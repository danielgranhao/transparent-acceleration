-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Ksnf5J5spyQtg3UEzsBmTBDujde8cxRs4Xv/oNqWsUbvc/xmOzU3vLQofn36Sx2q
xyf381+PnyWbgBHZLvo9f6+iptnm882CG3kpOHeDOgaah2jqwHn9sJDRTYP0P6NB
IwkgBCt4uneyz3GyUrf0ZnO/3Z7EPzCExwGgdsEoCEI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5186)

`protect DATA_BLOCK
lC06EFqknrhFyGhWyZQli4NLgDa762MYq/MBHpfQ0FA351B9eiB0+FXS5yhnN+5n
pg2b9rOPJw+U8nngXCOD7rea2EzPRtrfms0+RNzVw4Q6iwN+g7afTfBh7A1665oS
4AaDy7Xi7X7oS3YDVOxlj4kaCpVk6fDE9qGjeZpzfryQd393XOq4zsmNz/OcknLi
XyrmrojiEQRYvLmDeyVH4xlly76yWQGwzg1HR09gQXPuxz0OiHUbMw7Z0Ja841bf
4eNAvEqLPJEneWWyUjHBO4Cybe6asE0irYxKFTw2LLrdRov5thPUw/YOyBzU9By9
cDinn9uKOCRj6AjidevXIDr6P7GvZLUWQzrAoOGiA7jG1MkpDlj0GpLl6ZvvwiLA
ezh3zKtMU5+blIBF+MSG36XHCN8BDwfZRbg5hPhDfCpahu9yHAZEQTPJ8jQPqD3C
Ol50gO3mSYWQqZ2jn2GLlj7zNnFJYGKF7jpQS3LBo+wXwI0aXZXec8Yz6SXBR9Ca
tWJXlFRbVyDyGAEG5KjDKzQZ/VAYdF5SysHwmky/xWzciXJeFx7cBoBdYkOMF7m5
O2luFR8frh3N2viGO9H8B210Eq3Caz0+pydbkmAvl5IFubOywa8nsoYWUoEYRS8X
8po+dyP8wVgYEbTWudyDyw0WsBGXAaOQyj3JsxxuBOmIGoJ+qZamkDwes09YZbaA
ezEueUAGMhIOBi0aOoKTXfFydAJLAj+NFs2Ad2bvcuVKSjs54WLQcl4Oq1sb5TDe
j8NOsbrl4EAdlh+tu3T0BSqoUORPwIswdSpaNDnTTg+4CTRO0m2MPShNupWhaAoI
gsgFNf/iI+xiyTG1BR6NHQRnlRiYggYShg/FQYUYaK6+0TI0Fp1nW+1SlP5ntUxB
/n5rAKQemNvwOS4ijS4Ubzl4cayRx/zA7sM49jF6d7ZWuhiTNJhMnf87dNyUbi0f
/FdCotKsum+AfGQ2xHxEr8q1iDvvVoK/9GUBBHH1+6UAvP1wBnCfca2sETBQGe03
COj5bF9ugjWMtbAAGe/EZBm48sIY8Noy118ZgV+Ok85dE3MEpXphBJhQyx2SR4Jk
/84oX6wzVqPDYa0euLRIWYLxysBp9vKBsfZd9uU12TxCjib2JETmNgQlzqMJG6Wi
FsPCpFvh2lCBywww/HXYX13S5ZudlqOwQZRdrA1gdY6v03KuvpSqazdOqndBxHUt
0dMsiJ8UXPbC9yOCPNn+y0fvB0SeSMbzHBfZPE6I36rfNLQptuxeAfYL99UzVjYY
n40W3jLKDrvg39GZ+rAU3OfsbnivrOd0/zma1se4cXXh1gu21JTcuU7bqvP+TOZi
ozj7fTnQ5+aynsxCnMqP30Xq1/jywf3aA6zhrn9k4yzOJ0G5IJLh6hkTMzH4uaqz
Rh/grvJzDnlAlKIWoXu10CIkX3WZNL0MchFupxddwllDfy8QR/7z2lcs5d4lmh1u
smw7NxHTevSQ15l0s25SGuWbEEzWGo8z3fwMdAMir8eM4ow2tMSMK8Q1W8OaEMV6
mJd9JJhc0UnAnYaZEAMf5gygW+MJEEGVfoRuqo4awbzd7u5/elCcCVjZKpOR4MHI
KO1GcOV169xLivu9BxQ6N1KwYdQgJPdaWLK/HGGQoPrwIj29O9VeQVBCV3wmeUzI
TfJ5hHQn75CJLcBXWHKM9UoRkZ3cVhNjRGbQqD0KcZtVzWF58e2U6/O+g+/3ZQEU
/BtuUInBaMDMpUaeFWGGsAhRUr1NctjyFa2jbCBQpMYQ9PsAuwOBs2LesS9OFb3y
gI21zZPAYqjuFfHtPuH8uPMMHuSdd0Os0HHPs0Jh5BvHfTACe4KKvCN4cTLMiSyJ
9/PP3R1dcmS09eWj7jLAwnEox6aB4oPIANshKIJERz4rWY80XIG1uAU1JSxD0CJQ
gJVv1FHn5FFVKHk0Y4WGyZkJgi7HwfZcuzuDUaa7P2UnL3s3FJJKFPzLddTVQbeq
8KOfnUw8J+Z+W6CoxC0cf7GGQyJAZdcPxh/fkRoH9rLHrKt49WC+svZSpIrU74Dq
Z0elmlsVqqpRQt6fHNSBJ+5dJNHbT4jHlAeqqv714Pkxbvub05QW72gu6jwzryfu
0Q1evN3K90IQnPEC3ZEGdraNlYUx7GjJBY0UJgoxQ0knKRBMnopRMoQecohnn+Nb
ItpfKAJdOtiyTffPwD0EK84Amq1AzjvvkI9QQ7/pGUFymZH8xx+Gs6Pitk+JvoOg
sfwhWw0YqnvHvuSOPoe5l1rn75PWZ3LdnJKUhM+6kBcE/jcD39Mm845B6nhpl5Xv
Xd0JgUliuDsbTO+1pRoJml+Kgbhe93m9ASZnshUyRSuc8xIeQu12+ALV1BbrlSY7
SHxg4FpFTgchXdPGpHU1O15d9M/0me7TVzpzfDDnUSoGU+BT//xH6M6PltmHeUBR
rZL/Ilxxpnz5S+hg0XjC3DgR0lo4XB3U2FdferPIOrEieW2Ml+ZXbfsL+gbB/+g3
Kr1+aTzM1pSHZfrP4q19MvNki0eFy8O7OWGGoBtGQrUgjpIBdg8VJ5GOc+LrrGA/
OjOdz0jf16RY88/S16IPXbzWwnfJRF6SexonXWTNPreUkMEv1spew8HDBNd8wEtW
R9tF0Kip0Zbsqw8tiz1VLcACc52Vg8M/eCUZ3j9Q15vkRI8hgUHctfFdyVzB2yLx
zZPBweoIrm43253KCdJ5diSU3fGbkqKR0Chl4RE2Xf3Jipnnf9Zx/bXKtODylVXn
9gWnf2zP2IwWB4drzbSnHVl5suwUBe17xOf8Mwl6J5AxJrvyEWaXdqrXBgb88ZY8
FJzkbd9EePHRDhkvmJeApkQIWW0d0oNVjh9NqWOHaDTTiEAzan3R0AXadYUqoVgi
yqq82WqzcPM7kWK/olj7xYECsjyPihpCOepf4VaTCgjG1DrSBJs3EZxAtwUkqPVP
CKIngQbigmATcV4ZStRisU9VYtp4Se4WQ1M5A0wmeD804h2RTt1iltupKiRVw1SY
sr+ZU8yItxu/bJvklQFnBslYu4+XCDKMkNF9GdL3LFvj/Tqt6j/YfXUOy2aHViZB
IODKn10rlKew6Ua+4c/Ci1wCw1Z2PDvXtK67BdjQN66c8dG17j/s/AEMw67hlFWB
0Gv2qdN8OWU/Xdhe6qiJ9AzNeOJ8CdhHbzGnLfCJWwaBl+5RG5a+qwcDjjK8YKR7
v6/DDpATMOWqh3jmRdAdv1fMvJIAj11pPgLJaPx7ggksmc9bq8GiGNa9JnqZ0Xzh
YcWsCTGh1O6K0E8NaKgezX66LF4TS6hP48L2pKFQRqu8zqUwVdrXqCUS/4qLoeyV
b/Subt2gUi9Yq/mMUH7ZPx/PkfxBA078+gVPUZaCIwpCXdeK5qyd20M1NNbAQLLm
xYbiuT8RACkJSQfrRBY6CDEBFULRAxYnQNlziDKsEqcoG5+ghaXy/3Yw+odOzYEz
e7jJYoCs/V1O8Hip3mHvQNBeUWTOXRBXDZgk2fRetdQcWNW1TATTCjDeoRscsA17
NmSb2GzvSUhmJ4JG9CFfeIm1zazPsyuyhdlds54biGDcEHemhSBQ8JGM6aI8u6Fl
s+tKoHkcmPZdLHug83S0nWOfmHHJgcCoVeWkPWVzm4w85Zgj+V528LIoTLJLGQhz
XiRk8Q1abPK2ar1eTb+SVsK6QHzF/5FZd2VNy0iqVIKRGWJxsX/32xMlOgW2fTig
Axg07i3QYAI4KDv4vWGAXVCAA67AZZ+U+Frok+i01ExH9TXNZn2wbF0ZplAP2yot
+FDowveXkhd02UsXvR9zoHkpvGeRbt5bAWDt5eRMQWRAvnHj4CidGiFCaZmMm5KM
8IcEc/D4cucR5a36klDbfcn1wjxUpnqSjr0VADh5uGGgX75//e5BiZH9oqBj7n1m
UwfeVSqz5R9zN/qjPjDK8eGp4ReINQiAkwtRWeXKI2z6n5QDz9cxk03Hf1iD6E9F
69xdGszsK9SVTXZ5uOyGOA1P6lBx7ngBhKwJROT0w1+JGecuPyldk0XF0/mUeoK6
IRznD44Mj6JnTvKUbzFkbJu5Jn/8V2O7o9uCXCXXshW6tk373aokaEv0xloPJeAh
nbqDmv3UwmL9qTuTPGGqd15zuSzqg3UdZ8ErcPISWYjmVVvwBg9kHGhqRBZ492GD
7O3PALHpAuIwJVNhnsYfm1SBI0BkKudboVKG9frBVgc/nxeGEH+FLaJLyunmZxsw
2VliTcRQ2ZVQqLXQbCTgQEg8cpDcpz4U/0NFO0Wnkh7IJt+z97LoWwUDdW/Fh7u6
7SEaqfGsQy5y+vkM+Z0vemQ2SK8RKzQf5++gGIY/hASFS/cLR3VK5Ih6U+iWuDFP
C6HelzqaCr6cBYB8i9hZZXVnE9iQMkWgVUcJUcCkAHVw4SZkj0RYNHfqesZkKtqM
VM78FTjzjxrqRBBmKG57cYFvKtuHbkWneZy/cXf5Wx4ulKN+xL/tckooJ5tQQiXe
RA+6aAYkkh6z2K5Db3ohmff9dzxDgzbajpTpDM7AP/AigCZCZ0O4IuhUrGLIYcrV
JmRe/DLGdyk/0Fotk+2791nqCrjqsidzJt0/St5C3TWchjbL+ai9OkxnxMKsh6cq
qdHlYZfr/+6F2hvKKZ6lQY8bGtu+7MJ6piAxLGSqSUhiDAY86uO6LjYCP0eaV4IB
rpQoJwN//h5ZRZRJaYS7ElWh6QGNXg7q/4ody/BxbxDDXaD55IepRuIioZh1vtW3
5Rnh1WcSKTcJgJGcFZJmyFj5MhmG6q9Bx6lISMQqHkPg/saObwuaFD2suDZYkmz0
3vHMoHRYUK1lNe5lWEdquPZ9Ojb85HJiw4oWUpQbNTpX4byBUPlrRpUIyaxgsVgR
Jw4Y1gmZjEa07hQWhY/L6BkyobDP4X2+AR86fJikzLG9fk4zqZd4wywd0+8pjuQW
Auzbu/25OwOoerkFXigRSWe6lV8oQ+V11t6d6tRlucm0PpbKSKaG5b703Zpu2FFN
9iyOJgy/K3ZxCh1IA1XZlQMoV9KgYYmhi9Cz3Wv97fGu13ocz8k4HMB0TB99al7r
Z9UMS6OJjMVtXecy+8GbVQv+ACTOEhWHyz2+PV5tvxCpKVFv33juaewrlfieqUzA
UqJnLzTGGSu2DrtPFggBLftzFyFWdjnD77levbEKKUOtR2blHXjGqbSqsvE4AtkL
HEoqBmXLryhdcNtIzt9eGNzybGlX4+7pcrBggXkLel5CR8icnkj7zxYwvMs4B3if
dhKAMkryl3JWDIm492Kvp/vq4C24+1k1z/HYE98b+QxnnGuZ3EiESI6KT/ZYAnpV
ytIXwml6sx0SN6+ESQ5FxN7gP9mbWJNnFpP5UcSsUjDZSGaezqF7EdT0prJwMwOP
lK1+Qzl3bqjVHW1nYXkxKa3SSdfOMQka3Lo0V9UDQ5aX3sGkazv7VTsLJaVt2bOO
uGMBuJc0DTy57svcltMCp0ygWuiH1vLy64mfC6c9hO6bj6UvNhBFRTv5QKdTzxyc
ejAbITMfhSeLQ1yECyPPjOlPrjMxuLw7kvnQTAJnDZ31t7TDCMWVENVU+YiR3+fh
2kw6mkFS5062pP9NjENWc1Q36icZlT8VyB7ZSzovNKH1St+C6S0jf7Vn8ofOhmMW
svBEfJ0UrjrkCj9CMetzHebmYw8swc0OIqFZgHgv+yIl5L1lLS5rSJLZg5Pftgc8
b8DFziQxph56OFIjVKpe1DJPJTcobuuOWVOOFOc7tnLFCLuNJCq+7nLXFxy4hrsY
vTrBlwxGXrHc4tjJ8OHUk+xunFptxbFuIgkS4ujCJa6mPoQGVw7oMb+BVUyS3Bl5
xEDuafe0ek+PKlMQeQfWkaAj3V5osthrS6ahGQOmQx2FwEHo1FOrdRqpBUdxHJxh
VPpIbF/KkzqciOJzXkTUueODDnpIoXr83doOYxxVK9BRrKEF6I7cz+V6aELiOBx0
NUztLCu8GEfQzCF7SjpGBP9pBm2UH8AvUIa6VDaFvgO84PIaviLx21df7vAxbIZp
oElRFVGnicOqaY/t9rnfXulYNtYVCb8Oz6heaA0ZC6U8xPYAkd6vu571cJSP0xqc
hP6z52amVoaXFZH4M0DtY5GqynD4ahiO5oUGEvO7EGVVGjjtq9cTt+DIDWhlQ6iX
Cg80JtBxoebh9s4HpG+ys1/vTrvD52xrgcUxv3Eh+ZP933iwJ2BMEsNlr3PIRLiq
x0xc53QrO/wZ72gLNeXCqrzm6DtbpbCYkFUN688vXt5M7R48OqV25QnHGsGll6Qh
A80GANqR8PvbwRX1swF/UjfRaavm0ZF8qmVdaqhGtVQk7fV8MUCIJ4s9hWLTF3Oe
7ZujYCJy8QX1caePjJc06EfXCZWuywLJnWnMeviM6ie+0nhJizuYp8UA/nNPlA9L
o2VD7o3lW9GfIxDuWhmTH588KEUPAV0n80NyPtRt+eMV/3Wdz6YBlRUg3Lx0AEeI
FKPByVOUKwjYK8fb4yhjaBq7GpRRUsGFkgwW+PeshB7wJyHvrck1BFCHZlyIC762
yuVSL8p7gFJZY1qMmO3nTb/urFdc1T740pOg2ChE/N+5PANSkyVXOpizbJmt51is
H11uTsx5HGmrVMkXK6EB1pcKPzbuGcfCP4MnK1ku4iIn10b91Gi+eaAm1Ap5dvyx
0AwUf0kNzwUDpZhr0+72aqP9k/Gw/baiwb7jUujF6piHhl6YDTBD5Ou+c0zMWjbh
AWA3NIOf69L4czL5l4FoTK5rf5NG7uCP4wch7z+iwrlJHOxWthId0V0xO+UdMyC9
62DLWFv4xRk8zrqCr97x7eM1X+R6bUzUeqy7T5p+xOZ6z5gwLIClilO1GmM7j5Tk
t3Q03qFUcISeqCo75Ct7uW2t5gFLPyviIN+gFluAmU+d5F8AQGzAIM1/ZdvNKnx6
gSzzVryYNaxZRM3mPXvpuaoWVKeld/wcZsamYMfQmIo=
`protect END_PROTECTED