-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
nEF7NRpuxZWv+rTV4ne7OExVkerydx5d7ui2uPy26kyKv1TPiS5VelJE8eIKZDmO
oNJ4ajKD7JkfgOlI2HwaM+Bx7aj0tnW0ZiR6cOce/l3IAjysSr7G5L+I2P6aDdcU
fg3FQnJ3yNGIGMgE+5O25K3lhpBdSlChfO5y1NBLpvI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8848)
`protect data_block
WWYV8PkrTY0OyP1VXa+t+S6g8nY95WMsk2w725TtRndE1+xyPHwmLzfq1IGJzqqk
xexbYWIMUz4P0udoOYBCM56cXCPZR3/raEu5O5f2mL6LuIFU8d8xLIQ0e/Oeic/z
8ysP18QSJzT/+Zj0Tn9ilBk/krUhC3U/DGRpBffyX/QMM1Wf9JWl5ca76VotR62D
AoqTUmKha4iMyJho3XKg34aU9cdQUzGip+L9fWWvdHQa4yZ+qbUInEfEa7+KM8m6
elxaWWqs0KPR3Qja06DxQK023EiPjQShMRATKhmkdfKVEZ2XDSStEiL2bcsrou7v
3eG4hywS8pUJeCnXYEBLMfaO8XhOlPkLj0dN45JfuPrEDEDQqrpfAmy05YwCXgku
HgrOJ/mqDPfK4o6BzZO+0nZgOlKq87tyWs+Ez93oI0M1seLWgsT+ke+inSyF9f5v
JA2ppTrEhXPiSknPf99L7YbqJsS9be1swOIOWt/W01Dfy71HwdAXinJU1v/T1+QA
6NTKc7BzuzmiLfwCtml2RPWKve4urcTnDSsMdOooNLU8ZeFpnt7y14oIeD2lWj/t
Nuin4U6jijwYbFqfXUfTWMW01bbQwJ0rmCYMS1pYitxn7wl9p9/ieeoXw+6o01VE
xcXFIzHAiTXA4af4VAeh4Zx6Ht80eVdS9HUYKgFkiAsldTqPdG7S3TbZM4VjzRi+
VfvYPFDinVY7pNtyBoPiy/bABnppAiDU6dbZF27gmV8sDLbWT0wwca+oiF3gBXh0
lbGKtp9FBrmzJWfBpX2ylGTzkTAZ0mMA0XSm+8VUW/Z2uDQhnRjKoImYa+4qmUVA
CjgBq5XqHDfCKetGBYxhK/cvCSMTOCY6IFWhacF9nWVMj75VuqQpyz8DBrx+v4io
PMqGSNWtIuiyW3CSi9LChsegLsik97VB7OZtM+T6p7rffs1HuuJMAjL4tQpkx1ih
49KGxrfEEChS3HeY4WCBupMiu0H0tiD2f5gJKuqmT+UFBoGF0CUw/fa05c/6A8Ct
CN/akOTjLuXKLlCVUbsEs2uyKxjdqSfnocVRCjlY2axCd8PePIuUGbgKTUE90VXa
x1ubfSayRtonZHOsGlWA4npUREk/Nnqf43IQyevy03n+6B8WBs9FZpGrzZAhbqFs
ezAryNrFE1ocVgWbzT6y4iQu9Mj3k5AMwqGHDy7OUGHS/XKHsCcnIMjEe0dBEwWn
zxOod8tK/Mjoo4M95z6Nxdc1hx9DuTDW3TmSTfAqvZ9mCC9ZFfnJ14hSzrWXkLWx
X0ATiyB1v7E8yLiIUjUArgBj2i1rAfPqKmJL0iVWO0zk5/sfY+b/PjVgZosadcKA
UJXHhGIBm6IBvKP7qVmR3TCpiEMXw0hnU69qV1OIMKjT7yuSzL0PUUjEG8rkOBRd
CNs8IzGY0T7M/danlvDJLHWScGQb5u25Y5FrRXVPStjdPwdQee74dGAMie/YVYsw
xrXdY4rrHbt9Oq/yUngPyvgNwg+vS4dCftkFPTcBS1RuBBqQQkUQM+BmscHZjHVn
8NV5VfPkL1vn7EP6MnGwu4+53LkvPkwt9ydfIV7nYIlB1vX4OLm5u1v9jhz5VPtn
VCI8mAfHXv94M98yUMRJX7F/UyGt27+L4uDJmzFNdoN0ENNVXOh23Ttv9x771SFx
LMI/1htwHNXIdioIy+eJSWU/N1jgUMeFDmhJ+FBSX2lLIW2rruYyxnuEIsWWp3GN
eSdg5WgXyGohIv87HTsOfO13aY1bQ7FFY8FphpOz2vWFJbMT/RYt+RAdxbeMQjTz
WQ8wkoBMCTsILlVEH05kfenCrnx6hxk2PYQReIgta2VmbV7c4vzyrRJK3sHo7Qln
47u1EwSwOoyTWu1arAl2AuHT6JX3mavLGdzcQ4Y8xgpT0hv2rW3xRLy2gKU8kzGZ
FZNe/W2/UQru3RGDeJdvFej56R5gEexPbMr3Fsa3WAtmiWyR1Mk2Zb14nquKGTmm
8g8MDjtRZnyPSXf+x4q9ds0nktwPJ13c/8/vEJIZQ8uhihkOdgZO1Rp8J949IbpI
v8jMo7F9HJwwYLzFlQIlOgzR2264fzaT91Z8oq2vhmbpbAYK8zxmdCuGiw6MOYrT
gcsROe0bTMuosGfkNPZr25pGKrofjoW/Iq6PvLxmgsETShPGFRgvyM6tEPJ/kXWb
4OqwKUZJam0r4rOkf+H04YfF3Ib9B72Jw2dwexL0lQHJBKP0WouMWLAL2HIPTqe8
2wG8sMoO91o5TOC4nhmLfP47yXucBiKEMLTGIYiwSXV20XbhKsc6nN/mzC266pfO
CkGWZDX91YSXdrH4Ma0VB2DRwOFXI2S5hhypuJed0tnB9smHlAyobDvgstc7udyh
8ZN+4QR7G5rRty29BwZx4ERrqYWTSL8bv2cVDqzTFLIL8nSGPJxbIKLv+rnWt02a
2LGDfGudEummaLCZTejwIl/f/CXgeq8cxZMrRp8DB6PowkVnUQd+e5APTCGsl672
jFmSjVceawqWv4Q3B9t9yWQLXiK7lyDBio6PHj1wiL/yQv4wUz/h24T9mOYW+7T3
giCJUc7ORpIfeMObAMeL9gUd2veMiCPu3aD/bVrSaBhUhGBXP2Hg9XqmuYR9WKZE
1DviBaKyX8OCIpLpdNWwBjlr/5A9YDNMVXDZA0ceX0LfIk39kIKMjQlNCJo2YuSb
mxAE/sp6vJRrriLUduxpFyKFiMOdOeX1BjiH35X3HZ1OQKPAPbY4hEsZyohDabId
Q1rWhwYmDpv40sYwnoGNzma84rjye6ovSG2+VInaEFVhXgrPG6XKtGBidzzSR9oG
RWGDeSJLw1qN7q/CApf8mEOdMf22yQTyhu08/T5JTW/88iSO6wz04bxCwN0Pz2to
74mbMxB7aZ9yn40wLhTM0Haj0CbJw04e8xgQkEyD3weTzFWQNZje9CgHofZBy2oN
RBEAxkkkW1DD7veOKknK9w0B1f1qxQGvKXjUmBg8aJX2rtBfjqDuxBz9sUwr6YQE
HBjPnvSpJl8jUC2RlRh5MGX2Bc0xYlAMw2GFOimZEMLO8oJrScBr3BJ81Ahve88q
tHaYUgbg1M3woSRqwJewWZCvY+01TYP+b9G+QXoz0d5L/MCQTajnc78IwrnixRFq
CdarCk54xdKiWX5XklOXLaY91raDRbkiOiMHP3U0sRNi8bIVnO1x8EMJtEgyKb8F
cIBrYGlg9lHMqI4PvEoBppik3c8iNqw1dRJkuCMTZOKhQ0n2YNq8ZkwNteL4B2AP
RBNKUlmqeegHNAA8s2TXqMFoVWhGLQagr2sZtKYGoUNz77PJArMCfJhdlPuXTB6N
AIMIZflCRKEUPu25FRaHT4IMn8jZqzRIG5oPU5qW6nXynl9YEjKGpRKnOZPKnHKl
QU822xzJURvewUP6vazQYA/+dlh+aOLsPbdZ8P6UzW4QceO+/PZ/0zVvQs5LyBe/
8jXoJ8yHmzM/hmvmTu2adXuFuAmdoS77CVwcfapiOEEMbTFjvyiz0HfsbGOz5jPh
+jen3KvV56IJe0Jc/WH8gZIJ3w83NyKBdGE56EM1uPoZT1ZKAF0suKx8gKq6NY/v
TiZg4oTDR1kKGjMbjnHc3nEZJUgsWJnpewLAtXwoIdvGu47oCwpzBdyq41aoc1Mq
jwJzhc3dtMJosDJqnvCSFBe4/nnLpM2T2QfiTvSR0i5mlAkP/o2Ol3oxXV8ZCkbk
GYtmdy2hBm0S/Y4J/1zK1S8SjYGeVpJfA3U9FiuUS7mcMIRGbacTb/uFlLmuq6kj
+aoWvCVBcl/+k+rKsNUduPWXfE55Ry63e7bXPQ+dWGo7AXNM98KA7wTSVyPfMEMR
q6y1R4zDjqAI99SF/MXaUhFEYhcuifFfLHV94kH4+tsBDZWFYmih/6B8VPBwuRRb
LYTbJlbFzCMKQRx24muPpiu0KlZ2j3/9qOHW/0prtqkY7R/te7KydsiZ7VCiX53u
0gYs8uFdtYxyBkQvqRowN97R7A1ltHZiOVA/rLnXiotMUURtgAykTR0mL/VI2rCm
ox1FKrBRvwi3YN/oQQAHsgqh795zcG6/z69qSrzgTg5XPQo39EMPGGdRc0mtBzQ3
uQ4469+nuQuMcOH/xpRFTihuaEditNwRcDvS80NuNDNoVmJxCkvrkMYrHnXsi073
thqLDaxJ3SI6+AK7acSKiHfsx7R3ICobgDdESjz62U7P2aFetpeo5MH3LOxAmCNJ
ZWvyP50gk5L5gErWBbyZhrDn1yLTKOcVQzmgtWYRWj9RGoeplGkzihVcmb4enDkl
UrMA1qRmSpeLLbjqeleezlas95X33sJUGJObEXPIezXpZutU9YBiGHokVdmfyFZ5
gMPVoanj4hyjuSD8HSoJvpS5RtEBR0Vr74s9pWV83Pi/09aEAmA7ihgTTS1uIJA9
8HAEPKCweXUw9b6XMP/4LaxXc454J13s0NGe2vJ46lJ/w/vmjzc7s4HU91ANWpYb
EmZkKra2Esfn31BKhVLUe9dFo/qTLmHQFrPliYJFqx5Vj+4NVKK/g/JTFXNt0hdc
LLEWbHNYt9/yAni1bbyMGocUnr7vYrA60SMfFPui5l+mQfV3quK2lGAj+1pURX0T
gH+VnK9ALy8KyjNkJ25mqlqstTypZla+zkftjPDqALKtzsftBHTw1pKBJFDjvh86
1t/mgud+m8vyoI+MBBCD5QxfpagPRJ67U675XcNksl4AIBUsXHsO4wzGCeQ2kaYG
2Gf0t//8TEnpW+w36mzBv7o6JoNJGzvUnUUs0YfVMNjdEWBYjw0vAtRBmuiJMHtl
kjomsSZROzWBNaV5U9lVdx8DsEl4Jq4TBAe7iQxCka2X8JkpeD0lxVK/yoMxrt2J
qkDxlhfFUeXWmH7sSf+RWaYERnJyLJOL7YI0C/XkXmFy6TWLbJeyqp89WoknuRMC
gsvXZURLdKQ+SqUtiVXR7PrZLZFa34QredZVB1RqPxkkQg6sTC6nFwfwNyX7sm6Q
yGjFqNufS2Y4IEd1JQI/PDrUcxqA73lcJCMdeFhSr0v0lUGGXs/yjREIs89V5GbC
1L7Ksxc7OBxo2BNGF3u4QkR75t4tkhEMVVK8FPbCsZqtKyJViOVoMIZzWLTVcnEc
f7SmsEnzSmdxCHXLlQDj1lp/T3PKr6L2L7TlwOa7OBZiSYmKnn2HacjYZll2ZXCN
7DDzxj92OgNGropn60MHkPNQvXunwstT4aF+sg7OhI5Bq+MWngHpQGFmQNuHmHGf
daye0i6QW0o64rceKWHUt4HHEyDjCizYd/hHh8pgt9qU+hh2DB+MHye4JCG660+O
RbBuQpGhZitd7U0fBLfxqjjHm9ZUzRgcyjV3YBjbm/4eTBQb6yFqdnihp8sYMKQw
0jGrcVU0UC78n+NITAZ2EAzLeZL7GiymjTczMtYC2Rqxl0uSIKL2bYUCiehEXZXG
ZrRx1wC/rHBj5+FM/+ICx+0nW0JCS1cgVldShPnWXyr5rCSUEWurIdY5q7AkLxjn
vdjyP12gSU5iVsWf9NUtlDuJfgiI4NfLogiHoDWz/kxYkDP5c9KYWIeeuII1y1Mu
OdboM8O6B45HlUVgoYuvE01qzrlDSmsCy9knJL5F1MInV1YcaNkCIdq/Q1qt0wv6
h0rk3rUyor3NR/i7kF16oY1wiTULckcT44rjsG8VyD4c7YGbIfSOUM06mRk66r+T
YYNGP2yUpu9pQIHwA9CHr6jGu+qPxGxtMfPW30WNt7+VG1NVHM19Tsjhxf5jw1ge
Cjeu8wzXpwi1NNHJ6rEPd92x1LnC/4E+ugigE1LjUG26UC1TK2QvU5NIqdDq1qw8
7lFtCTgGTEnqOcKA06LrkeNQrvebVUuT+jeNY3KbRrltkO6QAPQyoRgGGU853Sjx
dh1/ub+IV75soXZHxr6B2iefqoYBXjnwoUd+zCAEhvm4QtG0p40j0XaERGAN7g+b
D2OfCcoZwWNWg10J41UeCXBx9wgLSGj3StZbKEzgK/Z1O2KCa7y3m/LMXdNzqzSh
ySWYl6q1k6PrBftwnt1kNBSzGFvO6BGfG2L2pja/lWOMa/68sc0ed9pVOUHZFhRK
rKCFrTIyUYWzya7y+0inCMHVRqWVFHTJiv7VADZYN9jPCauaqKzD6YIbWIPMm3NT
/jPT727xxoHsbfq5YLF1WbE75L9lxLZwrywTSBrgEAW6t/T5UBeoHghSk88j2xOm
RY9cJi+l7qXlqtL5mfHEsm6M66DTXAe7Xh0jKTsoaouKXZE2ZUBj/7ILFKlL98Xq
xRb3vRxhqq7Nuypf8WHHAMuLWjQWVJHHce9U81avHnQHTddT8ZHpGE7RBgo8iq7i
xQM0slf1E0lXt0N6fEEYzuu84aDSQxiPpBKhjxVwsFBK8Z9dmE4xPNS/nGmxzu7X
zGEfcrLPtd48u/v50VOMtycPymAEy+FN2zthh+JcJPrUK3+d7+w0z4ExsNvUoC8F
ha0T+iy3fqf3ceGDIbtNOwTppWMpLSZNz2Ts9p/R9duXVnOqHJ8yTpvBubILgUJz
pkcq4ynRVoEv4ayzfhReC7ldxb2iHg+xF33RzLfwQf5slCvrktqmKbDmzjct1Qar
xMhliUzAYWAMNhL6L+aZDZ91Uk7Nq4vDdT7ePuDLBW719E0orrc/2j3dZlug7Las
WT7e1IPwPrryhls8OYsGGyzLZaGgQ1xydREblI29+uQaWSdFy+6x0ko4zFsW8ru0
0CKFSGq1itMLVaULabLxVBOCCeAtb/np9Bnx/6jz3cpTW9vvZ6VXODD/kc1lsUQ1
/jNU9amlfaPNgPCz6SFY+GqxNQdqtzxynuyv+w4Fcfqnu48X5f8LvUXEu6Et0im7
4kAjhz93IfDUVW8crxQYrRxQ3inlte2KQQCu0qGGLcMxeBgAjvkc6GRwrUYjlXO/
GOXOlc8g4SB0cOnKoH9pPN8B0EeCkqOH8NN2jiFGppRfqCOtflUvIGa08WouBp6m
COx5RZT1OzCl1ElsIRF2HYcqnsRXJcR9NLJCA0TLLe7CYo47a2BAT7XJ7VQ83Pye
dyBM8xvWvG3pwyFtIzNTAQrXPPb6ZRpmyRf67lJa9JtyPfPt7NGnP7eWC7ZZwL5U
z4L3llDF2BrSgA9o3LzrM0zg9waMOFNGXsH1lsJwX4jt+3KrZkzHOaoG2Sg/Z8+J
95t160Qsf1bZUtnngOYiYQEiPz2rvt5Ic9rPe/gNzy0LtAQ44qmXOkHlOkQ8ydAk
kackYt/gAlTIZksrYOBQz5b1+IZQBloQVURhkBakLWgc3wyPR7WIOB+Eep5uhsHs
gejYBN2bpKQgFZsxCZfyn32ElNX+frTfVjyjmKEpMXhl8XIDlXkd1cDX+rFr9zae
SLZFwviR/eAQbBSxhT7h6M6Gxxgpb9OZvV5rQs2AHibYKpRgMphZjyTGUVoTy5HI
6hrKM+y3nryj9c02nclMKdNDpAMpckYFj3OJB+Fn9t9G4FY+5Bpi2MUUl/FTA5Gf
hvNcK11ZJeWwei4zOEOAx47qElo8piEN82rz2TfXSzIKPbOo61liB4j/8LWCCNC0
sWYkNIa9fvoBS5eS8dwK9DTBlqGCenraqQWv3l+bWR0mRQwHp8wAq0OyTOx0d16D
Zuo+N5nOqo+kJ6rg1lcnv0gM3md109J4rHH2DLZJYuMVvB5hKrv2Z0CoiSV/LttD
nrkwcEY5QplwKuZQoaazD7fjoIdCOgHBRVkgegtGO8qo0LkSjDs5VKBIkX5Xb8lM
X/qmgBIQnSbmJ8hyWpkIAXMpOfSLN2uGnQQc/R5GPvneLu8MFqpXtui8lq+Bqakc
85cwXLUe7l548EeL+xOBEE41OE/IfSVpDkNrBIZK+r7wNZdjYsEtiSKmzTezqDoc
sEJwlWKt77mCEcIUOAPmjXPUJ4wMHZ1iub7suCWHpPtxE3C7wZ4LOfgGJO+toOsh
DVadIlNBJq+wHShKFhldfn6vFTiYPd6MuukV4lqqaWmnmx3PbFywU0XGpk20dADU
LWIRwiv7DHbwtq2ur8B+QPunuysh6JM81oBXagxHljhVHUvGRoKwdKAPsRCFt+E3
RNMYTG8O9KcxNgKkG4KZz/y5YfiSkxExagTHd/9UlAPlMgVNt6jgNZIEkyxbDYf2
iXNETGRp0JQqVRe58WpMse44RUBGlst5F/L2EQ9LmUbW14s6LWhnZGlvC+CY1S+t
W9eR3aLXJRVG4XNbPFOjJwbWFi4hmES6YqrB+eQcmx3LI+ARgxJiTXeTunJw69l2
N5YeaaUA4NIAeEjo4n0Se6YtZ0vsja1RSz9ck2XRLUplIPU/rphTuS2M0lLC0y91
e7y6AligDzp2gI0P1rkJrAVEpA7gSJ8EthYCwub5vXtu7j9d3SdOWuZUluxs67Hq
AlxY9FKbsKGBYOBmqYwuXRY+AQqUdQYi8GnAITum0B2VzPbqrx16aAAeJRixsoCL
KwAzKVeOnV+7yqBJhKzEC778ZkLuj+ez54EE3Z01TuNYTWKu8lF8B23ZpDS38t5e
2TmGX/Q7f9RGlCRNTgKn03fkh93HQHJvjqhYjnVgFhB01OKjcHaUf0Pq7yuyrV1A
9vD2E+owWminQzOl3lDqey5eMTlmDJMUW8PifpIBVoEL+/AbcG97wRXE+jciMNVd
CEbZXwoitpFmEJOpToeo3g2DakIYclYM+cOTOYpuKK9eUyAxU84693UGDDVG+NEc
/T+NnSnTgxkjm8GK08+GJqfqhOcZy0CnsiXrmOJUQszh6vCDKq4dEbFehZoBWQ1S
M/WPeqFN+fMTW7AvJIrBTewRfuKX+zQFcM2CYzgx6pPAqrdajnMcyxBbvTtQZ1PT
SJm5/Ifs2YMmujY4O2BkFHUK+KK+zRgz/6NYtkzhHLh/jLbE/7ZwetLsjkzG9SfV
ZZnWzbKYSbx5ajHByxLuEXuH8fdjxPuHg8+uGhECQ7Ss5iURfjiQJ1Atiy9skiY1
T0ifywEGOjxTlwlrlQNPzXvl/+kZaRqQGxfPcMxBVbZeIG7pI4sbHyoACuet/HAC
on1LwWTwqxFfvrUB1//Kv7fCAR1JqOJkPgG2iHH6El276sC+K1gXg4ba3BxIP2ba
4g/W29eE10jUF8qUXNUsbUNJsPOWFkiXOPFYXWbXAv8dKi+7wHTMLwB+qA2tEtXu
pERKDghSjG6UydY/s+YITUEPnkNEwtYGW0Dju7YkG0D5A7gFDLbnda2bWKJPgPIx
93neCKyhh+/hvXkrEjucL4TLeDfxPQGEgB4v50s78UrugKAjWAP2TCsIm462+AfO
zDaDOe89T4MRDIkPsjnERPe4rz22LXQbMjXSb/cWy0CnQBhX/89p9y5LFai3a9Mp
wuIhvA8y1iZUIb0OFrVo3Xg6qeibpwiBGdTPd8RRgVCBbWu90svIpJ6Xn+K2+WqK
ZKeRylpwiUUCc0lRZ5giKtLxlLGZHU6d6gd55S8oXLU3m2teMAjwBeFxSLz4vk2q
boamP480p6zfHUJQRuohIg+Q8MsNaRE6xfmU594EVvWqPDdGYInbr1eWKdxRGsnS
ggH8PBTO+6kBZ9rVVQZypIfnDQAyq61D4mbNbwyjGgX/Cc3gcIzDYJPOt03BtsvL
I5O3YBUnI9wLG1dINPLRNKm+ZN1afLxVVRezx0vWaM63AoFkXJjAD6Ts8wUEDr2Y
V9qgIZtl1+m5ndwzq8Lb6J6Rr17ME5vN9hRNDHPbXZVb7H7JZauOWdnjiVNVeCpY
qiB3tPTCZIW2Agewag/LAq8p1UVZRW7jeyTuF6drjntPyL49z2iwt8k4v06YNuew
FMnsqtDuTeGh5BKh3YPJvU6gkDcniOI0CPKMYgo/Ui/d8E0a/Bw0hI2AkRE/7hgd
/hDhKtKuetkK9JAc6Zro1b1r2IOIoh/FLzjbHKNFeMvx0wMkbOf3MHdAKkXQeexs
+Z6CXDf7I0BOGNWMize4ueeTTc1Mk8w1WxHgslH/iK9827JBtL4wdeVjBrBDmYkQ
NLj9xNosIlWjE1xLTzdJ0bmk3QswLQtXNG4paf808FihGZbEWOMkQLeJ+V5j760c
KhPGKi2s4uVjvHDasMR1fslyE3jfKNcICkRq7WYs9AB+Qscx+8FVMSlaw85CXidr
UyRzK09Vu9GIgf3KW/n9Cl7xAIwP02LPOkgSXYbpD1uPeEgVh4LLG33uL6JBlZ0t
sHDeEywpXAvd4rOPNe0TkakP7W1K7Ao+Sw3uwH2CbaoJcf2tZtqDipUR6SDtrRMA
WHW0owZZFxLJCYjApRsxQJfxi9seBqrcWb4hjo2QEGDdxHdNuvrJjZBqmfYkgTES
wyKPXeaTtB29BVRP4ydJzPtSnRSZo90n+7YM8pp0qTwt3dr8x1l6B8umUmHGouEA
f1eX4m+F4nBeftyeLugPkRzpghV/wzq2NvkFYIwfflV1lZCS91ynwLHnd4IDFALq
HfVi6z0MK41ljpSZZbcMq4SiJK8+kfjXkOjYzAeMaA4yBiQZIHa60QSsScBOd5kg
7c/TAiRHhD6Dt2AOhvwpJog6wxF+GV2+u4ZqQ6kpTsr5D9IVnRkyD96P9alVNx4+
CeCW82xJgLxkb58VQLVKQB4OaRpVR9/+KHnx1/CZvLS9kuSlkABqQbqw9T+IZr8I
Pn1uJzZt2jqxC1XrE6IN0cYRitfskEDvDlfj9SB9wcNlsysiZIpDSdT+EwaiHKHK
68Ci5ZTasIHEYya6Mb5od/1ScoqnD3MQvw3NnVhSwVa5f8olexwafnbmksgicYhm
NKevNIIxVITgMH6H/oaNj1TbBG2lUa6YQ4oRStZmUdxk1Q4q0L8854blytsDrVhS
HFPsyY9xXr3FN/H34lCzc+4pIinRWqWWsTmBqhzG1SOMjbKzZ97x9MscPOr2yTvh
+oJbRZDaWzo5VcNYzw/AAAbbbxYquhFWJtH0E8h3c/ahbR1JNSCszp5nFnrAhKc3
7RpZPyKdkfuAU0xcWYZNAT8TRxkMYkIKp4rN/o0ZZoYx/8JWveRcaz6+KnVj2px5
XOTvbYZt5O3N7ufTmxnpM+Dt5v+DIh3EOgZwgJemfJE4+u1MY+e66bNg0VkEZx5c
OCwRxAucIOPfnJgm3jzYqWcfXNXr7GeBscroPYHrKIoK4KoqBHF+ghmzILvsa6bM
2S0YdjFFITT//vtzoFymIPQztS0HgPjwTbQodDr0wYqHbUHKCV0FYemgWKcSkCHR
aDkHqZO+g5lbOtmdPDBruStjjuvwHS7LZ5GqOjR5F8xa7l/5xKR7/+tEU4OmKhQs
piGAExIlN/gvLdT1jP4FjwWTGI6lJtLa5xC9ZmsNFA3eNVV2aMrivuJsNZve3IE5
v64UNyED8AvbRPH92eaKarUz0pfu3UaiUhia0sT6NmXc8ih4bpUDaTSSGXhNbg+n
5+/gq6cEW2uSeI4kcEVLA0c5D8OHBXjuauCpcbnhi53VFJQu4GSyeXh/Xjdlz1Nh
s5Jup5frPtvXHI55MnQSlydtq81KKxa2OL9iRMLb8eZ93H6tSjJvSsEAM3NY/Jpx
ZrENH7IEUV8hTF2DJYPfLGKx96YeQoeAtZhN0zetifDVkbO9gq2KaC2vx+aake40
oUhCyUd42vUDxpLTiuLTjabaY6Li2+pLeAP/AgCg+XGy/hCdwn3918AV/KFMb9eU
1yW4R0VOvqI27PfC8RTw/jNFZO//xCjfiFlC/swWXfd4fYG6xrmB3mT3SDblgHmf
eQKy4Aj1zGZuvTjaCNxFF/njDFYHb8nPYN4aBM63j3mFPuZ/f9Um9lXJe3NsgRiH
Fm8IAK24FCHXx9utfXIMAQ==
`protect end_protected
