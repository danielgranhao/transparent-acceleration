-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Hs7/XheJtBwDMjfLaRcJKRNIlTR59VSal4vAFDAdvcXsy5dKsRjIcMCop+M9bw8qNpknrWPcngv1
qUOEMG9bxGiRYh8zjsZCWt1bjgxgGcZkkj9/R9nzOMwLWkvuaC3iNqOjIbp63h/7e01i+AKBMkVD
MnANdYrEkpwnrnBI+ce1YQSW4s6BC5jjF3VRIrUoFEuEDyrJhE2GXUKzHZDk/Y0BjO8TzXXNhgkc
KLoBQjVA12wUDt2hyVl2AgM8GrGjWVpcaL2DB1tLrr0gT7fIpRnNPmaGyjmGr6k/OlOhsEF62jlx
w7f2AjQJ5Y5rp1scxjzGSzl3S4nC0dzG6sv0Pg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4560)
`protect data_block
3tlkhj9sGtO8qhropUgrwDXAB+BEy7EpEOh5wEaHsZ6woLE9Y6AHjgac1H2NUv4VfSG16B8CPY27
U9ZpiXO5JI0EwIuJ5778jdpik7LrvJl5ktaFmk4Wx2t+h604Q2WpJnypqUg+APF+xajJAV2c/sCt
ulL/uLeZwr17D8WkJkUnssOF7rdjoR7bXzLXzWImVBBWfGbNbGO4wW3r06xLyiHU2zbJog2Z5Orv
9cuz2kaGiWNepYwDxg0auuB1pTiqzsguKrIhi1faQFZYdaT3hAh7v+5S+aWXL22E99YPCKqK1fOU
rGTVLPm7m/tSVA6wf5Hf4Gw5bIfV9FJY2TzD0ELQbDdwbONMde9rfC4isyet8Q6Yv78HlacxwfOr
SLVWzCfQ/+Oq8KLmK4/Q2QKe8aQ2gQDpM+ImDmAygysC9PSCrY2CAMPiN96qpdkPDMJHcb6rwtmw
pdnqicXHInKa6TfZwb+1IlSs6VovIN/pyX5Dbj59YRZ4m27kB4KjCuMuycanqPqYWVq97Jia6HHY
CJv2XyshyxBsX1vCKdR5vw6OB917mzqALYyxvgzEjJNZHSsEvKf9HSg5Yac/P08wrGYO2YFV83ek
TxVRiThPSBgFfyGrKJ8sl5Pi71F40nBndPWyh3grp2byx2GIDYcZYzZpgpU4x4Wxtz/Lb/nho2jF
C/O/hfMhA+4hxm40/kvkrLgNyutcLp79RWJCQzOfofIUr52lyIv+RSMEorsJOC5OFgMgzDZryWLZ
9L8mH7SGYd/AxdERs6tf65YEzO2/yimEnfh+b6fsskdnIzv7sWkCE5Xp/uP4r02CkLtEBR8BXLuP
XEBCdmPhAI92GBO0TGkRqdmCHQBUiyg1CjRpPZClZfKP6E1inU/14w9rXDz/repEvMpYhiaxHnmM
csjLmcfi6c3sKwpoChnE+dgfgfp0VyFjAB0+v2NpaLwb9aGOwwBoHOCzfLZdLBvuF5cutURK57Uq
S6Up0xJH0JIjgohUd5aVZs09aPR0yCejkxADaFEwI40FEoWlvxXydJ49WehsnO8J19f5Ucafy7eb
AwuYkwERKXaoo1pCQ4S+tV0Eullv5w4A3CXpowp+6IL8ruy5F3yxxilY2ykNj2rUO6g8UZJ2YvNU
KswMLULAS55aajHGcLeAkH7j52YhcfF+Ex3xRPwVtSuvqa8Bb5GwLdnHssUWqfLWe9v3TxQMnCKq
8xwr1bDB19eHq/qKcKU7dv6u30UNW+0EEiVggVvZzaQS+sgd60Oql++LPP20a+LkUerO1CxIuoor
STZpi+b5N5e7ZHR1C0HRSTlOStQ/8aW+M1AYyHabaGNXLnxUU+IYJw+66pfhn3TEdRtZ7qNxiMfW
6jCTQoBDJ/DXHg4HFUj7dw9tTSim/BdmOVZ55XXHPTboNJyaauqc8DzF1aS9CG/aQ+31/7r7z0yO
0h6pVwfTk/zjhUL3IRlspLL8OvWQWj0orDimt9idrZgBJk+wlHoWQv5zB7goHL2PEy+I7YtCT+ni
lkXPeUDXLFQuN0KlD7axmhm1kUWiXXnXnBa2aXx/ytKx8ftXdYhDWM4S5sb1XeiiJj887cYRUT8f
ZSK4ET6S8Y7hKnPam1fszZysiV0g7P8d2YYhVRPI7gJowwaBCmSCmPeeneywH0szgltU1jdAacq8
/TO3+LnITqtk4s6Buuz3Y0KdQfzkbZjOF9zdq+iNxLQlRIHcSzlmIonROdUEERPqlP4WODU5DJm6
O7e4i06iYqCnjAp8B11TL/KTFCEaId5vUtcNufUC7rGTllzu41FmrvQWh03xQIVlf/dsMyHshZrx
04XEhEPSYxMGOYZWqW7PMWplqjkPOQa2tHIY4531rygT8Ibhd1W2w9GMvP2uTZ4QX/QgjhNFwGeL
2hSFmF1PGM4cLf4huJtCkv/RgRbn8LfiJfhQNnHfr3sjXoHmCPgcr8H2WdJSzrQomaDDlqpgg9uF
UYkeTgsMiJz/wG3x/aythsMryRNmUxPTDdyVccZ77bpDZJNJu6HXQaoB0wrbE9kVHzxQ5Lt7TVNp
Us9sq/oqA0ViAftOXwB7r/CiXwW3I3u2IwaRBMvu1wmaabIU4VaD48iVkgTO5+J9EBGFom5cRqkV
vMymNoEdnkJFMY8AWyww3dDma1itnnEsY0YHtBnMVhL6utaKvLbZWIOC7nSObSNmI4qaoWuoGn5c
LfdZPpvHm9DFfJ4CWnwJNzRrbbZy7kjUg1lGFvbvh9mBMy+Sl50JbGFV5rpnGbUDMzd9qv11pE0u
uNKclmdoPGBTU1nynFTKheCQGZAClqnGWbpHMRPqaTKADFjTx0Tyss1Mn8KJfPHiC5keb5Xc3HgS
ekVD67x3y/zuLN1xL2lkJnPLW5wTxaIUsHObLey+EoTRCrvCRoDM1rQMbV4+HkELfvdNsCS1JzER
4NPRIHKgyq0ieRKaTs6T/2lC0ktIuQS26NwViwArWuz5UhRwDfTzmdZRoCKyVj4T5nUaI01Uvrub
PMd2dhn/xmqnw2ImNNMjT09rs33EAF8wiBew19Tpbx7VRgn+HnsZU1rnREEjRYpYSBnZ7FPvKMaK
sxHNHDavrns5gkt1FsKkgx+PcYgj0ynhqH8wVHWju4wYiSdAsn38R3hUBSHL9UgVYv7vsJtaRQtV
sbem105yPtM18IkLnFw/V0vSA6eNE8Y7QiLZRw7VK1cxL3EBKM3531nwv3Y5WHehm3KB5c5vgLgO
YRFJu8GkMuMqA5NP+WxSpoAA1epqQSJUPew4JPKSGBvx3b16TJIUCaYnqPE9JA1/0E4nis2iQ3GS
JF7sH4KRXTtQwPv/WYFHQt2cadETdLmRIQZVs124lwahclbDziNdR/TdH5izmGVKRsoxqw2tolMz
xwLJuIMYBS3nHYfZ6aO7dxbcWWPVcBIME4uFrP0+LAoeGyn8vAs9jzVwCUmYQw2ptMH/3m4M6MT8
fDOiUzL0n9VHYQSEAPE09BuEA9sCaWIRjjgQpdCAXDAH2l1vkrj4KKunBvfikUq19XljjBaUgwVj
1Gc9JRzPeqbyYa0bDc3uEmn8eSc7L5PWe2wPM1yFxUwUNZn8z4owbx29yjMim/HCm1euAXG5T2FM
4nVHUf8h32ahqhu1DJ4hSE0yDYqMIPiNfjv9QdXsfQLuLoqoxYRiQmUpAk2532JGnVf+Jaq8nNCe
rVBORyrQAEcBMzP27IBxd2bGtYJInKNMwjU4BpZ1O6a17/nNnh+9TAvQkvVq8yoLmCyKCfjKdrdD
LiyIL8l+NjydVxss8+NVstjKAGdiEfaiAxphYpjW+jd4UngzVOUt0eaATTLOAGz+1yDCEi5j1Awq
TEbS6dZBzstEK2CH2mqRQbRtoXmet5cO9GR3syJNd8WdBo52W6qm8taRY6zPlG126qUQWjIgsKnN
4i+lCrayrSvahSePUPGuPgg1b0L6pQKNC6Dj5LaPlWLE/iuSG8s0JSlOcHcn/z5Jql6IYcOtTWRl
64OsSAG8h5a3MGd0t1wzpcGOCzkOyumU9ZFkXdVqjVQKqxXkkJR5cc+mk+y9UmsDvfFzyWDiVSAS
kAD5kU9AIpzHAc7BJETaUvwgSV0pysE7Fu6380Kr+Uqv0IIvWqEhqAvw/m+jII9kw/t+WA+Qnvci
iWHwlFKUG2QEyRZqKktd0cfGBmO7XbKp9b8DmyONQelzSHJd7LyALScj/5BLGL+PdiBJS3twkJYx
dqSGKNuuLoRLn+5T+8nFnA+0Vg2RG5mflVStvo1+bJ/Hp+ftOB19eFt/StEN8wU/PoYKzaCKJE3Q
4yBkxBSqAwgUQpe6BUcJQ6AdQ3+ZTBxyr5BEQvWp6Ttnh/a9TlLrduRbsFrs3OcpT+coSpBoabi2
2I8vby/5WMz41tzvQ8RxXD+SFzr2TiTFRtcisGSPKrDCPJ0Hw5Mfa4d0UbkD9Sus8xSNFSpagx2U
XBWcvscgdL+/wqxcmrvoygC16kWATO70eElJkcr29Qf2KAPv4DAe5LaQzCtEwCc3ngmUI6EwvddV
W29/9WsRtmfVQGOqlUr6IBdYJbjcIVrval2eqH0wLSPRdbiXQcQHo2/nMShirTIaF0npD36tbgKD
m/94n1TvTO/P4Oe2vHMv5d5IRsf1lXm8Go0OXDNNTYvztIO7ED95wM9GSdM96HtvNnhcO7qYazhs
v8esWJsyIh/45k4SUnzORZ7TdvxTlPZzVWFziHTZ9fLhuWsB33S6uQOY0xHQiQJzxh2z1ekmHw14
hIL8Z4nEOA+3LmWeeXF3wTJff688ELeWBn7ieX49nv0L+QVwE46/jPUwzAHFV1f1BOF4YMD9PV2k
5v8Aix85lfTWgJ9WGNxf+kwKx/SvGL/fZR94PRUYjVM2rO3YwxqU/r1X++zU0IlpJQd5L0k0rxdv
XHMU9c6x0zVIqtloHs9HrVUt1Ow9/qEHzopWpPMcz6xRWhO8axmRHUnpU+HR5fG7Cluj2GoF3zU9
rFAgRqJvlhXVQ6Qt/Sf3qLv5QCq+QkZimfcWC/awe4ZNDI6nX0cX1r/4Ye7H5lRBTJulh6o3fhRq
KFZTEcCw4wDiQ5ILB7AW2LUlk5Zcp6cYVE+cTiwBBTKvuh2ttOUJAsZhtuYxPuQ1U41WuQ/uvy7o
5fp/4B7RUe0xS1qO7HGYyzuF4UaaPRvTPZQWDTi1ZYCrYazC0H0rZ9vJx5SroSH0bLvr/wPDThmL
IYImli2Pvc/YSVNSzSwMW1kDDWpEUB39WuDZk1mfmGkMs/M4yFUGHnQZa59lXODjJfbpFOzr1QmT
24Y1oSj4JxHk12zDpMmGIV0IsdK2SrKEGcWKXE1FHEGOiE6+xsjQ26xILdUBzyugDSvIkVc62K8x
GsCU3lJ+UcAbB3SZpsObtpGxoJMNF20YU7hrSJxoPAMUZgPRAE2M+Om7mCPxD9O/WoFKXghL9Ccw
jWtniUkuGwjBTI5YMGWiofouSZ1Pk0lB6/GFs5CfW6ZOG/JenCv82bpdcgSGbMxfWbXIZzJSbSQh
7YekaBthxWJ61P4JkyZ8TNHQKcun6Uk0xalcAd0EKe4hp7MbuEYVdqjwqBU/ZChwDTomYDpBz3M/
d7SUUvgkG0HheUQvyJjZsPqcnxqhX7oHQTGbD4D021t65KBwAN7mxXC97S/3F/rLzwgTK3bUgbQ3
J5ND8meNOA/l173qqXXYu0kKgJBU1hB3aA/ANL5WulNNrk5wYVnzyCIJqTnoZMM+AsuHNiDnRPtL
yP/6XvMW3hbS8i0MEpg8fkRuqgBGG5/ebBFqHJp6N7ymO9rPo7+jCBJt0lda+GKxP0XDmLhnsIkP
yhBdgAPggo21E8wfzL0uUvjBTdVmAMV1zIICo1LZDAdxpyhmZNzEh3m76Iv0mv8NAYKwNN78CE5M
uOXqzmKRwNe7DXMjg+FQp8z65blIU8Df1ZfQLBuJi++JwBF8OY4A9Z0U9XgbB6CaSELC4MD5mcS0
AtetxD2vL2X9/MKJGKDpLIQCPWR2uHlwrO7adAs4rtCD49pzSZg2xBCzESnpwnaYg3uqolLlM7zO
vM/lShK5iylC1ZuZ71mLHV6P/8wG3OJ+XfkqTehgttgQ93UJVuO5qg0MIB0cnVROCfVSqmVNYpQL
OYCSqf8/mjPByfD7t8b3CUUskApFHH/Li3ew2o5Ub6ZT0OTvBzubgU8tv7Wu+NFkpFQ5I7UXjKSv
8/gC2XZEG7HiSHbZlcU+0cxyQW5IktLMga1hqJXcHM1m4v0+S8FS2zbEs2FTOsUoUGp7FOIqYkqA
JB8zzreE4QrWGrgrzndlPxYDODmio5b8eG9IVuyQpN+sLVAFJ9ahK791SXNrvRJTqW3+6FqCKn0M
awH492FTRxHigHx4QY6/LD0vuqN4s78S0GeaCz6gdL4Z0xm2MTDsoWnmPHoRlPLdKmWryFvwV1JG
lOapmcp7BLkxkIqX/pP7HEjRcPxoggLVOJwZVCdcVlPhMjgEIfqz7l2cGNU40QySbk2Ocm+/+JCL
CUySaDxTnubYNtVwOliJ2gqmRkeBzTlOxe4G01Tg1P1wYi9FVMLteFOAp9phzDyoz7VhJYurRxcx
`protect end_protected
