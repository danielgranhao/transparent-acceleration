-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
2N/ndj6GPwGr9nZ/CVewxSBvOQm58w8elAByQeqZYyoAWICkzauODh0Y9a3i6mas
sMGavBE87VZQYMlxe7qt00sVgG7QcFGpeb96DJe94v0d/qK1ue4u63a83MJ4maI+
HajxtFAvw7F/jUBVjKXEyQ9HQdUlDIG6AaqRaDkV2qSL9QPoXYZ5Kg==
--pragma protect end_key_block
--pragma protect digest_block
P+LhloHX8lcSKrf8EN4yzSXTptE=
--pragma protect end_digest_block
--pragma protect data_block
lb135y318X3viPEeAhgQC93kOaflQpar7iKoOWBV1e5Ud5om+zPIv+nc1mNgRdZh
JGvRew0oUnDlYBAI45CP9lB8pkvVwdyiN3LbWuOl0rAcdufH9SmZc45Jim/GuhNT
KKpEsdD1AGLaokptfTu2IcteZ15w8PVzHtGgXMa39nG/FJV42DMIhNWLM1X7gnpB
uutVi3mYpOgzCv+clNtXxkFskTj7r8QMMs7NOO8rIZFeK337yNFVPewsd5n+0EP6
81Zm5HJRRqs+5QOkkU++KbnGgaRaa+4+2BlAWxqrcYvCuF61cnHW2UoL0KEHI/kJ
CrPvDxZXK4rexNW/WEi7zOO8rJ55FILRgOrbPbEQfpWYVURvbGmhD9F3oQ5IGct1
spE32T1eNIVnXKPfP7IQkl7F1b6+4VspCfmLV10lKdspzJBpdeWt3WRE6x1cUawY
5qhity+BXU4bdl55bgfwG2SrkK0JQD8WxZv7Ao3G83ibPbgqC7xGIgfhpkczqS47
Zb2Mhx/eH/KUODcJ4O4kQickY6JdcO3V7QjNrwL4weN5CCMfpzMX3K7SGIG7qE/W
Ey14hH6tqjeDORfpaZyHma1VdL1ALpuKY1pgQP8GYgGf27RIf1rE1Ojkog/wNakg
sSeAm6OWKJh9kqgMOHBE0mMAuV2/d6F6RM/yTyEGcOqOO/f4hepm7PHJObNsF0ll
ejPbKPOoZV7/09xVgrUAatydl/DAyUJHjyEuHZMiKP8euiRMisrRKZhvSh9wfwOo
A8h2r+xuvHUFv4YuajQIX5vnF1aJ2SUTow7K6em/xjOSO2iAbzddZ6fLK2rjS67d
ZZqMAYaYYC5SOjThREjDvwdYSQx3jUMJZXKX3/i4VEJayr5PUh/aMTJ7PTsetZ5R
J9rRpNjneA9M59NW1YHoPWPU0GNMA0IKUjhTMxRnnC4HD2wKfgB2DWOhWtl+Bdqr
MY1CCizuMDTS4E5nWAFZlMcPAI4rO1htE5/MZJfmpgylBkPW0sL0KFY+wj3lm6AN
jdmOkLSFxce5PB8iiRYMfRRxBGIJGfDJuwfHTIELysNCVNDnByVctfRLx/YQpnac
4+rAnPmOY5Thtvv7k0Oqj84uFiESFaGutxy3DbWaKuJx8X67vgQ+L+5tlNg9SiDu
E3ETCRlojv4PtjBMQMMaoooZQhnqNLsXqXNEU2xtVufNa+Ai/Uf4tEuU62TIgUYg
lJ/5fX7/cE8zFN4k0rd0DymAxxraC31mxBV4j2+aP7w8111l9UUky+7h98eLWO+k
3A9RbFME/ucsoOYrAqvvKf8kZtR+daD/IJob2oJcfZBOAAi5vcj6jBdY1MeXWVbd
8L7GGOrBQlbpgCwlb/WWERLyc5q7cits2IMt1Vr6HJZRNzUvaP/2/ZPEX6w5po3G
PCHydlrNd4CPvcXUMxb107WUNAPELWjzIFQ3OPzQ3Z2dKoF9vGx3uE4BQX286HB/
c8r13pIqq6X4v/o7j9JSwQLX/FWtveQhBqXeUL9dc5TdP44zR2g+nww/2BW6vTYQ
yMHkWA+Jr1AbQGq23MbURjSxZvLtuXe5OGFnC1ZRQWknUILNW0lDrAFRrISA3r5f
68mKHC5yxFYlrPf9zS3Rk1e0qhGHkPyMrC+ZiKoYvWd6Egt27NGbXUwudhzN4P2k
99xF9+bx3Xa9QS+cUKjwfTkmxuQ69XNKbphMVQjhZntD1BUS1O6Tq8qW2RZGKBoJ
MyiEh3dXn5dJsSs1XUpeCajB2Z6pfs3b+sA9JosA8B/AGZqOXjgS5SDTB7PwViWG
f7w1j6cxoeBRDNuzjR/DrY7xSXKvAy13GbmUG2uPcbWq3PXAx6n0LyZvI86+fjjW
soNLn+TBAuXKGHqv1Cebp1EP+c/9e9lg1E00X6LE5Jxxi7b3YmIJZuFbow/QbuDQ
nanNuN9la7K40XW3uV/qvFn4niQXhJMYzzCyRxGEDqRbC8+u5tbaXgkzgTOXGszV
XN2yaQET9irRCOaQZq1tIN9KZIqs5wku3Y0tzMlGzrPzqf7p1Z/sWVGmpbMnoFDs
9LKtYwizx4a8SufMIQ7Q5pYTurKk7AjSW7g8uFOgE6Lx8GPZBn/vBGxUw9e3J1dR
1USqRyKIXx7+SmuyjqznhiuWN07eNp2Gse81mxWuhjBUlQEOElYmLw8lkyEDuWTM
954LYHaikykx6nsKNOyZlJKvn1fiLFmnOkIlzrq4NXqWQOMB8O88jjiDVYrgv81Q
vSsUe0wRbc3a4IpUm/2poHP0Xy11sLYjMVvDuGC4Ho6An10Uq8XqyNJrHnUThVTq
bmN6w+JHQJobdORZzTY/ZSdHpHppBC/jt8Ko9n8+Hu4fJwReDvWEUXcydAIM9JtZ
OKwUOPOABPKGfYULQj4bwNoGSWhBoYewspIyl+nV5xvn+mhVWkeWhBqIyDFovXuo
CIbJhI4RWssQGUkmdSKq+sQTEXASrNX18ZmbEKt5kviJqf4uq0tq1JiMlrtPtIs+
+xmOH8UW2EI+Z9XvDNXDRkQ1D258N1bJAahMndoeoorJN/acTSJ8jiOj7QhMmMMc
e5fHHbHOZAv/v6emPjTpyb2oAETunHVoWZsGB2urzjnBr2I6NnjnwLPJONosj2sx
2wQ5vYASKGGrmlVq3qy3mjnQlWRJJR+HPAyOL+B6FeBboZMUIrsa+VqQg0t6vgp9
aIFUsssbveSG2OypwZra2l3B0KcLg3Lki1gyrV22OcfRPkjDPEr9JMiYW5Votsr1
/gaOBWDrT/mmTTR5n36zjeVfNxx6GCCqJHKe/TO7GHSceFndlt+e1exGRtHthfIF
mBnUiGnNRHlvyxqo8hlJgKE63fGFLLtHPobKFZdWBuzhv2yTs+Zlp5xJcyda1LDb
diCQ+KOW4gNbTAZySvRo9vv1aMH7q8x8N+63RCPQ7SdUwifMnuyzzweNaaPOoKP4
gtjo6hGAY5+asn4MwreORSwg3P+jex3XHqNW00q0uj6hjdFsnuzaK27QiOfkSfrU
AiJQKWLhGg1XFCl+gLqCLiDxtapFMzUwieo36/enow+6dii4qv8iju3jp8bF+8U7
d8OjfocD7mYB7Ah7JA6oaCEGkIZVn6K84lYIROHubMLAqc4/3bKRNXRnjeiQtGB6
GfxMxM60VgFxBJfcd2wsDW8h6OyTH+yOroo19ht5qwR3m7eTAeBC6P2+MTuXEsCy
BfH5MbAt1Y92tvLgAWVE+CIac/FYZ1V2tQj7tY6nTvOztVNmxBUMwPzwbz+N0VVA
6ksE+HI7hxFfpbUW4pAFRGV1qKbMBrKzx7y16h/8BS1EEIOsmJLr7gvKGNo7VvFj
DPJ71VZ5JoAZIk4/EnpLFLUfAMHQ3tAt5W1a84dgfjO477L2gq08BTE7V8gR+eep
GTSjCawE2D9wfo3/q3mtNrEIXs1ki/sXLyIUSCTqhTEZ6JD6FPEDB62NFJTbkUt6
aJv4rDS8JV0DmdLfa6XEHhA3bAq2GgBiAqkmp6XTPwMmPd/4g+vHv8OcmmKyKKQs
h7u4UefV+T4LnIGzn5/UpOEG9Tv/kfnRYvuRIKxsy2rvmtrPrBf9AI3I2tcJ6onK
6LVJ7aLFh9kEnXnzBF8wm9rSZjjT7jb9cavhNUZGlVscT5WbYSJSST5gEypNjJkv
g0pBkCDfZi0WciBuNgcBIRm210QvNBNXl50Hnd5ZAFQHmZiDliptOTs/ehXbaJQh
gQUy+XBOmC9Dar79G30y1eTsw+3MxMeM9xVY2CSZ+zFJh671Q8LVQV18aYHr2Mli
jfYqNd+FOKOx3V9rd7N5Vuudznip1jhkaFzMLKM57Q8d7ZEEFqhIwFZNYjkw5IVE
jwgKQXKMINW3uLhN/6F7UExqrm+mjY3fmgdUr2QUhLN5S2iuHGiLM+Dtbc9lmahW
EovyvtYHeLFfca8DACkCqwzLLVYc5UPnIwDDDra9uVG3I/GmUNO22FugAL6v8qyV
4qTDwdL63sQQeDRxutlnTdH5jwM2cyKzttcRskaKhFZ7v/ZlqyMSgwFrUh408Mxc
P9ccdozvpN2rsmfKrNgAcw9IfeFfABtdSeoUvNBu1U7v4tb5mxZWjTEEjCp3KqKZ
B1RyQZ63jU0cxeorqRYyRikQMEtAxQNujku3v0sfLQKlHoElWnlWcLY8QQm9vK0q
/1FlBL8HrhMssG1G8U1zgY0BTsjc7E63ESKSyl05IoLZLdAhDLKDSoMKq+QM6uFn
IJ3yGffa2MkHxLdfk5KhLNyHV7Zt1nuqHOGxkEBVpQO65DTiFEgE/Bbed8VNU/Gn
sffxvVE5lJ2D88LHIMwMD8WdBu/dHpJm1dZCd+ZEIP+6obwHMQAuYfNH1fE4jfgw
+finU99BD8euoySnwY3RE7xelJ68h6pao8QehUI0OUj1SNhTRQyuaNk7h7rtsQl4
+qJ+3t4uX/xBKW84ZNmNUyZdHoA4PP+Zm+Q0bnEuQQYzp22FCXGl1iAurlP1cR75
GjnqOtlXg5El6rMViqabBpKw4bsGeYX8LCrzUOePz6HvJ1eDJ9pQPgR5N02yIjr1
dhV79Q3raEE2HUPURax5Sc0shTkSD31vKQV8phGZp38urKrs5pvJw1lStmgWnrkg
wHW/kNUpwOULvWtpNeDTpQrq9cdxaVtM/Use7qFUjc5pKtLGgstdtN2/CjQxbEow
oJ3G9GgADcKmFk3/yV1Wi8LZOWMAEfgurJKgn1P3n6BsoOmJBb+bgiiR3guXW77x
A9FiXfXOxpZJ+Wf/jotqXU+t92C3gRdIxG/shwqbKNACbtH35H01KYTcoJqsFq9Q
dVjdh3XZIL/y0cBfwWhT5UMtk0rpsOPxJinq8A1VBuvo1KN02O82e/fg76cD0TG3
jnGNsDMxZoS7NGsKX9nxdJuykqeSJIhe1dd1h5FWJPD9862U62rrapSlihk1XTmc
3ZAVVGO5v5hqlaDWxg4GKX4A2GMlCc7+EPr7KZhFUkWa3uiJYuKmH+RCmAIC1hAo
cdvDsAk716KafHw89sPlSc5VsOUhBXtxavnqUwscokaC6DrB9IyrJwn1UZrIxMp9
W3y9kkvLWov+B0aYj9BC8D/bUui5mBmk8MMX11fwbd3dUyGhO+RJVMhf+myhSkFs
jOmmd6PendBGthZAqxWkH+LaAaStAjES5VzHadExCCwiTwT/mNXtdr8SHIMJXp2e
Jp+cyDBwUPsDCIguIoN0Tf1t+zuW8dTHj3sSOoyo6697QJGwPZPs2x10pUzzvIS8
S565BGuVZ9Cny2HlknSM3+/stIAkQPHcfecLlDM3Mun4WtfC6+h8GwEQ/SfOkd4h
hLE6DDWvgAxHMYPfMtOOhPICyhCQFXMh1g7l5h1qwScrgpRHt7AvJwAMOialdS9I
dHpMJQJHxhssUzF5U0zdcHeoLlpf0kTQTi99yPetnAWd3UIPFtVhbGAFUFuP1nsz
BNLfk43J3uzo/OrrafpOlVFkJiCCiPwBNljEqkJh73+PadiOauxk2KrbbnEP3rPC
vUsmsrcdaodzyEwqlCYQeFzrZOwsjgBXsbpk0P5ycVQQLJFpsmUeVrwuAQm9hGXO
y/dPKdKn0ZdXg11WGZHSYBIsyUFuIgybDAUvHxVMAp7bnpDHGfAjVAJjagiUV/Xj
ZfipDluTDqFpkmW6fka40Q4fVNFqUEPxtiifb94U10+ihi95Nk4NXISsviInwKSe
k3l7gk0TbCjz8tL2PZFJsYCALPfTTPCxk4cEPRsJd6zossYIsXUlZUWEMgdrdrpH
CkgYr6B9ai8QRNTsB33s2Z7Jq+kfOE0S7sjl9R4wiOsViJyMW/F5OPegk8X7Daeo
NOH+r8Sp6AhZe8dkJmRKEvwHnp8bHzsZFh5kgCSowR1wj0/qOJGaEO3S/vfPPaae
VBrCtS57hI18r7I8JoL8TsXVpuyASQ7Mryaje5PMWoTKvhiL2WVS2/On4Ufk0sko
CYxSmyd8z3PN9tA6U52frIYm5ER4U1Q4YTYfe1n4VZQWgI8vt52gzLGFzPWwtpz0
bEaCTkQZ7JBl6f5cnzP/qk2WJ71MNymcSGSVCF7gfIYy4dTWJhFThhRlgnCi8jaE
UAEhNpkLBvWlIdiaPN4ybZWa/WPLTdcjqJ32gXkO1hcsxJG6ka3AqC3CUvIaUpvL
jV9vaVXq8NEguYy5WyoKj1R6J1uQKYWnCf7NYCRlDvDQVBxS+CEk9wxUATdU8WfA
MuPFtJ12ZhzVRl1n1YXmcBSIy8omQ9ULgHi+3K9Hy0l10Xp1N972YAhArHyn5QUY
254f5QElbzw5bdiibiHL7tVsdwLP/8+yfeG77fb/ONJS+dMEPZY1RqxB3FYC2zdb
q2ornZoJ5Z1kpePX+pBy3BRa5jZVVqjJUVqTccENJZRilbFXsOe8HCBD2Zlo+CP/
LKRTHWcZZeiAnMHB6v91Q7Fcxh1PqVlgdnGXjNxC9DBLCruJfGndUBqrVJQxKWMw
eGV3dEWLzI9VUrUo9m9OqzIO3uR61+lFeDGBzhdiWJ+kIaKpcbXJ+YrB26M1Dy3T
PgxPanS3/Y0s2yiqtSDNnQZo5ZCjjByRs/wmkO+6S5lWvZHTa2+wqoNsmTsLnj7O
0uhWTh+6aFxPZhBd7A7D+uiXkUb6nOietth+0I4lpgTLQvZPX8F/QqL+gGQs7dD2
dn8ulVy5worvhMRK2aw3XzKKURKFK2NCA14hvoG6o6A8lDdR1CjIHrvjxZuhxp5P
lvbAc10sLvyj3Po8inIuwigVr+lCDpUAfn3wiRwZXkbOqwCP+K8Eejp73E+CkGEK
Zl3dv7uCcgXNrNW8en7xV3hkr7XGk5YtQrcUMx46CCLvjVCzrRNBiEHBZjjTLOC7
fNLW3xmsQ1pbKmcAZOtOxBHQW/t7Dz2GmRfVuq9lRx733xvgaTjgSuV2pRIr+d3C
mNS1k+Wv0foD3UMMwFic/Eo9orcGhh97zNahGAmTz/OI4awM5+95Cojfj/3e+li/
K9l6kzMgx7QT8KeheB+uumVvAKl980dPmR87V6UGux081Bo5qdmWd/EkRAol3SI0
SCLpJDzpjx49DBJ9dPnab0x9Xeu7TapIDBw4URBZbF2pNH1YNcGjY8Z7EVp8xW9r
Wm6j+oz5tIy7lq6ONTtYX9h0UNgrC2fdiAsTJfS8WfWGgIYBUiybvUe90juEu9z7
m18M7vmgdBObc66b9B/zbq9mFFkJXMb8zF8n6c/CgCb0sxs5W/06CMkS25c1bj1o
v3N81eE4w8ObJ+1pFBgQL+E7gbgON0UOan3f6Zj6O1aCEZYKu3UqlcA4iHAiCY0A
phq2v4NISvFbE/l3beNZhkVyOBx9mQUmPcRg/ajpTP1A13G5sNwsweLejrZe9g64
dMlxiA+wQtZjLgZjK9Xd0uK8yknsqxGwAxbILCgZVf3/Sx95b9b67VUPOPZZijjp
oFIRmgPirzlGjBE1tZARQHwI4X95/jE1iOmyLDEwIBbkGOhW15Q7ZV2KC763Ugkh
MkNwhtYq6bSC2R49XnCLKT3XKPyBn4Tak3BPCI/V5IJ+dLJ8igXLfEMNys7pFvew
aOe2ACKnGIlTqtqWCVXB+AzRzPt7erOsur0/v9M+jEXDG6OKiCTI8W6H1MSyVwoO
FmGule7NBiGz2eqsQmd6UHKRqJjpWDopIB65agjgWTU4hcChhDIHCVNkrtcc0zTN
SCUtx0t0jQEIHBw9VTXlIXRGO5z1jtjtcmYmTMMt33B0V0EGktOsQwuTherxovIS
pbSTebjp26jt+t/IxiZ3EckX89QzPkyorqKl2uwyeD5Vl5p2/0c7mCkq2YvhaAGX
eI555p1AWLNXk3jj59bo9GINXnKA9BBkY8Q16ClNSyhjoDMYlF1k+U7eYNb1pgdP
+VP/iN6a4p3p+rYO+1rCPphiuviYm2IkdwrLC11olb8Y0J3Du33yqxB+KGs/p5uL
wzgdyejr0CHP45uXli5mmCp0M5xLBZktdiptipl1Ps4S7H12Sn6Ion8PdgwUr4aS
7hFdXXDMgWJafffTH+E4aV8u5XVKpb5hTJdt8ozxdooGQ3gZUcjD3gQuJ4kL5yZf
E+BGV+G7DtnCKcHnPpRdw1skDeLMh29iEqE8m6MVCMgI/2OJVdyq6iJCmQcqXeeQ
FVHBykQgt5LhLF7MamAm9XSXEqGz3krswlfJ3gMZUL1fAvD4jWqsF6uwBuLmFPYC
4tIY1RiOFJIAEXvx1Ajyh4H29Cvfi6QqPfWgtSZQX+AOLdgEC+QdhtoLs5AirVIM
Pm7qp5QLf4mTqguZxrX15XVj/U59dU+HvP79L+Hy8L5JQcewNicckAoQcPLt0RN1
VYTSBqa7auzccWa7Awa264TCIF1veXl9C1d6gBeK6rZSYQOQ5JpDfrDTVDUJ1B4H
9VrMxHurjMmkecfRumvAJToqdLZumc0PewEqo1cmRZDW9f21s7oqsO078HiW6dHE
vmMuima7XPE/WjsbdUXl/QKGbYER6Sxyx27i3mLY0ktX5IlUtBzqOHLjhJ0jez3R
CbB1worTtnh1j5HnaQcqVFWj1NWBjhxfrBBo6RAOQhFHk5oDklktiN6M1YeTP7iy
OcC2+v5P/mAb2ZwzZAZ35KSTdTMkt8vQZd6U3sTIYMyduq9+G/lUUWBVnT6oHG65
TyOlvAjVL3oLVy7WCZFlzo0ZTf8ujDc4CWKCZ5IcdG4PiqGs8AtmiC1OZ71Gno0r
PVuYJ27Mdsug18FK01HXwBYGyLFTBe1Jk0d3T0OGpTutj5HBlYtYPn4DcErzSjHt
zx+fEXNSLneSEHiBymPOt1YPkJW+cAVXcVckSfmZ3fdrdy66TxinNwzivbXhlrXr
P8J3ZosxR6DXdNKIT8xBB6bKDkGFwP/DMRSpEdyNpqkr8vWpgR6LDCdxV3jsVZBv

--pragma protect end_data_block
--pragma protect digest_block
zy7CMhSizUuJMtUM/LT3Wet6vMg=
--pragma protect end_digest_block
--pragma protect end_protected
