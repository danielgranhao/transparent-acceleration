-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
NZWgatKpzvnwNazbaLRrnrASXDH/KVd0xuoBTy1qZ/J3ePkIjSGO0UhirN7gJ7tp
/4tz7WDKfbnviWtwjBF37BLX8yZw/NjwErs+oEqKStRXZCRRBEa7MuZaqZo9GW3x
VekDHJgpmD6VfNLY2NRu9jFYKHsqLnd4M+lbuSK8Jgs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7559)

`protect DATA_BLOCK
rkJNQE0zIVzHy7v0UvONyK8QXK+sGooHM6J9d+LQ3Nq/SsWQt+DphDHDGKZURAn9
0/5o/46nInEj7oPorsvcsDp9h/zII5rKYzB75j0c2QkkC06UAipV/gQEztrmQ4S6
qU9UTeXpiUfnmdYmoRcRHbkrhsR92eSjqwk4KfwNOOKDBvf52R3vITzIAKiHd8m0
KbRdAsE6IH6jdoo1YJonl9keH5FFbQAWNvn3LA1qszFpI55adf+DfXA86xjNR0iI
d7kcPgmaszX1s+CTlPRewyL3AZyEQ0ZtRH/N7QXv3FR9tkT7Bm9dpDtpVjqD73mt
MvhenrLXbnAzZCY731SXzw6jmAlisI0LvENkbpfuC6tAEy9gXSIwTogNwVmM82Uc
h6Vu78Y79wGPXXuFagrDhWub5lQzOAcFGmE3jVnVs8tm4cYbdnG0wzBYcg/+jkXV
tXH8Y4gBrsGCSBmqaJc2l5NfvydAzruY/9By7YQjhRLiKwWkD2VYRa1b/Vf1kHqh
lagC0ftyKLY+x32xvzYu8VFWwIm3tZ5XyfWKwgwPB9RIE3WNM2/3Cvn1SFWLeOiz
ZDbTxsJ7qb0x1+o7X5UE/HVoLlkjveT/KUQ+4wvP3WrHvBvU8ZeiTQKkPWNpfInq
o7r64itVTTXKwI4VpSKFg5H77HTIBzdiJajpxhWmh6OkYk9QPRVn/YERJJ3zIL9W
PFXEf4kafzJFhF1THpv9NhHKChJinkexr0dnHGknaLh5rLPKZeW6sXg+7uhu+JyL
6MrvPdVFff+wPE9B5ntLIP/tL0QTiHhk2DK7EJsEFjPvyqJAc/ASYPqzC+oxBk70
5TQoKiZ0/d03hwVzq1mcb5BDRc9e3/y4nXC9njbRukqrOxU1xXRTBDNJ5eMHhsOy
aACUZ3sZHk3vkhztm9ugy7z/n/HJHVlVC8klWMgBBQeu9L3htS5kqhf9kddc1dJ3
QtXodkHl8rNPBU3mPrF3XVVmwr50XEKTrJxwpH92xD+9moMIdYXyyQseHvlhxv8+
9Ja/iy948GOEBFbTtRETMap0XVGEe5v6w5uuHMEfvzGThncIwYTt5y8PCshuot2Q
+dR4gwTCbtjFppv7rn1oDMQQxeYckuUOLfj3B/ha+cC2lcqMt1mf7aCOjoSnXZc+
QuN0nEFU4wTAX19WfyvsMwYIPRTBjaFVVJ/0HnX4eEMW4gZzGvZrFf+7QPPfg11s
kGOnP6NyShkvPv0hfc3FTQT6G72Z8PObdclUpNVHVjTnY43TkjJZ90tC6/oZ9yDl
l6UVm7lYFXug+KuE36mz2KlKeSIyb5oGJ+SyvptY6Dqm9sZgyf+23YoalG1sRtRk
58WhSbiQM1fO+BpIB9DtAGjOowWwJBuSTS/9aVcEwyabe5FmrvKJ4lc63560nVoW
LjOZPezD98/G+pf+i1hjk9aqYNeDTWF8bQLrh7BdtmZBWSbzM5i9WGdB1av7jhj9
+heb+I+3PcvTYdHdKJ9PCM1SIwfQuaCglVKFDY54oJM/xeKZm4tSrk42Eho3Yhyx
OjFSZaTY5axz+wumQW5607yXS7FLsohHFFG+S12nIlvZyzC5qtNlxqes5rr/jBEO
MqSFpKgYeYB2nDg1otIvjfNFuUs5JPYV4PhS2S4BJaexvynF2y2m2mudHPQe/nnv
r82RejAsyK+x8LaAOL7VgNKMJEJ4JD/CbUOBe3gP0UNeH5NdNr7p6hzP9BRXCKEU
317d2vyoGQA4KTT2FbWUKF8kxYs+xPjywxiXLXL/m+Bu23Cd0w+mVBq39W6aiBAh
cotKWLQQ2C1LHFQhXVdw1nv0sfvmn+LJRG5KSR7J4gH6z5YqlEXk6A7DmE60U4uV
Em2lAslacFpiBammBB821idmUempmI2yLaJdADcz+wllIXn/YGFt8nA8GlWpJmTE
a/u76AP6jZVi365kDvKAQkNHdybPY7kMiNnE7KlAI9dcWkEvLwexBxfnZdrfR0ID
yO1JCt3jZUVVgVDYRxBoIBtfjz1DqA6mo7l4SE3vNgetQEJBnx0dvY8xL7t0VavL
KAxszT8TdBa/b1M3akEZumJoa+GMFjf/leScfxRR7mxXPUcBMpD8moOvS9zX69pE
a1sSi70f6mMGOK4N6tJKUoUHVKQGYEpe15bm6uk/x1ZLfvtYZGICff9p9/w673qY
XiTYm//Y3ibKmbQDqeW/fGHvuF7lUIZ+vEKS1UzrvU8S5Hk0JC8EgQVULrAnHvJq
f/iKwhi9pvp4Hs/ZZxhYlujSreU8jddX8XjJXljN+0+r3unWSfzlz+s+4nTHxXNv
6FCL0dR7DVKxSlmdiBumGiZ/0wzG7e6BAeReMt333DL8uT0W25aR6NQeqgVoJhcs
WEAeF6GG2FBG7gDi0q4hFSiRVeVIosX3wcanGW7+fSfY8ObcNrD9Hc0ZmHMdDWJs
J33e+9ag0Ht9Qh0t3VCEUzE3Giz5HxvW7o0fbcyVZXqgXirDCRj9z2wHkJnsXFXY
V9oTNyUZozRZpzdW+qp8uRPACtuI2VKv2ResvjJzTeYQna4FTg+sB8HNNdZlvFNR
ohCOlGBRegMUgFE3InGge/u0+HIVME3dczdTfCLHJ8HH5PMClFqEiRtYKxgLCaVH
CQTNKjbl+ooFC00IsESGBbArTthJguz9IQ116+OXaZLYzdoIodVGwo0xtBS7HdeM
v2Y06yQMN6rf5Zn0BXwUaMHRcOJn718FlcO4TKu+duE+84W1ukFbVFJLc5iGrGN4
TLY82PGyukpwdrH0nFrzemXv2/WwHFSvlTZyQIny1FXhHT+QPAZ2nFgg8Ek8g+g9
yC+HDuUY7ohZ/i2Sl0GwFvUBtIhNyFenmvOZLy08fOvx5PFkQEXgdsWRYh7VIJtd
WRgaawaqrzFpJh2O6lxyJkYpu4QGsf6hwhoD3enzXzKa8D55tJc2qyXx8vTsvoZY
ioWuq962izXxUMTVjOJ99ae0KNhrU1Xi5YtPZqolfrA7W7nTue1AkgWqLH7XNcIh
WF9SfP72Enyuh/8N5vJOKaynfVQTWs0+HBBLdma7o/wXW1JLwlq/9UWIc9Uja9DN
6IcXQ+hTtDFykFbCyK7C26L9CLu8taVgtuxjr7rKTnDbGC/j23X/Dw70PN5BXmAK
LhPJ/dyNG5c8Yt/3quO5wP1uUm0uL/E0qHYDr0ei4Z8ny3ghzbceEuSAQClKFsrc
6HR0G8yN60vRbq7n0zV7jn1CRI/YQQyP2Wve9p/Vjxu96uwczcR04qlej1wp9BXg
Kibbo0+k814J5KKkNQ9hP9dVptdWAz6IPaw0mogipKBpEx98Br4JsMiHlNz1a7Se
C5n/iCgPIKBi4csIinR19k47Lc1lov8h1e3inzTWymkex9CM1SRvMXy4frzy2yQx
g4wCmCUXhfKIq03MqXpPn1b3CiUuNOKcJQ0K5T6VcBhhxlhkdshmPazclOUoHWhK
GIIUhFx4fzHZKln+LU8adUzvmbWgRIzzJ+2qHOk8RTQ1dUKCHlZTgSkVBNPjchjS
JJ5AOKm0Apj7L29RT1z3qTG/urighsbCwVYkD4aMT4s3qGcsA7Vm51PjqREjraAg
bOX5MB/itp6U9CEVJISl4xGiRiPpubs4efE7R0TrEWapcjkeotx6f2jWjqxMd28y
RWe1n0H6dxn1tQDbzm+q+Mo0HQBa1Mo8ZBnxgA3xS7zrs0hcKNuuaVLwnYXzQpBo
50QZpwUxZTrSQmW2qNCnl/K21Y8bZH4nM0IT2Tnn6ky7otgH9Xu8orO6/1B3G5rv
qSMpaNSPu/uvMJdlmpWYkdziQcwLBuv5YwTBQzBzQmXZBz1PGftrzmoMPM4tcNMz
tAXYs0Uc3xTI2fp5PGkP/X9XnCHvntg5mo5/cSz9iBZ+NXZGnAAlHD16yXceoFpN
TKDYTwcBtS1oh4y2ZlrXkedwKQw5VO76TndSzgy7Lmm50Zy6qFhL38HKR4OLJRHB
z3LIDAdVx6Q4eGwn8XHgnr/sRfKdJOiPlyy0oyrpHb2ffbdHCGpmtHqnxulGGZcz
zyt2/2OXF4GVaXEFzQXrd3bPhbdTeiWFtHjIvU4Xg5fUTN25jOurRX4VLDvBxm+T
tfT2jAH41BKCL31VbcflVtOdg3NXcoaSefDcWiH6hR/DIcIAEW+Fl48MBu37KVlr
g9xsZT1dviJGd4DXEwrjcG7M07DNHcKt2QkdxMmmpQ3O4L30yepBvi/CNdZRQz39
3LC7ohFDJY+oyg0PMtagQwWjgUJV8T1hTDTaurxL4uw105ugXNrOkA3i175YBLlM
47J2vxGHMNzFPAGhPJEbph65zDbSlfnsJ/moOHrW5py7CnsgXFMDgYZGHFZvg7ab
Hk0uk5Hb6uPfj9OyIrViRvvMnR3H0CXzGXaTjpxVXTvZwBrPzOpJGZ8lh3kk0e9/
SEXDswxZEpYpzVkJ0/V26kF5qgGw0Up2nlAO5A/7x32r6/YTUVj8jyJZz0lY2J9P
ozESy2hra1DZxhUKH2xAc+yWRRgMmsiaursC6NZdHCoKzPHkjUlxp1OFyKT62dM+
IQsTyc2+5bcOsg/Dj9sf+x6EavfzY5AQVnAuTi2bz2a0gfv0ZvRwGMOTZXldBU/I
FqEIhNdLM9oHxG///povhIDLomVRZP3qCyfNtgL7WtH5i79DtdCM7tWm76r1WFFd
Nz/Ay3ZLe66KR4sLhqEDU/X+cQCvxViLSvrnm6w6EX7GmHjwljOxXlkdBEAr29EX
vUGNZoveaMAaf1Qw+0ke+oxQNihGS4EwsHQyNFOdcCf6SIEU8jH5xci5W5O6yZe3
y7nLv2WnFt+FdKCzzIgnzq0GafZp16EIPB4B0yFxls5G+jRdA2Xy7Nor3ThAoBZs
aCB+9SkESSGQfJq6zaDlDUg4MzoU9gePk++g+EW+PSV+hJlMtw1iDghApxXqeTfL
xEYBXYCMAv/UOdcvubI4FPBPt0YH9Ov8uZSsyp7n0spVaW2LItRzl++i4CPSMedT
Qfez/XgPNa2cBddlBHT3yqJ9Cbr5a4WDGaBZt5dIFHog/BTFNuNTQ+P4uriqO0II
84ObDTtkrqKPHCpuu6bn15U+ok8mAbFuUGzRTLfRno8312eoqQ+lpDrJxfxFERwd
2sPa8+0RtAag+08VZ6sUVZD8FuQICpUpGnsNxy4g//2uOClD6DvUE44nQWHAdmzW
dRMoNYgREyyoZME9i1PgmrnIfO35egnS2rJX6LoOE1We4kaBgilQW1Za8N7TxDbY
vFJy05xb4w452ONQxyijfGQQMr8x9bv87asdh8n0SZGZ5NN3Ukx/NWD2B7v8hUty
X+ilENjiGPMnvdGfGsFCoqrRWJSfqrTiPWH6eQGSfWWlDR3N97CXDR/wFzpDEFEj
rX6C9U85J+Z7/Ulf4+Gqaof9HJnkCcF5NHjG1oRrppk4EbDrUbREWcMN50FYb/jQ
yw1bOOC/tkgPTDZR7NonV/QjEqEdHXqzrAP9CjUT9KDT2/KBaJewCDlRepwyEFQe
USv5SbmtMwEBkKzHF9IL6FMTxK7fQsz6VmK2O5yE8fwmF92tRyeXnAZqbCoh6pkU
O4ln45z3Fx4hzN4mNMeadfxoI7n67lCON1vlCTW58Z/2q4KJKzYHeDl0xUdu5vTq
FGEsBM8ejmz7Tj33Awr6TOrJSDjNEwTKkrRiznFE4uKXpbZRAqpa4395Spi371s4
T+sE2szPXpUAheXCZOxOge6LIOjeEzqUYA6pNJHQ8e9g8V7TCxMM71IsM8bKcsJI
q/M9mAG9/4OR8ZfegqdPgPiUkh/t42HnirzlXQyeAeDXRBRyW/ROpA/4B1OJspAn
tBHEctnjAHFGuHOtmdLD/RV+ckSwI5FGpqwE2jJYxSJim3mAIdFy9Qy1Y1deQixw
1NNcKOw0KPSYSvXn0AETposU3yeOS/hMwBxtejvuS22EkRPg5gxsHomMi5RMFyxN
sLte65iTnbVHy/ug9KZ+nN5WMVCwtMKLnKXWUFYQKSaJjO0K+1NcD7YAseAzWmzT
GFETq9zVNODfKr5WOrm6uc5L3Va4/cUIJQ55DH41ReMIJ2pv3edoQVTam0VAoOVI
KHrJAVPQq8khCIHh9CZJCuI/U7/ZsHo3hDlhHBosIEuBnYZ2GkO+exqod4jwN1S5
+fxcy4k0Ip6b3hsikZCJ/tPg1H+nyw8LSXJTwyMQEIhl0+9D7XT2FEvibJXulFOP
Ge9Q2Llcuf+sPlDMqFkgU+srkTYVzhiIDGI3lRoj10UDj4Y0k7r/9cDLBMs9S3U9
UKZfPuKbxm3gcbge19FXGmstqjAaCOtF5GiGbXP1UyqevewhRHJ9mJ7qIEvcK/Fl
EJCBjhG01hG79am7p8KtRyllkpnpa+vOpzTRz0WmyIST7oPPW8iWtKOGrtTW/JAE
X84OtXX+ZvDUl9hkLfFtGxbtxPefMDz2hkls9XKfhz7UB/pt6oWr4AgDekT4NPaC
78TTSqvjndXGQkVEBiBCP/O7c5FMUb2SHtTwWriWciRy8umDRYp7dTfui3zEp1ys
G8EZDJ9YlnAPjyrSztjLPsBkc2UnuCpCJjlYNR3JVC7NOxIZRR75HA6oeZpGMEcM
uclEiL3f44ZYejggLJsLCh9s6CDNUygiL9uB/2iSR7LsjgP6LNufDJkeKIKryLeM
w0K6KEajWQQ08cigrHmcqNJ3LRP9Xz38lQXVjGmXNHpOU7bDEUIeCSQZEsFxi/6d
o6oPdBMxUJOmH0LrBD1KYPMM6N36CoDU6gQdHL9WDM4fe4vuZ/mEpb6bkqIukXFi
6YyXzoompohJBalbgsjXqfMTEATZch0I7PnmtJ2FdRS39ykvXa0tXFwCAhv+v0R4
hyGbPaXZLXQK9cChWAKU0SvvqNtHmga9hrugciEr29gfHgvh+SHe2oLFa+9zh9k7
ZFeGLlK2yTj28zRalLghnHh80zNLZVW9Kw8BeP8Ula9FDctoLJH0BNPZ1886IwgO
dhsIMBhgI3DFBvEoJmctTxowSSR5xj3UqrQc49fT0Vt9i8i7VY8kfrp7v8DFQ31H
qZA1v+VWR3ZhhSnZkWRe2I/anTdeL5YYRRpSDYCOayDuAUlds8Zd1sh3LKVkIFKB
sSbwwVEi9yrWwwz0eUJw2+CSvQRKbF/fntATgiK6Atdio0JEFHnPbkTiNgDsyWNY
g2tCAyj8u+lmb3xGuDezwKad6wLVhKRmN5CWQ63n9+mfn7a0unJLcyrAuJAMzzUS
Q63RDlxnDhSXv938shGBWC9c2kZI4rP/tTfxVMtK9dMvztx5seEKx/3hC0RshS0n
ryaf7XYF3TKk9I5DcX/cmr0BroueeqguB94YE6JtoEwlidX0He3Hp9gZ2MrvG+ph
Ie6nK0XJbp57YzW4c1uB6LS+nUYI9olwtwzUxvmApYzvvj4rSMkjtPVjHTWccZ6/
rRycDjriObI0oUIWbV53QvtsDfPFNEiG3wifNyV3HsKr8+/aVujG7GP3aCFVeTN5
eg5bKWjI3huf7M02V42lGnATUw2cKzRFU9v5gTYhflfoDvf+8+yhSobEzQc+wJFq
JhL/RAjj7Ebk5Q2taCI8EcJgbf3AbDkw4KAI7UxIG86wVslDTzFw/d7U7bPSGVxn
Hus0Czmi/pLZdLpc7teVmxzDy0jDd40jZ47DkFG3URAXF5zhRfDheY3tAp+DFoGd
98j2mjmrS0wt/NG93gZrJuyV6L5bPc4SxxwOIuTShuowl6/gboPL4EGbueRRZLog
H+/SSulhLzd36owBD/gKawFE4gzEx2KIMkP4W6nerZrO/lShqGCA1fgsRs0xySct
8RdWJLNSaHk/SPStUfaTHGChJvL65XiJViMowF6MUzvMndmLsWgd2Ke19YecWBPw
3zZecMXx7o0ToJy6N4N++7TXIaHoIb+S4wMRw/ecWr4MqpQHDqyAWCE0XWF59MJ9
URyDOL/gSnS2lNedtfyqn0xJVMyMDOvZRHun830e5Y634S0t+FQHF98vpb9hB+Oy
tlwiuuXaxl9Ay8qHiRGJhKD7gBxR2lRyaAahXJUgtbQ6JoO0v2xoChIGuRSPQ6Oe
6urY3RYe6LxLPwGvC6FVA0UBfQ7oHbLtputB5lByUpgFnVyGdjEYYi9shDaDCKvz
MuNHvvvOXh0Z4oQahVUnpmlJvrURPaKa8En0s+j37FfMEzSHJTF2oBR0oH4pPNrG
uAoEaGaqA801luqsNMdQE/u/Xu2w0StrWxcpEVyMosLIoFKljXMH2VMwh0zWt7hF
ABNSTrhD4mMie1QVTz8YQXTVJuC6YRi/iH29bhB8aBG3ZbTqt7Do32j/IPf4XeQk
mNz7sNmPLYOI2jCrTnM26bOgFtdcKF9kUUIERyZTGbJ04YNJ+uJ64mw2peoKNlsa
XKTqy0RmVwqlvpk6mVPlaixfTQO2upASAFCAb2eI8O5MtBPD0FT5mi17mPIIhkK/
k4+GNFaP7kGrto8duI0/cx65rtAB95BlzhXGDFntMuPwDFsf0H2u1CKmLquEvyQ+
0BXsYzfG8nu75zW1tfzVmBhBrQ4wvMTBkK+GD9XJyjMCgQ514LLjrMR9S3sGG/U5
taCyYPvZfDF7ALIET1aMQ6HSNUbtd25MB6N5yTtLTJ7pI1XdJn0f9Rgc3lvY72xK
5iUFfqJIrzVgu/4+pePTp0EEVktRaC93Qkd3gS5ZSFvAtJjDK/7KfAq5N3tNemzJ
5jjg8AYbbmoQ+Ed4b3CWJFpAPOitLEPoB8BUSZ9lE0LlisbWxH3uXyS7Ru3YnZaQ
NSvjat3kxPea8XnXxaTzy2uFvTnzfIodkRs0KH8PTzhdMwDEYGWUxaEYL3nM1YsQ
9WdKLThORNoJrub+ZTxKW0jCR2WmLfVYqYjPTo6eoWQ67AWprXDr+KgycFF+8+rt
Bt5HJ589de3ect8cXG1g1fhzCnugZXZ1QGFplkeUKopkWmSvNedZnjnfz6PZbXJe
zPzM6aLvuEQbbDiyj8bDk3CF5ZsAIWBVeL25eVpRyxu2Rsr9hlk6Lkjo4HynO2y5
J5EN9N482sbSHq9toD5KqWIDwObrAiK01TIcMg0lxejpEaUlIjVaekYTzoaweJL7
BhC2nOb+pNi7+xEccySZHg4rjijqbjq9B2vCf256LPJTd7u/eznXpDUZyLNMw+s2
fd5zkxR+hTzIFJyWf4IdiRkZITsM2yy6KWDyJOhNEQvWcecuFzzzmZ89P/r87NtV
Z1FpXPDNTBi7GyKcIJKby4xPSs3uDgo/Z79OSy9zC9HNY48WTQMsJySDTRe2Je94
5YO1su7nMdtvWnmC/Xv1EAQuYqi9Ez053HmHsmYy2DPK6Vs/hzyMctPHr6ZDWERM
UqlQ1p3SNWB5kjtq32stMhkdwzokxWY78p+2i/uA7ayGJ0LA4W+k2blt0l82Z7Kp
J9fmRY9rTxIg4j0V14xtdfJ+sleyy4ZBNTu7exOHyCDpMTiVuXUoJCHYibL+mtQF
7DiwahGlekGMMWWmWDZxVDqjdxUueR7TIhuu/SadEd+3RqnxY4QX//WlFhtUISJM
exbnvGtTo2WSyR3d1dvhMm0j+NG/ejpF10rW/R7x5I4v6KTmK5E+tP31V5Fp34XS
70xIJdw+WuIpCmeEHWm/3hrD44Jd3E0mkKiOW9ESnf1zetf/uLQlzI6L6N/9bblN
QVrsht0tcupN0W4+DBiJjm5hu83Rr95ow9GGObVHDCQ0Oyul/vYpMumTHIG5rz1N
UKZCJpQirwctdSa1dHfvGhgJZb1zpt6YcblcuAnCjeS71JcVdz6gmz+9u8KGqHTt
VirOQAGwrYs6y5K6HVexSWE5pixtzjEbD82Gg9XfzTIVwgOAPXYXQHICSM7lAW9/
CV6meaU4XNBRYoq9NuBkEHGMfrtYGhbxM02kEXthzZVrdnisPoSJNdKVSbHd3iZT
OJkt0mBmZoAIXWoPjREholfnMQra7+vlBHoCbfQevLs3vday/tvlh08WCLrx3Ybe
zNqL4AQzKhNx7X/k2jrl2GxzmNTtF1A9vFtcF5EWWlRTZaDD2tBTivLEeqnAYRhU
BXpzejtqyq6F8r02E5YEb59OUe+wWMWg0CraxE7Ps199Sfpz3Ijvapbc6kZ341mN
`protect END_PROTECTED