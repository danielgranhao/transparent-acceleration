-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
cVRgHCfpNscHuCjzgMFPtfC4rbi9DqATd7tK/XV6F/i6BuaFUeJrIkww3/50gCeutF3XZTE8AO9O
LzjVGX9JFwd4IOl/k+6Du/jAOIZjWnGvjxlaa+HjezoZjc4kGFiPpBkWiklmRCSOAQQFkuRnh+mb
MTavl6lse3gwcf177fk71a5mUYdeO4KXIk+AgrJJBbiDh1HcwRYp7j/czJU866H6bfcPyzP7Rwz/
dsU0rbDWuFY+wPh0yQJTqkmkVe0fc+0OFpVpda8AcCNtGX4rLYIwKGCCWIISWwEQmdLu8U995rAi
Mv4mNBBGCzpeeqwrBUujiYTbYVoFfKBYi0TTHg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 42976)
`protect data_block
WpZO4XVmde/cmvIuDDC/inIdZwx8LueLngum6DIH4B9gks/ZvWVaiEpHt+M6aO8Sz26iGIa6b+Ff
0sk5MKUGd/d4kjZpG+42UiceA05VgSaYzkFmHDr9gUSgF6zRzwyBQ10Vv/iHz1Tw3R7M39Mlbr3M
++yt8XnaeTyVshZkt0cUsOq4h1HWPH22Q6vUb39viruykm4MZGG4g8V0AN/xbu1hOdsxlIjoqo3P
QoluVlLlQE3CjCZ1drU3hMVPHh38yl4g9OuLl7XcC8ZTG3QMB9nbejTBVPra/eF9ZqQ5idCnaGci
u8Ax8S9FLcq1chn+mQ2CZWxRKAyO94lT/VXKPbrt01NUxKLTXDl/wcEUA84P/tWxelVPvw8N0tB8
Qs1pO3j/n/sRVddklEU9tNpPkVFKD9I4Q4m0Gr4VX8o30AvlyagRMcHVrXOrKEu+5hJPaW2wUoIe
rXgyB8DLiAlt1LnnlZDZXc3KvkhuQ4zCujvS1cuL6N5D1zMBwgYEfwd4FT03eQV1Eg3AtaeA2KgG
2EE3PqkgQh9s4/i3RcpBb38zQxJYCcnD3Jg6z586t1mJbZd0a2MD5Ku2vTAvu6BTQdBpghP17j8q
I+NpSXYOHeKptW8cnFqSYfhUKfryFGY7d2LdyKyuATjTX6DwbZbw5kOc1411y7boUWBsi4W2BEBk
+68ieY30JMob2TjucFaTaR3XnAKrewqQqjwjQRZiPVUgicdKkUylsp4lOCLOzYwZLntqvQzxqrqg
zz0Qnn/Ogw3I367xESorZd2bfvosDRiBOdqBXWAySvISfbp4RTxHc6/Qb3ju7hjZQL4wj+wwrTvO
xVvDLVbbrcD0gHMZ613MpOkG5eH94sWp6oqSaI+bTvpJ6FY5rTHN+uuLI95Qpsz644xC4r44oRkj
eGWkVqrQX0FT0gtZKS5pV1nb8PehB1X8c4dIz4YElg5rOn5CCqnrtP89SQYGB1DAhE8hJCYRmEvW
NOO01LG4GiMtqAfKpxTWoFj6fiJVBbwSyE/fNNH6/ptWDlZizXPYbJc8wCIF96kJ3L6UB95T/G0Q
Rvb1XvYkyjXAozvRur8ELXbTTYbAVk/BaDNMUV5lK/cBtDUcKUpp0oVz7kEjuKktlJ7A+Slt9lAp
+ht/CUNMFrfFRSYAGCl6x6vPKm1Ahn3ecitbpDCKsgrB0gJCwFXJikcQXIcRgiOBAYtpzvSusvQE
eprhatls6x3VSEfczX93DHXPVcrkymLDvJGf6DV6fR5355M1wLoqu26x0PwG1G2b9KiDh68ivPkK
kkPgmqE4ovuynhIR1PgPfiGzXrNKV2QTur/RlmFQ1jalmWFGQfbG3GM9ysDMnZxc3OajkkXiLQFp
wACwXbKbWcQoFHtHxxS5PHcYeBk8ZY8cZO3JVh3dXTmp3nRvsCnuViDM5+MR6XOcnEpVupIELmIS
i9IsN9aQLbtRvCHCaskJ0eTKE5W3xpJ7kvP4W6EMhYe2lh3Jqdj+x5FGoWxm6A8IOFZd0NUpl3z8
Sbbp2lW+IyT5EyBwIecK7i1K8rZoE1WEjXjHrML9pW/L6pFgX55KhLVUtbzZcx4esr334Fpabdim
qeCHNIEWDqBPf3PdHx4pnDuX1m68kCuEi1ZO8z8U1X6dZNgbZrhzjO3wyCByZbs01kefVhL+L151
PPmvYsM+XlVClPBuH+W1ShaV7DwwduEfHERJkh7TJUskv5yR3zNYl9E/Y2vDJM3pQsUzGFnTGuZN
XwCg+5FWoOW1hh2b/lv3df+gaUyqxcwSA1BGj20Toglsz+LrGViG2S2SUE5NPBRJ1WaNbLhLJjeh
lZzVtrpYSC9XpBuPWdAtT6pLHq/XIUxlrpsI6ayltEwtlPi4EvUdh7XMDZAhOB+aQPA8zPjzET2g
y1kJW2+ZtH0AOXzTrK+M2pnjTcXpPbEAy4HQkZ8x+fai9BBG0S4z2NNYS12misKwYnHZpn0IBYEx
LTlQ0zlCRGVkbOLxeobMW564nvoBDCTx05Y43ft+Qo9cNFG+QCIjCqPVblIKidUWRG3SXHe5UCrk
qvYGvsj8d1WOUneWKVJQ36dvP7kL50kk5Vt27ZgHNst4m/B74NjaxPSrPKJL6p0k56zoqP1e/f+y
IN6ciezYeA1Uzw/CW2PBUmBeIA+2uwzmjsqcy0j6DtKfLMomDePj6JD3PnA47WdFVvEj9K7SNqiN
mVqhh4TDlXYplV2pEXlcH3N50r/FyZsq7HxwlG4dTyIFFaeqZl1ZmzE9xGb8CBu8ILFqLrWqHdjL
5TpPsRhLKyDpIHQFSvzAGPstqE7k0v1SP4taXyp54AFCtMp6KvD5jQjacEGSjazjl0irHD21eBRr
wDDC7v8XKF6JnxfQwYun7Tn7ScVnCdNfNnQexZtpkNZ6GpGTiWA12bf+tE4hsyWBBeWn6a0J+TpR
71hpIoeHy0HiwW4iD243USkmQD9D8W6VkBXh1X5a3adg7FYyCYNUYssW2Uk1JfhD/QubpXV4jZuS
+i/SkP43Nr4bTAqDK9v/koiliwP2DpQAauG6zumRIx8c/OfdOvfpWIjIuu12kvaAtl+xg6KTM6Qq
GVSpiM5Y4H2k5SGw+lV/bDrIwD7lioO8HA110VHkf1msNu5Bd8QqFMCtaKOIKA26KtcFnBcN7VWv
M5ouW2J+DaTPpj04a0+vlWZkLzbGHP2VHTTAMq+DTOPuMi6AsIQTyjQnOEhyIzjditVs+fyvws3Y
1pSjI7FcA3kyAjD9lFJU/8IXPWPmZHKKj8ighxMMRWlV3Vik2j3nV+Yehs353mgAYImJdGAw6dJd
bDbr7fAmT2VNJ0Ms1uJlEOkqfhPHnVucQa2tH9B6+PvAyvUrMaRbfiOs10byM3m+Dsi8BkD/Zuyk
jadUZ01TiII1fc/kGz4S2tEc3rl5W6q6VMyJao1tkCFYcTJtJoQUGw/mk0Ca0w3pdAWvVOZFBXwX
eZ2vsTaIjjxYyC8LmFSSbnemHNOYjX27DPPinJl3qxoj5MiyA1xws5oEl1lyaoLJRSAI/7y/5BRQ
CarxV6jTWNZTQaIkdg/g6Z/SlTroKRZMr2szljP4cQTDTMLXCv+Ii6/sZMZKzFQUqMxRHEDO8BNk
EwRs7rIydAtLMGRqZvlQHxB4pa/biLEAddSOxa8Zk77jhbJGeY2Qd7HCHBZlbPHgpc1+P1fMvGwH
1/6dj5ywPo8S6ld0U0uO5VLpdmsQ+ZNUqCsqCpeNMTlKhconFDUZ6Ergus1Or7L92i6T6OwHlQv2
Fy9THuoBbp6D4LOKeur6VLMO8mxUbN/lyx0KLjFNIRwO6dNAyk67mBXubt6F+iMajs1qsTjHce+U
82mVQyqpHjnJrnUBL5WBvAPjrrkfVyFFpjTP99sX6g5vBqw5yQC1UKrkhl2YBn+EfVRItPi+Lr0i
WAV1APtIHSgHRdnbhVys5ixlHKjS4HkNj+GPeIcE2nvC4BSxjUaaUlZcxJ0txmcc7oqHkQIMhj+T
kwnBxb7ttOAiXM9Z5hdCTcuojuu2ugOV4X3OOoQWGNFD4JX6FnmkXH6dxp/7cNfWU1NxmNMrBGdX
fuDo8Cva5wCNlzZTsph5k8ocOkMfU0b3uSVDiKLCozU1LlNdad3xWv0AmD2dJzizFk811du/dWdq
TeLt+ds9YIsUnBcmbRqMLqePLoxWotMzSmUmFcOrlRlvtkHD1OYS/uJL+Uat2pR4VVuwt6qWZCWv
tLk2kq4Wvwdrp8r7nE4l3F/5OI36TI/ShpCjP9dVwqhuC3y9E3SGiGTtKqOCSq9das/Z4Z/xorEd
7TEaNLoYV5xdp9d0MFLd9vJDhmNunMQSqmamKl49FlW/9x7Sr4Tq90IzhLffYUUFxAwWlydBSish
08l06mGr7izZ9Lw3lp2rsbkadLT/EQH8bN3ptvPuneDsIfWzp9BAA3RiwyWb2TJPtpUH6l6FZqbF
8BPpKFKvrlkKxjXCOEHTc35GLGkgM4TeRnpPx8EuFtlUmGaJg4QAhPFNajCkPalgeo+ocnrjfJfm
syl8l4Cnvr/YfFDzOFXMhDmBDGgMPZ/QRn7oo1EMVsEe8GsSthn9N1vrjwLbBXacxcKC2HVoIuSo
zkWPbkwebMIR/3bo4Hf8s+EBfOVxZXgESz5qihRe6/43N1PD+Zb4vRd/hso+Ls275mTIfsRjpmbc
UU2k3nl2len/vNZi2sYI28NQmPIGEMxJ2xC6fJ7CyFI9kcrFDG8JbSKStsiO+iCZZFwd1SE7JIsq
RbaptM49nv5zefSI3srcB6lyOjVCoNJIixL0aEBpa/2UE0Bl/0iTyj/EBBiLT+12PhhfUaWq9WWo
NdP55QY/Y94HnyUjAk3bmDzj/CGzDo7dcuCnlGcTbNxqxGor4Zr8C4iiQdxH+HGHzLPvQuSYlJzJ
Fb7UtHNpCVdziWquTW8feoec0XZdV4Kb2eS/zaeam0MtRkhhkx4+GlpOOK3n/m3zHvPvBpkK093D
GJr7hFCrtL8U4JaGsGRS09eVjEj3ZdR4IfI8v0Yw+RgEoLv1EsTX81Hdank/Trc/gayZ51ViP4PF
C4C1aAceyfru+WNSSpJK7Xrh9fz4WxgKB/r+ld821/ZQNT8S6YqF7rYYidX/PTyqm8B3JRZXlZog
wrP+54OMkG5oKFp5Ly9R6XFWNef+rx/KsfB62R32Cwh19T92rnIaG1iwPWyXFUefZNayhapMg/+W
1AO9M5Lr9/L7NTX5CriHPm/4BhC6zogwm7sxVr0z6zjxmYLP/mhpR1vbQ/6b68Q84aNGs0Vp9Hhz
hKGYH8BqwbZHJtP5fQSJF+S5hwzV6Ed7jfSzuZon9f6aizCGoBZjF5cir1Xz7+98Ck4md6DIu3Hg
IJg9eCgKE3emtIb3tg+Yo/Se6qkHy9yI+EjkcHkTCLxMQKLq6Vv9eNslc3D3OMzxWJQn/w+F6XbV
nwC/feVJgBRL69sGx5rCerxd5KKi1DNfByiit3R50TGQmCOW/47TgRxGd/ldG9DWrQq9yIm/iVKq
ENHnDAZxT92kxg6xs/shXtaCjrpKnEpab560hAN1JfbknYCUsbp6+YRKPP1mpbT+C8uaJipETyES
mpUgNhqyYHXyJ5DTnqeXZIiIb+kPtmdMpjwEKsSUVHW85hzslbMXsEXHz0byG2+Hg3OkuxGUgMmA
NG1pfQ84uIMXVm0oCoJl7yKuxX4J2xvpQKtY84J9gqPVyygyew3FoPdXHxaPPP0iw0C5RDDh/wmG
o7NV3DCs4YC8tRgwdVHV8D6CwNrfz5Xhb64sQCOyxZM3ccrtt0C2OyITxNTgD+EOg85XBSQwAM++
CSzoyw0jnHd+mter9kKXj51WE5KMJp5RprqGybFyfR25DjZvhjTpDIPwMIrB7wTAtw99XDsui2bk
s/p7hqfZRpzTTR5Hj8HZWSXBLHhlpboQSHToDNME4OWS7U/AqQ5lxkUn8/nPaSnNDvKFD4UuGiy1
FHqfsBm0RwiNsKtkMFfaIKQ/1f26w13CisWC+bk/eSiQFud0v6WZtlbSE15pGsiCBmqZbwHWdM/o
AJX3Nrhb1bHQxJ5HmpgamxMvN4VwWpltif6r9q634Z/DZyMJtsJ8tYXn/fi9CB9dlMraz3DWGKuW
TCuhmSXdFdEu0K0XkShKOPXPR6tTpGAgbEWNP5vdrn9ZUGkQp87nhdABdSVXQJkkwz61wbQnzdrz
jsc9sW7cp/x2FfGxB2sT3bdSBP7v+JNNJlAG6UfpQ3KGKx/ytNIYvid4qDqf2BjVnZUbNjcTwmDQ
JVO6zZdzRKUabS6gRx+ZgFJ+BR+/LzI/kvE7axa6aHZWrw0M6lIFDN7p0ylpQWy58VcpaE/7agzm
6IlTF2N7VY7K+7MHNQyToY4rzgu4/Kah6yr98t/5o1flD1pbX17C2JMhbz8ckb9lkq8++3xI0K8D
d9eZYbFVl39PrXY8KCvouNWZBbVong40DN9GUUr4M2UDkZ3kG2jq/H+l5fbTGp4b6QT0BkVV1PmJ
81RSaR7RbDnuZ/tRPxC0eQu44n5OVxuXTJMzzWbtLeNBUrloCHJCzanSkBcNAAHjkNhSqngF4lB0
mBRzaGuVL+Oq87RSDYwslGM/Sr/CCQ1NaxPa/mLM6q55qfjJ+USEUuP1zgaBTeZerbO6x4VFmoJw
wm11Ul9ttY5sjDqLY0PDNtW0e5Ge7hynmgIaAHXTofxOSFFZyy5f5XdPqVa5+6bHSMcuJEHmIuSn
ojqFzrB9ss1HNu6uZH5Hdu0K4u9uoBc94ieFn/dODsA/k4NV0xso1kZpT/J9zUUPWR5usB63ZPc8
t6tdRwHhnxdM7kuA3/UMS4iNEg2kGojz6ga8rbmtDYoG1ph0AYDU7HZz1WkDQd0aTgv0RzFZ3r7q
3sURzRXxd7zLfYzHHwuqoRIpfJ1VT1GcpVpfipRZ58iEHk6/nUdNfPZ0JEx7WxNzRIR4Tx3GA7kK
xAykh6F4bUI9hxZ6dBb6dLITBxM40BqbBstwr5kWyMchOR5Ipwq6PIxiZI3xXWxBzaTpeApG+0zm
jnVo8u6YpZ82AtuI2zQHKV1GP2wp4mZj7ruboIiNSesrCXCi+1G1XpLza+NvtKooknq0G3yBT49g
4SgLfi8wGqUVWRm+kFZqAw+DXg8522MbmDz7KuNT6WQ6KeYIJiys6jZjKZG4fvDITDfhgIxiZpNp
2Q9ElNi57jt0MtlfBjCeprNMht+gVO66G9tLCwOQYWfFbOGiqihU+xmjhhtm4o1yaOgdzLhGNcLK
wpJt8zxErWMq+98sce/NlGBq/rSpkp4oBnLp9bB/R+sv9rTZjU4BZA5k/Ow8bNdlMX2DYFzCaSZm
WQRCSyFetgTqiGEBz5UWEPdvOKTbc9zJd/PlrVEmWb99jhQiyqzk/5xP0/FCBqy5OWq1oZKBPeRE
QBoIT+noka7N6OU1Js4gVep3XMTzF4LvrPlyxsQ4t3A+dAZ30V+0tClEFP3FzL21Qk0tTYXQnI1r
lBjmHtqaafSEtPG4i5MoarFK15DnrOjozjN0Zt2TQAhuc7bjksbkmlbQbJ65wm5YXiNf/fRfWjI2
mpuzcMA4HtUJGBARzM5crqvkt9bTqMrwpPQo9WUVdY+seQ1akPQ7BVLD8pLMeBzbMLFGcbgcJ9+o
HTTV+Yw/I6J6naj5DX2k02dsWcBDvwJ1xr1aZhk9BZZ9Rv3XMP9E/PoyQSSsL620dMqaUYPLUU6o
NuJZLTbGk/ZlS4+mn5PdmHgXEM8BSxvCoyRWlly5kw7i/wOeWwm7w2oDpfTDwwTYHlk+tUk4hLdd
AxAjJ+xxhtL3guWfGK9p7Neg/NkKPOMaHtGaRZeREOdGeHb+pcfKYs9nxsxC9P+wUEU3zctZWZn4
PTTU/ZIgdxMh8iQAQWSOHROY8AMC/aXJd4/T7qXBF/hww8SXCyViIgchGy5YGFONF6L24V/pKeYL
DITgDjuhLFwz/ErmnPDlu0F+nPkxmTRocp6VQ4rmq15fs1ROxKXy46i05QfaZnx9OUOrNfI+Mbgs
JLq4n86D6FlgUiC9+qTxOsm3HXdQiuYB/lEL8nsMP1skUyzF5QigWRpzXWDCuKTklfzkS3PjQzXv
qIjPKf7PWIt/xfy8nDAZBK8BVMb/JeqTX/mqqPyzxHoWQmovOtTppS7oVHKciPXTDO/1HNlpEpGz
O8zsbD1yhHGQod0YEbzmi6eQkAvUQbZg6K+6WSnjt6XhqDg1k2fImaTtMxJQKUTeA8ERAT/MFPv+
/yrwMDk3xZyAxm8ZY+ZDmdPxT8AB5B//+JrgfXRVmBFqYOspuelQloVti8YppfAyxpQ6bUWf1JvR
QMqlC/cRbQvC3MursPas5I7/JRJTPEOQzxQuIAGoAY4E3Bcp5pS1VM3CODgAx334MnrG1KYqYn/0
g2mbGOIf48otTtLtp4dPWEIp2EcC7JpLThFf3ZJRCF/68/YWxzMVh/Ibgh8AE1AhMUQxdSdH0q8g
HJPp4VfNPa675uEVRQdMSkKnP6JD0O9hWpYr/5jopY9PnP/AaOuX4LkZoXfCEoYidDcxAGBIrP6F
0cxaD+5lbqhW1jCvSS6ivdnAtSMQRbSDR2gULzeJRmyIYVrOtF/PXFyJDRY4NLpkNf1gi/kT+Uch
hULIzkJ1nzgVRH38f4nzt3iF2GMeGpLKPvADlosimeyFox1NukPBQOCcbwiv/JkVvwtADwGlw24b
bP6FwsE+GnwL5Ug2mwzhqGlQHDvsJG9DMuZk4/hf1yZJdsPJyPghaBuXej2oWuNPKwUsntmt/7Xq
U0BqOUaWj+QpLc9jiMut+WcAcyyo6mFpKbEQWkp0hx1/D2irs60J58D5Ujgf+QEdCJ91BdJ+8g3Q
xf8nFDbaWzvE9R4aTQcsfKPYInTnVaDAfx5xH0DKpfv3RrL/MQR4aGgxhK8ZPkaCHiPwd+0swVTR
KSfXdRQyPs2oQ2v+q72FZeHd5CWanlzyZ0f+jBMhywI3Pjjhfs0qbjvdO95sit8bI57NEjmqLtEl
8azjKKQN9hrYatfhxZGbGXexNjc/fnrVv+4o7LbWF2puetOG27XLXNlRvGrM/UZ+OPvKFHqZjr+E
lBW/D5nBnUO6YE4OhvfKRQ7H/vi4QZdlNwLAuZftbUz7OB2xS+DZ9Ws5mbf1vS6qYIfBEruRnsBe
Z7Bo0lXThgAMrVZIUhkpRmy9zqU0+MltMs8iAmvENpQ+Y7L/hEOzqwsX4Eekw3ZuHb9h0Mc/Ba8E
qV5DV2xvmQXBmvk4SjYjQDMntvfq3gd/AlsqrWLNWYVJRAEkKwHn+umrNe3zz1J1JtigQIEGOpBN
wlSF8DlfnKwsEcBvcQkoExJg6ZMqBolpiP4smyt5y+MHutn3HYfHPXhi8Z+t03kUJdQNEfYDPrjH
LnBcUu9GsgAaMMuBzsVci/2R8BZ62khTD4h1XSg7hgxQgeZcM4BFxO+eOMqilPxQu2R6w7J3zxUo
ng0bcZKBkXoLn1l0Xkr77/c0xiTGJFwivG11x+FvTLwAw9WTIGywzW0+4myGFfKRG0xzXXoxL/rP
QB0TLoBVNcduNWlt3HyWlTYoiToJOdgtZ3RpDl+Adkf2ewi4wnb6zsdwOarA2O+cvZ+KM0i+Niqi
nTBVA1vr+OsGP9nfouHWgDY24yHf9vemgM/VsRrYkN+8fZLLCKAxXrfhvCPzkHPI5QgQGANI9yOA
LJle+ZaVjJnh7RMNCOwmtAIMtCuSLp1zbI5Tc1l0Isu5BNQzbuwz0PqQWf28392ZUsnVUJenPUpz
pU0UtN5ZNIFMCp7ahA9vOFI2sXuUjW07cr3GWnb7+45W0SzPrUckA0qjjFi/2EjzDtq6ksUYJPti
DHPRFSgTBbqM6QjJqr77ZdTd7DIxxP++LQUl4jxAH0fSPIqvjnxIN6/3gSG4mLAvXwWU5KIVy4Kj
iA7xIUThBh5rAT5SROQqu8SBcgNi2230G7KvS8fvfWtdZsilS3E3hFSbs65VqFkGudxQwXxTy8sz
Z51aifJtHWqDCA7S/OavA1tYh5r27QWmvsk12/iZapR/ZHEub78F0qBMmf8E8/n9gh0ibQAiElxQ
SOztrYkUodLAeCxAIYIsuBinrCeOKXo0oBP0cyb7JWPpr7+PKtsOHoP/at+eyrAEdmbQMVO39dg9
oAbkQVkOhkQ2SVvV6wr5WvI821mfPGJKIqBBEEAzLClYAaY8t36Ak/qcJUWsGhP13ER5CZ6W+D2a
TS3BxJer33gSchunMv0XRAMP/PGorlykdpBD4ZQ1EJ4DFtDofJTockjdbZX5Z0gOFAwYrNuE8fDi
raXX8LWzOgRS9L9A04xgMVmBliCQ7ur56H24R8ZL929jq2EHlhOW9hW7BcbCWl9c+epJnjRZv+Kf
/6r90UM1C6a3/hqp/gf/S+SF5Jsu5l/UsJrEllXa5ca9YARL9HFzGZx/LhKdHqnFQlvdEQ3Q+lp5
q8xYV/TYwwtJDL2Tjkkya2bEbvRpCNfiyfpOICpoDmFRQGADhJxPgpulcjX/Cr8TTrcMwd5UacDZ
RAQItOa8mGB25lYD7C0v2bKP2IAGmyhGa+ig6+Hz718KWUbrbRAD3hJGsPUfne5oZWn0zun6toED
M1ZNCConnFFQbGD3dkPXnSPUeA64Gs4VwI93X7c/R3twBEiuvRUH8m6/WmNE79rRYmWJc78nCPqM
rBmBLv35/GyqzjgOaD69PmUrLhOCIeL+FSX19RiBBmwHc/LcS2Gu15b+H29l6Aa0IedwMNmWBWKA
uttP01luGUCOG5ExjDxUqncRkt+tfubrgT2jyqL1e/w3fQGQKdnfIsbWHqPGjvMVx8u0PAFlnFOe
EiziiosuY/0xr/ZY7EcaViWwuoC+U6xgtgaxQXpPzdqikcIvBZwlzPwbpNTcNunRu/nCU1yIK2lR
q8KJZPtDThFxhCDcyZlcKs9fFnXLpOMjqORCQDA3eT5HTq9c78t1/g4Vri6oXKvNIix62V40W1qa
WCP8ZxujcbOIihKS+ae6iS45b/BV3GmlgyaxeNOY1YsvFnM1BI5o+niDDQMJtgLAVQHSkf9KQjkL
hyYRvC2RAVVfL9B0F2wf8Kxn2HANjbgpW002qOLrI+UOK/J95EP9c4Fb6wO0c5Lgg/d30oFvsWCk
MhDWW3PoI0JkC//TNy5L4hUycJKJHshwOBBtu97VaigNNr9hVfOu0CSI1iLP0OM/ckflXWj+BBeO
8vQoithGdUAAoQaVWI8bxvQhk2F7CM+VHb4LqJmicP0VZHUMQXRIBnmQl5nAp76EYmCj/JUxmM5Q
zCF+An7mlRaSk0kdGw+55PiDbu4GG3fnK9YD+rqg2wo4KfNGcGlUO/9KY4TSLAVcaBX1PKLJqHo/
+GzMY0sYsRjt7wZOE8eUGuUfsK9bosKj0Rv7aM2/VyFF2kcmne5RSeF0gt5mtoV0p7kfazIWtW3L
dVT1hcDQjfoc2Q1/q7a+Z1EpKUcupVTrSIfrQIp1jKVtohPTeEcnVpspb3gN7Pb1pHd2UyNN8H99
N8lh2mwipwjvqXsxlSk3/sEd9+f7xZRHN49VzHV0vJdNW22Tjn+ASqJNjT11QykkoRlUat5+VeOC
pv044ReRcwytRDRQ3okzFoaIq+s0oL0o+TS5rzNO/5S/IByBkYJ2YnQEB+GXPY3YlOA6dI9otMV7
Mxy1vMkaB+046gtRKhup8+Y8kpaxeyO8CQcwIvqjYL+t0wbzoNAipWA0UAiUJdJgeyh+2Aus8oPr
yv4bG84BgQgaQNUVRnLNWkKf5W4ghLXm5etL2k0RRJ+7wC426f4GqSMGaSKfgyFK71Fo/69FAppw
eIZJOy3pN2Uds/CMoeihNc4yglyP5pdmRfl5qWvba+z/fsqMqHuKwXL0uE4kchoRi88jGWFC9qZQ
ZgGQbh8e7SfXm+7/YFE/+MyUhkpgrCc97NLfXmsayTJVBYE3k6Kxd6qSxNQ+yAc2Syhk4KC34vNh
s/whiG8IDTd/1ebiZJ6A52XSJQXnUlieC/b44mu5j/xUv8ZiCFwMF4Rd81/1LxBODIZC8kFGFPZn
Rg/jQ6kLAbYflpDVTlhOPdN2Vsa8CgcCBXPZ+HnL4QvZkj3p/Wp5nwmyblAyo0dT1xTch49tsXxz
RdwePnukWn5kndX/fEOSCWTj1R0dv60oV0xdbX6Hoamue2H/YVfMtUELLRXFVibcXgpU5q16Zhga
gKLK2eJvVWyEOe1r4NRR9YnH1PK1EEhJMwrCtmLBhjpoH2j8ltWzwIztVMcVwZX3/VpoErWvSYdg
QmU25GjvOeNr6n84yqslkgueUp5GruoIfTmpevZOaif1XX9TjJyKRrrD0l1JpVQ6brysG1FvbqG2
WyrHtSnDlHCYAb9Ei36aR4l/NdcntoDObWigb1NimQSFifyMTYEk0Y9yZONQ5v72XH6yFBFhm5zz
OW8fV0EBkQfMxbTI6F8chEaPD+pQevCGxxBibr2CXoTfnUwvtgZ4NNP79gGgP9F7rBVabudjKRlh
MqX0+QTmbK1cnytXASDrzOmQbSpmxfVrnPxmBYKwHTpOqD+3DDlGiXmCjn0Je7BPEEXwPnHHRsRW
GP6x1ZYUtdWR163rKwB8PEWiNEr0dc06pa34hHd/l0C7ctaQmpDYnjhfqrBuZIQam/FHH3+GzT+8
cLEsnzKTKgRg+kkSMJRD3K7x9dJ6Csd0vpLySlvmfXeC1hL18gB3LidmbcGRH3U4o3Gdn0VwNLqZ
d1tRwK4g87AeWYtRdfLeVstEEConos+1hS1UncsXQirPJaDec4wPjtt0A3h46zc4FV19WSZ1eTIe
wXkFVWnhT7zYX/5w+5je4l8MvavbAIss97hCFZ7dyfwnJsr/elan3Mx2UDWYjekFcGV0hVt/D4E7
Whzqne/YOTX7KNwj7Sd9LccZWEIOKVxJ7Nog+yCYhYuNlABCFOtnOKHedfJ0i7+5TGa6AdbwxZ5t
6yaT3VBFWK5c5/blKAwD3pl4huLZ58MyZOq4izPtM3ITIML/61GWX/kVeNmkbHWvJiM8r7XYrAw3
D8n8XvB11sb7YAC/QrScDc3TaFvC/LH+dJ9j8PqMVbNge99l2RYycZK90HQunBb7RXCSU3da8r4m
K1bAbiv0IcbwAydB4Oekh2cKaIAIYw1lRBL8EFqYfROixpi4kIEbaxKlWdakzOw6Nem4tteo2qXg
/PoASyoF9HwQkiv1ggg0M87WTSgToU9TjOQIkSt/U9/dMPelrw9Jn7KvIs+NkCmTCoQRB0Nd3Jdd
9E54eYXhQ6WJ4L6hK1/xnj97csAnpwYUAf5XO0mvwUQO+/+4N+EPY8qTN7Ru+sDTWETZ5MDyte5c
xbPNRjX9o9ke3ec+/Fc0Z7QfkEZn5Q3Mv2JUmgwd4HSSZVI1KWc37zeZf0uW/WtZnbXjt1XxSDvl
8KwEGKLwUHu8C78kgn2f6OCf3UJu7ASJOJJoz6A9j1VQpOnZnoJX3q3TlxX4qdVy3uPdj02mzGd0
WVlFITcSYXcuCLPTvWlBVUe56p5YjO0jgKnQV6OEOVMKQvslbrHikQVDjYzDVrLIw8NYdLSKRTcp
HSAJ7v71qDr1hBdpATuH/OUjLvP2h+1uIoWn8fuZkonzJ7jYuPbXlkpxZjeCbmYm92Ij7U7qQx/s
hh22mrmZz12VvZnZ0GCQAJUENulktUml/mvUDnTA6qezRze3H3hStbYrgbF/0yL1bTB1SW6cyTaF
36lAu4jny8Yiq+K3XK83/LPP68ebf3bQ5pOicEOZkJvmfm4oMxQBQ7hIjZMlb6miVkYY0hOH1XD0
oaZLMivaAuKpC6stnlo2FfiKaTkCCIj9wGsCBsYn3e0H8eF1WfKmiaPBkVmso29bPxx46JvWdlTp
Ho8S9rA9+X0nxxSnZqAkEvTAA5/v0e+w3WXJEPQMNT+FyuarZCkozbTceTfcumM1Lao3dZlpkLcc
BuZpw5VvFNIMg0sEi17cVzeSg3iNL2p4lCkF2Dbwa3lgRxUOFHF/Un8s/QjPOoQ5OBx/D0ujuL+2
uEMzzganZi41qLnmICMHYrtjc7ONjBuJ6jC1dkKJ4wNMwoQQEijPsWl8XaAmtxqQaMnZ4FRCUu7e
gp9aBfrNnt1FCZjDJO0yCb+cAEwzR65kjHzYRTwcA3JiSFQCBmdBkPXwSy+4L3RJ2mTfQMDJJ4wH
kZianXeOqEOKlB+hJuYGoZWvp303F75ZrQ4GAPa6FV1ba+v2Q3mv9VMV5BqFaPD9wyDL0mxsQJqi
nwGT40wPTIuYYHsyq74VYTFUNuQT9b02/XO9VTHU/fl08tYWINtR71EYKnDNY2qTNGrryrmado7v
xO5EwdIFAEEm5mWFe4/XuYsEj9QWVW5b5TXwo5InY/HK2tjCTQ+vcPIE6Gunawl0N9dt6h+imxgO
2mKiqfT3E+1oY+11HxP8zFk366QKmROqzT5wjhpAunveRnD828PzAshll/G8NR/SY843LVWFbF5P
K+n/2K84ACJWX2NZF4eUEQFKdnryBwYysHxVBy1uYjQUdZJl0qCoa1zcYDw37v4LZHhXz0eDe0AN
Kl00DMfxUQCwiJ5hOlJcSYnI7UNDvPA/+oA1JAs7wiyo/RvV+IrLvIH/EEZtXaLU+bzdKqGVfrQW
UmCRQ7qIV/RiCaU66BZidswqy10bJjt0mvBSUOQxHfOWK+cznwaPHH4J6nvMsgKuQO4A9HlvGN3X
C4V4SlJYAR78Capt/MvfYuR9d1hBtfy+DSCK9qdxBT4AoCVkkjSui8rBSnk6aCzU8xOd6mCGsLXy
ZBC37T/WeXzhxTxrs6sw22/L+vnpwsJFQmnBxG7ktMbBwsjJq1j3OxB8IydcmLF72fdvO9Qhts3L
wev6HDTROiVgzlwn/c3ny1q2MxBgUaudqh9+yyEEN/7u3tfQmbaVjQnQ3KZ+6w6VrTX1ZbU+SxKI
3NwSLBxNl+Xmes4S+S6NK72/gIxVVjbGkVzJ6zqohistUT6XsPP2OzGDabh6ZqCCh37ApVZq4CqL
uz1g9oVzH7NijHQ1VHJOKcBXKcS17MRlMl0+mUcNBqRdYKgKqxA1F1icJaRsCi4QcLq0u3E0b3an
8Ebojj1ha8iyLXCOrSC52HHeuSqRx/RrSPeX62lXzs7OF82I0hVvhovSESvZ3gVAC4WvLal8u59b
nOC5QTgt4b+Px6fb1wWb7coaxuZfaltr8fDZnIHSx8eY4atcLuK8oOH6TosJyFqLgqeOsfjWL41c
xE4bkYI7ZPh++p3RrhOlI1PBLXfLHc/71rIhihnbfQiTkShpftrFTHF6IeF4E3CQblQkyOjE33AY
Sp5x4dz54Exo3+dJF0YxBhkgXBVHE+ZGWN/4rNA/4SXv7DR+Qp59kQ5QSQIYehhfPDINNjGUbHi6
lm0wxfcQm8E5aImgs589Ynvu2SIee7hxbAb4+5hdH5o6ArV5zmnG5nnTrhba+Go56yN+8H88v7kO
q8MF8jm+p+YtbZvMl2WkQIdLFwr+fsmmvLdcmma1S0h8xlidt3vdy9AxXTsGGsxn3IoH+rYiK4yb
hsHdBiNKRlqbf9n7lYTbEev9tjnLtUFtRfNtg5sranx7bzNUYbUldhyhqsVqs/z610beE6iOTM9g
cD8iy7tGda5lCnAZvgdY4BU77d7ksCSUAROXFTTUB6KJRuxKAlQCn9TL3euSjbKlIuxLw8TDscA1
6s8rbAqhvGkxmLUbAZf2RyG9HA6VGqOyoy4if20W4ova3Ecq6mdq9bq1Murc60SnA/Ud2VbuWuar
0XPDEGuZ/dwehQN/sv7k+ZJifi7E/CSP5zPRUz7smwi4zk+zTxUbCBdEbQTZoCKMzVoW62G2Xplc
s40w5I1Cf1oow5Bli2vPkUtk8EbZpt16OxBkSAyyc5J1/WUnx2xPbw8WN2DFQUXi2ieM8bQzlHUY
ZpdW7B2ezduLsuR64FgkEJFihOlFTtp9og2O87Yh4RxmzMf1tQZnRjsO0YVwAQViAaiuGb7jNcWM
1n2eeICy+SQtyHNM7qSgbiPdzQpV4ofWpzJebddfWlsQBKstNXQ9Ce6jw2LEJx+Xm9mpg1w6OAms
8Uo7xxUpXQKfm9S3viY6s+M/caz6/n7yoPeg4G68sMFJn/Xc0k3qtjFYqbueD06JRh+3tHdmJevc
Y9kc+TbY5oyv+PTfsgmJU0kOkg9Gksl533LVXAGCS2tLT5vcJz8+kqvrhx5slPJvqAK3P+/El8T3
JYHtt0PekLqbmf1k4W6iWcsm9dl7rWF4B5nPEoNYjIBwYb1Z7Pr/Sdr2chN0l6ws29PY7P3T7fjQ
QwHUlaKe05sdAGaTJA39uERWu0O/SK+RZGdE3ozbBEe1rGs6hjtXy+oARsZhOufGGG+1JvCUsLw5
XW7FPSp7gU6fViQ0S2PCXX1tKez0n9TYbzcIED/8QaAEfQ52A5btSg3XdO23aYlsFHUxCR7dHjd2
z/qN53n/BBzYXsfIOL7gCxAhM7kOTelJzpDm8ULSipRpzU/2+GxyCq5L0cfg3iWTnK//aBPrOMIP
F+DkATwLWVcqrrP/wiiBabHK/9RfLyOiMqE17SlHudPTVrhmFWJl8TZkoeif66unEgBU9pZDANQ+
tilFa9Sdh2FUdRcHdiD68AyZVt2aJFwLqK5GpmttAQXK6KGJ2I6JD+6Fblz2Je9Fk34UfJBEqwec
UtglReaB57lC1GQGkPjnPoAYzfCQ84iqGUgSI524pIfL2K7ZUEWrsm/m565V4zP/9aUHlqdGOypa
JfkcY/PbLoXNr0XjLuqrMkC+7dHZfwHA6KmAqgsuG1GQeK4QxFhlbOwdUBTrhatoRxADCmpSeWG+
Y1jZqVGA0EnPkA+QaK8Z3i1vK7xo9dRKa5LCKUQjysXQhnsBA0RuTqu+9QklcqYjKtFgjrg1thTv
9gikXK9X9eSXfAdI9pkeA06edokiI3HqpQJ3cTZRnqL5W7AUndJ7Aiy9ur/CXD1xfU/Zl9PtzPtT
AN63p7z6WmFAICSxPYjN+QAu5WRHfWPey46iJ9wdqyziXipwtSEL/sIUkVvEoLdXWO7rzQAlgklr
emJBboYqYgN1HtGA/jFUuwKwpZb2nKRR1k4lha/ocq6Ob6om2jWRiDRjALJetl9khKkz8e2HXjNR
ktm7n/9jrJ3C/inDdBAy+G5sv/Z28bsv/uZOB3WV9KjEvsZhghnnVMTeEtmihKY9oRX4vySO985/
ALbeh3FZXem+4ADKDBVA5hoHxMRLsYqsIjIKN3A0TLft3HaKnZeaJoio6GcxqgZbIoE1YfPxEt7B
qv9bkhFj3KFCiyJIfQ7HegqLzb9H8VJYU8Z59iMabKBIf2SUZBT3sI3VRusTpd3Nyf+zbsW/h8uu
5HeW3ciFu+w04/WF1hogOygrM+qfP2znI5TDtIOFfcUzhYO+SK4pujBauYxBZJqf1kpksBP7kDZS
lfjHWQjbnaKbgY0MH+B8XQIQcK40N148AEdy0Ed4dVbLntfJcbAaPG/mPV/ptW+YKO4AiRV4E9Hu
wRXPzPoCLCjK1b4X0nWa5ATXSoiGarwiFKLV0GOplOWrarhHNfiFhl3GJJSL8GVC3OEjhA0HLb+a
9588aJ1m1ttgS6yxZuDPKKJ76yKqXswRoxDEJR19wKJFPWjiXP7JmKSDiYVZdBmemXsXnPUMgeRa
K9/RzUKZIXLRBOr0fnf1D9u8g4DZuhqEqNNGnrxSaPUobAc5n9MtmDTcIRfPFGUb5cfvGfQLrfvD
OxXctK2WAkTIxu7UDyS+f6lh1PLznxv57RzINu6dAK54CYbUF27tkd78Qnsg7hDhs3100hnk+iBi
fZEsmAzYJaG51TtU+dlNoZuq2AVJ8xaTDNmlspOJlHjDsZdKOyNYQN9NNbFpwdBf9Z750OmrKCQD
1VEiDO+4fTYvi2sQ6uJ1qO82jnho2QUt2opqymdZ9xsIh/iI/QdnOobq8pIRR2Qa7jjHh6GkrIM3
rmDqAren8QTv+ermYkkIgZtBZZxmC/JyMRiKckWOBRIhsDZYsrOr3ULC2bD7v5J/EC6LCs8BZsb1
5JBf+IN8ft1mpxRqvstt+mSA1aWxGHnxyT6NwWT8xVt/4B5s6bdPhY+2nSUe9sYWP44xp/VmxQXi
Me/KeeRPL1RHJdKQYXc5J7l5TacNSuYyPyolqCRVRiWHLoqQXVosgea18A4uEjvdB7BQFOgq2T+u
8dwscs2VP79hqgJzfNEAtxL/PET9JZax7RlrKmhAYG9zKPHNAseYFa3FuPEvkDFBQUUJVtnGmntW
EqmD5R7UVj3CJhwB1W9z4Yc5XFdiBBZIJgoB3rDxJkFX/qg9nqR43jdw1tnf6a0CLWdpHnEOvxUn
lEPpoRkWjSOyBmowOFLno5UCQw6AoLwO5BTg2x6I5OgXBqaAc/7JdFIDAHasJUMrSqJNlX2n4S/v
WdmYJyKPuFiWYv/gdPDJNy36c2iaKqZstBK6fYiqqU4Ox2C5nR+IkFc/EFZNyYJanTvqWiLa9QPD
BMHLN+DmsJNsBhTwsKaW11ddR0bQkpQG9eZ4WqYfAbo1Ap+S8hi5JujB34iCBe2abiSHf3C0we9z
dykAUwDHuRBkhXA44xrMTsdNvVp3B52u+9JkJoSQ/51AfwwMRzkBQWGHajJK5l1MZAngxIwpJ96X
YMKK5vTPZFfhjQoETDCwr5PONL602dWnxRXxB/SD1gv7cQW+bC95bcvr/EicucYI8XwTQNizBUTM
LoT5hb5O4re8cywumHcf9FZoku/UOuP/gy6UpXYEznB+H/o/PVRVl9WX8U3l6oxMRYE9iFeBeOsb
RoEFOlQgwnHroHQlXLoAih4qSPK6gNmoiej3jDphJ9zXzY29wzvw6MRjgLPNcLOmVvvwWBdtNHOc
QxZdMu5eHXbKtkUKEgWB4TNtuALS+ReNdn5mh1Qj16BsO/UFoamR64bluTM2gHGUyn67wWjpvke5
VrTILMUNVobgEwlraYMiBSu6omsXo8qR1PYNKpeJbYaEfTNzRluoYnlWEf4u5rpjMGT3CCVDN5/n
g9epHyLaPwjhb7vXaTh4GlbwM2Zx1fydZfvnv4VH3FSA+tDkRlKTQjN3PX+ZTdonZ4HHG75+7WaF
1gjmTjEesMEZ+uuZB0RDFpjzqvIHUbeHPQ4KNZDQVVwqDYxHOBCgJgD87QCojra5IkOK1QvMDweH
LOHAlILeAe+pZUfFN3fxFhwrzzWgjNs3aHTnxUb6ZrbDRjksxG3tg1Y+gTkblX8ytCtTFtTx2f/9
2MnYtYryOabKrbwGCEiGyZQMMd+pZcsT1pwc57HQ2efYBVMqztViES/TV4D0ARSCd2B8QevrgISK
3Ao+sdESrd3JkXzSqI0AzfOClKNtbUEjwHDJ+R946x+/dkir422/3lg+fQHPbDFEXMyYFCTTrs1O
RILqVX4pmDH39sisIhPflqco3kH/F6XoOKgKf9r3MwBP2IcfG5uQDyyF06g2x0bccNeofA3s6+ZJ
veuWqSl0DoxF9SEaDUafmGS59+bh1+mbiiJdYSgX47hB3XOw7pLLgLLtN2+WMrgkhWyUnV/vyEz8
TwfN0jHWSpc7dohMOmrEAI3gfdVOHSrdCwvhSuMv0wYztBmsoNfbs9HkQdBARiDd6+DxvLJeO2Yu
gPBQiPeY5YS3rprCFXYfzzFbMl7q0zNjpJS5E6W6fD/L8A0g+3iZOEvvzLhMUeJjRZuyGtTxqE8Y
/8z4AmI/xzhudhwpqXYU18NWt3YeobqZcWxtdOqvn8emrv8jtZ3svGbxXNXKE9VBFy3QFJ5mptSS
2W2p2P6E94/q+uL7stR1rwjXREjpLKjetVL45JnhU6j+tLrMa9/yfpAf6c24pkUhCySCHi5A3SiD
IC0F5F6negO3iB0+yqqJl8pyMbLT3jHFDS9lWSJsA5j8TTIiHWVAp8p8InsTshqJaTlosKIFMGoH
ZManWO8JFBi8vlhDgrxSCsHgtT1COrBmUclVR0RNXcC4qSj4v4+txfBF8lwNDyKZE0SGE/LHhiWa
g6gQN+2FjwMm+v+R41hQOgl7yFKIWBq21A2gHoe2gfvBgWtcGSH++Xq2cgRKOJ2EQM1G6GADoh4u
B9zbpN3hQR69fOTAP3TZiXKnnc9ObRU8csh6IYjOSJoR5CGWIlni7eQTKavcM3mcIVG9qfULkLbR
gRr4lQ7PFH4dZEU16LlYFcnWEGh/y4VpBMRuNATMwv3EcliGOt47gufLPFfmrijHPvyZCDCSV3PH
BhBAnuJC+oVGBIQ+jIXRapBCU9pNA8if/Bto+kRoCh6wciJUG3godbbuuXU0j/tQHrCGKZAJ8JkE
Vxi+t3qoDQqBuWQTXrxgyjd43xMFhDIHgJQKFU20EoHZOdO06hWZMNLDgOHHXqzrp1/TWgAU/lcS
4Yoq7TwkSsN9b5QhqJ0dCvpvowSuusAke1w5s66q1XGajyzfSWCRUArWYR23sVyDPq1zvtqNqyKs
/4sF6XIpgAPW/4zNczCTWY/QSrx9JlDRB2jM1Q/idCrg3+vWx6fkyzHFziYly+efJWLTzTeO+6kL
JTlUV5j6cu6pUWiWRu0Evpe15BzBcVcp0PWxrOMAJrXAGMngPixIcQ5cj8cT4g5FA6bTq2OcEbql
Yj7AgXagNy9lV5e+P8jWqSybmaEwdQK7go4ZfZWYeXjupDILxL843W9smnADd0FALIMvUZYD86eo
hEIkMqQxG1rAecWfOF1f4JhpAYzKc8Utf88EF0ZQ2+wP2bmcaL4PoobAlnBAK8RaWOpfdu1OH9Zf
Qj4z8QCrpfiRQZfdqeqaSSvgxQcbYB/gszMVUaqRwuTxITxEFPBxH9vwa6y6vDdANmIuGc676E3m
GX+Wno6gBke2PDzWyNxqK5E19L81HV/JEbXOc8pDkai7DRFI1OW+VzKef7TFT44CMYDAhUXsxx5Z
pyaY/pz268CKsknr5T+q/vfo02ahO0RSgc/mWoWjEHE+tiCTi9wWVzvWvarJ2tJl2SqLMFzSg2WA
JGVsA0Y9v2pnN5AbO18624WiLABpeMph2bbu2Stuyxbuv+fd5e3D0kD9eKV7ENsinxgmWZY5BGlU
qrLM90XlneychA6fj7mqgJm7VnUVe8Q0NdsXAUUEmb4fH7NTaryY5di7F3EzXlm/oVv4xQKi+Be3
2Yn10fkaU5PWf5cNz7V+9x6S6w0Cb/OFJvcqGR4cePgM9gdSOe6QRVCLDpIXoaIozfVmM+Y71+Yn
X2w6cLaTcPfIKmBArlPMC7GE7EOwNFwFB/S7UWAZkJpeOJMFDiU9GSfYgrlpGcNHcioxQft4AAT/
tyAlyLFpqGF5pxxq0RXtjvnW/+97RkP8foW9asuf+SovflfHGZ7nNV/Rjpix923AVZhzvHczGISE
xxvXWyA6usLpY1TiX3BqrYtDqixx3mzPuzXUMz3PXP+LJeyWAVJJ9XaWTU3T+nUMQI5eqP3TopEu
hRP7wzTauQkeGFMnKqw44FcS6jKYhpU4IeAYnyqNvhLyFr2oZe0aDqeLGhgmWlJyEVn+peqqlrv/
B8R/rxySCMXpL4y31+/5ApuWhmdlE+0E7k9O7158YturAFT24CVmgzw2K9N7RaOZjBeQswJAaHkj
DJ8W4iggaYVdevWNnuyu5Xgp6fQZyhOK9OWXEzivR8KbpuzuASAaStmyFb6KXBXbcMi5vR6SBOZO
XPtKkHdiGQGmjgJNKUzWdgXSNAoAoh+hdG392htezg2ZK/bAVkW9D5FwE6ZTyNQjGdQ8TiAaAlSx
J6xr/6WeJMTl8LGzDokAsl4Y1qyqmHbAbvkNTEOXX5EkhdMvrl+vzwkhH8irQfFkdAuzcg6g1olY
6EmzZBi1MhuQMxM8rutWtZqZxT1mO5XGitfAdRahxFZYVQbXfzVgGrM0jHMm0c3IlOeS7sSZF48P
Yk7yrT9uV6diP7FZZ8XzF0+cSWYA6sbV2t80Tfm2GoQtAB3Xbe3H6wtGwGUCVnpmRJ4ctV9tImAI
aTPAKyjKUbEreyOR4a9sj+9o66YV09FnW6bxeTmljYHV/I9eJzzv1XL9hx04nsGJCVWy5nHnJo0e
xTTiYAy9Rztqa71ZTyD/sbBWQdZb9Py7JBl6DufcvW4BbnL/Umvjko7LWqpE+bsFfzsY8lU3oPSB
QVmZ2ufonfrKYxXkfa+I3uLy8/QxezyX8Ez/AY4tlZQpjuO6Nf+ld9sQJOYcjsEbpAPtbfPZlwbv
ZgJ11JEhr0hZep96f5Py3j7Cw79Fk7FYy4CGJRXFz83EC1efJKYV81nTYQ3jDWZkXQo924GnpAgD
qu+cGvOLZ0py+I8DmJgzYsNrESzBzJtworn+rlDVma2xoGqLg2LCuVHYYEFhJHilcEcTL07/edk5
W79mzUj1+b9dOP8JB9iZGPW81OvjVvwF9mO/Rfhby7lC7BNKGGdIeuWEYMfrEPFLihyK839BkKiz
g97zaHRrbYRMBeX3xbAXPrVoFsNvVWR2NSAbv1q7dkBOVNuOtxTKaN6LXdqooS5U73OyJSks+VzT
Kon2Fga2R2mZAwrI4SrfqYrE18lHSAEcSnW6xh0rB4MQaWqxkwa4bYFiMMaqXcBep2rh9yES0GKf
4WYJwqFbdWdAIEekA+0TE7QADJWM5fAnSeGU+CxAQcjwUWPd+A4Y70Jjd4ax0uySNzmPBSsToxkw
FtiPRvdzNNylIiaL75A7eZLPLb6ZmId/dA/IMfp07otLCq2dRwrFt+UVOTu0QLsbAnfeLlhhrfHh
4TjMZlr+rmIqp5fqMitfRr8XmB2b/wHnEhh0kr5R53pI8mHNqQWjEZNDDTjJBmmdTqQLYFOhLLiJ
mSXdGev7+xDPMWn1wvMTfzeZvjBnSOUf7DTXmFMoXq0pQtrRdLrP6GGXdBW7R+PvwSSiqcRAjeaB
OSj0kZ6wgCGjvaGKkSHmhyTk6EkrWLt9RbKbkcy19P2VeW/p8nAtrMxeSdHJsl1oVqjKizCmRGiz
tKO7GLrbY/U8vODE3rMDxoRiH4U4/v4W4fDlSI05wcuKp3Y7/p3NpXjuNv8PlZCmm8DbIb4e88nT
qztbucwW2iYIi4O5E5+1Lf3JgD0/up2u722nAHHBFUjI+7cu3+AbsHyo8cE64wXHPB43+vPaAJWh
2u4X1L8vyk6/dswqBxqSmmUnpdfqSwRrEBC4dVeFejFS9TS3m2Sk8LP6XDUoGO+TrkhiYiI7/EQ+
joe5+T/LVdM2/+gUwau+U4h/HipU2e8w/5A3fAKWpa7RUjO/BeYm7utWAKenfPkxivWa26uXbze5
2QQYwRK4vVcJD5a2CfgijACzwxS+ousgfbjWm8TfNPmCC5xhdkCDY3UWmYhLyD1aNELtf3VgCoMI
cY4LP+4WBYdJm6ztZ9Ijl39SnlA2+TSyHgXDuUOjqXkpca+R55oFIOYqcbjCzc7rm5QRDIc9drpJ
9Cxwn7W9RL3ryAR14cV7pxNQ6CGkDurYb1tXdCHg7OyU8M6HPGN9YYgcDqvwB6tDpAgxglbTXNC1
lhj9zX6uE2gpkXOR9drCKD/PXU3rhsw2kI7XKmgRPN582A3lBb/hhT7N5zYgvE8bjnQwOYiS4MRD
P8Cb/G/pfrO3ns7MoUr7jR/naZPbiM1r/fXi9Kzm8gkjQjYT8BgBS7E4ycyfga43Fcpd9/hSuA9Y
NtguoU6a99t+ubip4epkJeNnQaua4eQo89eGcgUzWiAiUjHLKCAjQ5Mm/1TlN1cQ4VvTDLC2Syh9
kt1+Ax5coy40AmPDLCh4qTZ/moZVkiza1Boa9wn5V97vE/P4OuquDOUI4EDKd/jSG1TotJh5hqWw
P0uCB0Z88vQFW8JuBeTdF0S2EleLUIZ8pzQ72OF3gWSS/e/nRMo3Ye9gcjVRDWVsjaZ30EFEbnRM
fBHqHtEvISMZMUuVCHfZwGCooScoFpNeFxNcl+4WLJQ1npzWKZmef/Hyoj92e1QczWm+Iapl/106
ajs/YnomnCtlvk/4Jn/L5UXS0DqYHzvtvKCG6OfgnNsQgI0cB6rF3gomniEUAP6l2kobSMVjmrLb
hVb5l340JUCWQVcaClGVX9dAUFuPgc+FH3iKOc6YjfRuoOf1OGLUIaKGx18MMUotxeN52d1w6HQR
BAFVHszfhUEGWw0+L+NV1WmTRojNQOd1AZSrkzlRnnQgwg9JuUWsseAuCvtMA/OR7qz+EE3f8Nax
8NV4OqJjwGhNFI+wqohu4jLbXqjIZeHeIifCb1zGJG5gM3Ka2102vAGqKQ3JJDZZlPmvXmqlN9Dg
qAQ4penUoPRBiWTYfcVLSn7rXJwYH9wzQObe4y6lpbPnz05Iw4BZBGvob3C4Vy8pIfukBAREe9yk
ouIZVScG5tNvqSWyDVa4QPrTk29sxlRL/2to1LQ7Tjkfs2NHUzE70YuFr7uWz66gNS6J9Qx/mVn1
8XjbIWCXBHcwJ8l9szSZGDl/YLVhHm0nU93U+TNvVcvlENIdiGPh8LH0Ws8OoYTcq1e3hjzd3MA+
DZzeo7MQRfAwPgKOlXbkaHnGJC+CsHasFga3bUdUbF6B2BGyvP7PxsZ63efgUDwgKkNZAXCSImHy
f0lWnbdzEAm89z4kHY6xU8+5G2eJ2jAT3VT/TYs1yBla7S/hG9bHwqdq7W+FIspnsXjOj6wXwx0L
b+cnkPUGCs7cdTlQ+pDgDuUt/wGlaE+xMBxgXexf3eeCl5ZDDu1ThOmJXFpRrDHJjHWy858sDjpL
X2qifEkYLpXNoFGPlJK3VNmC/mi1jCCtNfKK/hw1UrgHC00MKfqa1ApCrbYL8ohVETcZUVUyZj8n
wxEb3WCOqOe4xhvFdiUevP+agMU10tNOg4KFait8Ti0EDsUjfZeu5NhTKn/uUY50ytv0sh7cC640
eO/HHvquEEZ5yvf0Nv4fxAFebG2SlmnrxWx4Fs3vCIfXOTRqAW41y2Ibr3uhBL5jRFlZCdMfifEX
JBAKFilkB9nEAV8m9R4WDabXG6PMeVnXC4ZFWOsWHTRPM7/XF7gwIAzOeOyIFlVzk1CY/yROZxx2
XXLXXgDYkhzNfTy67y3xAA8/rc5cE2dZg8yBqPNNRZEWkpiWm+HSA/5TF9RSKQZo5EY1uF8dub7X
eqkzWAusQD4AKi9aZ0L0XE/EfVsDWZyDIfwkAHPhij1puwk6T+yr2+nYLx6IXEBllV8A0Bx6KTeg
4Ty27w1ZX1QBw8nF9nJgH6NXS3/e9bPb+EAMH+RBrGjFj8PxmqsAxJbGszArNo8VxxAAXGhL+ex4
fE4R+IKX/Dz4DdR22o+uyOAVbeeZMsDZ9Y8xMVw+srxPTaE5FZ2I8XnT1jx6tl6pxNFnHV95dQoE
F+HBFKfeIBuP+dXqDIC7Hd06HJYIBlZd+7mAvPkbZdjuIiYT4KCHw/Ckrudnp23JdsEd2APUDJdt
uPAwBTiNdvn7BTnFH8KOVexrVYCDFsRaaGqQQRn5r476TrQx93jsLTWyP/7u/yeEYRgQlKeSrXeV
q66TPWZLrs0zamAWhRWzKmskF7GkBlkoeQhtXyF8O0/9y9zzFZyV/TANgh4UqEntaj7hmwsUtYDD
GBG9FyUcGhSGtZJRctYwXjTSSfzifW+1jzyybqT9DpCqAlyFXx9rRQUvuFPnGJiP1Ub6DYetMvTo
Bt2OjPz13WvR2+s3q7ftO6vsMJzVPfziW2yuN7/ivp0ei00ruJ6qmdSyag8VSS/T3mIb6HHDba59
OyGXsNUN8tvqlfqjQ8MPSOfsGgnOjjtiCBTNnaL5592OwuG3ZooOaHrUn3AtX9MvvYgR3cc8i8zX
lZlBFEiTdPktHSyu3MglfQ2gG2PLSjJELgEPBfKOhYcTFwk0Ik9YxQTcnq6QLkfb33A6/HB63wwa
/NWuxJP2BNVencPeKH9HswRGExhqkBbbepvsPMihqiVfeWEsTvtDG9vH6bGSaTE+ej/1K6jarykm
X2pABzmgdeO/d75Dtva28x9eM4y7EHBunYHtbd8Y5TZZDMaM/Y3hKXU4CEkBOnfysJbp0TBlOt/8
xkqMr1ee7CvawHuWRDfAJCszKCNw6LY54Sjm+6YK8Dd0EgrR97VcdHntRhfFW0Zy27k0EWMysGf3
c4H6oDVCQqgE/O8AMg0whNLkW9AaB2zxOOeaKnrhJsyR1PkNVI4a2aw4bkjqNLY1k5ojiC8k+0/a
brS6ZZ1/6zkDQWpGDnmNYAsTSjXEBeqrzQo8J2/XcffvyEB4iFSagB4VHRnHQ0dlsHA1gDUUtgK0
ykckabbG18rn9evOBNHFkwp9+7iVocAEm2LcIK1Idym8Nr1MRB70LvUTwyW0q/h81puUuaclcRro
enoYxYId7kG0NKPYeyv5TKr/KqURy71kUSsm/ow0MOzKjmrXMDgq7ur5JGnbbeS6fi0nsjiOM+8t
LrS2/pOSt0OLM1vTKZtr8DDro3JtMlEPDuTWdHHZHqbJZ+ips3S4Lw8Q3TsH+Pn4ZwB1xHSfFfMK
05sJh1Iv6SwX1QDMYp1GsMvnh5LQVHlGh+ff0pUp1Du2ECsRe65g+3gmHUJdbXDE1MzcmeMbwE9L
6RVaoTOkmYOCkN4OgtHkf6A8IzEELjrC7n2gFVZ4pCF4jkCKiWW8BxcC5AtFiBToDSX7nsSzrM43
4rgTio29XE2OQ17umwt58Qn7O7cnoZBGLMS9Vy9ExgJXzNgi90HFbmrUZccauZvJWx0zRLEv8+ug
y5dkhC9BnN8Qoh7iDNkNceqEX/HqiGSOxlDyyNF5n/uJOg/bb14sPOKd1EDcnmnc8sXBll00wY7d
RTQXwDPrt6rtPduLiXH/izEQY5wJJp7lCtrcZzhp0D/ZXpwDFuTFqgrfTuRK2xn6EQkMKTEJwKdu
twdNyi+ECRREcA6YIznq97+xBtVobK7PaNAEkfXbL34RYwTLAuPd0JQzbDhDWFyDCH8zOVq91EE3
LY6L9SJ+XjwbHMOXpEGbGQxv4Ozi5X+egBoaXx6z9SxzESazxihHOloEnz5KyDFBPZvp1dajifDB
ubTVxu5uapJO2Mv4SCI348m3ds/TkVyo5oh86h3FNyX2yWbPAIPxYosivAeuMgpqfsHn6CBdE9EB
mmF+ORi4Y5B2zsn8qnMrZruCJK3TovFr2jY2XzvBO9cLfjaPEZkf99DvjYZYcQ9bxIdMs6xRf3lm
lEQHpIbTnyBQ8KURCgf+T/Bko3EDawCqgz8Fi6Aae2z92lF9oE40+uQexQZeLR9hhoywUCUf5Cor
g+/F0M6S2qdk0/UDuTJVpFSetPmQSoMrQwYc0OvjQMpB3eHiS+BBoUn5KD0DwER5QrytK1BE1v83
JYSeHO2kdhBhw1JBOVhrwNarIwocLAixH3P2CUWM9SpErEs4Y8zy86+QlecGobj1wLl+bXtIqaCW
V8UQ/1kdYAiNGeLzUY+cjNElN425hMl6s4brc1PSwAFQ++9dXqJQMJ1dEJgBP8aQAiTVVFUybNOS
6eKRpPuqPZQZNTG6jpd8FLWGK/+WxOKis5fuxWxZ/0hhv53popE1lJkfyqtpSDS7NIg2XYEpOWD6
XlupPJF7/5Nd9Nh8mgeW5Yyw1iw2EXRa4lzgRN+NG+oNpS/o0T12oyGIYke4ootEk3cnLgludmlL
kFI6dZD+UajC7eQBsjALZJIBemBxdQXqkJ/iUUmsb4LEzFeYeEcdN8YW+jNHoYxmpLdTMIno8SBQ
ecCrZHsDWCp3Sp+rUZJUrka9nU3Xcldq6CtcAZcCq9ROsZHccTVIZ9oi7Tq7yKs0AxlKqJRobrGF
52q+5PfL+zldlfc2Xj7JrRFYL/i+NOHkzE4Jnf2QPQ28P6J7xKjBYgWbOFBvdS5wM3gogQGaVmio
kEQzRfoaJfoa+mnLHybKF4qqqHRYNCMz7+BWXqkNTlEu0WUd1TVwJlQN5ZBoDBWOQ9PmdlDGPb/n
IenEuc/+JRRL9xWcZYB1mUl2HgbQdD3yuACec0QMwYSu1ckr8O44MP78z+/JCmRxvMozN6oP8GW0
Va7WCsXcVoXvH0wYn4QGnRj3zZ6IPZ8Jas+UxhBMV4qFL0ttnBAprkzhp1DxAyxwA/bu/wrcF/Ox
5zFjD+cYWRNw7IzFwM3eLmIKyhO28UwEBl2rrBngpTQtU7ajtC0RF+OPeOk5nP/PvQHA84k0a/QM
PJi0MFtUQjdHw5C8n4zvvhKWsjHd91Q3RkIO/jUalGMBqwZSuIzb6aUY+eQ6Bcq7QZe9700uRuU8
XmQhKg4A6f3aC1MNzBrhBBHdpS4CApCHyOvIzYXhD3A8KiI4hJWXQ2s833lQTzIMwBxq4awkvLbk
f+XJ30IRcCp2OGAbdiRt0RPxZzfTdnlpQ6MvEkiEghiwcb/vePfJw7vxBsduameSBKeWTH4Zm40x
ED1NXdlyzZ/EVXqQdc52aAJqKUUsFqbucT59txWZY1kBb9YtGb+xGwja3h2yA/SohDjdNN473hcl
qOaGl42t/rthxcBW5YbaqQEn6YyjaB9vJ5Oju8s3paSSyxw4K7EncKezbrH6IS/Hy5R0gs4og6Zj
CASWIQLlNuBiCLTrWBtoqkXyBLO5ekc4xk4NVCRsdTHsXnrnb2iWpWc1ImFHUCcAC6VTN0m3L9oG
zg9nlA9TYBK1NLr1uW4towuxXffEaKWkjSy6ymBsZegz8iE4d3Fwn9tshGlEil/kkbhY+dZqKIyX
zVRwWyu0nc/ZkCleoUYiN53euW4itNWHuwmwpYxU4VKqO4Zrq2U/H89krbD6b7AlLpYkeKHQHv9C
ZTI+7ighefmA4FaoVP5WW5BYhnkSfR55C3WKs6tZ9BfBrn43OPrD7eqf+LhnISNCoSvlWyImwX4N
L6rcCaYsCwRc5LnYVmjLzN9cmARwFeYSSUTv52NAoq3CQgFAzbSyAGf3bxjELdjyOQgo4eH0b3nB
KgZ0TAPCFEoBYgoRgDoo9Jq6h3HpEWl5TAKOlj6Bm6b6AuwbNVqLb7oMS3KbtfLdJJPPRK1IqpwV
MEs8/+XghcqiPcM0u047RJW2NFxa+RD1kBr6veChjrOJFjfSXo4bWvW6vilgo1Im/XmiTeRdY9vX
nL7zvkJ+Eyafp5SBP1F22L5EsX82x8UHEvTY7izwGbGhisMEkUbeXrvt4KhFIUw6Y8B1W/pIASbi
JyORwrr3fWilNa7QVp2eh2tApZmmIpnwD0kMHezOi+Ep2Wedh6kic7LeWcLpWspj9y4/mhinKrdY
cE6X1yyXcanEQoMSIpRR7/v2Q4ESqv+1yx2jANN5/i7WIT/v119pBdvBAzNXfAM6NnpEx+S14TNY
GAS+an2GAmZ+HJ3IK5Bw1z2V5qt5AscvfXOb4iiG6DpBWFqfR2s90Ds5jCPRgrDijc75lvNL3eSM
DyGcq65LB1NNwARoP9ojUXMe0LNHpXFZpBdWktMvUmu2XUEjTziZ5g/PZw/sW0afB7DdR00rIXUH
D/9+/1jOSLs/eT2ELq0wiaYbpAt1CiU1qm1bfEyo3smfVny1R1a4wP9ol7fsmMgMFtTnc/2ynZfM
X50tw3qxc3HUv9HMoi6xFWk0nLH65OYIr/By+XteYX56H4NRZzHGsZhVzNM4N/zmAiHp1Zreciwh
fOt8L/LSbQbB0UJDelKmnQy9cVzsEEUGYX99toDL2r8BvIzA6Y6e4EXRsOH/MKgrew2GJwBbsrye
aensXglrUaxupxte111f7Mg6ZBUgMn3SaJrOB3cPEgBQsCR6GWWyC2lEK0iQu/WCrWTsA2LpnZmF
fSHcVsB3OlxNb7pwIl1AYDTSqjv8pkWLWFPcaGwqTRF9Yuaf4/XygRnjdY9jfdbd0F+6vtfvDEjN
daRFdAB5ey5vp16/17QE6ksXSO9yTYr9fn10iSUjb7PvJp7HttAJzoXQUUcB6kuaRYHGzDXY2flz
ej76NhA/j65GbUSPUUYzF2a4Tvry6bhF0NO4r8R+unTno39db9EyaYgPL4BcwVSQEInbr4pYTJB+
lt3l2RTE5b1UaT5NsqyKNMGAmrked1OnoVpRJTFu+MxtUfrP5vNwB6ix3CPexWVsvJBBrDNTr1/r
X+fQjrYkNc+6U/dT8b48RPgMhZOeZICBsxxyxAm79dOGFltuV2MysdOwxRYUaWCO6QaVOKS1Rfgk
9xjogCdXMMl0oPNHzrcWqQzZqjLmMOY8wAYFY5/cqVBE3wWGeSjTteM9xj4QkApjYm/Ms8SEw6ub
u06uqeU3LXRcCEYC3yNrhzrhBBU5WDW9GHYMMGBffvVFwkmMdstRsyPoYGAdbbxidAJ69V+tfT/S
pT31Xxy2XR24P1R3oUlDsBfrVFGKj1gvygpVj17kMjMmcSnyAcxUM1HfURpI154b0h5mksK/V1it
+A4+sXRKEVmIkgs2vXIFRZdxJ9QHUuXk+lw7CAd27sLsrrS8mOlpZPUiuKK3GmRXfsnvrV8C5i2s
Gs7gy/EYiziJUUeqcNbzrEckjgcqIR5jm7DB7eNxbwcQO7qsYR890YOx6b1wvDlF1Gtot2S46HvY
r1LUP8BAw66HmfdFFJLDJ3IqV/Ehr4pZ2rm/YoWgBYDdjfvmdE3nbXdXsF36VY4zBITrREjM+5la
1/zSq8l/yJMULEZTcly/omwQtBsfoZ/lPDI/XpbhM2+HZ0lIXoPO2KtX6SpW4mi0wwhAWqW4/+f+
lW53Yk7pIILapgmXYvZAqmLqPkYb6cfGm7+zW4b/WGZB53vcfRkxg5D05ECWKFJmckKzRPGaCldc
zIK20GvTCXbn5rtWiO0P2LqmVGt81tj4vXmc6h01BNqpu8CznTB0aUCEMmdf2d9bszwAV+Ox+M0a
VVma3k8obHfh96Ij2tQ6hAjqd+/F81qdaPVHX0TCxcINGvP1MFDbOw3jO7DcCg4nCeyzz1n4S/GH
yE2jrL1VXDT4lcFQUVN8MjCbo+KfveSel8jGPEFwx769loE0XxppavRpKT7dBYTWJXO1+IFnt6Yv
gAZ3VlKITux1u9KdLFKVVAwe8B0ckQJUjmc17UWIIDlogVf0hEenhXPNDtqIZbNrr+atUwbE0PBc
9hZK3rZl6u+7KAfzZ7Yz1UjOa0VFO/yamCNrXCn7VARjD038T1SvOFf4TEoFbUAO6ijOfMEPXhUU
lPUgMq3h+/hou0eoexAC1y+SAqStLW7HD0DDoNTjPHLbCRpFLlLHAKwzmezS7bZhNn6de7xaxX3l
s87uhQv93coeye9LzrwcYgi8eDCYnScs6T34mAdxuM2D5Fk2T1ia00YYpddJXsfLxmxZjHlJ0Txs
xP+fDsZJsgzYtyoITvRbhUMPdSf7kqdodd/cV9WaG0PgKqY/8XTiY3XzzzM05Nleb2WkRJbNJvM2
xaFenzdTCoqzSDRYKuY206DDgHcLF6rQKeOxh7Dya98WJivHYBfe0PRBMQ4shhzjjMsKVEe3nA5D
yRhcKZMHOeGgwFdm65mmcoRFkzT2Q+cT5UqISk6Nm9GXfjiQLzrvZHBJ1zaUzuN+zL1VuXt40xgn
6/00hrId+vNp7aqWAYZ+3bh5owmj69QhI8HSBgkgIm53GgMo+ZebtSqs7GUQ9bsEVQE0zKNIwmlT
Qjwvhf9JLZlC4955o/v01yHI+JDv1AFHw4aYJWcAfnZZXNWJlKptkMazCdAsrTqaAYKof9/guvPW
DIjTVRa8LRx8ab29+dQLNUxsjbKc62svk31n91I9oUcu2y09V3yvgWQM+WVXfbUR3LMl5YoI0DdM
/d1GG/Ik112GLA83v/YvOJ7Ri6zkWythQUBPtGAkTRILgL69DxsRcixR4tJmZYDou+43Ee8HT78q
PFbA3qo3034XZJ+61o2yPjqfCxg+9xnaZH6flRLMc3E72xcpB69rXneDEpyYSkmqXGwlfoJxq3v/
fEYl9oZHBzH5meIOlNWMiSZ37mXr7+WG276IOeTek10DHTYj0Wo+U4cWbBhpmznHy+YnR+mAzoE9
0HrfpLrWFa0gBUDLv6yxCAiKZVMxg8w+VCO2IKcJAZ6BkIBk9Gxn+5BZzlmkcUSHN38bac2+4L46
k1p3Vb/VPda3p9wydePKsnblFyK7EE80zn4Ng9a52pABdNJ/oxyc4mdL/zjtYg6l3hqq1FOsU2tk
4Fq3gsCKW2AP/g6pGuF9oWJb6L0YV1xsT2wgp3kvCxFeWg16IGfqmkik0fzKyMpkPaDxQCqOLZbj
YsQFOmUCu14w9SLbPjEEQ1UfqGaWw1lCbJwFNwfIFVIh4Bd1oRKfFK+hAgoo5Uw501mT2q5XFpHU
GZOcn0eQPCm+z6Nbpoe92WbSAJ/7GNQY5c8ZX/suqeURc5giwi7fKdqNHR8Cwe2hNSK2ZB8/pDhB
cLVXPuIX/kMDBz3xfwMQtrnoWuoiydrnK6qwzaScmX0iqlcah+nbaIek6lFx7sEfUHFqaZyv7/U5
5lv+eQVgcQUtUnLrHcYBpNUMUTKRCJzL3fbpnnPBisdNP5prmZsXI8ejhPb0sSLZgKJzhPNNzXnt
MRdMy3ihfgcN31S6RNjlbIIOkBycVW/FHrlj5TH3eTDXfcgEJO98IJgBYD11pmX/ACw4yjo4q9IB
iMKKQtzmm+TGLn/7W6MSWAgrk4mkLmANYN9hXaCNqBAalGbWgZUSETtCJQLsMfkpmU3OQVZYMlBH
0WMELloymNyTXOc+8CZLgMnoX0hrUexbuQapiyCI1CBngkIuyABPaRH8wWRtdcv9E3Ur6rqUHq4j
BvQg30kUBdVyFqTX62UwYLWuemrTQo63ZXeg1ptmHk4LdDErqlD+KhM8ABRnaLs5QUdAj7QpY4y8
dvkfBPhnEVwbhwQwBZ0Gc+z3vVV5GDdXUgwedK5Vy/53BkGhmb3TOKukkMUPvdthzh8Sgq4wfnav
ry6S/COEapsJiuhpkmJbEyNlP5Y93WD6WpcMjdnqWdy/ZZ0If5xglT2mtI2q0PzNz7vlJD1yZ30Q
ymHUiSUPAyIVux39f3bYRTBgIPVhCX/lvGDfy7duBPJ/gKsrucTbeONDkEW6EL41LTOs2Qi3CQFz
jUt4L3H4pM5h3dbKBR15gifivyq6DwZM4oYK9/qcSel1vOCnHvTQbX2KT74TbvdhMKWoJTP7XJN7
GanZs3b1XsIJPlLIqY2u0dSAsiNNgQfWoQA5Wc4EbraI/n2FQ+50MA4pE1SSW2PcwGpscM01xVCS
pw0aVQjSpSzq+J8EOuyGVdQMjsaQVRhEi9+lfQfbls66e1vPnjLCnEnsJH1wqMFYjm8RSvJ8Nj49
6J8lS/iWV9sdB86DF+b89EybTvW4C9GAUqvfAzKiRFZ+OhfX6U22x96w1Su5GOSGCP3aA2qynlfN
LLCCVOa01zq6lzRpTwJGTpKX5Z6M4AmXUUofG9JPYAnNavph8FAvJ3xReyRgkhr28z+uv6SA11fB
uXHclbV7X8fqI7+D4l+N79hmfUzKaRRL/KoAhicy0/1LSqJz/gk7UqWvUZLEFgyoN7fuXRdme0wp
zxWYwJoOtH4bapWqci4qRGd8vRfOJDpVBTOyKcKDbP7KI9+B0kiDOxGHjlsVQK3fnRPLxS3wZjcw
Tk0LLvPym5V+Qet/ELuSkzdC0oJg5VI/d0EsKJnqkfZ5RM5Ewg/9ALFeVPJRXh0jV3aIbZDlH1zQ
x+KvgaYhicggneIFUCO22gEOgh/xzxb2LQYhhORvfnAIh4cZuPWCnbFIBNs/3cD15cKHewkQrOaU
AfwYbJNlj5+mYzN6o7K1L7da3mWCL9lTTZx5RoF11RrTsZRuVvL3yiyFn48otwHh+iGP1CDPueZW
eAJQQZ33N5jXYUBB330UUwZ+4xdCa8Re367a8PLzEm/TNWUlOmoeynCqKGhWyT75WqTJo4Z2CPhT
lqI9+KLFN+xvTMpGbqG3ob+nm+W3HiFC8v6muZI4Ta0vARPEhiecUX9mTgtqmNFPOIM5JbxIbzma
G9+q6uEfTjZbyu1CcunJKjZfXI+hiHFU0OQBE51Uak1JOmeXnX2XUNJs7RLVgcJeVrqj1Wzm/AhH
pYJRdnVZi1Cdat5JJ3F26niWkTbFOnyg+wQfEB+dAFs9ITEs3gCMZcBq+cG8JbBQB9gYCULEc4kM
AgvTad2xBwkNi1MVeJPhbYnu64Zdi++X88Go0qr5fr0+bpCRW6HTjFrRhSZZJ07/E0ogD1e6YezC
17I8Y7cRzb+6+jyErgkcsgcFajBUn3mK0ACJPm36wmiS7RMkd5ZCQR6cTtN7oi8U9tbogsrc2Lb8
a/s7dKvl9hu7XdnyZTbyCDHjC/jsWbGqT7h9fCGhibGVV8Yf7BPzQ12iyKtMgmRfepP0vomW6ime
7fJ5/wYSrMzICTBbofky6nBJ+uncN1j0WE4pAwPZ0jCFeytjLJxwJXP2BUuENPUL9/RBp/eggWOW
FnmqP31u0Pu5P6e7HIYj+wkyDXYTuY+kMmBBbsrmyHhaxn7fZq91Vr7xPl4ZK1YCc/xxKAfe+/9u
MBaZ0wmgWUdZdGrmgeoX41V1r7BSknmVYKcCHdvYNXHxyxnbrnmlThuUIBHi0Pe1+wc+O49gDK/x
16UFe+dN7Xfob7uE4KhQv3lKY0o4InmD0U3levH9HDnO0bKp8Gc3criedNEA/qtljGbNcrnBnP//
3v8h38rtP1q70Or8pAj+y0T4kuZigB/6P84HeFCaC4fSV4Xv9kCik1dNp7K9Iq18jXpsM6GYkSAG
5WJPpjitspEphLRbPH9+gM2WG9Y4s9582dVAtlBexCRzpUDX1FbggZj8NaC+GdZbaRFo3r1RY1Az
h1JvycVclTYW51e/xyO73PFcd/PBLgmJWHnGLB3TGRogStNlevrMb9nxBONncOilgBqszNmWV4oJ
Qo3or22xwjzGsRhrBAcHiCEIdi3rD0UE1RdO+/5LXulKcsSpv1uABZRLTTiW5TsaicFrdBh9QB/c
FF/zfugjQBuJug3oGkoX4vrOv91S6rSCk95F0eIhA/Abn0ZVrWWZ7aW6UNLCPvSQUaLF9E+Idpmc
0BXqzoWmrbreNE0amARf8vgHowUjxdmFOxPB/maU8v0Wepnp6Ze9sZAsSlM9zztDMedDUdiSTiYj
MipLOhg6yA8twvBuVGl7jFn6fCOdRQG+3hyR48/B4i5NQnZKtCNtmNFi6fgT35MrsFhYXEqACOuR
SXSL9cjlPBgOym5sHyl+2QwQ6Et7QW7MGGr6IYp8wQzHmm9cJ+wi4BPUiDRelPUhRgTUrS10bema
JgwVG82A4nHL5E3AHYxj/ZpzxeK9ollqZetrpd31iyDpdTDZvi5zbi0N4Tx2WEKfvd46VEyZJa0x
nPX4mBpl3N5MFPEvi0h3Em4+897wKwnkahXYkEOR2AUlzID2URyDwHxXgU4h3TKf2vsP6ugPr+W9
XT6EOc1cupiqBoBshBk4nUyEcLYbmH0z8o4j0jinDYiz06QHNnoKG5gVjcDzh53u8ywx4/Zc12do
SbEkIR1tmDGVBMpf3ZHBNDPgxLJF4kj9fNLVWssLv3pFm4ze+llAIpVvR/R3Y6N1i5IYhn2/PXVa
yitxXZlISyLkJCaqHzKeTGREYdYHZAa3RQ0XOI6MHa2cR2hOVR+PucfKB+UZftOxdzJX1VZPhFjz
5LU7MtZhn/Cxld4RvkwMYXtw19IW+UtYlqrCZ7rppY211bq8/5CKuYUUDlVgARTDucCDEz7oVkDM
y6rqqlPWQKtiw0zkka8RxleNyHZaPyDVZ6K9yPsb/GIKaNY1fkbBrlO5rk9sdaxCRFHYuAmroHl8
uUr7gBH7LzoOYWQ1qx0PDWHmNi1bXeNV88Gb9n6T5g/STocaOTBpaJhsqf5BkRPEU/n1d7pvpk/B
ItMkez6E7GK52m+1SD+xu/h6tBDR58Q2qxKSL6s80OH5tTZltVm2WA94hPT4fT2TF5CEs6qVIzzc
S30O9KaY3mKDBbJLdGYfY6Gqi/D/tkrZfmyWNEzOoWvr5HAY3e4NNM+CsoHFZYrZAPcKfMdraKen
fhdiXh1MddQlHkAhIV4bAkXE9eWfHyJJclcOk9e+3enE1hvrs5jkMi3oJ0colPIchrtPOQUjCWTV
H8xOZNeOibj5DUFgxRrPhTdVQbynNDOvlSiKhyPCSqNpv072oXAwN3HpdYS3o0R9x+1qen1TfMg5
EVwe6F68TsFy0hLWbwnkkkLzEmWgPe0cpLGkW+M1mHV7HVOTeLTfgJVn31vbkkjwh+16YRjoAvJL
R/ydEmiwp2Zcwm0QG+gVUdqlIku64MRKHM//86priEApKbqQF/pfxiLNTytUxgSoiA+EuOllYt0f
+qxU1ls7QvSJQ3AWlTKQLB/Xn7ZEC+rSm05608/ouffiKD3izqdPrqv95q75Lben+vEnTNLqOLtq
yndkVte0bjTtbP7u8YasX58kJGPsC08ZDWHlzIgyRGds4Ui2j9dxEPp/ru2WoagvkZMdrhuiVJAj
VNntv9ZPfcmtyLKk55jqqINO3/OohRCspG8pnTV+4gTCTZVpUvbroV3kC5vSaaRHxfsaURQX2sk1
A0WK1nrohocny31tQ/eZbtEOgkFXQqv/O+W6lgdkfASRP2tctSiVJ7bb6m/n0Tt4VUWaxqL/Zeg5
xC2bgF8o8RjF8Q0ZxhC7wqy6oYDlfz3yRyo+oeYuu/B2nP6mI+NrqvyfgIA6t7ADtSWGSC9jxrvw
qoABWKMjiveTniTBI4+t8gZn+pQ6lI5KZ0E1sRMY9EnAfwZ7RRNNErX/ZEP4WgspGvQbhcHl8Ljf
TmLVEGOfK4zBhPIMOMZzh/ZX8jCf0EYYmwi/gPh/ptrK/uxcZSLUvwAsRRk5UNW91kUKYimfI2ei
Okky1ydcwbzPCiiuB8p69A03VyuZjnA7XmMEtUF4/OUGEAmHKaNYCSwg0mg/BKUWrowMbAgLDffp
kbtD3uljl8hapXXtwTklBm2C+v2Nd+PtkJ+Z1tcI1v7WmzIKchnkNn6S3OOEn8TI4NnMoxqQfqri
oCKbhXUjeQE4w1arXcwAPoNx+PymC9AaUK7adHxfxHKvybuOdeU2nMI6/aEOmjfoS6BxaFwPNFAJ
PUfGnitj9x38KeDBdIWQpI2THO+GjXoYjBr2e3SxDurs4oL0ECEGeTc5oGMfhy83Wd4dgGL7T6Z5
xgFAbMWXUbQDEk8VFeqsFezi1cXLNRWIserWurSUp0c3R7gF//8ElRq5OiaOKrhk50T1MUW0gIjJ
LJNA921fQ8xb94ta6OvM7DGHXqdqv/4+DTi3y3M/bRehPCUqgSUtAgswoSb3hd831r8O+oJ7rxdK
cB7ko7hrSrnDHgD35reeBiWKxJOeNrq/o8dLTFDFvX3XItOiA59RRKeT4PAneYclbFVlIzlnptpX
khl0+sg8GUQoi0TzbIxn3Slt3UDVi/q0LFZngndZD/at+aJSBnLONtzmahA3/xHvUkrtDec0W4TT
5Xv7QgrjwqMOaOpteSu4TH+N9lUTnC8vtjntz9BwVhEXvAgRMiUbVli7t9Kb4HhrhwxiA/85D0i2
dkKgTovdjpvk5R7OiLbURJ48XO+9KDswc992DriuVugr1ddB9SmnPErAszmkn5NV/XqfE1UTqLKb
nGLrvemJ9n1KtWqd69/qf5udZc+aBFjFf5X3J7kKJTFajKJJtWKCz0reha+zN2ojXQRh13bSpASO
uKi9MwdSHd2u76c5P8qVWZLVwfXEjBv+ttxHW77iG4Ano6OUN8rAiqAVfCZT4TZx45cAHOeZ3Rwx
wQj/OEujkOOqEviCAg7ai2b6Yrjk1jDN0gsI358fx5+HrGnXr/g0fAev+q/vICOa8c306W+dzaJ/
Rhhkw6adzUcSAEtlPVOy9VgSsIe5G7GfbMRovBwXXSCP5765K5W+7NukqRvSApfJy0xwZ3CPKkNy
mwFeuY1sCfTwiOz1Hj2DYT4eop3gRt7gfbRyOXBJohSE1IReCzocPrjStr+y7tfxEgIJFQnsZZ2G
oRJnPK7hceRZs1bIFxJX9R4W+btYq91ReFR10vroHC2Tu2wjEgVEL4zHrTpclAAsIxkFKVQOSvuJ
vzCr6Z0OGMU1JDA10qL2qFcGXmVLf/B4IB0wM2KyeeEJUMqUjhXakvfCQyTnds8pdBH7dSA06bl2
LkPreyrNNx3KWf8/Kdz9GocfIV/4mQaxX7RQsGq6y+pilPmbwORbNucOmeAPD2bdO0l45OhC2mIR
amoey7VO5y1N1yImXf2NETEruKTCrzbA2ghnDORQu9QYdHB3yiZ6JKe8K0elrh3NESrr1rG6XDTV
L5RNuUdUzAEDEy8PtJlob+Z8jppLiiAQIcGjDudaigqm+jsnAt4C2fHcUbqwhehnoIvZA7yKIDDF
r8QQDPZe7YZGbNXyYw5MUbcwOc7abqPYcEw8dYSBV5p8hktLtByCbKuTw5/dTQmuPo5YWA1xjlpQ
cMerCFvVMag44138/8K/7rIXA8bHxK1eua+w88o5b9a8pt62Ttfr4lKozERdqntum4b9Qo38SN+t
Vjabwus0M2GABCo5r0KErVZMV5X4IjlpeDWPotlJJpMJIYuq9NMZmU9NeiUZrtddK7+++6CRr5lG
VwvM/MBSLAgSDptUq8UR3OsiX3+c1VjwX4ye8bhXOf9lZxHZ5Pjht/SSVa/V/z7jpkRqOaR6RNH4
2c9z8P7SaPPC8Q7Q/wYkmW6p+WN13sv1wQEhxC4X84hT7MLPFfxi5YFCoJZE19c1HbJuug+NDiKz
0dGRnF4erCUvHTUs40JOyUXG608KNqs02e0VIcZJL/PdsUsIC7KaRXgIMgD3ROGUGLahN99L8Mgy
jyKdqPglDLrxaIJkFMXVD4z0WmGqEFW1viENRELrbG24qF8e2WbnNIFkTzHktS/wf7sMe87F+d6E
1T5QitZVzC0bSpfkWUtSQnD2SguRnECi4YjkEOu5fU1dlc0075KKeSLgEnn5w6LT4gu6WMH132sm
vf4r7+CQmmjNcCCg+Qmi0eVk54nQGBuGFjZoBfWUkBEJOI2QqYifZToMSjvaimO4krmTmX7A3+GA
IVjkE8WLWDyc11OF4gopvId+1sxmBve7p3w8nvmxQpYwHZdzr5M+LKhSkR4BpNoF0nFdc0Q728PZ
fzCSsqwGICKuAut7M6a61SCEtSruvNOE+caGqXCKhcuykfp/UHob+DVTRiwT7K3sjyg+gJ/aE+jm
cUUJnKlRNxLWFEkDgZ9cMTPY6SeORmVDwUq5S+8oDqIXDz3vzImocPZs45zdWmXL64G0uDQ8A6D/
PfDzmROBkS8sNJlAN/qyV8RXI1bXAeZrYd/VTcYi5qk1itlmK+6aDVF2lGlgt3Qw6RB6zrCnTPay
D8qOOvlVUeU4FTcBc7kJCxezpB1aGaN+oSoHxklUDpJa+ZYVyiscAecyCNTDvVtzZm8R3YX8CX5l
jMBGILUTZKQMCXO+09Oz2o7lhLssKbVqz6L2cp2nDGdG7e6iQ0pbZ5lf7exAoVdE13PVto2bXmjq
h559i1RkvFIqJawJMDQuC7DR2796Q5uTkmo7NBUjrmFNzDmSEenAad0f0TeE+w7UwJi0yb4QTUNm
6i0cGtOLbVr5zmzeRMAuwOTi88+dVwbW8MfEqYIGi2FZbzRvHA29DIJ601yJWh0ZqO9C3NwKYBKS
CEIL6Zie3pAv3/SkLSCy8To4uFg9S12MyP6NpbVU//BPVBiBq32ERbzHHzOGmPbYEU0DMuI1Ouo9
v5wGXKguNJxzJVYr5XI6jPrULBXZMjrFcU0MrX1cF98k0ryugSFIpvV03ggd+1olpt1TWBcGulTt
hIusxSYvFX0NYYi7G6nVtbPQMNZE8GJ6hl1Kr/rnYXNphv8WYSEmOKWs8bleOHKtjg8wmKITf6Wg
9X/aaXZoJfKIixbcp396Z3Ek+emn38st7ct+MYyLgnviVILhi+KtnMeouENPkj+pobRCkI1rb6ZF
KhE/6UJz32U6rcT8VfeAMyHcNFZDvoNswwYh+3//RZCifNxHsu8HdbbAMBPY/lRYC0++Ex3tfKq4
pof0CSYxRZd7yBHx6xHmf1Sd5ADO+/64ignaPuMNM8xEog7Bowt0c1BUd8hUFWAEAjKaFFqO9peG
aOfMoJrfnd79pdacrm3BDWKSxkmENWe608TSx05Shxj1pYEQXl5VBY2Ywmu8ZhZwWNtYXoY6ByFn
bggyRetYrrCzUF3sypzzJfRcI5UaTaqAUvhmrkdjQNY62ItN2FZYNIZAh62lJKRWYwW+SbucxED+
srso/Oi2elhInxsNE2cbzVElkKqHTWtjteDqGSUyyBw0Pr5wMGNpJ9v18xwofu2kkFO4jDpzcsVI
HOmyzE72y0jW8m+lCaZzoAVK9NcaB0vZpwV6QCji5tn+kO2K4JKKxyp2SuEXWijFw1RyIFKY8fGf
wduG1ntxoLV2PDqHiAauFRy49XftbOR3GlN48EWJ4gCbIduh26hnDenvdmUlk0syuLu5Y+OPJtRX
1aMZ7NuOdAhJa5r8wqEOh+QlxhhSZ5vCb0/PGGkNGws7OtWQA+UgBIcnkqS0fAdXACxqfwQu79fy
jD9Cd6xs82zUuZIhznoBT2cnGt2yUBZQ0ygknLHPj+W27r8qVeaRr4WmrrBEhofbuGsprmV8p5M9
1iMuewBw8POY1IvHUJDY1xdg+UfD/e0v23u/K+Jz45cTiV9alTR46fMS6Ezy5LYRhrJLdNrkL1rR
stwu//yg9weRv3HOSGXFth+wW/zWCGTRcDKNu1lAb7vrGON/xxxKaHddHy6ti+7E20Fz4E4Umn/7
KRvi0sjusTzFvKg49v/FgNPN4bAlSwcTzPnxZ2XfjhgATk+BqCCoXUaZppDHES/OHAdZwMCvaiZo
p8bihVTU7KufLizt3YRMPt9+qca2fB7kdXNq0+xj+5fjF/2g0ja0AYsRvozGMTkqvWwUn+mpC+9L
irR2xhOTmcUrE9UlOMeuPO3ZNs8CQ8UEsyN04Ov/92Oe8aAFuunqySxiuo6mhvwrC70wrSL18CKW
pDMuWac9lntoRzAQRjpYGPVdm4kSrn+AdL1k63s3InYCoqVCWQOQtmQtaZeV4gwb0DmGBK2mOWja
zv2+Mico5seQMJ5hiCouty/syTdDDDR0CqeP1QGX4Yddh6R6mVllY2lWoPo8lKDBDaZV7WkhIJnH
P9YiTVuEO2zWuVSgMNAreKcQ3t1Y2srj2+KcoPPuaBO8waLOyNygWfgusYgOLiETdfgFL3Yf6JPJ
2cBvQpAqqqs14HPfqjex1fVMuQOzyPP922KBECZsu/cjTTQ6ixEsvS1B8IyxKgJqtRthzACRq6Pf
ov9xxL7ae1ImZ4LI01VL1+f/gXstLUj8H+ESjNGKqXmxnF2nN5Fehk3PDPE0B/NAJqI4KFJtvZcg
eDRsPS6ZlqPk6ercDsS2vph6WJ6kKWsMuv+wx3FZq+XZumr8rXoe3HUR+mef3TeNGLjx29tGbbM4
zt/xED1cWtUB2YGFBVsZPq7QZT73q1MF5LemL+RASOi1ImgeyfmEsrUoAXbCJ1burzCR0s8zuBDf
2NqSYK28I/AkUrwVYbkzsrsAtsTuG6sGWGFV4wETJVxothVk/dIolO/1BNQHkeuwh77l/zxlT2I7
YnLYa2c77C442FKqXbBBxHn8L2eDN3vDD4Ykeqtcmnpw7HqXTTjv5qPfJTUt6xXF9L7w1x4OSWJ1
WrfmV3sj8rzmobiyT4gWtdma/VbfhizN6s+lUF/Eg3dUm2sNdbhbY8xNoZHVb6cmlgTPIEQb7MsE
jeTc/XTPRzXSPyZYbKUl7Fu1TCX22oY3JzbKFj5LAcgSYTvQXGypvqFwkqQ0Ij3a5Lvqsk0L9yOu
2rfchZ9d13+bzM588L4TWmSlvDzT7vwjAxv3YVZjmQKbgCMYWfZ5H6BIvxKVAwbKvmF8Bc8zbfAN
vbEua8d2ZOSbnCGVunWM1+xB44IPOizYruWHbrX1o5N+/0tyYkrq0CNep/NHguG2+DD+tkOqXwIm
GVbhmR0pEXBYAcbDdzChvGPNPP/RVgh9bxqbw4JtaBkN6//yuLU0Fa0njKvx4Duy50Cep6KRGG7N
olKahDJOibKAgbmh5nT/XhoIM2uExMIp/xvWFYDHQ7iOuAPenaWUchQ8Vrqe819KUDnq1evsGcYV
P3OY3MbMYzYYSGHSDCr28jMGliFUCt6mObDugmx08S72sT5EEWhrQYfVQPeegp5DozZ6U4UAcvo7
yLSNxKaTYLOuNIeg6dW4FIQqJAxMUlwsJOgElc4eys79/pr2TkK0bEyTEpzF357569LiBUSoEpQz
lgqNHPxROvnIdQs7VdWyd9y8UBWPQJSSOs6MJqoyfmqpuTlTMDJLEfgBFj3kaDz1fiYeBuQ14wJi
PWJ+vCU1f49jcKGu1AmxeYqtA2AjXsHT1G0Rk1aOE8uQfZW9EMeW+W5SEdmclwlef2SyjOoiXtnc
ySQnabMs++W7oKPzdDVOtm6ckoRSsOYEP6zlGXfsGdiNaBocdxVi4qoGFPfdg2uhCzPQBE7Hgp1P
TWiXUL1nQz6R7CxT1Ytfvuexkfn/Ywnq11fEXxdSQdcsKH3k1K1lqFhymEahCpJ2ckZ5VZM8G5DE
IKWme8V5rAM7+wJsmax9RsCAllifirl+Vu5uOs8pvRlq4VrJ3NYx9R9yBxU98DKvouAhRcr+6cPK
b2xZQAES9c/Ct13eLpjFWxzdvcdUYxI82IkdT1lh/pD2hcEamhocBmuQByqoYtSuXkFQtYdktnqp
r1US7ZmqVSUQIL2E1TxyWnhj9r34VXpyb4W+lU/66GRdS7m9MYgctHBaHtZSoUIv08YiVnI61pjb
x1Zp0jiu6/IOooHUA8zt+MnaV0MMTMv5Z1VWPP0vVlG9cn1SaeSBMH4/zD494sERLnSZTXpT1jH4
d8iIbx4K3kKfCO8c1ilwPaU3GNcQoDxkVGrb3JKBGL38fipvOymV1lfMs+2iBhPnKQJEx/LRK8lK
7nx9T4WwiE5dYBkBhzR4WXR7b3QvpRNKcq6AV29YpqXcojBvEjePSM4mk3PDPVQ4pm04wbaTblY2
RAWdiHD0AanZDe7zl9NEjnzu57QdoWYmn+T9STR5AaSt8zzXl4+R9xjkFzR0tGBqHzTbUn52H3RB
WkDg4CL/enA0atWzggAqBe7X+hdcvXi5nxhGpRKlU3FxR6zbgB2nczgEALPG/p7CvBTS/dpQpIz1
UBi5n5RrEQJE/mlWbWQbycOMLR5SgOkYLoRazapdVh867oQZCJ09m/Su102N93wD6NwYrI4IYKxS
XhUwj/j0gOj1UoX9tsFczr/C3HPIPx3vGeqASGFU4oQS4IlcsplHbKtOV9XASyPrarwPK1X9vFfa
tLPtQJRTbvHYrQlrjo8QA5HsfwIgA6Xqe+zYoy3KVghLUlTr21n57MexUlGbEPEbJKd4pQAfsJFc
LxMiH0wc+VxIQziA4g8YZeQqAbEME2JhhFyy5pUKdRWSY8mw6BT2KVXLuxtyKFFugYnGSN62A9qg
Any7ltU5eZtosglXgz5cLgGCtQ59GHcRr8O4oNvELzjulATSU0DmbaiK6doIG1gdBtcpwY+a16kI
sc7zKgVMqm1heF8KHkud3SmOaiXleTsucKSJbtizZ+OpJcIH5BndRFI6/6xLSA+ChrhJtP1fyJ7v
lBzuahhUex1B0LE0mYqs1QCMizeUrTW3DVpXo0o9VNmwHmVO8SGXwvT4YNsAADSU49T3xN/L0eMl
kNDVN01rfZEJ9nnLCTHY0klorGIijKZvRb3OMofPKBRCArQ5uPHB5cjAkeulb5RIEsRy3p7QHn2E
JMjfeTn4+X2LRDBwJDQuXnn1I5v8eEBFnn82TlsMkLZy3TPz1aGUCl9uB5whM1u6NbKYe2R5TPGN
JyefE+KMeDHjZcwYbzfqXXtV09WKnBM8Dkgys85qpZo7+vYTouzq8V0eAVxxFlNPikO9fg6Y2gSA
U7+GLqzxkj54jq0fGEApqUgKPuk5CNzp+hZ+ulpkR1dBfgZ9h+5QdVhXkkIfiJ9yj5beFvVUlA2P
GElLgYe7ix0XSe11o9UNJEi6r3OKTWcLBu+1uFzLcSEqldeKl3tlYiEUBj/MQjRICPbUKQnuiCiL
qNcsP0lpHhBLVou3D3KI19VdCEjjRXHXnlsRLh93InLz+47FREMly3C/FEFuHPia0suu/tHdXORk
n7RjelHGwMe9hKEd0n5T1f0ZnqSsDnDtibOLz4UkuWqAQ4BRojgBqbC46HHs/7+uokyyxmhlrcy6
8VgFs0Gqy5R1r+X0PncviUua24KjcRxf8ukSpG+qLagRBVHMYsiejtCnlvvzecwQqAQBvJMGcG4r
3OjTylnWjZC4bOPq4f8x7BrsYavVMis5wsIYnhwjv0d13swtGcNaR3TnXcpq8j0F3ljXPvd9Mk2M
+8UQgOh1fdj2l89ZSLOXWlNSebAOwrFwiL14JisOoOfgR94ZeUSc3G2bTEGvdrLynOCFU3HhkulH
jj1Mh4UHR3dIc/KN1Ecc0A9i1Clxze42z/SUdRQAKpjSLnlfuglsigx2UBJZjTJXEhwcvLIAiml1
8XkhJ/B4S+ecGYGSuCviwSHxuQa+YCa52ce8lW1d9uF4BFHL0k+8OgQwVdkVPo3FGT9VD0WxSh7R
6GS8raI4BNPQUh28wgP3mZWStrh0uXwyaxUUOee3tMPfjKyKtpvYGvqdnj/2H5t8SnkmlQ9cfLCE
915BFrzcNjAcNaYbAOUNkiUzoIzpucI4+t0degznQiDmg61vdN36HBY5PJl4Tq0ooQFuYrcvTNdA
Uxxg0h5HcN+7PNf/ALhFjQWUufwtv4Co6UpLitER4CzARfy4cb3Kvrht2ZS0PYN4GSSqSunyv+nU
SnWeQp7YrhIXmj4Pss/+/Y8ABtJcA28oj5cESNGPboKiuvq3OSv+kzIDsltRZC9v/LOCyKPN7TDP
qD6lic0jnkGLHfypT6N2qB8yERAiGMOJU+g7iIeyrIBShLPfvzGHM1UAjM6FzgzFrL8CUFdaMJDU
Nhz5P/NKw1g6QHydIkddILnhpV4db7mLckG8lr2voAI96aCaWnHlwWmTmpACbhH0LSZnxD4TC8Lw
9wL0+wCkyuOvRKwiUcofL4gAyvF3xey+1WHWDEcrYh5VI969BONJ0OdF/jhMMBKg221xf5TdjFuG
dJi56UnbBP9y50R5tfW9aFLQXpLG0PL2I/Ialff8meS6BvMGAxAS0+Vdp5zmDaxwmaVuTqiMi1dT
VaMBY9OXst5WItL5JtisKSsyAnAwEZ0Suf7JL9mnYuhHNNYDoOIrY2JKElocycSbasv5DkOnK9He
z+kwSm+HItQyYTHbnXRERT69yVZchaoClOq1TMU1NCtAc8pOiXHmuBuoPGTLNhqGAOLIaN8nJboO
cA2GMeM2cuiTtvdXB42zXgCdk+2oqTFxmH6y4Hwwi4qcOEjU1Wbs50VmHo8N6TwDKoxphP0APciD
4jrNcuo0zinv85Xnj7/D5cjnikkhooy+mH2Wi4Um5USPOG3zVc3D4roQ1BXhWukbuyQuFSao1tV1
MiXFv5/7GEhcdkz3k3b8NGnlJjagDuyKpzVFEPH0f5LmYL+yu5gcruhV7bEx9xbSJfyQBtUifVRA
WFLXCmNH+07bRr897Di48USRCEX+U7Chnyb8MhPj9Iqrvon1Ub95qDBB9C8CbxS/qt0Wlterq3t4
F2Ts9qU/Si2rw1OPh7wnklwx0k4vHpHuOAzYJ9mmQhXIloV3GTFgOrzfYiHCJ0aI87W6QgNxRXQN
KSv1DblNPri6GM3rMXPsRJJY9HANpG22u91NTWi03/9rPg91wdftH/O5f82W+/uPZTmbNmX/J+Y5
4T8GsAkMEyxD/+teKIfiOBDuRx0ILqk0f36K70iMMgbQsqYZtRfooEnq67U0KPRa1xmO3BdDO9QP
YwjpxVUkrLbZ5gGuxe/+BdtVrhkdWMSQ7RkCft302e7l3cM0K+QAbKgIlRFb5EAdjHwIMgJwucC/
B5YT0hyec3m9J2uNkRISSHLq8zUUGNxoNqm9ccaARi9UwH7DdmGwRO0fO2xhYqUhaC05KOVecGGh
NqjFACUYfN30Fz6YUM31C2aK9n1inXblyWhIuQv4ElYs/J8Bzzhpnv0V4tP0kr56wCwhHj9uSmQf
u2419CV0BcX/DlS0FtiFH/hWw3HjFI22W353IEtYz1QhOlY8rWgoWHp11NS1r4JYjmQnK5uTCyhF
K5h830tGBOGB5D7jb0WbnfaWT0T4towXOoi8rTrkwg/K+f8uFlMEsc+qy/2NguUHTbRWk9HiSkQU
E03PLPRWsC8yVYALG6vyEZmXYbJg91aI5HsM4oncKGq9/LE7XzgmzVYOBF0AyEIOF78DXOtzS+uR
5cWfMhZy7SXVPOk3w5lvo6XN9XU6Q9vpGJYg5L3jNAoXDGcYjoeagOFjJsdiNVKhINBIB//CpQnW
JOJgZrmhS5ecLW8dXocyhzw64S3WoqrwcDanBGSa0FQqxINlYSR0ekNU3uhFUTfsqqLnQy42KOgZ
auOE7qdfgzs5INI6Zp89KgWIXXJhsvkffaWiZzqJY8FKzvN+yB/UwDrBmH4kD22QWAWmHvvTIoeI
vE1jUP+HytSF3rX/HW726w64ckJzbV/552DX4fCoDMr7yxQxRjYiAoBRpXdZLe0guqccnov6gskK
EDD4si4/DQHQTQGhlE4as7ZTkmH8cjkuvFRqYbWaksf1T3HdQ11vVdENJcgCAkrTcA56ThlQvh7O
UpGYM4wmuPC1ftcldTdEyAE51pWZG/7wuxN8i3vxxx+o4TkdQ+HcKb9NXwVqPCtXfOjGi2KjBhTv
ZbAHn7P9h9Ugu1dxL/XUnXd04MNet4lk70ymp79FeG9IfnE8qbJe/NYMKgdZ7pyjbMPMXRRtpdvl
y/5Yt5VSN2qB6xyZVZnc5Oyzbocx/8ebDnVkXGy/SOCWAZcd1SuA4lPTPSRDlhkAClS5dY1wS0iO
bG9nEDwMSTbfaG//TWLeNcPto7cU4qX/ac1HX+Oqo8gbWsN0+njbj/Ir5oqD2eKCx2DJVEYycVV/
1Km4NkcjhSL5f/trCNtrzk9wBscImVi9D8dYfwDx7Y2OTlcIvhB1DJzQtxSJL4Y9Qd7LNRfvl1Db
yEpSZGhEBdbTHkgbv1CPr6vgH2neeVMNlPk8+29Q5Aiv/g1kK1EigAKr0HKOcKyxP8K3s0+YkWAi
gQVrKg6Bf9wAAGVPRoE5ikU7gvKUC3BFWJqwDMlmQoDuMPtu32sAg831VJDvbOucCnpsp2tNC9sr
/Le11hqd3GH1xNxkFc1wBvDHlVMxtzYPbFJeCJcbL+tf5a5t/pwS66T04futhmTeAzObmV5VAqEg
Y7N1dReMdVGknB9dkT4lzno3Dfk/XFnr4jfVTGTZzLP9WzkLf2nWzOfQthnDQ5eYm4XVXJLI51qI
qPEMdcd7lb4i6FwR7l82ucp5YIxrff52mo4wKVozDyc/kf24LpjGm4IqtQ7bqzl5yXcMKfnjbVSk
AwofYyhBz0nI6oDHfMUuhC2tY8BaTVt9vZphpDm6SjiwrRZpQnM0ql0Kmrga7eW2Re6q1IpS3tyl
ywCfGuoBiGvwnPH616jIFjSkf5EgLR5YLAgKHmfzzBGuNWfY+KtTeAJwlPYohVCgR/aH9Y/3PzQA
T4HOnkGE8iV3CDeBddmqPPvFEEJ/t1Ez/43LHn3bvqtvF3r17s5aUvgMjOOBbuf746thBMQVR/HY
0G5oZhx5NyuT+FEwls0/zqke5lX7bo/bkmT6SyMwoCOIgpISaJzl2UEN0ni31jDFq8eOF48FZwaq
mVqIT1u8mmf8wHXKS+S5ALw/BBN7tEbQLoGhUpNEtWEE0nGPbb5ozKNxvTVBmliK8rRqYjwjPVYv
I6nbtcVZUp4T8HLEpHm8m2qXoxxRWI3SlmDKGnj5YNiKF7HBFD0vSagRfvGXCHfZwPJdXfdyY4rz
oB+/7QH3m5+Ozispn94W8QqASmFgstAW6TOcQAa9msLmxAglMOo7BfDqMImIr9w73+M3NZvFygum
60lU1ndqHvWdXrwV/yHttxHbLjj38XgX6rU4qqfLgIjbACAlzXLZ8y0qk+ODy2yR4rv0QlRx62LR
DYWZA18nLT+Ol4NLjfd/t8pNQarMvREreuOtGfAkK7nlh/WYYPbipKXsJxj+yDGrxXoVqvec1AXL
P3B2KthRQ7mnLo6EQTIyKgEzOeCA4OA1fqknuquQAD4UpWQASDh4Oa88uu+K1KqmUGf/OTgLlPLh
3uc5qBnNTgt/o1xuCK63q0xzRPHMpr/uMXFKpWxkx6Xw4x0yTP4/d19xNiApTSwbBmblpwGE6ebL
P2MaA6s5oIrNhqXYkS5se5jI38ctRf/RmZioxKPkHHGC68PPmsVRtdoof5hd2lr+lhNHIQpq58KT
S4NTxgtQ7XMN6ynY5TMfGRF1/JmGTmoFBsTtGuvVTHwoN8iKzC2ugXywq9+I0Z4XHt2ih0lfxt8k
nfWtfSs5DLBntrtMVrx+NaI/BUDIusREZTSIxtdnbBUg/rSG8FgZSCTSe9tR8XSU6IiZ/wFxao8E
PQ1SxTIhAOaVDDko0UbEWxiwpU0FNUdpUg8QVwRsx+tOLCYvRHcGJ/nLu+V1+AndB17dLsZeoknI
i0cz7d/0vdMDLYdIaQJIdG0jQDuJuOkS/VuEw6sFgfr27+Q3yWFxPAkvhc9Z6x89LMmwtzTygGvv
cPAKQNI26O+yuzhSt3z72nswp7F4GWl63KT6bwONBoOrvZ8pQ54LjG64KTnOCFbY4qsQKIAYkskU
gGB4rhDKEh0kLlTxj0yPqiwZCjwssgGRDx+tkv16ei5PD91FlUM9WgTtfuVRJ0nc4ZawMzktMaDJ
n0IeWr3h1j5VzTwpQp/m33FGOZaIg/wgLKvxrZ6iUXVoQKvNTYeCjEKvJS8SLhaW4zFe1Hp0XaUd
GByg23xNrACXUDk189I6SNIoyPeHKCI69ooknQbAL0Le29hy7c3OYcN/gi9q7tTmxBhmEGzcXDX6
h1fbDA4IH/34byGfjd2vyOziqkiL/xgP6x3ugoXG2+jZLhi2gNo4Z0Woyk9oct/eez2p7JUKbdcm
x7RUHcfcjiw03Xpg3CsOww3L+hUmuNnPwXox0+W5nIMS0zKiHJpyrbC6qOowdcLqC/RK0hOPJ09g
XSNi80irjxwFNh09+PFYCsCn8vU2yFU4DhiVIIQYYv7f+LMXsJEamIZevAoD7JT+Ae2FPAqNr6Dn
JP7wc5+JANdnSOsLBACytJLryxZqZAfUI5N2eAWw2jTJoQUfHKZPLSCA3gGJeI6AvVjOP/fYRZKb
ZDypToYv7UL/2vKfkC5Q9oL/R6HwlhhZnpmlRgz1m0wz/q4OwCvt6wULI3+gymkZxIyuUHIHS034
oCBOAovxeORJ+vpXHdfZeKTmnDRUuppRDQciwiM/kPL1LIF6HF46PzODX6ofS3mPQYQLTdxICuYT
LV+6DCRfcF5EtCAwkC4AWe9RzVF/G6/ukNG+PpoNgiNvytlClU7oxkvvFpYkH3ECHIfRycyULyWk
pLL+oP7UGn5JBlBTknS29ReccqXqvp9k8R4c3h9dUbQIc0SEYt+/96KzVfOoFGxta4wnNT3wO0Pr
N9kGidFVdAs65o3ReN6IPZreOqOSg+R3eZF/W8lIyYOMx4/z8bgmpHb0LrgWTL0euOYnch8ubBRJ
Yw3Ly88674Dy71r/anMEck37mq4S7IKJapWFQA8dujIrk0NnjWxrJMg1okaviw0bu7tzyXMuCyPL
b6zsrz0wNvg90EIOJTusvAI6F0Q7N1RH8M7NSA2EIxsVbBoWPurtaWlhFFijeqdae31S9r+1qzWZ
/ICYkASKeo7Xwa3tsv8+6eyn/rm6tkYgJy6gB6mBLiT5F/H3trZZ8NiRqxcaeDYW4HwGlXYBLAxK
Ad+aMOVCSjyzoVq/nwBk6ZV04Li+p0ouTggySW6HBLe6VrZkm/Yt+NivhLvOYGdD4yKeseo++nap
wePvBxcDxTJTxY8wRsGaW7KBKIDZ1Ea8jCd/HLhExgAzzbCHDqA6udrCbBJ8Tn7D+1SX60EaANAV
575AxsvpDKKqE7LQ/gVlISjDCrMSPZvT784YWpy36qtTgpk7ZHaUxI/uney2wi3V1C4JwD69je+U
+DavHXI2Pqip7Z5Wb7lPEJfp1F9ywCVmQfEgmvhAzVmVESHqlRj1kAeHcESyCNpuqNueBTnNBDEx
OJsa6JpkdB1joc5aqGlJxskmjjALz8fUY1V8Jg38v69YkQgUInTpGzK6n03XxCDLA4yNe/q1840W
Q68C8tXl76xuFwnM+3TSxORkny1L6Zs58Wnij1ZAbvL0IWH5W3WqdBvNCoowswlPn6sAdcDP2P2y
13gpmeCD/RkxT0Kt2grnt5STm10uH3BUWfNDpiAG3lOO72x7vy9XTK6x2Xg5lHKqSk0zAg58p6co
QPLkRqN9VEoel8jxJNAlyUuH8TflwQFaLVK0Oxawo3hn9YlpoDAQwG9RYyWmXHL/H5pj+Iwzm0tG
wtDBW6K7qg09kHr4ZrxZxtPD+q+6kioPkOaaqSYO7viYikIigPxEpONQGh6nyQzlFvBlpVzyBi9H
fhUcgXklTHb/JJaLH6V0Qbj6Ke1cpNkCd9oakkVRXLAx4/lvHvSGK+dbzSTE6UD+Zj7KnhGkTwL6
eTyiESP/tmOyWNx6Nee0ImlYkqtHJHfIgE1nPghQ2+p7VbsGj4hlw8suGhfsxLa0Nw1Nu8lJ3I7p
jWuZQ1fkSWzfEtrB6sNP4Wj8SOaejQ7Z7+xim6DtCe+3VIWjj1XdyhluPtQhzBVcApV0i3zLNeUX
UrI2s6Nvl/2PjRXJUzN9eOuyUXcQsd/H3WO83EvLBpr4lLdYCw1XQ6pAs3d4etIyNFtRU6RWidn5
66ZmS9BttyaWM6YaizQc34E8nIetITTZQkAMpB3y5+xU9Qt8JaQIcLF/AOY/8RFLQjsruIjGbfEh
iB550EpEA0XIEj+l2GgAezwhElnEkcKGBKuUUIUUqW/1+vsUNcWGAtNY9LKM6PkhDR3z+HYiMFpt
uJOA6bS00gVq7QUyr3tBe3PoqdHz6VWZS/dRZbxD+cqUX0+pSzplGSqMeTVdr1D1nSK7YT7kYtOw
jN4+4SbgW0sGaKor/frMzesu/SU+Vo6RXBmVuJkFWt9Qm5NQQclK+pYwQNBnAtEtJwqh2LSSKA5/
/0VGQ7w/1rB/9nFT5xlQiyjI2cFxSjet6fVel5vfuZpV9WJjhZMPay9DWnKTVoXHamW9Mvy/N0B8
poIeA3p+swOKVrToORJuo7+4RBje1YucSzgzfBvHAys508c096h0LflPAa7sA8h9QlAfyync4WSW
QDrzeM654jC8IUQP9t83oi7Zg3fdhCx6zAd9gFH5/+W87/CauUktSc1YHU4FAUzCjO5TnLtcC//x
EfsEEDPCIHR3hfAsuHlRSSodIh8i1aifBkBzhf99SrXQt2H/+AiRA4zSjsI+lIGb8YkpFsmXovdy
uix+bvFqeTEqHgIW+dv66xlv3wCR4Kz59/cZrlBRfAxt3mkOnPS9yZR+eU/sPO6ZkI/0X9jl3fnG
R1ZkRh/aD/JLtwX5xfXGkDAPrVMDXdFJqWNK1x358d4oHZSlJs4cG7lr3GxUTTEgWIF6sq/igobm
9a5gyi5te7RacvRgALTIkYsz8OeDbshzliN6i80zzDAQs6+3HVmIXAd2EIcwcNP/1HoshpiHLOdC
NShzcvd8sm9rZTfMaiXFBsj+0v29OFtB55KSdsM3hghR2l5Sd/pglStQFc3PwHDR8SZiX0mGLJt2
B5I+9xx1hqfNQ/0PL3H6aPTzz5K7h7uk2SQnRI77J7obJvIdLSDynZybvEnIE6KyV76gIqPULFhe
5Me7H5puHCdzvrZYDKXh/zQ19x/Nle6W/aM6vljyXSZbTOezLZ4TA7irXhLYTBCxuDidTu1B5pv4
VcmtjCbK4wS+9ofCk76Zu7H5eK/jnVDWWTnDZYdzQgJCHbzM0elDd0F32ssusQcgqRdpoctpoqbl
4HzFv6J9YARo0EdIAmMjNkaEb1qaEJ9hhoOCMtuMq54pAOmlQSXdwGmjokCe939gNQVft1Vdtduf
ILk9GecHUaEXNkOKRcz4e9QM+xru5mnGRYAXKrypOaWuGd0kRma4hgkAoUWEwYulESlhOYleJd0+
M/KfPu0zfODZ+nYpjrrNO+oTHojSPys7NUbFdUUPym79kkjpGEo8vSZ+gtLHGkwLYOEiwzWtirTl
UXgDQmY/z9SejR/q8qKOM6q4cnuUosd1XT8Udmm7m1+pqIN5a2Hn5s5GRliwG8V6fROuMldDLyZa
D92bYv/QxE+NassNTiMP1HR8Zwn6TqdXAHI3BiO6UoJTHXj1v3uORunPrLZgbvXdz52KCYi+qCxY
BCvHJOZQvh3DMRzNw8KGR6QbIgXoW7O0XUdWI1PAAGdQzu0o08lyhMgnCYyX8cvTLYt38UZ1B76D
9yQRNvjCPrq5n07bDPgtC26E38nwHJXH2PGoQtm5jPrg9XvpMEjdKSxECiGDLSJtfe8z97dk5x2Q
WpWG/wdpsuvB33Hl71QsmdW+PAKncfyr5+d4314zuK29WgkJdiLgOTUqq9QkSk45cmw3Z9V1tkx1
MEuP885/R7X3fmxrA2FsUtF8IQ18ChskoGi5CUkcrPRiHGV50e8lCwAKmnS+YXQBTP2xHXprYlQo
tVSTHBHcI3NKisG1+ZywMJ3qQEXeFNhpDDGtao+zXwrh4pmJT2DDclEz/bcD4yrFLKYnv6oaB11R
lV1nzMsQILPy8VNvW+UqoO06c5rSWvLz0EcvDMaCkLUXMFBDwctGRVzcmpU5rbGsAZQgAhALhiz/
qgRjLpMdXU71+vEbYYnHT9JDnFXPHEIe3WHht3nOW/LO0d1ve+Zd/9vsUpS4ODCuhyxEH/QBQdvI
gWdo0eDSGChGP5hfMVINjOjGxWZoDJ6+22UN4nyHLSgkfDq3mY8+4libTl0OK4eIx2FckK+74N9z
549qQg1YjCeSFpoZYfPSrWPPql78Se2g3No7xtgJ6NGQgJtqlwHvWxIsyJWGRazR6Q9Z4zEvpVDK
0itkNwlchl6a0fSruMEVErwW3E24Qfu1Xy/iYm8z012IXE/p7iAP8wJkbDPQWEZQzRsgaALCcQ/0
ALiQ5aHxKISmXxEjQz9njtOFEVBeDO0Jua/QjntrFXjNJG/g9t0wB+79Dat4Dmc5S/BND9BAoIAO
efTbQRlIl4H8pei44AIA/1BZbgkS3jc0HvxIOl3n19rOum9ukyIOHX9qi6MfFMOLAMI+0kvF6nH0
BjQOGvVsVCJ0pNPv8VCs6c2s3AC+1QE3TE0Jkdpqx3dr25+FGyr2715qkAYk/W2exLIF6Z/q2qIB
aLMfVGMP7DSRj8GxySr8t5kB3vwsCOOpZkFbEmzp/wfAo7WvcvmhOWTp3hqNOngoiDLAnkVfxHiX
Vr9HMRoXIPgoIQWa07Dv4SKiofHmenk8ZPr5J9FWpbIytBfatFEnahn1mRluJgOxQ1F7OPE4Tvv6
agzOqpdN26rcLMvLBIUMK2LOonXRDTGPwsgwdkc0qtjVZTzUQOVxzzIBd+w5asiYCQpI6xD6VCUI
xfwMoth0UhOsJyD1cv7PHy6AnRzGuSwjDoonLY6X+2gQdNmwMMuVSd5CEaD3/VtFMMNCWZZLL+3G
jYnV+dLQ7y2EB+Ly9aAdDZaN2vF1EBSc3pmH/zHl73KaU1TZgAkOBuD8nj4xZ3ni0OZayLZsh5bQ
gs/i82jmFvBXRmS0CG3EmFZMnIFIcfuR471t6lGfknvjx6yY7t9NTxp4rP2/pc8TtisNo3nd7rbE
3beXdYD8YKU/d8zKyMhLEcrHvmKD9JQ+24UrxmZSIzvGbQv9kqqYWY8bw15oinsb/UK8dQ54JTyU
1yDqAtQoy+GtQs63C4nCax5IR1zy+nbAP7hjdvn7DWasQG3+vsQwoK108ygAsrBC88Dw+l7W1XrY
8XKZ+RPDn9HSyj+qwHSJS4UHbehkAV1nzFx3lPXyzwZcHFCP5B4nRcnKSJGulO1+Ex7fjvBIfIVk
3IrTPUYhIUe0pTKfP4L1IJ9XmDLUi2EZaLGT8kM/KAPSjPJGEXaVs6t8ceFScxf7xUP3Ko8wWSyD
WjIrac0fK1fq4XhFcomkDoLaKCwOaQLGbeN+OTKWOeysTXvuPsc9j272fVekLrHe+ar/BATBtwka
VyWl3/rupjN1TIfv2mGeirO+beZw8QnU3DpQ/zyXT8vICcfOd7/Q1ej4YvwXHsemMOcWybcQydYc
Mt4nbc1AVyl2R2yV6SfGTNzivwIDaXO8i15DO72MeXTE8f3FFBel4J2Q0WWiioxGQR4x5uCGsoai
B0Sg4Byas/7ep0qWUMFqgezRmiGeGg2eDNddaZCxjt5RYjtBJNIby7NZzStJADMzyuoQtsnLJzWI
xEsQgccC0vkw2oF3irtBBYBe5BcBhIMj4tgEeNFarhu9bvstA0TgHCHbjP68ABcUwzNSU3SHMAlN
LrdZwc8/rBo/O4OVvf4VGUMdkAUIZqcVaxdGD0PwOo7SlmBuCFq2/Z5BXfNO0/TG09PHXgqFz8gw
mBlzFgZVBohyBOv+0pqbrfwRZkEYBYynllzxgtoFokZekb+3IisxQPl6ENFJgtHEwGOxBiFOJJp6
Ho6jrm0DySkAD3f05jLokWS0Hq5UVVW8p92RiJ3P3PR/D7a32HPB+cXYUnOPvyIUDhWQmeXLVZRA
sVlQApXn3XTBz9HeDGALDUnss69XRRkzATpKNxngWj7S4paio7PUQsXglSkg/t0Ghj5fQx+7xmgv
iPfxg6E4Th91yuRqrOYY/hXCRjdU4jh7tS6o66PtfS7/g3gqqOCxJFztvG0ZTYAovtVnDqPwrhVX
DNkHoa/6ZVgjMaO6AlK9M4NOSHckKm7RJjnE2BPtU0aqoBhV4pyu/2uijyKKZmrOnjbo+F5nExGE
50T3bdsuCofdq5iX8AntiHenmf1NiPWlQpzfp1xM4QrCZIQQtoZ/3tNKiVzopRFJXVEH7oGh8NwK
nMrbc0Gc0wgexV1ZhvqyW3L7Gvk00fpuHEsrAdBsrCFFP8aKiRUpgaIMvESokJa1EWiyCjzGn+e3
JNT/Q5EtoNwr+9D1BsUbutblCTgQdXKnuZaxpYvYWlYFtKA6tJWIn+Hbpgh/8tfl45Oqr58Fxs0x
ZJJiYQbXQST3/LGPbUEi1s6Y1TSon7SfKGvR4iP+0UuYGU+La2TuvasFSAq+S3cemiL19MW6NUyf
qjm/u1lz1vvJ2HFFMEdRio0wzqwfA3o0S2RvQSdRcd7ZZaUkPkNp9aNJxxoY7TkdmxsB6M/Cufd6
O1pTKbsn0Ht2SQakF0Xox2uEwEzWdy6/x4fluLF+mq/JvTqa3f8PuaHFPHLiZ1drbSGBZPe03s0A
3gkFV0YYNNUiI3/DL64tbFl0un65Mp9xFdYlw5dVw3kzTukhk77YoQ1Z4NzhMtKtTpdTBAGYMlV5
7ROfE1eJeVOW9C2VF7TgIWXW0saPh9mnMQtk18cPgh5Dn93fPOH52kSW2erzk+jS4gplNKUbc5uB
JXv1XKwog6M/tweQdSGZX/N7HuZsrcKGe/93mps7xLGDXaElZJIET2Gc9dhZg8IIc+ggi6sDgU+h
kViHNuT8mPpkNgMNQWnKJtWBQA5YqnW2ORVtpVCAwsKQ9kDTEZv+tpGv6YadWiQGoPSzvHD/etF2
Eg1+4spLOqP7JJpR6YCA5a1LfpFc0/gY3IVWQUwbSp02JVNS/gKfferKzWGyx813zU8mTDYPdATX
QV8apDbDHNgKheK0cmIYVgAPCSBX5dClAsC7pR2z9wbI8d41S2/2C9zExkFH1m9axhG/+nF2YyHx
IcSbaZl+UEdushZmHdmKg0FBJH3+3ISls1V8uJGfKHVWEdXmWkp+PJsnmjpz7BaU5wS9g/IqyeP5
TcmBiP094Je7fcQIKOEXqcxmO0ZGW4JpMLpd/Y00CvwGyq/VbpLVt9eim2TG0xaJ/DMVxiCEc24M
zGe7M8vnC2CDfHysFBwH2hCImJmG/lD5hOyhnOjc9G9FQYkQD10cVQ0Y5gAicJiYwrjUMiDyhPxW
BIpqePyQQeNaTezDOddluTYBWO+l27egzhtYsqNmPfYB4xyV0GMi7nsLs9WBmVR9rLGou+q+MaZB
eHfx4cvVjrPZcNYOwmBwhHP9FTet0pmP+RRSPN3Kv7nh/JOgL8bJAEFCs/rIr4vlAtlfL2alZGYq
KxU0kzWM97Luj4iq6q4+4SuX2CHpLcABL6Kxs9ZadR5RTzCqC2HcoVYqZFS41vqnu8SF4/FJYYyz
BkDI/XN/b9D280mGnBM3jvf9kBz9l/Xe1T1uA8YYU4fMALSvPEVI1GcluI12CQr/QbwUgAPJzABP
OVycvNYlhU6aHKRJSqqKm+gbDT3yPVvS5qgyFyP3b/yM7JgTqyZcM65Tm66j0vy06lnDMpqWL1Nr
REQfKw+1zykBIs3WV2SxYcUcmCRk01dp/YsF8SnMHBk2uMUmcqUWs8KsyFtw7SWCiwDFEQnX+5XC
WtiJslamehXFY5U9C5ENxYODGc+8u5lTryR5D4bUwKr9rXovS9NW/fEXYY31IaAQj77WkJQ/UkmN
OrTaCgOLPG15Q3M3UbeDhwSNZazhkLVQ2UUzljzjRmviAKqNhINOZqdUPcjG/66sVK05YD2FD2ue
uRx9iph/ml+yP5np/ZyDAqtKMPBY5uVa8yR0xinB+cX4rhz2st/kbxl+xVKmkIhHfSeBv9eRUvnd
yquEsY7X6fHOo85CBJbCejBqwNaE3vgKF7XE8HYQiB2PDIe5TpTqeiPiGZZQoCmHQXb1gMYiIwlk
i2BoC2yHMR96vKr2MjkIRV/izKSwx/Sr8A7AZVkvgD6rN4p7fX5p4ft1CRFTsRh2G+i53W3PZNwT
xYAobJMZ31IFYTIcB8qVzFyZP6yGpuJikugquxAoCyfZeOIocspEEHUTvVGQdJKBBjA7kVP9gNgC
73Wmmm+KAyKXm5wx5YDT2U6/Tr3biX67Dv9dPz0p4SR926Btby7/c8P4PBNMg5JxhAOEUrmy+XyX
NsTYZoQaz+XhqNeTrSi72+gWDRuRb8VmGp4pmoP56PIXqCO26jo98oQhtZOS5N47MUgxVuvJT+Sz
ch9avpmos1Uvrto2l6Ob1Uht2fKJ3z+PIyeWDVPU7uUHYLlvYUSm+GgZLxyWdPQ2NoPDHd/ilB/w
spOdaQ6foOvnDtz6XwHeuqICzXqZ/5rr2A//yvx9SSmuUnKX3Oz+cnMmbiYVcR1YcAlCis1GQ2Vv
iZzSskgZE56uR1Z3o3fn/Y7oPUjHotxmvlXdTP9elhuUVCFuXu5lM6p7xmfxzpZD0ftHJIP5GTmf
5mDckpR+ASk3WCgbVN0NcZ8WbHiYxlXRTvcM7B+a5ZjNvdD24e3bPi9Ml1Q+70zP/pYucmeDfrOJ
Rb6aIY8qkZ86J9nlS6u5okwKWh2TbsYdNustP7Tm8UEOP8gHKB49MB9nYgkImOl1RP/ZMQv9f4Zc
Pnd6ZDa5A6vMVfkfUo7gvQxNnMPeblA1PtxndOIfjZ7RhphttGmOrHegT+xsY2Dxuq8yF2hn2wyK
NSTZzBv4mH/v7TgP3CvgPGIhq3lTLFYU0Zrs3PrY3yZVshr11CtjzP30cYwnIjI1JvK7SF2Q2w==
`protect end_protected
