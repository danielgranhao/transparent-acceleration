-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
8gVNGI/+S8kGlXP0kgXz2iidyPSXw4XerVfHenfacL89EQ8UJ3sJ4GWM68ff/BFh
6b0ZCetposYuMzR63W/t8J3MgTEXSULF7bYD3LBKzuPuhKuoW89CKM0iQzoyPF0D
taaoYUklUL0PTTZ+YT/5qqPNjH5zbAzbRpMrn8OSrV4+Vx0TXl5+cw==
--pragma protect end_key_block
--pragma protect digest_block
zrmPypDzOA8pjhESd+der7r9S+k=
--pragma protect end_digest_block
--pragma protect data_block
ZAMcmRTw1gc82qVNfrfqMxuVK0OtJbCYedypkSDkm1wOE8/jLxhiEc3md3eZ58TH
65izkEUjPjYIYY5fELW4z3OlAtU50Dp33gfiSmje8VzLRXs0J9oWfOBP1byz5YuB
BTu+OD1FGLBnqSiByqNho8+Rq/4O3v0LsCYi1o8hv8VrCBsWHg1hAWP86Gl9jfTc
mjZqT3sW6fhbebx0M0rsKOnhRlEgRCiXYEKbY6XbC/U5Gd+rofRDq1YHgKERtA4o
/30fVdUoKvMO4ivwaKPWagGA95Uu1VDkwgXpDo+u1qwArCvQWBODr/V60n/bl7ds
8jYnGSG605ZWTnuQuW9MVy/BGxbRA/C87Utc8Uy+54y9ef8qhyO2ki7O9FV3pJkW
FuMbAekodxtM3eg743lFafcfiogCbPIKYMaotSc85zqakg4K6Du30gFlhs0tA2Yh
S0IZ6ButETq7rQ/c8uVfzmi6pVjAMlNJLXY5PDouGUwlTMnd84ltpL4QdoVBaFTb
YMWC5h28YucFcsh2ueEULwaAfaD4+FEYC/+FdyDorKw6TiKzlHQJr+vAm3BcZCDS
GfAq8d9LgH8ied5rlgTP//Q5PwbyPDuz1ogieWpPZHJyNsDvi4wsReUya+qUQCwp
zLgjCw0AlWDKmNhn9QoQTKlMJ9NA/DozdyGpBu4l5WQQQSreJHs31tX4zLma777T
CCHcYe78MV/NeQ4Nd5ISI71B4tonWLIFGd1VjUNsCxha7SERNSLfld7YzdjrKiHs
QzKMFCOAci+snUc2nwSmYKU9ApqqKbouz20hURXNm8CqEl5A7Ytwk+HgvCaY1X5v
XDfFZskUQLeFh0/C64h6YfALLdyfUDaUbULQJsPomlPNOWEbAyWcfYj82ZcWUs94
mxuA5JJE71fCf1RZcJk2X/Ysar47u1psj/4/QGUBKcNspl4O3uowlLlAlOY4oXZD
rzsAfJSkGhWPqf0bR5a92fpj+Vyb/B3ZfrUIBu1nBW6F0qWAy9TkcC2kSLa+goYB
4wp+BIKQs/ZXOew1gnTWldO0mJuparjQZlDBU8ynfxIj5xI6H9566EN2gvREwRkg
Iu8t7wgWMaZ7qAEeM8k2jd9J2JApBc39Td8wQhlGJccR5hsAvhpscQjKupk2KATX
diyBCGYAReEDrTNmYRIJAg2TTr5hmW/lPUutKoyzQmPwoMRJVridN+q659c6bRqx
2MoB4Gy794kfS77gkc20osX03O6CW59heYdUosTnSoYmpBpkZdtQx30Ci+CmDQbM
oV3w8yb+YcV/uW/TRh8FsCED1NmagTF/dTGtPhv1R/jGnIV5chSy1AUkqet5cOiy
sz+oayN9ucTERH5EqrPqeqYOkpinaId7t6JLa4FRc90YwMx/9yFfd/w3QD7uKDZI
Of5pJ00Bcv7Ryu/wnq8u8KRUe83pYiT6Zk6PEbvsv4xiKFz46TzWuNveFYH7Ywms
dEdvvJiKWj5CsmLxdPleaUEgBJ8peT5dGj6p1c9g+HXutSHsvILNFEkHKicADEfK
Ns8wXFRXHt3ZqlEscXDmnJy6DQnoTfMU0bGSIZPS3HEAGVn5ZtWS4J0zeIrI23XM
zcfa4uGcJ2rJ7tCDM1K8fe1iW5zXGPYIN+TApwpdGGH5AKD9CXLNAcHTkBGSV6AY
Td6+PJAbe70niwbNUIO/Hal7l8uPZwv6N/xA9CSF4UcdeMKQdovKXZCkKsBCt5Z/
EZtPfrMLF7PV9je+OJjt9EndgTl94gY7lCJnEbecU4L3W2/rj0Vb/7t9vP4MjSwY
gtADZuXJjF0H10XxNBjX7R/OYxDy3Rm4uIYbGXiCBFuQHyoL/iD2H8NY4EyN2bIs
UwPikE3tHRaD1U0P2Jtf/hH/DTak8xyF0w/566SY/XjrpkzOgVY1r20vh448XJGP
VSyRZkph2/GEUE4om+CKZIu1icASLJEBN3SlrjD5ENB/+KuGcOHtSRLmTc1XifPH
Lzy3h5BbEsoyvlKgiZbp4iuNQtLr7Tv2NYNKHlG1SmYhpWYjF73pj0LIm3ukjOl+
DMD2BG1orv687EWeF8UJ4p3ce+54iymiKH1RG+SxIdJfXB/z+5QjcK4tq3maVkC0
2EKnWaZbVYT1ErmUaxNp+fLEdO4DTrBsQWi16E8C8o9YplQ7b3FA58/iQsVIZskX
4JgC4HAi+u3o98QHV1LMXyWapT2wWCWjyWtjCcpxfQeP0sqncmoY3RLew4/tcmRb
7rb6cmTbaMP/3wxuJc62iFjVNnD/IcooonoIxZ/xC2I960WL8wt4yjckEDaheC2H
D+HmbO3gmC0Kww5geO4a2gexRB9I4AQmHkG3ti6uMzRXIGL4rZLp16z9NCGADLmy
4PFqP7Gm9BMA/b1nj7ZF6XgIWV7AME7mlLX62R8x392LxFYJAuC4/Er1IlJsLjbV
auMGlqR4kYni1OQPLJjhzyKAsGi5mb9eltRHak+q6dUFp3xLoQyZbCFwoFWqra7Y
ahEFzhBtvbDl4/tdzkpR37UPSWRgDx0FggBQ279PXa+DvH5HayTUQwolerqX6Oaf
BFpmVFuTnnRljICkci+dyk6zv/Pd0ZnbnsUuJ1JFaVK9ol0bm/XA2eK61vzrUmWQ
01c7f3GmCdWTPZNdSgXQUkVDAZPFNt0HOX6x1X0SjAdhHMlkzM2FiSYyGmcwDPmZ
UFazgtujprdqUb2ozqy21GCAkzZtvLBfOfajR78X8+hvjT18WETcfm3mupjo5DN8
VI1Kv+NSDEei1Qo5VeolmmSxudndqDolJ0UsQ3NtE5as73wQtiPoabe68W3PEMLJ
GdxLlQnlbZ/vwq46lS+6RDMyWbZVWfcLqmau5WXJGp+Dta5iS/3AtAF6u+t5qfTd
QAZUjvHLOFoQXUmPf0/2fDE81hbaWBIFQ3FDPuAe9NOkpoM5ZCVZIG5SFcdHYLvz
rmy8Q9WZpnbo0Tu1x3ZSwhDSU7YRrEHBdhQeXN+pnkXp2hVvqJGIHulG87aUReC+
G6/jQmyO/JGrqZdayEwfOQP0P8nBVvISd/RiJu3YguzO5Vm9uqXDX5qZ8qPuq9Ct
PpBUdnjFthNN9qt0AhrTUXrg1j52oCrarUq8JdzJWxuek2Cgy2GrzEcZu163WfG4
pceW8qXg6oKc3YwiJvICCe16TmAJJXDPHgFL0+9DFrJde4K1G6ZxYpuDQqqbW0Jg
rk0WA7XWlqDkEMyosYu5L+Lv1UQQ/E2GtSiI4I6pcV2bbmv+RiJuYrGYRMVmaW2T
tkm3NsiWq2Vb7xEJDUDsXzxVAVFgxCOEzGAVyR+WxYnc1Kb40N9z6Uh2WJGyc1dH
/3ZDnx/ASFhlY22UOteHlGtxYDL4CyZFXHzfIlWbck7s5LXVfpXpgLmCe50RIqEG
4KKxdk0GPxFNEHwOz40FPlZG1q9bbIEJ8o8TybMOZ2XGJZ1z/jUShF2BPBqnFIIK
6cBT7l+XiWKqJr/wgwdb4YOiQXS4W530B5CaDS/Z/+TLU7BMt0mAZ7Kz11glLosT
azCYS4bI4pHyBCq+s8RCI70R3p7+CmyQJ18RDeuuiBpp0noaxZ+zX4ix2Ew/Qjtd
C8lze++Vd7973djXOGbkVcDMGJUyGzqUDduf+fntSbErk5zbzSXksdcD696C8tUi
/ZL/cQO99RcWbrzoPJEio1U+KBI2nQRi7XqECkdWQwH7/nVGR5BT9zf/kFZ/N2Ob
Eg3GzFFcbNN5874b5bQJgywwUvMCZnI4Ni9TiUq79l7RxP9tI3J5+ViSipx5UNbH
GwtY9V/Wy9CI4zvQzKcZ0BIM8XiLekb8yC+EI/EOimA/9YO/lO6SE37vTcy+NacZ
pjpVCWwUoNh1HJl0WUXDyddI70h1GytRUzwnTvlLggYYRgCdUk42F4nVLTJXm+zh
u+IXqFTbg2J3Wg2aB1a60J3y6TbEc1FQt/XpwF7NEPkUJTGSOQoZIhResp1NqZjF
pPBqkNqry+xhKrPJrBX4bvMGc+2Vm2ROZeKRVcGIeXtGU0HvMULwJsHRIgWnAuNs
JJMwQ/u5/lxwluG4l+uBSX6LgXQKFhW5s5SGvfeCUMA6wZrQF8p+NIp29HpAwgN5
rRSencs0xpdKlDxqD2J2k6X0O6B7t1OppPr99xvy/IYDk9I//TkOSmYN6i59YJNx
4E2LsJ6qJ6jwSIFJXLFu3F1fN9fc8zenZKYaGFA6O5UREyO7rJMgg7dCHdqJpVPk
hvuaJGbH600ALwHZrpUZOdKMF4rJkmPHT15CMMTfrhyg9PU/JWmO7bGPSElvK19o
971zp1r0WLbltanUHcRbXCxIhy2s37tgRdxGo6W3aJh2MFjUvWD1iyQyWQLFgOOI
C+0e1lEnna4W+d/Dehx7PCiRPL+sRAvI+ZcHTGbSIusVb+eaGthRBbUQAXeeOY3d
R7IbXgjG4JFn0sWHWaSFKZn7W5MY5hplG9nNhXmJnGRsQYF6odEpAfRHXfqJM5F9
cJdWN3lQ/WNW5HMZdVk+1CtI55zL3qy8OhPrXhltesz+v1yr/Zpkz4XAqXzJb6o+
YWtUsSfCa38FzjxBcEt55cwuy/DuVoZKclTFE2RekQxZRlUaQSFCw+Wd1X70LKY6
bxyT2ljYRZhbaCgulOiFipj4SiEDfuTk0UWemh5JX03FqcbY1YRv8Wtts7kWYTGg
WIyBgGDvChU1FxGt0SIW04VA5lAvdb+lzNqRZdfl9hvzXICPByfQlvS2EINQ8ZVG
pgBdqz3n/UGBhvVsXu/wzChWYlAfvxVf8cqd6+rWF8Bc26istb0TNQf8HEHTk4Ip
cXKxgw5pCRO/WYMTVr5PNs9kLEPA2yiAjoLfVX8cXBdxvmZtEqJvfoe/4ds6Mz/P
2ozN2jzRl62ThUshZuSSW9trMD/D8iOJk6nWEkbOZNh+k7IFiFnerqn/6ilaTihZ
30eCo57lw2yLutD1IiP6O1FSKjymLBYhktlA7D0fPkyF6hHOqYnuTQzm+a9ZyDNe
kp4yWOydyxtAAvSNUzbjxaJX86naQVSszczSvBRhdFh8UOCBMYVQwJtuo23D52xs
Huvlb2L+2nb9odbVmbK5LcZvVunuUKcx4MzGjN2+Mw+53Lu/xuP9Y+JPHoFugkqi
uf8PEIOcCqfq6l5Bo+uEr3mfF47kYjh9qAh0vVWvJB63osZv0kjuISRakPY7egVb
vKx65ZaJr9+xFkAcF9LMTloBFwhZUuzoDM6VKimKznEdQDVoyowyQINcxLHRFbpF
TQVgmrAW2qMymANhXAuEVCKtcG4bKc4rgrnmKpm58YfcL6ikzkURfLPZe4zxba4u
Z3534nupi4UQ3h46FDznZDGolyOtySpyNzHQgq91LZ3qf1ZKAnq1xf+uW76HjmB4
ewo7/7UmpwQmFhN7cFzJV02/Ag7fhNO+sNj/eAlTwdsLUMyT6vz0vWqbLlEPi9t7
ht4AGsP/jUUjURs3kE/19+6Y+zqeDvbhr0razf8EIIkRv/ml2B5jSkkerepY9REb
/Vm1ob3j7iwsjBb82tFcV2e2kivtr1WJaoV4S+lynJ8WhgDzLyiY/HTU54lcKMBI
ZHv6AzpkcB3vCLSqAIJpVtVBR/wcd+BlMLICfTUiBl+OuATeK6xRWwB62uj8yB7c
D0hAPOeSjCP7TaTQYCKIrKsZC/LAOaWOPhqHbVozJ/JPLzSdZ5skz2Dyaxw3SGas
s/cDPBOsRMtttwOB3kf0R35CD1GsC71He5z1ydX/mlRH7shVKVVvOiD52U1XWfb5
q2eOy245ilE6V4DEDXPTdYlK8X9ei9tq9FTDPcXDCJRvwA6wkpbhHyIQNvfHOEJh
OOD5GmwoGWD6W+ECuLZqDdrk2nLVAM4N266SqmpkGrVfsgxUBBRlmgiNl2pUeIzh
bLGZWw/t1id0br+f4I8asKk5WacV9cMJQz+cCB4YuDagXdcXd1Q1vWNYcScRexxi
2c1pt9lD75ralFj+/JCPTYjiwTZDB+GTsbB8XamdOH05IIA4GSL2WfohryGIMfSu
cpZRHIxoJ1bhJx+tp47MI+1Gx5xAUmy9AGOm3X5KupV0HsZ/YrVCBjtzoguhqE98
VSFONzNoZR8AHLCUu/Pjjd9wlyWs+cJtfc0jnApvifXJyd+iWhoRjXP8A50ZSs0u
XNIE/Q4ql+vlx5o+u3PLYuTAERDtpniy93N5DnL6rGnfEYwE7rzBwaLjE1uhC1Az
aq3kgeDRH92T+KdK8xElCJzF86KATBpv8Qw1CsPGL50KHw5dDEHQOcTs1alVyT5v
rLU6IToGp1LpLFcq+HkPR+ioDUSSkhW1fC6rTT7CiJnZcMroFVFDX9aF8DpMSPRU
6+zCObGNGpHysczW7hoAxKpPKHMVg5a/0kK9FHjhJijqvTG7tQHsBzv4L2PrCFE4
zwz+yOBnpnwCDoks+AVwJn2iycXw1tmvmaUc6ZuG3m3jtOVkuaOQQLphg1wdxSUG
XmoUZDaxLuF7fdC2YHei5uJI7sp+asvCxdtDK1D9NVLa+bznq6JidRf5UsSBYbEQ
wdP6/HfXHtTIFu8lqxlC5jERgm9LdTB4v3LwGn8uCIgWalsqtDus5kaM8PW3rkYc
aGpC1xNZztJE0JLbWFgKlg8+hGXovUmdEHLIbE5QlePDFmfakz2MlD+ZLTR+7QBt
aFluXsEnre554IZ7liYtXfdNeYLNS0IYkSGm4g+7bHAsigw3ezHUXLmD1UF5G0iA
7MhO143E4q7ySgIZcaQ5xsjmHE0td3kYfFsZD63/pqdnssIEFxKIrffLiVmuhQrg
jAnEJUMjWhge7DGayOGyVLj+TggYt3Iv5jFjbY7GaX/zFP7jgcKm+A4mAMqLqPrl
zyCRI/+e0T/JB+sS28GYss5AJgjtfOUtgZGTKKmpo18oAsOqLhiBOUkbtINu0BgU
aOizM5+O9KEPW0G3gAP/YJlOZ/8/GqnH0qlkyCYmoM7z6J1jGH9tLm9wTd6ada3X
iwKejPOWBbAr8CjGzPhx/UnzyS/gsm8nrhbb31saS5OCeEMc3dxR4a4lxsyvKOn3
EfKdSyo918XUh8ASVXZwETiEVw/xiozgniHRM0M6sZ4K8AEEnbo26rKdid2izGhm
A588pXZe4wWDj12dhRrPgx8k8b7QVUFXU4koNTsukqIw1m3FOAaCSTh3bmB+AtmF
sUB/WpWjCl7clsraRWTcv91OckMOB0U7ZRIv4p1cYD7OKSD0kFG43Q0hUGUE21cA
ngikgmpaz3MnuOtg5CWbBnHg5GrCxFej8QYuZ3br08Kg2Jn534E0THHUNF0X8NdN
FdsDZpGq5TmNCQWwCuV1ughtkdS5EhNZAWfTTX7DrBrW+8MzPGyDNt/pn/avaBLB
qJh1GD33F8gckdp8x12jY94epIlnv33xKDI77H+lZ/3v+YTs5bGXq/NU3J98p28s
3o+sgmMMdfg0mFZmbEicfmcwKZsgCK6eyz1heiuDgUczRuz5nHaK1+zmDiQSfJzL
xpxdqfDiLPvWlhEwyPhB9zMpeM+zsj6nIced+OUV2Piyw9tY6YcHG9BISWcPzdyb
MFZP3miPJP/EEzT5Xv2THUx1blgiIU4NKrm0/sCN5Epz23AhIKmy9bJktwo7WoTd
l3ZgE8nSgasD9Drbys0a7ebzlKZQmPDBHQJ1Wpzm82OnXDJvff2BI+FyKX2NJBXJ
I+TYP2BxARw0C+l+yXuu0onv1JvYZSrJaC14ZEXblv7+Nzi8RBuI+aAwh0PSSZhb
1YQ6HJouqUYCju9cPzfFqiWYSx2cBhBxywiMp+amO/kYiV8JRQGnEu8j9Gcf694R
zBbxt9QfIKhH3zzwQy1phTY7ev9AAIS9VXaJbbR5zELePnXsLkZCXF0m+AJlPmKz
se6rW75RnG689A/X89ROmim8fEcFLxxyLNgIAwJ0OVgTOwZ4iaqG6llzeWT2CMeW
inLpL6aY9LaN/DFT6i519hyzRE00qfSD0N8QEyNzmg2DxT8x/o5pZQudsbGgfXQT
zssMgBqprMazDh6kKt5w5fO+zNz6XEHKG2LwCZSjnL4T+NFBD3O553JNYnyajzlp
kBPBU7slxoFnCTcszueh9FTTOyw5B9Xp2uyryfIjC/TIRGLAnal0dTzuBTkhyXD1
733538HI5yqXZXOtlACgJBBN2SK2YPVOku5SX7OGmv82W4yBTmQfT3SVr+1AmWsw
x4CAHgrCqH4jJPg8nTvMCU+SwJEpc68aUZFaKq8SMDCnebUCo5JeRpjzPwFTgyus
g9xJzWpx6m2OWLZ/n5xMP14vFBhYAqFd3OUqTWcIqTtEZ+m/W+yK8PI61FFDWp9e
eOU8P5rgx3xof04QkWbdvbVSsxioH41QJPxoCb9NIMmZ8hMX1nTTXtrP5hKxd9HH
Gw6AAiiryMOw/wkwqD8hXbyU7Kfico2gX/5aJZ51qJmdfFZCUjTefLhY5mSupqzz
VBF3+HXMk+moSyYG3rVgpTYl2GZH6kuyQl0r/fiFS0z/bNNmrI2C/WZEFELW6j5u
hZT7CioIA90enH8yNfjhz2d7pNyh8eV6XRd5i8P6tIlfzX8Xk9TpMaKIDPfYbZrK
NGF4+BBC147BbS+er4KPmbng23i+l7yfj3gtfyx1iRtsFItrzorbl8fzCjD1a0zg
OkISCIvBwWC3sCmukjoqsNsKBB48iVIunjhDiHwO4z6vVBQSZbb6oCOVdE3Hhwgn
iLt762VTn9i0Z/2kndxPQQ7Xe15jVYTULHgcPpOPpcJmYxVQp2Ipy8jkHWHLZ3N2
R3iaZP6khY3fEuID6wt/+8MOEoY4u3YQxSi7XEWNUFnnJ8Krbzzvc6GUz7cUuEzi
OeCvqCnbdjXQ6xfgm8tEeZ9f786rDLygNNSTJ4NeS6NUIsHiwtY5ZT2JFJi51SFC
VWvdhPTfkVG2zBzzjf5AdG1M+czeQZ7HbYBVxDAGgt10CdyihMYu1OPquehht9AB
cgtoFiJavVzQCRO9RQNjal3drsJBTbjY4RpsnOkskkcwgMnCGftqp58HHfdd4Q1U
nZ2gbDl5pCb5xCplAGpzIrIhK3eNhjGcdo7BSjLjrEw224JsYGLjECCOB/I07LL5
WIyglULUpyveHwZTHBbrtuBAhduhdsDe6JYZ3SUlxPxbp/TRjJrNxrwTTVh/Lrnd
iCM6HiF6/peK3QbEw1sSODXdrooDtJ5IFtN4Edj/kugiMvzMZTbXIQ1iGdHvr1Gk
5ELYwAWnaKN3D0b5e0QmM+eYmYezp9PCv8dbqHd7nsEvVzqWtvoB5xooeJPoldkA
OmU9wmAn3p2QJsnM49s0c5logmOiI0JikZFRm45PST3D9AvifUq/n4Jz6ahA9lWs
R6QM5wEN0MIlTJRxnsBChuWwkWSw93caIlpAKD4aKhNY1qBa/ESevX4TDM7U7uIo
c7iLT5GuVMEn0LClYWF3vLYE8PEfGDL+1sYgT7/UJ8URK+ijGi17px3dMGzwXTiW
JzCb9WnZL4BweZWesGAeEol80ikQz+X934DXYl1Ty4sLw6YFp3r4TfY2HRoRTrHs
6CsjThTLKmnWGg/KRs1fBzf0n7cJEn3GEhSIZsgwwLrnv9ZOkwKZtN4WC+KvrPVY
gk3h1+AWl7r7lUf0s6bx62VpZxrn2yugQf5xV4iThlaNDnJF0lzIyETfLas3DRJ/
vI7mDABub9rVZ9t3Rvd1oM2Y7NagBM7+ENp833N3Tq/6R+2EdSBpHMWYq+Jhbg5U
lePAPUW2LgdcwBrwsi08qV/7ettcz4LKR/02MSxh/8Js1Atyw0W8GrCtIi3siLpk
ZmTFx/2sndsu+ZuHR2LVZaaxnFzxi+2yY5RgDRqhlkO051+LAvDgJrdbg736DZF8
cpkXgfrm8biJ7UNtdmtH78qYz27I9zTdTcNB5JpESqsR+n7jDM8kZ1u7+iAi9tTZ
QYKUrJmrla6VHmDUnF/lU4ShC/3f2n3vrxw0d8Wj8FoV952ayS/xiZrBNfQuZhLg
hCSVErVMcZ5+cFULubHVG3XdLEHxuCrB2iEZ947TAaXxFaD9v7goAoPQ5ZOjUx47
CIBJaA7ZVGPdJ5LjAInY/8pJtzy498lwyCehCbklKjOoEiDOsQTYVuvwwhBWtCNb
zbObuyVWohGsJT4pIc12fDhDLCl7Gh910Jd+kjgUOe4c8vxVzJd5tSkKrrXdup+i
HugCc9enppj2zAN3zfcSaLsHdSC0TehSEbLs90wYarCH60DQUArReMKErcmNDuc2
Zbb24NcOlIDPxO+xHJuwhM/+gH0pqAecypy0L9RyYMw4ZQpmm7giATa1ieiddgc9
W0iyn+Q5VcDg53J2fr4AE8yQNGPTFky4W6QgiG+/k65XDJc/hfMvy2W/lLvYJY9f
QXblyRhxS3ih1wC+UOyegw+C7T01zZkuu2qi0P3z1ggNa3+uRZUedV/1ZJhaOrWq
v2jaA45p+dCDm0cEO8PQ+togVSxJzW9w+KIE39FppoNmEFMsrNEC5IbW24K8w82g
6DsLtTLLPfDm1GuaNVoWkafJr1Kb5qvnKHZIgW0/Qp/UDkuCPKfErqIzOFbESTc7
bl0cD8pCXCEy9iK2JNoN0GF3mFS7S5L4rbgWmOyQ2nIifVakHyGtYehLRjgSFM5a
NBnjp8K/A0evuLMk8OhlnxHDAugZvThFtnz01Tk7eCamMRUR8zzJA2KLoMzxHRsQ
gE+Ikv6TAfyK9tbNikyA7XE8d6hMEw+MXV9lOyTegGJ6/XzpH/KytI7N6R359dc+
UUESu7zF6mHYLp9NCNsyKTvF0Jv9ON4kZDaGzJEpiG02IGMYkCPK1elZ/FjNUXag
l6Wmp8cm46E0c5CtgcgXkMaV0P9xapON2vL/t1ksCd//iIH8gbEwVjrMXGbcMhjG
ojCtSkV+kloTVFUoK7cqq0dN071mc9D7rrWzMwGnGdWab3Jiu5oWoYv44f8McpRO
w1/2r5VAXTMgw2ycQEqXNQVCRg463GCmafpP1kTBUcHo0mLiUwEu/xCCwBxiA+u1
2Qf74DzrJvKMLOn4w+SSGHj4vR5jtYic8HGXEzUyOHS1n8KHMXo4UiQnIfXMzNdE
dsBKP+FPPRVCuJxjcN7fh4cct4mZhJuW1MAZ9ZoMnDAdPZgurahU3iSpJMaY514L
np6zkDrSWu2UMv71gM0pbOUQqC70t8zLEmtfYKo+lIirQlHwp6TkZmco8FuFUdTX
FwbM5/Jxjssu0jsubHRz0XqJ0OGZ/VtT/BM1z8m0wHSKAzdeXvi2f2sf9ltibmhH
G/u75KXFvCM6FYi7inovBiAgXwpTbtK1gpYwrrTLi9/MmDMRADOhx6AMUWHGTnl8
9WZHIyoniFk7jY8S1euQ69Rm3ksQFp0So9Yz/Gn1c3PpqptUi6E5KFAiNEn8uQIa
NKyEatXj1E4PahRkAsA80HvwrKKDa4hz11Ebi3sdza4HmtQyNIR3UV4p+UgexEhn
utWHJHEX37qr3BNUzRmz2Xfw9fVHIEHSIc/YWpR8WNcnImkCtMjkB92O1Y1dpDGa
LAH+nO/FlGWwJyi1Ithyryp9/CT3uiMkX5cJxhuFUQ7b0KCHGeEkz3YHLOr5PSZY
+6VT3eERR813cFt07LQnfe/qPcMwbgD7+eAw8K1rH4h9UNbmn+6Ymobu9iYyuRFR
YK1UCCEPeVp63d5iefue+lZrZXxyvmwhMSIezcLQfWlqmi0lLKko0gFI41zLHIiv
vNjOxFBrKx2JTeSpbSW4tpjgDFc96IQ24MCtPQkqwdL9pXxdWxj6rVJv8xbLzOUh
4bdOgDpVAL/yJ1UIbvGIJmjSbTTdbvt8iB6+pzdQEcsU5/RbyORjX05quyjYwxiF
S/b/CuRYzZtZN0TljcjXfKn1pka+4BQthWPFqV3YbWC9hbD8Y1JOM/k3f985XU/t
7lPw/2qNJ92W0b1lB6ExUdVNwEQYSW2K56ijaJb0afqtIHARmR4Is6FCj90FuiUh
+gkon5mhj6nzf8gcp8TvwUtkQ9JpqNsReVi1iBvSEoMZzrCrJ7/82vlYXK+DUH8d
VXwDgqCzhp19V7oT4BVeLMu1nqwkq1rfgVfYFh8yUTtAbXOOxweLIQOP2GQ57wXl
WZl5HfoOnYLFDVeDQ3kaSsC04IzEOL0xy15wjii6vTueJt7QlCAFqjGz1Kyfv1M6
A1a7bGpEiYK1kPbB3BxvTMCROXUdAanI+LzL5XEDkTWQ9GkE6gfKIuvVxMlK5fGs
kFYmjdQe/3FKEloLOOtq7P53ZQm7NMnQhdWDa0zNcpo2CngYj2piywKeOPxO3JZ7
Ook8d3i4fUyCeVafWZQllfE4XKqoF9u5zCR4bhwu6YAEjsHr/H3JNwPZWVpTR2GM
h8fGVcAQQDGSxZ4fCrYBpZpE4ssACj3L2ST29JPOJvjTw0Jy0uG9U19Plh9hyWiV
kw1kV22sFunM/0cAFJLfZTkauuZbCE7LHwqV3LH8zoXcbID6OajsV7KQm4FUwiPM
s6gIWYByD1ZoEenRNCt83+MFaJXFmhDg5JAQFZYh3NHorGaMuMFuUYdYm2TCNWxg
she8rLqBOnYLVKdiOnG69diIxflDm9HC0/uvFi/TRvhIklqLD6Q+iCEF1Oh6R6sN
7DqSh7SGsaL+3yPNTfcy6wE3j3IPsmi3nNR0ljDoXByPzlcXVa2OegVvSvt2FDFF
1Pxtphnve4De+WHUjYepy/ycMAga+7n6rN7RpkL6h/aVUIpU+MIReRNWYyBBJsIL
CgG/0iWqcUB54wUBy8rt0slRGsgnnY4tv2k2YtFcoApETQ3hd/7fqJGKN8lnJ9+b
knUGkdzGtKqHT8GqXCKwpfvTMUd8dn7T5C48RjrNUaFkYMDtwhqwuHrvNVMMz2Wo
jjo4xAqHvSHTblKX/F2KKVyAFbfb8Sn0o95BFVE7NqpM0j8LvGb5BpxTLwVNXgPi
u/HZM+Z579tjAwWxhG2TYke/1ShFtoh3Tuoxdu/JDvMv0zvMST/DPSegWagFn6lt
kR7bT923H2nPamG2wwA9LZaGP22gJRyIgBplTBmP866NYeXHgNIkr58iOo6Ad8bQ
ClEZW4dgvL+rzu+PV8qFR7eGJ57bIl3Cw1lPAQdwvGW1Au88t+ZmWQqUegtJL3tP
zMhRTTSvgvQGS3omjfolQEq9JhHXIX5LRbFo2zobNd7DkEyhT12ns7icgw1gYeAI
5NOO3oApclffkDICcXRfO5b+qP8EXGEi6fc6qRtQBL/aXqxNNggwCAWTtG9WBac6
TWISLZEpE2cpa0gNdOr1dpGcRlFabMoSARrY/2v/suZnpeK6ntdVHy+BNI1LkyHU
Kg9ELxWugSdidfli9RQntR0Koa1j8BazsEFOBVJAlm7S6+8fYIWW7AiJ0fYKxV/4
XNcjrnduagTzICQXYsihs7MlkMehaqIsx8G9lgGnM2cnSJG2mTYW0vUjsJXH4hss
H/yVFld7ZFw57MMm+shZjDwzphm1eR13EZ9lScaMxWoyTDNAHcKKNMjUYa/VS+9l
DvOl1ZycM0TcUARWKmypjPiT3darUkRuisutUHct7aAqh7+b29qkwwM6Vz0YBLNo
vmw5vEk8KWRPHBsCdrrheA1f1PGAyEH+qTKe14pdceZ7nzfV427d3qYj7i5RA9hd
BePhKTq16XXTr2Ig1KrulERNnp90Ls3YeoFzAMs8XuFl0lMXM+Ft+246qJf7bP8v
cTK3ROhU69w7ympLDbuaHExq2z2yIdaB+jm8Bqfg9on2oyPUal6OyWfExJQPghFA
/zNZ89dUQpNiX+zSPJbx68Y0/wLphAqW1Bk+q5Hhnf/vrQgu/HOB9slzud+vH48h
JOSrR0s5q+mSHYwKlBp2Dlq6NEVVr7sVCCYIypekukdtXwcmS1xATU9AERXkyiWP
Q8cVMR2ClETzFl8A4zbGl2vTnoRu6xQdYeAwefyPuwx66+V8nfeMOHEFYw10En8l
YNvc49Sj9SArpquV6rstbVsT4xXWBIMFJZLWOvuXBO8Vq4oxVhfuToiDmTwCoOMj
OQ3eF509dc1IBhSBW3Ds6nuE5rK7v775SpFiZ3uKihuJkKXWiN5g0V2KAkqOdzmu
u0WBZVFafqD4ypBWiJZsowjAeneKQqDyssLbp6iGb+ADfLSm4BSvFxMBYihFL/Q+
O8TTsDsCOGLd8qN4hOc7qWDYdwD73Ey1lyoXbm2DigSK76oLGGYlf7WIuRjPDfFn
WABziU5pf1YtWap72dmJNtfNT8D/yClRYn+k6hV5DrLBNw4/5CV0QVNcccnhO8tj
rb8uFsm21R5vEgCC4pdNIE0NvEHX/GVQNARsUjULKJlh4Y7sPt3EHziJwFq1GgBC
I36iIYm4BLcL0wAvzaQ+GzPj+y59yy9By/EaBHRYXbrCjLqf08OzOkjbTBbbGzCn
2o4QcUEF/hBbbkzIxFuC046Nq/ALJM7hZPICH452xGZdzhj9Um4SFgqN3mhkdVpd
dOFz2lSKxKtHVjKGIsEegO8NgBSoFQ1pBgBaCKIoW0iP7hOeV3UPP+gc7xi/e4io
mIceFxEcvBvnAmDwrsZzzTwPZDAETCtPGQIhL0bHnIo=
--pragma protect end_data_block
--pragma protect digest_block
iQhIE8DVyrrip9mftNDYiQtR9Dg=
--pragma protect end_digest_block
--pragma protect end_protected
