-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
JyToZ8qdS2coxjL+Wkq4hN4TzPKCMDl4KPCagV3rXUK1Yl0mrmhtzDUBCKKzw9h5
Eb14WDlQ+sBUm9PBeCUJWjLy8+HmpJwKgaaQQNgcq7ZFWqXKSjqb4BPknfkqICBX
zwwyNOddxk8ZA+mWDg1qo4rk+Wm45CVDwfvedx8onNnr4ecjki9pUg==
--pragma protect end_key_block
--pragma protect digest_block
Us+m6t5cAn2u17SRPGxktPwIKQ4=
--pragma protect end_digest_block
--pragma protect data_block
zrq8mTWKary+sF+Sq9e/WaqSe+6k+GkhKFt8zkiXMeSdyta6ZN2gYPYCW70zj+K/
sa8NApiQrW0kCVBXI+Ix5aTiavkhd2aI+05umBtunTBDwdyudWYiUm5ncROLS9DO
3wIGA6z/1akcOdCU4eWm5KUSb5mhmmpWCjuxsGu1YqgTgykFmdvxMMtAY4Xg3SEg
IzI25a9Uf/xKoTI9+Ra+nNIGmEjKpsBvyOATpN4mpIMX9ZWU+vxwDRBajlfE/PR0
UDQ9K8cX586qnxaNP5pAYIy7hWlD0uui/7KdApmYrebDmg3cOPbRGSZaCS9WuSbx
khUG7wfIA3f0L5btRk7DqmZhL1pkyg+itja7Cq/jmu79ePPGQ8osWRihzqNxiuho
kfqXXPRgRU/bVzuRskhJdwNfpRXs8LTlBi1KLIOv3TEYLPCmRbcQiUgMihzsSLJe
y/Y+LSp02Tqrp1ARPCw9fDKbZ54JYs35PHV7icB0++okZjzlduupeeYFAO7uUQzv
E+HcX7kFWm0vNYMpU8MzMuAy7w6MERvzImVfPMHJOSyrfzu83i6b/gSzjhoMDSM0
E88fr0K6mMpgKcnJJIqXm99p2FHYwowaXd8sVq0cyssPdQgJj0BAwym4Kpj4SSmW
OlCIPid5dyfkEd870ErjiL+GBbX6KyWfdAdSl6AsSbW6yvRkgzV28ngjJnDjsCc0
S3Au1tHPnORoIi515jO4C0DodQ9mFeFrc8SA/u8snT4VXiEZa3APEUaTNV3CE/99
j4f03hXh2kGPnVuxXy5/R3KG7B7kcZB9kFnOvn1Vwi35F8a+1IY5k05w2JtymHFe
uN1Vp6zz+FTC5H/JwP3YDs95Oe9v5QVU8FnjCzez+3LPHCR1EXyDhKBfqav9ypq4
3N2c0z4Q+hrVKzifqU+7wgVy2gCRXwxV+vzcANVjIMfG+TEKosHWWGvOvxwc+iYB
ytN7wZ55UWQAmTHETuBqj5QIN9OVMye5enten/hZcLZxrRtP+K04NHcnx7ulnmty
eP8weiTJqEmrz/FMpo+/R8svpUoZRvNeXGh9K+Y9Sb520irgGCJ9VA98SKz+OEHm
alAnaSpSPLaimNpFMnDtbytcHQrfcakBZvbSr9PA6BY4+E1aKVTFMl+nv95TFyZo
oApRhsh8Y0rwuRgYmySH07HQt7gBC4DpVOdbJracFIkg1vevKiIZTWAqEStoBmb5
pZ5kBDTKdFeeeN9eSaSU5m7ZkE+lYco+nNjsVrnrZEejTBbSXWUZVoF4NdkcKQpn
aNyOEcmH4vtt5yJiDb7YTMKl3pGYBgVetpw7U/TCkeYbUL5yuDSQX3P1yhOtU5Gd
EcbafmFkRPGGeKyJ0P8WSYko1B8ARJrZ1VsDuzPfuEdyTK/Z6vHD2qwZ85bUAmWD
FmFUjv4+W9j0OiU9yHCGdiYUbsC6mxd3WkFT8rsI46yovPoNdq5V+orLX7xNBHM2
EQFQd56wKxg8cniBegWiOWqbUe+dwxSSIwUunV2M12NBC01EgA5adLHD+sDROopV
NRq/l5hs0cDxHbnmWtsfXWY8ULJI1fx+u8Na8foarBNFfO5+Ge7KLRq2ZUlz8dCe
XGUeZ/xFz27rYIJhllmJDfNrJmBmxUO9YScu0a+u0opv7UnVAH8X2Wbs0hIhZuhH
bLY+arNB8dFQwQV6bWIwf3dH8+5i8wE7cH6pkFT+7/2je2XPso2dk5qb0frYsXka
Af6qtmAsdeUhcKY3o+NL583NN3qksJ2/7gmN51jl4ygvIHImDWMt01ggo3uTkM99
pKPUSKe1qNRkMZylGv8XYkyy9FCPe0zuHholt0JMDijDIfLdz1dUhxYRvz816CHD
1D91PT6Mcm+afJk7noyMWZ7zzFFKrBicL5uM+i9nYwu0sp/ckUjmqZ90QysSc0Gw
KmHfEInIZ97BQEAnJLNwYZohiL8sEK6+inPQGHrbgPczqHFrdf26w6RbZg5Tobe/
zGmUBS+CW4ql4JXV4pcEIsaFNeZnUKk+M5cCLfu/HkoaEg88Cd5xrflCZwyznV69
Flsrjj7sbgT0UdzTFMG0iSx5SPeEW1HILzrk2S8vhyShJskny9c6jAr2st4Exv2/
k67ZZbObytYZa3grYv89XM46UJUeL11e80ZymZD8dO+SZ+IBV5SSbLbSrjVwVKi+
lTuTFP617g7d4Th/PdakuDMQLD16VaiMyI5PDSntdSJYYjV31OuFWvK/DpPV1U7R
1w/F3eVA05M7T+VwjwIz7P7ch9p4us+nebX1Tt9iecsreb89/Fle7mVu7CbnWsVs
PD7TutT2XSvYmD9kP2XqxgxwAn2B6conciyeJGmWEHtxYK7/x5HNOe/aFhOEHcoU
BbmAefcGO7/2ZlMmifcgwAv2Jq2pC68DXLp8YKGZ2GsolsqvdxiwJMu6xF9I20/u
YbmD9yIRetxS3k20wWvbubd6TUOs4Ba28GgEkOOIk1EnUnqkSbWFiVQGZhSL/jyz
cnGdz33e2Bo7IPl1PLFA2wLapvj/4mFB0okwfJ1bYBdFcrvoMWHheYJpEvWYd+3h
6EGkCVoIDNFLZEyIpF7YvruC4aLazRuA+0AiY5LsVY8HMmqdtxlOU03vNQzZoQu5
OuaY51txaHbLYAzL7dzHA52aknnWBwRp/N9oebU6KnoGmQvutyo/Nn3ug/eBuJnY
LFHM7sg0gKUpgxU5wPp/GLK4kzJaSuLK7c/bisYEIoOuM12D/m8vZ0NPE+u0Pos7
Bp9AJm9P+o4UcHfd90gEJiM3b62DQ8cVFxWe8M1rIgFHJIZgQA9j6MFP9KYBOPhh
WOiXSY0qkcSdSv9B9R6YMCwA2XIh1XiTH97by42Gn3E1JCPeyv33Wnx4o8RaJqqh
lXr46XU7dvch7ZphG2MOoLgvq1ks0/QpZ2wxVWEPkrUN361Tp/SBQnNkPFRT8QVN
7HOf1r2W+GfSfuPMHZEmF3z0Bz/WiUDtH/+AZI/fkxLL05/qvl7hlbK6lLEFLpkq
gBFoVSB95FNIRg7nGaLSJAW4sJc6sfUCXr/eDhw8ZMIS3KQuwgzXZqLu8my5zBCJ
/cLQ4O9H1ZJ53rkoY73mqm9ELHBvaU/FyOD467f6RgorfuLMigfpRbWn6D/2uQQt
zURYQBG185zR9BlVHB+cgXSrxhr6p1LA5Bqqc7MqAYKWtJKrMXBTq9XO3jPXoow+
Uk9FK1m2CcLxs4EepRdVAqn/2cAJUvk5Ytfc5Zyq93mXUcD2RJla/zrdGPFEAm6q
jgaFmFX5+q9oTK3/PTOw6d2kiRASpFor4oFPS516Wf7MMPMWbtzlb5iorsojL8W1
eElTgnusOl2wU5YAngoWK/1Qcf4UvCZyzeyokAgQpMa3QS5M14+KaO+os/RJoIuq
FQeYxyj4xpGxk1gNtRj3mwM7mqIwg10OruLdWtTUnUxN/jiezuR18UuVl2X1PLiM
0G2ZzvXPx/dxFwYEVhWI6rsq84XEPUAaPvdGy6z0S7u02dy7NnmwRV+ETnNjCiHp
kzSJrHARrm3DFXSdvgZhxuRCEX3QUwQv7DN96bnuv0wmA34mEqntQQa74VnW/aX6
q6UxqNZpLp4uwbzPPhNwgOMzlLQG/I5k2972yEXD4RMQa5TUQRgXa3R+sjHyCTiJ
4mADCAT/CmVT5pz8Skznib3vgzrOcchQWunF6/1upUtEMomEVnYj5cGCp1UDZcBI
tFKIeyR03cnhUh6UAo42waHmpjXUm34P3U4Cw4Lr7pEcK0qnl+0Sc+mcu4Zby018
dzw+tUATQFM4zYP7qnFw2aY2ttpkyXTT3qhSsKqXS2DcejeCtW6pwd1iHUNddnqX
EhtgI2ka1Lf79LHC2oQbvrkrJ2rqtWlKt2gsa9fwD+axP5ab8hnoX3SXNwtFx78d
n/kGfPSKVFG3gg6Z+DuQqbDl+9ECOgD5pAGJonBj2988vYWwAqqxYGKhOnMODvH4
ui8fyWw7B5Enh/n+xQPnxmpm2+WBlEIYturCIF30MzmfKZRS+qJ+AbNs4YKIgz4I
nufcejOgy3N27Yc3aqT2+KFF/QcEqwoxPapqcZGC/U16M9WNoOV0x/wKRBQurCXO
42cj8QKDVnNFlAAreAtwYq7TjCfuJGkdhMeOV+FAr0nW5IKOq590mGoxM/f8nCGH
n8FL/hiBLkE+hSjGjMNhvacn2XmxG9ZY0t6DZ16RI4SsyaDvwfLe5KP9B+5izgtD
G/TzKf+HGfbd9rWuOji11eq6B9xh1UzT+3sGUaVDpAVV6jdglX0S6vNpPZvylsFR
PGUhhmgTbi40sFZG/l7dlCniWcf8UNtP9yWgdpzn82m4GnVY4FfIK9zz6RLHWAdw
nFWlJwOlso4aQdqZpCuwibFKCTvwxDED9kGk7XSxSgwdsRLYe1/+bzGqMOx5FLUU
ZRHx08NpjDITF6gr8W51alabb+eq2xJZFJSiGtipMGaNYMRDZ6b2nf/YsyTrmkt5
rrTPIniHbakPeGjKkJp70ydyGZOitVSyIXsCXgYsDZXzMfX4F49yx/5/J1N94LPx
tPHXJRpuhdac83pUuTu7wLeXIj3GFxrHp8jM20DRBGgfVEjonHveZRRISpOBRWop
YzkrgYrfMEJ2204vRZrQDDGKoRBYKn/zn+P6NfJqp8dCs0TJT7tKWH0S32ddpcKI
qN2VukCx/raNclXsn+gkGQSYLV2Rhn/zMk9vYd8DvMVH5Ty3UOv7PPvkS66ONpOG
MGOaJ9iNmYdxzBWrsLHSr0VeqiaumxVTjJWfIkpldlPvJgxrmXXO/6hYmeCS6N+m
mFy6zPJLV94be9qNbs2rNMb9Vmgi4E0UNUFsQoUNeyi8DFAqwopjieqM4HzmgSJ4
ZC4/JQ+C9m7AWj+3+MedNpQ3lPfSxXEiO3AsfdKVkBQc+Tma53nrsom8RvQchuDb
Azsp8Wf6DEPWp/ORUdIdJ8+KInIupSslu0/SqjIJ1AQiO41hbC8WjbhE7EMV/ZSS
Q14OCNUw3RM7k8uJKbmi3MHzh8VMq9gRI5H1sFsuAvDHi61zoC8Os6Te15uJc30Q
Y9Eb+5M4gxo52cQ3YYynRQMzzeCHotGkGrqOd5lf1HB1Q1T3gnGCwQ2to36hNm8l
yW6+eZp93wCIEyt5x/okD3Z4Ri/qnpsnhFUP7KsUaXiomxJG1eArD8PTwX/n64sY
ZXjk3eXUZKexaZcj0PXgpkNLDCdzEPLHpFDNv7GeuWjOtT+6RTNKYQ1QgX537mS4
m3dpkfOLoUN4ibFh9LCG26UccabxufqoHJBqWUw/a9VzXJJ1B9s46gOzPReE5Ubs
jvJhKVa5HvAFpuJKVVCxsROAXlje+/o0D5WVtJisOwPhMWHnSLlbrqkefBKhFBIi
3czzvpewyxaupkDsDWauQTIhFr8LXdkSADadkywL/5+4iNPREd+nNqe9MUlDiPU+
TnOB4jv7L7ww6k5YU9OskUCu4VqZ9UlnXK58QqNeZquDfOdXgreRgPsrx9MgN3z0
SesIsvdnoyD+nW1DuRS2AB1G4aLZaB2C/Iy3CFpEcq81KtHWmDawS1vPMWFjvCv4
Z0OxyF/bBvxG/idjQ2POeFMjnFxINBM1hG/1elrNCtmd8rYPFjUXUhNHj6sJtURw
jHznZwPJOb3K7QAVB3ZpWibxxZYyxiAaJyfDFF8xSSnx4fJY8JohAszzo+PBj53K
a9WN0lf07ku+WVpnr7ksDaGH7i924gw6AKygqTKVJ7WDWR68IbHyF4g3m5vqcXqW
DLH9m4HKY2dc6qGzPxfsRk44sQ8zCj/XKlAsFt1UZTHQFhiWjFvAvT4c+QJWJSxz
B0snT7xqynwgHwnuNWbHt9M6Z0xG2B3nsspRnwNs9YleygAadrPw1wJtxeDAELvu
8/3lXoRAzqOcpeeitRRVHo8tyVWEZ7m2dD2xqEFxHxPSSZQBm6gynBbVpON1wYOP
ra9CarYjaiZRC1URggOmkDsNtYCbDQ62BJhJVVhvYrPCun87YyMXjQ2w7o8vFXFn
gRt1JrSpOa/ZQMwQcT7t9htvfObrb5Gw90FBjSpftXdU6rs9LPJZjX/7kTxWPRl9
lC1mCnjnT3UrtKqLHNswsDOfCmdjHZkfO8gF7exrO2n+IJjcXvywLTSneLTku7M8
sUK+GRc6X1CWFo/iUTe2o5HSWoQGcHNrWwOToMh5VA0RXXEf3XxPnKFjexLbKnqq
C+HCyIrMJzEUH1/Iiqxokh721o9BAa8tznWQv+OINChxEP86z8HYpEZKht6TNdSg
vOz//zvMWL8IqM8vtP630eqhULmIYY5D5OaZdBMqe3zSJg0ViJURpeKrazW0XpwJ
IUbgLq167+FnqR0XA8kbH6pNmBTU8K8Taw6oXmdhoaIvh7kqAtWkg4/knL5nHw7d
uufLS2xcW11+psF4dM130Y15ct/CfLYjsd5t8PtLKzU+DrkAiPHau82RgsZ+5kiV
C3lv3hxD82rChVgLKIWL2FXsonl0lDYZdNEHiggmiFRHFDaSARhWsZJJew7aHoz9
9x6ZQ7u3Bc4ACA4SKLMmJNVGtZd0/MUH6Aq+aQvcFIZA50GMLZHpqwYR6v7ht8sZ
PS7S+QFSvk7nwAK+hKQqhAR/dlKh0FVMic6ldxW/AIKSai4UqIH0nKHj+d6YeZAP
pNIWlrSAQxWVs9IZuUQ0GRBWkYT14Ucysw+UrjjkzP4yEUdxcIiDTpGNyz3p7nak
S2d6o9p5HMnhKtAZ6E3pSyOqT+IBx3AO5VjPkaN/HcSh76xpgcvXqysmQs9q8I0F
oasZwJ2WmamtSqwRP++QzwVKpcTC3L96qShDon+PjYvIdJJb3U1ox1HozIZE+fyS
xlGR/Kp9rvTCWXHTNpKWxJ+S5uq6tuxyKT4upNM4rHrGYgime+25Ko/k5nuytSE/
srCu6C54xWeThNpBKTvLyZ+mDM1Ml3ojJXLJmmO8oRk5b4HfcIP2HLpBjKvcokgO
1Zt++7gDAMP7OvPluXxTcQholDV+0QpBwKdELs1h31ZmXC339FOJ271ipZ/QAdD3
jvCIbm0hqA1ocdvpp6lAy2QEfUJ5UyyCBi+eiTzq0f3daKSdHUhCLDDJlqoOqlKj
tvkhIgunpCVa0a6pDlM9+rOx6iIWTb/DkTnbI/AG+8SQFOhNeGZ8Itdopi4ezjbX
Jygd48mwk8J1K67VjKbpA7tVtn3bF1Ac/KsabVMHbzIYhxW8vvXnE0EfELU/mrST
ZhDdW68HKM8VsTS9mBQZn21KuFMlW5qMlIaoskvzzYeJsa1nenhy8aHsdI9tUWQT
G+FwEXlIxCDEmRei18yHhtfD04mPx9Ej2HzTk/NXi6ip5CvUGyI39/bTkvfQ8b9L
ITD83Mb4NEdvCgEOc3jNmxoEwAeatRIDM1qNZd4Hg2rNlBbYaLDxGACHglHhUi74
lnSiUQ3yeKQ6ZnSpnlm+v7mx4s87Xsu/8LtKjj/lawyugJ992wvKGahLdUfgRlrK
7yTUwedBeSII5hkcAmkH31dULOxM2JRpg6+CEMkCSyCnyaZj36rVA3HEEexjWjA5
2hxxPCx1y3bn9i7/NCUJAghKxxywYRZgZJstEUPUUz1El7C7mafzy7eGjl+7NP4m
Z0yLmFtI9EVCGWE2ZRgnISNz7t8JUg811N8PW0meCv/dsfL7CYaR0iANnySy0GKr
S/wIjwqcu/Cs6dahXLV74UEEL3xIMPC3GjH6f9AkfgQ2JS+iytUQ95yL0WeXLIp+
R+B78cqBjDOGeJdSKz8YKYSxbKw0oj6NPgQfhb1tPJNjHErvd+G4fM0TyCCa5p7r
opgX6OdlugbOsDUBPXxlS9abXdSmOCX6ACGDlHC24f/G5ZMZd4jT9EqXkgBL6JHA
+/j//03DAsZRq9Ix/CnaI2hMnqm/xg321d523+VkbBcZ25P+Vw+kVfTZ+gaGORfP
B1yVPdWF+1Kk5BbOHcixd4iOFUkvO6O5uGnny/kMs/ESKoOxQ9laTuSF26zLy9xS
sEodvThWixyZC3h313drZ9JU8LEayq0j9cpGkOv0K3r0zEfljeIPgvwGHb8F7r8a
egaptjVaDcVtNc/q5DIt3lk62t7k+QO5OVRja+a369ds9mqGIPAld/q+TYrpv+Pz
HoReHepYYhYfo+6v6wURxQRmNfxlVB+kd+Wd6A+bjIcvp6wryZTprMazY7zhIMO3
RQ7oskvNMoQ/6wjj8bQPtcOR9BTGQMreZJCKoGLTdT1Uasj55l/wiaAPRhw6c+rS
Tx3WyDZ4blyZBCeKXsvLiSMevPLcMYumzVEkFasrwzL78SM29g9tHuPgzYFuas4O
VMR/SL0LhwmVdkM1hN4da7iKWA5tO1rr+YYecl3+yMmhB12m2Rm9HGqIsEOwO9Iq
3EfPOuY6RTfwPUbmmPLWpmK8/k7Q8DL0k3F0H9CAq8+/XaYVUX8fWrOzE+QWO/8k
lzAj4jiBQI9iHM2WtHWcvLG30lSl0Hm0XCMThG/awaxbyc8n+WcYVaHbV+9+8dXV
WpoY72ueOpo/DbaKAqoUFv68D3YHsMOanSI+V4Pe6IXIzmGN6Cg6ao1US4mTWUPF
kqvqyNuv4MQZlxKMVqXBG5rPn6UxF1KOETv4gcFZfwPFFoF9pW2d2xSTv+bI3G3f
kCCJrBuuGI/H8QB9Anp9tXwafjZHEwGQzKXgN8vkXos24MtDfEF7PZK/6plOnFa3
4BoI+y2OXyhBz1nckDP3fd/aoGyhIBZCUODDXA3vlntHGeZwsBvSjVzakQIoPssH
7RYS+l5eEhY4GQXoBUVApYk6PCYGAQDYK5y6SyVSBJQ9qFX2yqN3lXyb9nhCz5Lj
o/Pu5XrZExaUe5Rf42AqccmJ+yqd6T0Yog+/MnCl3noh2SWDM46pjgYY/Rg4jUKn
yjj/F9Qr0Kmmov2ttTZfihUSWmNo59NW6ELA9OF1FEqaUXN7TYHJCifG98w8/Xuz
9Agz++lduW4l51+YHvRuczpGx0BLK0bE8HlaC/Fb8+V4d3nieewaMhQQ2FFoGvFk
yOLgpioMepqEr/XTROYdk9PybQJbUU7tWUGs5Uv9nbZUL1SP6ak4MCejvccLv7Ce
12plJ1gizN+ak+OeS1rbs3B2C1+Mz/yAn8PywZO8pyoGGJwNn/IEoy/XS4Oj69IG
+moWxhl8k0//YTSlqoYepm8fjWXYiKeIdWLDHH9RN63DsApS9n/yTmUSlRKRPdwx
5Z/pFsTfYuNthEbSi5n3JW3XSe9ObnFSdC3L+/j6uigfwBIad0k7uXvKjWjx27f6
oJhYmbWYu6K2ets9Lkv1RAfTahhDDSBEPQlhV8s0mYCkMLcitIpRjeFWcQm61J1N
u/s2oaAkfyHJaV0BKlzmOZajKhUgX1gQFeB5ZAo2AFvrZAY3+SFA89HixrJ27gkN
iuaY9u4CpV4TChL1ApRjkLuL7exl5P9DxGDou3fdE9P/5n+bxEmeBVzf5gjUUfef
s6bZ/E2eKouybW3jh4lwdpTVOqrNRUZYzb0MfrJ3EbhAQRnGZ5/tT7kxo5WgPJoL
dzxFiZgvayEtWnhnTqaGayUTeno7/HnOlxAECQXSCfFsFepTxgpBC0VdRQKviayv
E+sbsxFQOlP3vnRJAj3RNHwWJls8myKDhSWPr5RGJcmnKoi6QTFf7ErqHZcOjHDj
A2NpcI1KPYWfnv2pqaG3ZLZUjhxQl/NpMqIW2IAOsYVfex1lHodQXJzevfR+HbwB
Xrmw452SAKpb+lcgJkt7HEHWmDpAuqs640XBaSUWpQICIUK5LbSAWqEB94n1wq13
F1oq9yoDiqk2U9Gizqqnm80q75uQtlclCi8XgfG/avB2T+Q0lxW71HdReRubxDdh
DGC8TaW0fuUNIJXOUdY/hyTTNoX3U4l3Lqdhh/YOGAkGi33hpj9EFn0Pyom8nuyi
OJPteLK4+VdkR6Db9Lua+mZgy2rAJcx5PaZl+opXo18mxqvQscSf3F+RB/47u0rC
nQ2RR+8sAsVeMnTsXi76igiqyuY7WZduNggCXd2F1zt9vixep7saDyxHA/i3bHIy
462xkA2U+WfeQXV8E7+OYShToj8Hg0Y9YuuTurIjzcEiksrNQM9872NqQNXlvFIL
n9T2qzfAqgktK9tOMNaDUKJ2vDd6Jbj7iEYQVju8aOu3fJH+qHm+P+27c1esW9kW
ozU9kAxQCa8mq+mTMvEnai2zLuQtUJ/25kktO0Mgy7tmlZsZZrOIgf8p4w2yZjwO
HWQYQ0IWYJISnh7FXH/91LOOvaOgoJW0GOAU67jaems6gLLNuATYOfnOcS7uniC2
SCKKMxb6eAO6nC7czibScArCT3gnEjY6w2tI5hHSK190C5lFucB353lMOCB4bGA/
MGhL9w0n5m9cAG0V2WXxPkz3lWftf5xhtOqc+F5SBGyiZZeOb1i54BZ1Xz154ziJ
0blK1p+xmAHBoRv7OiDBtGy1fyHxvQMWNSkw39Ekz8116xxznC2JE4d3N9mIHFyt
MLawm/tMt/LTPLXY5RAUIJ2lDICVg+s5DNn3luJwUKYvq2W2nUaTPX3LMq0QwK5y
CbhyGoYI+QjCokOivMezvx/nODUXz7rGHc+2+jHFkiWPZ6FoclU/bJMW86A0OFYB
6JYk5x4+xgXlXG7EuJLgQov7Rv0u1pgVvvYGPx5dUulx00fnzQyTN+IWxUjHtGcd
Irdjt1dPa2xHs/LnNfafFAByAffH8c8jXYLlMTY78EHkQ7BLVe+b42F4bT/BPVpO
AS9EBTU7e/vU50BvlSyljDMhDiD/uy/aNK0eeGm8iwz1J3N+J/rLOfRr/3PEvAa0
Vn7tMWU8oFrG2mBn/4eRdGJH4+NEqq5amPwcNnk8304duSv2ep5zAOCddqF5a7ce
pbt9P+N63E2YagUHiz0FBHLY3stJ/0Pyx0QvBSRA3U1DMpg30AC6FNyrzbBczlmS
a8bwbYcVNzL9IbK9Ool6WOw8dj1/YkmATf8fse6Lmw+ZU6JDpuPQwmfgQrBQrE0T
G8tyiTYJt6Po2dzX1Td+mMRz40tNgGpJtESs3yV7Fcgj7y7ke8acwn1X9TmboM0S
otJ1NChUNFplnuz9UNMMM33JzsuNnUs0s7talCcEz9qMtqfllGL/8t3/Ug498388
XDCXFTTpPvttLSDBOQT96uLmGHyzmnA7b727LxAP6gkMl0KKwzTkFgNOoQqEWOW5
N4MAoM4N9bP681crLpjMXeggKbdncTTX6ZfzruArR3g4ZKkD5uVPyjG6wcTrqScu
5ID1JHsXSP54AAJse8LD14XTGM616HwSHPvGHoRcbPr/VxygNkwXwIxhpgQjSch0
lJL3JftLr0qqWVVUetyCRDNuXd5UB6Z9FmE1mq5ATo5B67tCdb4rVtWa3Syk5GZx
RmmoXt1FIemgk9o2IytMn/env9MkbQuP+1xufSBY9UEXYdA3dERjoMiBGWlpD+oY
fwO35UxiIR1j3U1k6yImFga31MdIUZ0/XQO8puTNeTK41CtXiVNnfs8SzUWsciyW
7W6yy5JLrKd11oGZcpfbL9kzGcSiAqYJCqJmPNhKpIkEhNW6GYE/nJqfYmo40tFD
YVNc8wxa+N+g8bVErfjAFWxSxF2xM8oXVboyGhtVWda2JpyjHl/yButROmdatuVY
g4SgTS+1HefoU8O+mp0ELjpNj69NIZlWIEg0omeKVHhkZZJfn2zkCpl/BZ6hijBZ
+wiVC5hmg2nh8Rt5k9mZrNVH+agAO10M0SVONf8/FyT/5nltLHiSfLjm3//qH2eY
XFQDa6LHMq2Tz7sTB4hr/fffrMrg4XATd5b0G8q6OeGNHb1LxGMsoXiMNZIpvPab
r+JtUGaKfryXOxURYaQo7N8764vjien4YaGCY5Q590Ofu0uQk8XyXSdLoUUYudZi
rn+sFm4GP0DsffBA4yyUJOlD0uGWg00jUCN7fYvIs6vt4mO/E2404IZdKmCPXzbw
Gcgz1ZnCLXGbZ0UPYUXFNcmBFyrjpb4VRaNSD2ega/8g3YT0QT07kpOBwrFdTcwo
EJvmtm88sauegpDn8ecr1k7W0sCsddc09c0ltRWPckb5PxehgtPMCeTrPsVhYqzF
SWytSRlUbsPAVwayt6SbQ02Hrdhy62YgYEACRXqHobHb3LYgjX+/V6fTQuG8y+wW
wF6sgoY5AdkyJ3obT7g3aIZ5wyqUgqzQcL0FmSSJ18dEme23x4yKGYoVSXlb/XCQ
lLk3amj5ZNBHbqKbabnV0BM8rAoKkIidRyAgUIPisq0vZKqmx3pvx8tEMiUzfftw
hCTM4GqXQ04FRFkftZAJAPWucSe3UXd/IwwMPk/NECh/S7xlfxWBBysm/HpsXB/a
7veg5aUOVGBP2jUCOElyAxb6/GeWBJ2npotqAhRSr94hLCJp1i9d2ux5U+cbbzh/
oLYh0vQWP6OXJfh9JKcuTseOojKo8tW43S6WZ2CrKXkOHKf2WGTGW2/RVy5/q4vf
qmNN526UeQyu+CL8mltSNEFyCjouAnlww+vBQoJ+2MYb8YDJLAl/KBTx53vCkAkS
9+bDH21aCIQPefTgqM+MpYvx32wgkSHsit1SDVYLQinI6wtapupSxxLMpB9FXfvW
GHKvICBE7FDPMYsj6u6ij9kXPPb2dxRzjwWEJPl29L79AFYQotlVT/Ncj0B/TdXR
St6eYlZWwpumdbT903CPjjX7sX3KXDQf3zbBD8ftC5iphEGawfP+cOX00YZAOIcL
lHWMbG3zBkfMVdAexj65vhkPVPPkzMugSTK/FuVP65h3xteGSfRTqSDltbO3IADd
NODAWD0FbDKZRlOTXM2p9SqU2i+z8FexCo5VXN+MNEiV+OtAHQgabt5MJ+w+AwRw
881jGDAcpGdjyL3hAAN/J6PrBmf4pDBB0WKNtCgc+DV82sOwwdK45hiXlm1GS3HR
VHkliPtyDsfcICNdLX+FUmfKABlyFglT3+o9u489p07o72IiYaY1DDFEUG4IZszp
K1JTkSTN9meMQ59cyxszgX7JTiJdbLk11a8wBYN9uxVeQVVqlqNBQX5p8JdL/2ak
RDp9t9RjProBbAgEwbNAI0o4sVllFU3pFFU2dkDXw9KLPJZosHtcpwGTrr8dgTch
1CDc/TKzmawZsfz/X/SVT45QqmfnJc4PYMZ1EYmJ7/EyDNK0nWMLqfOopOC+UTI0
H8RK3vEpJNv7nN9zhPdUjjP6OATgMUEIsXx7TAg7BH1AorjcA710/DMmA0XyNIhX
8v9ufKK9BeVwur5390Ld/FVMuYUbsiPAORI+9wtO1f/BktXNx+tkfk25ePDE00wc
bTat2omy8T/znotp33SxLxxFOTabJ4wqYyoW/Ra6d7xeVhMtjI9gVwTmDvYGtSB3
zZKxPs8nrEvqSnJBgeGOOTq0ZQtPkpb+m1Y7XcKeDAyU+z7IbsEE0g5r2KegOzGg
MeUgIEPdHo8SJU1lcpgsua27eqrnq6AwbuOlmXqNqxczvRPHrY1yLWmlvuLaFoXs
yrNx2mf9R7oglLNVGLV3hea2lylSyMbQDDlHAd99BZ2Pw+Xm1QjlgPwK78V15cJz
ORN81CPqBgmdlUAz4fILNqjQ+M8fnmdPck8eDLwOnTUVuFqMle970Vwd90LhzCao
j296CADwXOr4cB/kpcIU+Rn3Lvqj7VOTjzj92uH8JZ2WEQSfs6uZJ+RMszEAA+T+
/1QWP+MfDh32s47juMflurk74rYaIV00xCblNeBEu/8TE9bFBacoLJ3SwRChiaqj
xltNDyUqVfFsAjdL+x07joKZF59iWdxCspJcpf2LCL2q8tHDxiwA5kz1lmmHaC42
85CGSDXYXtrZB+7adpZ0sC7UgNy7SzYw7fDV4+eT814TeBvJNHtsLAU42+EIXPzv
ZHHerZ8pwUcFSzY/C48ITFlorSE/hG3NE9upujmHuJOCRLBfpm81uY9JusXiuUHS
ij4jfthRUjPLDBROF6C7wRAaQ96WUo6tVCrGvf7yYfDkJIjZvLJIdkGAlhflGdNL
XiX6YEclnwDBdusXkDjEOqHe1Br/o+lsLN3ixI7vd0SnqaZ4qZr0JyTEbGus6wXM
D6BveqIdahlZhDv0XMUsBF8u3G1XOdw77RAJACNEWPLKyBQM2ny85mNpyBDKh7rT
n1+xcQ9rLkmdskLdEf6b5ETS+3ncNkRc4KwOx0tAKKAK5PVWXgtVe/TvQ1bxMm61
Zf0kyUNsCTVoT845e9Jg5Bx9JRtzDg0B0ThyYL0QxD3sHJE21DzNA4Ux49avlwLq
vp/t4dImxgO0af9WoZahSSW3Z1fGNYofb0afqvJsP1mMKH0+yWto1Q+5Ixv5nouz
6+QSP5b8MlNGfCQf36pFQmOzpuMAc/FNIMBQWrm1s6YjfB8INKHo15khDJ/PS8S7
kaAhFPRbHDtZye3JI6SpFIq81zfJbSHS38Q8PIvioH4d4XjPuhG7S3ESPuo9GqPJ
ztebB0BYeJV6ja5a3NPO/VR9yVPOpy9Upz0E9sSi4K86qP7Ugd4cxTpXaa5+75Pq
p+MW+dKNNfcvkDUVPwnxeHOMdTEVeGnEwPYCXeKe3ilWDXhtyhgtvsxTWW2H9Re1
6Y4yOoAdtyrEgpNoNCN4MgDBKAX/0UKXhIq/wXnQ1aSiMMu6t+ndPpIVvFx9SUu9
sw32oiC5voo4gVDeU3d8SOBVCPZQEJV94R5z+3KNPyKasZa8/2sq3s3n80a424Vo
cnbAP7tpaV2o/1CRw8NDBJa0OQ8Rp/vi3NXjkALYS6EeYDx3P1jMnl4WvWOZgjVc
igZ3GcocCGFP27IHGeeA1v/VAeRDYaLNIU0fYEnj3VAT72RU6/IFtT/ZeleNi9fR
xVISC8EXQolDujIO/7vaV2rsFBRWLD/tdsbOu66kH5vNIPM2M2NOjQ4jGojBvacQ
PMsZiWbt9m2JPTUTNru5f0UlyB6j/Xewg9Glx/8/Gfabfr85yXS+Tk+FuETFFpNo
l03Lu1pTYEXRJMdtDOfu7gEBp1NmXlfS2727NFmXBmnDmvkxPG2gdz3TMM8/KhE9
8/Scs2re6S1E3QS6W0WZSvdGjzL8rKn3hF1tZAGXx8SZBKnC1ffz+PhvpH64EM8r
/6UZtl9MQ0/6IJWPUDy9iUA2zOIrsIygOd6eWet7BGoV7ulEh8P5bgpgZvlGu4wX
WUiXXB15bUIdqbJF1T85ThxeAodWXx0FsjNPkpbiHCZrKOtYjI/zXrFxZLSr+SYV
e1B59hrt0StrFmsoFty30bjCepAJ3tbVJ28aw4MmQzNTC+dUir7h83ehA+sUCaRW
1mq1PwefAUUpiOeUy60Q2wztIrchpBCebLCJ8sJadTcIQNpHhjBPyusC4+BA3V61
q9IpBmltODMdNkLAI0kPB+1DgAL9GglRR/d9fbSd+pOKrUMW3552EOlT5edgs3I+
DxVxuge1K/e60wksK2sIbIMhEcJIdbdXyxpulS7+5vxbghq7dwqdYdS1vpzZfq0w
NNlIhqh+FrKd9YSMPUsIL09gpbfOH/h3M3Xxrw2k5xiT+qbCQP6V3JSZd2WDQhuc
igh6hPcYaZ5Xh/zPZOuOKDCvsdniNN3RVTbuzLm/xC67SS9grhOf47PPHBq3O1NG
MlpLLadalO2DrrT10GSJVpfW7p5YhjnVV0QX5cH8YJF3bcWWjWFVh0uCx427AWM8
P3/bkr60K7unDqy74sPCn7K62fyC7xw+L4JVuwO74TEDBrURbA/WP0ebDSzoKwaw
VxNKsdbkPsLC9MqeivPL1/xR+6nbM4Y841V+O0cKR0RdjOoTB41SbvnV8oQ0mE+X
r+djZbzyVCjYPIKT6JxOpTG7R5g53/kXkWA+S5uSrGxluHhu258AsjZtW2PaqRtX
E5DimWe+4cin/NBc5XGWMChdJ+7o/iY1J0T+Lkbf3qF7ia+zN9doiyWL5P7XinzT
PJL/laZWx0H6/qk9kYGOvrlPub9D4MdaZ3gPgUnY4CoVaxDy5VHFAJzT9PEL/RnK
UDLKO8WrIsIkQn7YyKU7xZa4VvEcPGceFTTvpCRllhIQrLiKMp15kS2e7FJKjpcv
vM+lwO5wyhlBNWzysBn/S3hIPHI/sH3MqXscku1lHuVOqpuKaZyvmeXy4EZg0655
f7VyyCNQBIHn5OjFv1d5Ccxho/g4jpT8b3xOgdzJx+lLIY2k+AiJTlHcyXahtkjd
jywTn7OR2D66g8I73K4mSs1qgPReaWUJjzMXGkYSB1mxHVLTKAdzKP5xoikS56GI
fj6oQaD15jdXUkJtdrdRSTaW6noGOR4BHdL0BvXO+GJvU8376xAozLI8ErU1YN0z
XBsG2BZ+nlJ4D2TxfIBf/2X/UG81DnSgc0SYQ9Np89ZKlZo0tDztgT/0eXMfmXLy
eTg8rd596ekI0tq27qiUFFLnL0cHtxGkjSLKU0gveROMm1OZ9/NFz1otYMTXKsbd
Z7PIDOKvwaUX2OxwQMjzaWEmv5nshEEwmb3JZAPcC9IFrJj5ytitzHBcv2KFOBqw
sIiP86lml14O304D4+oUBtGTJhjVT2UqPR2tb1DrsqPVk9H/SvUp5IYfuc2RcN+8
B9C1+sHukl4wAhNg5mcrfWc7QEi+OAkP9NbJT5teqLfpdPoVGLCTlRNC/NN3+Dzi
JLuhhqPRJ0wk8zpm9IXmgy2RGsR1g99JWONfLT1C+PaDcSf/Sb23LLAsVZita58U
gRr0O79AN+KTqKCIVjJTyK6RLx+mTxrMLHpcbJRbHVMLcyOtM8xSkcT8vL7Ae7tz
7D0K4A7e5uNf3YIKUvhTc1DzkaIGO75bsHqYKTcMxelhj9Rafiipzq23s5wzTe7i
Fsq33ZTZCIE43YvXc+Tf9NbOUD1i4PYq3Dd6sH84np43xYHEORnZoO5d/+Iq+iAf
zSx8kW1xPx2l0w46DXKcBB1myPScEisyTY9G/SBx7cWISV5CRbshhE9YNb0euJgP
R+2NQ4nfuGCscHwrpnpHGpHBid6sw1jvo80meTNoeT1H+rE0x0guMhYcE/dOAXJW
axu+ZzuAXQYYTRkutPcIV8urYBMxYZFAL0p1UgiBuyq4iX08/OshXAvvUxxGlvfq
+0TlteDfLj9CHyTHo16J121ZCJDfasgxE22mHo08CZIcreTyzEFkUf9upkNGAFl/
HoZKS6jh23WdhuY/3fZMim8dfxYu4l7g0P0HDrMzXi4EddiH5iuL5yr19c8LogJ0
6ZDEEd++V96lWHmAqhHNVq2Y9K51XHFvAwCNO2rJZNXA1RBtpsJvFPdwA3836JYX
goAHb3GojLO0Izyb8v3PWNeqy9kqMjYjrJxV2haLYFN3dxXQ+UYvNkexcjMnCHuD
SefIpLlcv9UyX8QPOCVLESxR5P8gH8A8bP36s/woBMc/UES7qgq2CZtTmBg3I0/T
bMQ1CxPKCC/4Bjw8UpyiIrjVn6tGiOuwRV+QYp0lSQIFuTBuPCO1ugN/DX1Vn8+g
utZJ08Rbd9MDnuKYfQSF5unEjavMhez9kPq5jqBGqY99wTWjhIOhbfRiQ2WfSDVi
C9GnrZWjEvcvpZnwPfi3qbi2UdHngYYlLxikxuPolla07nFv1kgLZPJ+h84bkPwh
lFjmTasgH+NzR8ZYDantoRWsrQUdpmxkKUhv81kGwot5+QHeDUTOjxINcLKIFik1
hIEGHqF80IhZ3O/e1o3K2YCI39S62X/6tfJFlhhxgFW9Ush+BS2jcXQDeWsvfKKi
iS1KMqWUtBib4M8KroPPH6SKQvd9VhcZ23PWxkVZMUEMEDMSuRJ5mXWes1lSjrvM
nn80vkwqcxrV8Ne/Q3WylxP8JPy7JscE27uM5d67aHMxcUxMNmaALr+hb1mjaLdK
ISdrwAGtnNZsxI/639+uY5YAifOndRokDw3IoHDeIvr9WM4kMzUbMo37KGhJBoYw
sF/U2K6z9qdfQiMtFUclCiSv2CnAW+BON1u1JprHCeC5qJxrieYzcga5u8gQy2RS
DLkaLUFbt6dFdyMszNJd/042pZfO2HOFRaokAmlFwjX0D+Z/8uxTQm44+SbXzWxU
DqYVkvu0HAxUhFO073F0J+ySV7RDGylFTY+3cq/+q84waemWeDlH2PBCsnGIncqs
mWE7xX1t/j1iKTC662HsgxIDbVI70OB9x2d1FUO0u/IDi+y/QmPY2CPDtqykrVgX
ZZ+6vvz1HgUsWRiP7nn13zFvoGgSp4p/SQFwe1WNELkixSexKyrdkkf4lnGKINmx
vK7ZOebpfkW9lrH2dTrXumGSYCQH5Fgjuw7Z05KnnxDjRdIWRbkwpEuVdIjcHK95
MZGufZn7QC3l8lLWXL4SpPIs6v7esmZx0CCDYz+OO1ztvtI7SAhdPVHxkxZ48Jmp
x6RcFNJV5jAiIxwvckuGv6ELo6MD8hggD3SofGjISvTBrDRHeMyQxVtpJPG2J9ME
zcgADwiXoxs2mCL+5avX8ehRVO8dIyLw5zKS/g/XYBBuribpQCcJdd/hLVij5jeZ
qFvn/e/MZyvB8V/MtjzCbbPXf9Ex2LYj6XRle/2T6O3E4vyfmQuoIr8IC/icqoyV
sJKuf938fpwJISal53CftQ5B0J/OPAraQFgyLOY7dprbvjNMg2sxlI8yXXcZxBsH
+6yWL6+Yim6FOCLo5aJMBe9NfPuPOdYwdmzxvsHu7ke0QPLdK56MX8VWAuGZ7XTA
5KUldNsmz8KX7ARSjyxtmUJgKsQlM6SBEcDEb0dyj0c3C87dG67BFmJfxGiskipg
6lxjROw5WecWQl7PzJAltegWI88bA5PwwfJVwCffw/My/TAmKXlJ9xDF1fRWNMh0
z7Ny0eJ8OpKU5wnyP5Ws5XpoNhDcavXYigVt3J4KaluBncDxPb2T3qXx/Acga3w6
9aWYJndWmfSokVaTU+UB27mc1j67Au5qni5BGZvpMDnY/gRPpkY/BRKgTbf+OteK
1SppLsYUiXo9v8tGyBX9LKIfAtOpY4mxIlBzMIA+bTDIQlATrs2Asz750XUeetxU
y1XOtBoVo3z4Yxtca+Z2gNF4PhJTZI5wAkoLVVRea9kpKF3xNQNqUBo5hrPpCzrV
JuODg4HBUnXkZRXtO3WUwYJfjA8xdUcZlwy9yee69mEslMHlP1hYjUbgutRLx0RW
TCbEbZOMVqqQOVpOAmhvH35lTpYOxwGwjknzwHD4hfu418NC4SXcvEVbtN6AcuaB
00LEpBOL4F+WkG70Gp+GistbZiKQSZF/HRE6LnmbwMXc+J7tqIoGXlFc4a120ima
1SGS99xJ6rR548Yz/GquN7yeh05BbUx3P0mW02xbcKYt4l+aQ9K1ATpaaiXadYbu
Cs2ZWctjDKPGTsVhiOy+fVGuo0wuriGF32Ti7cbs96SG3tyBF0GZqqby2+uZndm7
crJS0itJpbPS6+Lo5XH7qdYYzv/bqFuYvZ5//peSdux/lBet30pVSYDB000gADwh
AdeolUVBjAvAZLKftByMc2jiIUtDB8/UaveAC979D/SAIw+107QquDsPpI9aor2W
sAtLn+DLlEtGKvmK3T0dLLztMRLPkBd8aDKfjgRikoJaUVaAhAkWWJS2aY72fqlS
Pn8cNOPnWGwwFIL+xV3nT6BZaApNB3fn1H/LsKkrjY7r/yPjSF+AdR1XmTbL6cWq
QLJplo4l9p6YeWeuwhyU7vR9RlTq2Vpb6z6o90QvZw2sggT111ZY/TvpqugsjH3m
CiTeai83yKtUSld5fFpk7ynSdiK2YnYwMLvSKWzemwbYF9B5hBva5j1oCILQG1tY
A5/es5HQ22jOmaXLDlQmj9ONBLUjjkJP1jSHWqo31kUaXR1X9fzkE/k0fY+JhmXZ
xfn0l1Ww7RqaVxjHJQKRR1Ksu6RGYjrRhxcLsPcCPggUviUEhFIcj1dBcDJw80nm
zkSr8KruiyJHGEbhWr0yLBikT2Z8M8EdjhaFMXkkuQtDiCgT3lh3EvLGNPxWdIK5
HcYuUtQUNz8ohjZfZgu7ahlVZOcxQE/nlIQ56B0MWV9oNUsjqU+aD6dIA6fFv7Y/
evXK/mHBaogRbIb/koXfcVIF05YCWw+g4dPINL44Qy8DAvFSmcfB3xj+3abWUc+t
I1ByFJyAeBWe96G49hSxWldkbJTQeIvL8wjvTDLHG1I1m0c/dXTY1fVwm/R7f15T
w/QfEUd1fWPBoVIhEvGJZaSUHgi7b5LvZD9GVGvk1km3HaGSezhGelZeR3TC31S0
/tpIo8cBY8S4Pbfa7Wb+nMbKk7p9jbkdQAIOLewURnJJPOJ/MTQk7G6xcMBCcL93
UpfVflK2nfSwZelCaUtgZ9Y98zQJ+wR27K3USqA8X5LnODYH7SPZ6R7XfxVGE/A1
6uTcBQXYTPPkzaWsBmNJl4PVf2ddGHgON1q7NDh3RLoFd6mM4DqigSsEkJrPCScg
Pe/s/OJhwupMSZjXYKbpaHx1Sp8S4WGCnwyGnIPVTrwsaDxFP5PM0cCLnYZwHgJy
sDlPOzztwXBYjlzq/XcVkf8DEay68JWfNuBv0IJG752ireFlyd5J/Le3TSrcxAx4
LMsQPi4CzBW1DUii4LR9924AdzrXGszjXmFCVMmuL0plO9E5Cfl7PZ0PKLSEjIQO
AI86jlql582G84FQxu7spwilp1dYbE3tVccO7wfBLFXoxMEVr5onHIFfTHrNRgxU
9j24+2fqFINXUgSR2I82OMCHdp8H9RZqdfS1piqmEYmvVmeQVqsZyecdVM8qGve1
sQx7iCuHOILgh5DoeuED04b1peiHUnsP8vH90ZkAARD1QcIdzrmnAC9Q3z+dSzXj
1//s8P7GA+HUEPiCRXQa1NLUjTwA91NWe7cd8zl3+FVuGo3SeNrJCR9xawOC6HMS
rcqmq8QwrdMRkhVp/yw8aRa9bD9d3np9AzqxaGTvv+qlJgm8786OaQs6O99MFuoA
doWvvhdiLPwudYcg628a8mzHQzsiwWg2S9dyCWk90waTobUMRPrDt34Z7a6aPily
GtvLMp3yOwlqzAmatOzsEIQIqsYKrifqVliy3nNDzP6ofuGs5kkrYr8sz+HVufvG
VHYsKkolPA/jxlfEOuOaHXEJ1kRV0oFJBRaEi2HKB+OgNDJFl7xgypcGyYIjcyzt
n9JgBKSJrCwEsncgo8GxNko+FoWnWszJnXbOkLWI5K9rGCxERgjlC5df3TDQWetK
2HpWgOzAbYs3qAJr3l6gScj/T6wS1MsyNYl/K5ZHizlHKsx1nubPj0V0MXnlHljt
/Wp37XOCSKlzuLG9iTMPhZdNi99ZJBF+CA1sWWgwYh6tBCmJ+hqkbjH4HyXTVi2h
TSMNTV7B5QSn1i2VM89hDDR3onWNvla4O5EE0XFG+LdHF90lWgdMljEKiYkqGPAR
FCNnaRuGRPv94ebf4I3/a/xcETr587eZnyANAs8iR2/H+HdMPgVwYHHyLV2MxMvb
t5CK4CNBVJ3xBGd/rhtK+Qc1S9y8o0YZMq5YQ3kFb0PwJePf4EoMyVetGdNpu9vM
itMaxkcYfpzYaWMlTVSnU9GpFWfp+0QEVlordF3hnwAiXQzKgpjNtPNme4aYuyus
p/1TyaqsvuDruyMsHX+iJw1I1Ysit5qtiwFG8jN+EKNhwwIxfnQ5FsBaUDhUYUxo
jFvR/FbEcZnanpZAjQ6oJDPn5MWJnk/IOouhBHkmpKzr3qmWxv9RJ9b2l3jfjZkM
Mpnn2vlH5iXO9IlJ9B62lhH4tYXYN/vmmlHDf6bMRDuITQImQf1n7EDC6m1GvvKf
ypfdU+fTAJ2cdLlzn1GgMYeO0EqbwrDFOqTgAlT9f8+frYU0qGZO0qKiRSQaAd8N
o4PMdlBMif98JHRJDFTDVS17gVF55fH6Qa5LwGVMAhgw8xcuuI2LdS9zgDVC7+wd
p7Gm1hXhJur2QNBrDBcZqEfnCcLBxjDTFYDXvsJbzIUQP+xg2i5lS9/FkPMPwmnJ
XHdlgMw+T172KAXSrGiRn4PkokhG7rQhBKyZQ6QRG4s/H0E9+k6NOy8dsJfc8f7H
7/XqJ5DSwWatq3KfXCS6GbCAIcq0WWLINUjLaTR4ofPm7mOqPqcX/dYFxo66HGKE
a/6B7erWhjt4rykaUhuL0vAk/Uhffv2wXbdnlUZQvbM7siyUmSv/n6VtUPriUS6E
fgicETpoIP3Zf3/EPXhRtK3ObDPrO1vwDAzIQkt9s2AXyZFBfIPyEHKPP9qFzp2F
lJ1mzV7krTg213dfP6QD794Ek197t6v7YeRcsdDrcg2tBUMn0jtrYHoVQanQRkMi
N115pJuhOxC+xwvpbpZqWFMgieBpV6NouVoMDqa1VBdImVvg0GlG2J3wPR9E1nF1
LnnpltRltkAH1D6quZagYsOyw9C5/pPVeueyXpTirRb3FiZPgA3C+QXsHEAZab1B
+cLNdvCBxDtYwMPUOr7BuAZgwm5Y4W5wkXCKs5qTbDDzTve1fxCeyG3wrUaB+/i5
1S3vGtuq0VyliwU5x2GfXJGWkdAa5ZdVn/ztYRhnEdR7T+aIbi/uNJYs/s8gXLtT
YELSHO7CGQX+9x+sNqelrBGHs6hazFJN6UaN1tL0YUSKgJn5Zyp/SYCB7ogUPNKV
HzkrpT25dp7xL3JhLWrqDmdyIyWmXS/+7mT+kWQp2MNTSoY6ZwhaKuV/COYHRnAL
Enf+uAK237v1s4cQngzR9ncd7M0ypKsoCPaf2U7bIX2z9Y0RYCGfyXY8/tPiO11s
LPeajz5EYXJ+2hwsB21Ne8FEjwRele6xNl6oMSoFrC55Dk70G5U0vm9qY57euvuE
ZQ2oCAhB2p+xfmFk0d3eHUTUbHVvdJNIQNrG76qcq45RIH9x5dFGp24RtQVK/INX
+5g1ZVmvbz2smnDr0Aq27vfvfxTkPaQtSgFTxTBeO2lgFdqElmQT1yuqKbs6PCLj
YgsbYm5a/x6OqGlWSwystVlbZuh2NiAUXqyDlX4ps5ayoqEcAo1LD9sEpy5gX1WG
aZ9ixpd0NccZIKK5llXrvU3zwhUrKk9qHc1ZKf7LxRjMNSjKA0gxmoNLnRhpdsQB
5coXgCZHyZtdH05NmIZrpjKfJDMs9Po6hYGBbmKaO0lcLFrhcBvNMxc1WEZCQtht
k45JVLoAhH9OZwDrkRuw7xWanRC9TlG/5Q+uBChAzGYEy5h9j/GEbdmSJbXS27YU
F6MBuLbIGUV6RgtBqIQ2dVMif0ULfmdfhbyQPQxwX4QOkLxsKYZ1G3ImAo2TtRfw
ofFO9ePqcSuOpSHWCJ1Qsi9UIrq+jQsgnhwLrTYYSgRjpn/QgTglDe80tWW0/qXB
VDsX2GqQptVp42dvuUrYPHM57/2/TRQ/WQHb8iNWHP1xdtxRK9U9EPiM0OWneCsN
1aJ6EDVchypwFxG9Iauqlpt+eGpkPSZ+pV4QSYPTBMzwNPIsNQUS+iQar+7DRwzR
jQjQZ4O/BdSNiNXS6pEa5QIddmFJlUx3u30sgFLDbmqV9G7nZ8WGQcdB2FtFlXBx
DTw///+IzXy4xfvf5H1IN3ElfMg83dYOsGrmVvG43x1Jk3psb7+xnikEF0CeFQbt
6KuPFZyi5CCMDhb5gFt1lN8kfxroR+CVRKKgcrARANP2IVGCBSrXN0738LOtYv0+
uQxMrY608p2aRcyDFacrADnTx4HBYgTIvCyZgdbjedgiUB4tQye5/jHjfU7lnk++
8y3whkFpBhP8WnncTbJQSN4R6X7JDyIn2t6zrKDL/c1p863k/1PiPDAKqf3VDBMm
QkHoDfIxb8rtvDQpGOMhqcSQaTbPhqFUdkaUf2NGehrhVI+LxgcjSQkAVKOO6e+J
04FCf9bTiFRkqxQG9y3CL29ldY8vecyJHjrwIe7xGGqGPW+UtAwizpqUqzKmKELh
NHUIi2/d3x3uHgiidMx/Znlha32Vn2di3MgR1L4cjtBRAt/66xMv8gtQvzhrdw+U
QDubYDr5uZK5exMYfLq93m8LRJuG3pdGjLnWNZ9s4MiXzu8NhIxLlXsbeetjKWOC
bquDH5z0FLbuJueLVuiMX4kj63Xqz0BUaBabWZEuSLYgqgUrUgxismck1wemdgZm
S7J3LqQcjGAvniWFoiCENuiqNmEeGTVdOlQEkeYMzbg6tv7NjqEnB/F8jL7QkUjU
PrCBeh2VCAdT+Aen3xYxru5zdPregOer1v7oajbDs+HiXcpHJEfGjcMT065LonTA
zeyePY3qcVqKrA6iZ9xjzjr/XT6otKzOVs4QfCTdUT869C4N8ceYRKjNensR8jY5
crs7Gz1BYCgSSS+hX0fzaAJqEf58OBeyhncp5aGk1eqpaSiuQjEzUsd+saDTsDxf
M+4IFmE1Rjz8jD7B1Z30y6y7SSIf1MO20KKjN/t3milXCrflavQKsGPJH157bi2v
fWX38tziV2eCBFW0PWmLyGKxzI0B1qfXqug80mOIfRIyGcqHAilKNFOZRO5B+HBk
cerPH6Z95h++B9AtoSClHNyivCcyJoTUfdVk+Zc5x3E8dNErY9WwQFy3DuZWGY7L
5XrJ+O0YXCkiK4bRiUW9mh8CgyPISY8Pcx69CwMMxqFYjuqMsgo2SW/cKdmMBFmi
uLHJMGIvIQaq+BC+eeZfc/G+WOThKwXX+kEepfgagQ9y3MxUHVkqN0OaO9ihskUU
e/vjgsdC+O8msi1c/6UjTHWzuuVKO70H/cOe+k0fF6MlWEWuyoYV9rziC+FmZB4F
OLBAY9fdLGgJckuXQMQxe+WTpjNLBKZvro5/oP/c/vwXr0lPc09IeqUHga915Cwl
63TzIyGl2HsuoGRAgfGDbMgXmcKyppoRtKkwBPrcHGsvpizaMXI2BX+S/SAbzhFz
q1HaEztRCU9O3X4FaPOU+a/isaIGDWcbGUFgdjRtFQvrHP1M5cnktYJiG0Y2GaSE
N3Nc92fZK6U7r4s9LHymmN/R+3qfIewagrFyaZ+zZ2R0yS/OtmSLA8CuoFzAy4+J
zvpiEMpz2aFtdOFhyyIt41YVzNlx1hd//b3e4KE8XETVjSWM+cnXXrlqhv0b3lS8
TsAyXA8/OrGZCM9xYBP7EyjebEE6w02UcQ9LV3oqc1nV1gnLqgQBIgPfbYHZ32Am
AMgWpY3+LJzlrZR/eTodoZkEKm+1E7dpyIFGJ6eksKBhsvgOx5RfAfv0uFKcwfNi
zbV9MgZwOlLF9SV2PaUdgt3uWk6lV086ytYMbaV3RkFZr2thklAnczhFcu512BCo
GHpHB8hPKfsM2omXnk7gzWiDvrmx//+RVlsEd02/6Ljk1XeZoFC+QXAbWEdmpkIA
2sRFfMII8C5XXEc97jZ64/9JOijH3QFezylA1zim/cHsJDhN2LRImWX3SyrdUwgC
0gyEmgIXtOPVaGpAa3Fqxo8hi+6cNFzMMl+7Mb25JWG1idKMU0sBxBj3iwvJbVwe
TSlBFTVnNGwHTQ5iK/WZ3tHjWbey9hZxWKQsDBPsY3gQKdyKwwGD2RzFAEBNbW0z
+479I2kbHDHft81KnMP3xstEkXucas/h10+C37mQdhTibiIpKEv/DrTzVI15ziyW
ZzO2LhBEc+weWIZ8Urk6n82hq6kSXFqCwoNKDlP3p9ek86F/BI7PpGg+4bG4lYsy
kpVgO0WreSYBPsNgQsHh+odMqhalBZaBl0GzVnQON5e/SD3ygigGFvzK8lB9j5m0
8Fj39X7lYWXYL13Pkbp4lgzHa+IugEmzIbYggO3v2tnLYxkCxZ9dwB4QPQKJVg9B
jUs8/EJpo+vMzPFvvlvtJDS7rY0omoCYMU9FgGMhrNUaZTWEL4pntDXRcj5mjW+j
8E3BohKtsO6ylgn150KT6yu7YS0YUfvzQ1DmTugPNIvAzjJ/vpbXSWUvlWRzezKC
Dc0gVIYXdgaPgtVew8T2DZf7KvABgxqjnM7OTNXR7pU9JMZAbm8i2iXuBi//Nz2p
u9kshVrrBvZKfJZedYQ6B4ZFZla+7O5+LbGiUZzKjIOjp1wj1vuv8ptQDzkIzesw
ATmwGftZAF8RLkDs03JSrMuhkfWRsOaXTrxYyZ84pmGKdvyzoER3lDpaf4W4d0ed
rR/+msm0hDjHcYi7NkI2BcGRcxGpTunm+H8KS6kMEJGdCpTnLbNVSRlR2zkMK18X
DdLU8i7uqBPMmoz9aExSav3cxdvE8SPC3QR/0sr31HiIy4V9K4Hsnkw0Lw4oNsRl
CbgTdAlZJYzU4FdQA0fNNCU2BYUoNEk8bo5uoJjiJSU05J7bo4arXeO15Z0oRcCr
nGxHN/wWp/Mqo/e99UZamoOfBh8av1HN4WPYcMIbbs9ECgfAHDx3cA9Xf0O9VZ3g
e20E3gXsgP2i8SnF6cYqU+8G+UKtMB41EKkdhHywJpI6CLiDA6ZKJ86GzgMTv7AV
Ul1e1aH1kTMBYUUq4LZphF3R8IqM5UkYFFT1FvErXryd1dRmzHhnvPV9rpL4K3AJ
EUSPDqGA2eS1tYHwaKc6ar+ByhxJnrrGfwRgYGkHw9RTpM2cy6gHuZRuynHE+kx+
6RO/8CwpnJYuukxL6NinVMvLJiVVSTAVU8szBzADHP4pBXAN6vaE/87BjkRgmZQm
mW5gzjwuOx28n7WuvbURg5mKbAZy6GPPZ1ba8A0+LII=
--pragma protect end_data_block
--pragma protect digest_block
Yf7WEa58fonB/J1zyjFnwV9WTDs=
--pragma protect end_digest_block
--pragma protect end_protected
