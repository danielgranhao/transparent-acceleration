-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
HbI9V4O+4gs220UNkf3Vpj9LgbxYgA7zDC3QtzHAJW4+jkJ66RX9DKLK98wRwB33
NqNnNHNgXBogIVdLnNSyJ+wwfu0X5sPaSGgyk6q1lcAg1f+iqejsQrT3pRUCdM/m
z6yFkd40whco1WTwgI77o90qQGgB23HTEtdltLCh1ww=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6823)

`protect DATA_BLOCK
kgEhCMI3l28eTE0po4eMjOS1PJbGKnJKUDoNDVdA8ntnlaBQXoFaGmKlvyMqq7G1
Wj32fwYiDGttzkimTcxTpg0aMyC84jUvAEIQ634BnElit/xtZWqJ4Iz5yBUzveAk
t7mMqKibk5wFFGh7H4ZwAyH6fgmOyM5Ee9Lzvx4Ng5blCPEgJIQpRkiM7ZYU69DN
bzM+poZd8Aaiv7w/M+0Q9Bxesjwuj/KvqNTMgAuq+MkA3NPWxOvuSbE83+bYmu8t
HZG8eCaq9v+GkIuE1TBBAVK933JZXynyKBKz3WcJLck67vuI0BHibc703jQM/q0k
d7BHiB6V3jt1eDpXZxuBHzd5XwHeQUsyDol7AyqMASIyh6s+BIWpngKgyYBsT69b
WeWAP40X4CC90hKAkCa58Vq7XdWxYO0lK0m083upKof7NigV6n/t2B1pr5c5HvUA
w4crATnoVbwuTJYxCKxFV1Ysbw/DVOMAUizt7G5Oyaeke7IhB9LyJMuNQxxwewg7
dhXpBQxue9THhiFUssqjSe9v9BWdAaMcuN/cTirJRjSE8Jxyq8p75NTBHHAdVcx3
gkTseAOuRlrULASqDt3hxLx6FipXY29mpquikJvv+X1M0m3zSeiT9qzxE8zJlBga
PejBM6C567DUoaXrIx/SbBrZmT4qCsYrVhNgpgPaUZgFp2i1mwjZLEANM0A5gGo3
qh92eYLrQEXMk9CMvy64myGX5/pplzlssSnFg5P1jWViDWEw+LgIbW6dC6AVEKhb
n6KXx+HA9et3XSQOKB9fnNeRWjxr29zpuQu+BBGyb3xyK+HBTqXUNS0bgLS8Z59N
rC6tM5ltl9SL4sohx+VqkH8eNbQZdNcM3MVHFmi0+nhRhxzZW2XQnGRorv/kcTz6
/zcm1qpGqcWiaRwen9Ry5J2sBooAZycTOGN3qtETdYUwsn5uaeWuOgblwcE8eqhI
C9TXvni0rAeLNmKqADaCrO3m5DiFrvfCnq7TvKs3cZRLl4mVbGx8ZrE0/Lu/1r4K
CwbvHtdTGuD7X2Gof9A9wGj7ECXAFU4lQb/Mj0K+GZ0ffcY2H7wE1iPiMKwxJQBF
ZlNCSsypXSDA1kMIUhofZsp0gzqNMsIx6Vwyzm5dIOMqYsUHlOpPIFc1F6sU09v2
LyyHTliXM0qi1DrM9RpvDYbCICadkIlZ1dpJFl/tP559H4GlxF52OP7SPDb7v+8b
/B6y4Fdo+GfOdYl79Awr4R9KGGnYzFbFgYiDy3hWSkmY+XZDJ8/3g0W80IOgnOEv
zTsFVRtDy8jE45kTuM+nUN/waCdqxsDQrUI99jp1rG0bP/Uq4uKb8tk492Vk6VZR
SRAxOiuLDPbrkR6DtJ+GANNp6G0OlcFqbQII+P752pdcvcIZHp8dgdfZU/hyzUER
krXqaSCBwQ9Dt655FUwTBS+Tyj+qh6an8uozMKipTLTAhXIs+Ze8C958AZ+KxQo6
jaCOQPtmXCa05N5Eb4TmYIjJrQ5j2BSh8A3RxaQuTkn+1H4oDLQtsfLWTAvsFA1R
Vme6D7M82zjMXNrukrioRFtVa/aRtdwxxDzhXFWTvhEStJ3ED6LwD9n2LpVsoVL3
pv+ZicbwySv7OJ7t/o5XnV4nHb78m2C9oeLS2c9VL5tpFlBGKtvS1CcdNDANBfji
ePBuvlR4Czpg4ymooV3CoZOePrzNGsBqqsfx4Euj0MPuOOzRMbSOgK0rsJFB69Lw
cmXqM8Zs9bsKAJV5AFIoXgEP++VTQU9hpIjuMHqrstCIG1dHzxnbxeFUrRl2xyjj
r/HjabP6k31UqIUXRR98RoC4yg6m8e/qTMBBzBWLLAedcXjmEZgmj1QIoTc9wvkv
ZLYQK31nFOotPVP0xjvihhERYD+Fux0WMLb4ndxH53HXhBS6wpo19FYam69tS7UD
v4DrDKxQ2/wFm1yKT5rqLTTtj9Ktk9RFABj8EmU1YGv/UeKHJSx9Z9Qa41G3hqSG
1afzuQgDFLSVjEZn9VjuuUSCbA5ft8xQ0HaUZYXMGDFrxuVey/isxuKN3/iiYOgf
hKBFUrtKQllJOHLQXrfsKuoOE0ETHUw4hclkjnm/C+008+UZxJrI53k0izhauXw7
EDI8orqYAX4LaicjDHXx5UOOL/mRdTKVHVtwtDIaySTIX/IbHqy/UBqIYDsyDcmO
oMsV1QZSUY2KvJ85HfJkrnJL3lbGRvjZxp+zHBQaung9H6BuMj6M4SVhPwBL/Vph
RNV8IFpgOtjM+9ezc42YmbTZfEZT+GcIxfvML9twbRJN+JP1SW0s5nd23jrJyjmc
i67lxHzLYq26KBAxpXuuxZiyhj/Bt9ryGllJW6to8NT4K8IIUlUCo/WQOZYrQ46x
471XjbTKwtpki37Ft+IYMB7vejj2Sm445W4S+97CGUK1TWBB8zO1CI99yliv4lbQ
YzxkHk52OsNXvc5aSsf8fY9tVGNjfgGJvap7ZgKvnQHivNeL45k2Y17V05tmqzJS
v2SaDzHkfktHg5bQ6VvoOhFLb91PBy3TXWDmIMJHZooVQmtpeNJw/l3xOoLgLIlp
B0oWjKk/J9A6WIB0xgUI/cHzV9jzdwYGAUyVBIYEOq+DCDL0Zx5qRBlkusuP0usU
LBFZtA+0cJvAMSl46ookt7I65X23G6h4XhVRny22UNOp0DIhH0qAEXj5nI6CxUNS
8VCEP0uPy3zzyMBhLgukbjDbkAMtXYqRwwR8vg0VgE5ZYdS2RV8LOTos8l7MXGNf
fpvcpF3/KEN3MvYuCXrj7uzTkb5a7hIo6TwwIwBttR2CuVdZCJqrEeVR5ChBRZIb
tAPPvIE2CtHquW5W1t4Q0TFNiTAmpTVRQB03QOa+2jdpS+Oh1xnJ1Sxd6pwWqj4L
Gh6ik5rqir4dxSAAq+em2PIb7ZeAWN128CWmvcoX6BWF4BTrb4GKLuHraxyIS0gz
C5JXHkFxbPdtpTT18RUhAWaFupOQi7BlsAooaX4L80VLQ9FRHoT0qcEBb6Bqh0x/
nE/q8bdlrnxTBJXhtyQOmxj+jDAUWp/VCq+LOI1PhHDD72/lU75GOHuwY2UryrXV
8wVh5C6wPsiZhVEbPwl+JO1AF4zT/C2VQxCAezj+u6kt2wksyKLErPMSbHoz7kWI
/CyL5/ynbhkb4AEMFgNWRUZHNR+PwNKhpj5ZzdmfGXT8iJeqPZyAWQd9m0HTzImz
ero9J5Qrw3tcW0FCOfCRQv5rVsEXcLzhHRiYGRcO1eu3DCpO06yeWx0dYQptrlpF
tYou0Ull9qsWFwDHE+CIuY8ZaXWyuDbploA+AfeTvOCFDApsv+qTOTcEmatuqN6q
EyBMvUlCXFeQAGDKnz8eNciPEQrUexzbOf/qea38KuSLIkZYYJggzOeWJ/xi0HjI
/Z2aoL59HNHK+X8sGrqpvUqF6C8argR1/Jfb2AfDHskKvDX/EwponZyCecr3YfJh
39QzoWQIxPAjw4c3nnSqpIJA2Fed+mUxqOSaI0Xbad0DYHcHcoYhtQfRiW5ovD4J
UBp9erVWleJ4wSqKiVl46UzZIP4f4dY7FFReZhh8z8l3FIl5HtysbBRbqUwE2Kj2
4Lido/WWjcNomUnw1qt+9mSl+bEclpwUFlt6Z18zm13bYrevRiWevDmjGA0s8h9q
5bwAkq5o6s2Tyw4SbaamJmX9+K43zd9/9vcMoT9juthXbGxPe+H/hZiWnpwzIeyM
MZsCyNCthJiDIz760WNksK1Us9aUe8s05z6HiHfM1YWYzLpOSM+NPjoyo/W5hkdy
S9pPIpGBc9P2+bzkA8IyPrn9mJ0Mt1TJeNIEh8V5Jx9zKjk329/86Pnydmi0Vxmg
NV42gFrHFqQR30/f41AGsT5IrSqjHSdZfKBoqUPcv1Rb+YSts1m/8DAy15+cNVaz
ceJ0AWPnutjLpUPlDtJpuHrXqWAZpkVDFILtwMIWuPyldmMTlXUbh5xX4hkWhmE8
5jC5nPOt45zI3TVfJ1lU38PwCirv7vc87CjF3TSotwvOXK2nKHT9oEws47iziMjD
Ln8UognIawbwAo4kU2QqMkMAUpgld09tYik5AqYPHNqQfvWJD/2PLMEa3o1ghEQe
Z3FHAZAfVoYlhiZ0Ql8AK0e8PFzhBVUoXVIyUCxymh/eAUzT7rdou2E8prOr7vr0
7cgGL+U+E1sywg/QufxfYFMgQPHdmSTco6/WpCiAD35krpK14JlQ7d9Sm/kDIBZZ
VBpqveQi3/SVz7iHOebNI4D2Z+Lpbhhen9AHWlFVp2+xQe0Fu1CFMV6SHdPto13Z
XNrzL2/LAvYnPlBTFHufKBzrlbSYPBL2COv5DNOHqob4nk0bSEmQfQNdAgGDQWvl
9Rx3vgeCFOEltE/qbhbmMXfypeyYYwOYK1YOL/pBFfR719PkQLABhJgvZiEQzelL
77ZonsgmfRZHSReF7kwxdCtb5rVsLZ1gxc6rvN8p8KpAPEdTC/wrTilJNZhgjT3Y
Z5UNRgMPtD3m8BiX5q1hEZNJFafYrMipz52KwD/Fg+yGEVvzPN3HXED1QM0jOuQ3
WaQpegZkAZdXDi+aTFaqtgrxdrSbo6c6JWm6rI+fyAjOJPzAmXwEaSBp82iRll68
palH4ilL2raYZSwHpGQarz3vnh5N+YKcHo+vUo9k7XoO5WQWoA8S4/x448EJYq6f
gKG7yljGmwpL8ShUJo/c6Ezih1jymXlelgL2GoI3b0LkpJ0vu5FUpTPzHHzV28st
t3ANcNR56dfuj2CYqGGYh0Ek39Ladr+Hwj8gDRCtTLiEjCPBYkHYfEzBs9wDsrsT
BIIgtToCB3bH0ktNxUikTiVTdWqeYlNqRDKj+p747CDCTQ8xKbkcrfEmwmTcqTOK
8K7t7CTPa6qWzMMF9y7Hw7FHJtSuUMv1+TW5A+DKRoYxWbgDOKI3whaK+RSkabHY
a+ixl9/1qrh9YJ9xypbpubjpBKhfROfUq+fg2wghLkPmHmK8vIS5BYNPYTC4PRtu
Dn8b9fj4wB+xEfb/uMwYRjkafOeuIH00ldEDDQk2V7KNtg3HN3x6vd125cxfYnzq
BVGSQnPLY2jw27plRxQy5TZNjxgRoejet0MMUPe0nY+7XeQL5pd8c6T/DKLBLt+5
keYq8vvn9CIB9seBKb+FUWfH88OXZzNb3x5XMxrHBdYM6GggOOBmRT2ptp7TdUTU
7+kqOm1NyLHelyJqzKpuEECE+0dRQ/INzWJKo8f9LqEbZ4mpJYj7Sf8c15e4qMab
FNkHfKvOx9MWs/LTxwuGRhun54+mTHkPspRU5myRKZxBmnA3V4DKKc5nrhpnat0e
OTKyS0ICV7XEq+7RrBbanYOe4SzqV5NDIGX1GVF+7N+QQuCAqWRYoyv7Jp17v+v6
1iX9Yq9L+W3pRERZTijUWfbfMbTaMQ5riuXSXNnrXPoAB5l6a9rK1YoOgEbce2Wx
AeYFpOSTY4160Dzcj2FZAvlPghthHrSm3A/j0OevvZfXOoT7aDlmtGEUIpu18QDT
6J870xtW9zEEe81AapwkIvJDY+Wy02bCRefa1f66hvgW2SgGlttMZRl9FgGjFlTj
Ouu3B7ZcboVLKbvolomQdBfupXBqbaToNeOTq0lOd/91x77k4K4IUexhNC7J4kqM
iWDGKJEaPyOtiCFxPCEJ0jWxlu39D1VEVegknWSE92dGOc0mZd86OIJotlj+r25/
edTffkRZ1ruoYo19O0aKwoURDpOo6B58/TTcE5gcR9EfBa8vW3SI2qIqCY3HB8zl
lEx5VXRlrIXMJyDwKTGfTduzRaBIQFfTHWYYFzOuVH4nec3ADNw0lofov9ffwCIg
mNciBAIlGHCjqI3zY7zgFs2zT8NVXtxjLIg78R6vRaOtCmLpTZTxEJEZPloTZhBM
FXmfWEpv5dpDu3AWQ2mi6aArvePUg2B/gWMq4lrkK2ZqBBNye7XkWi/c4rGKDqju
reK7kQg8kJ9224XVXATM6Hr0AC0IfRm8HM3DXu+uVjrSNrA0jOVVYJiGoBb1EKxf
xHq7Iceh0C/Xubiv2BYcX409NfidwDTCN5oCzn2a4bacdcSt3FbrlZ5T+G1WyKvz
IsMb5/XLn826G4jBvqNIfn72jSi+4ZJtrIeLBmq/AAZ5B83tLzWz/KHZYInaPmES
uFPb37sLETJCZt2NElHSH0TIZJntS/1PJozB3CFv4Lax+GMxv/uJ4OUMsZOzGlkp
GbJ8SjtUyqGgdIg7e0+KtaEJprYKAVwAb/ap6W6820wdjtg4MdXMahjAt8TAlH4V
hAegd4ovwX9Xg3K/VnAxP8DPkqsMjJ/HY7pnRgWcwlbhA1BjsOXaKM+YpZtH09Vl
Tz7JDZjqxtbJkW70PnZNopNhQMHNqO910ER8gv/0Hfs3B9vdWS59fgAZ1csrx6vq
s+bUeyAP2RqkgIAkuxEm4w83DdnE9S0hTNnxRX0jHVe72Xw2S+F4jIQfUw4GEVhO
QOJRKahNuraPd+vgtnAN1uDoOabFmuYo6xAFlzKXqiyMjBqmNZaYiD0vyfxlz/77
gGPC18Jj1huyfoIkXATsOwXZu4HFiU/484lBFH63foJmZ2GVxoWo2gTdUXHyQPK1
amAew3mWeBFNWh5gBP4NfcjnrwPqM0UW0IBY1Cuh57axJ9J+jghvb3f+jVtl0CZs
QzkQLNbMOwnP7y6/RMu0fFCoM/bjTtYt/UMQZMTHPrDHdPJiiPlg3XlNKD2cj3h7
17DP04yrDVvkSdi3swzWsoZztJnyalfrOSm5dvR06FTn0sleGWSfkNLTpImPKOVJ
YnjoTFCB1hVKTx6oArEYUMJS3k9ErFCtoiXXXkaJT6VWaVYO3AHAmeypspqUveC/
HqhPhfrLEx8MFDs13rQd1IUOi23FrFBDsp+42dlJUZwyzRh7yFON3QwNVt63Pfzc
lExW2qEnPzx59ZSbK+alxjfwsIZdZ7eexDK6kHQFc25zcvCHkb7IukYJ6h8zndf8
dQsgz/S3Sj3U32HIN0KuUn5NQOQtgHWZ+N4BuwNzTYQzEPLtccxwA9cMDKUDfGpt
sQvb4QZQtQxEH/u2LJAlQGXAdRED0Plp2I34Tagob9E5PQZ8Qb81SOFaBXAjFTKz
Yj2Nt+IxTLx77jBExZfnbRvZ08xH19UnoUbFcx0TzXc8ZeM0KZS6j1IEPge+sf8A
4XcYOv61gBUNi5iYLr4uGYR57qjBLDX7+lekAxkNhAdZvcZvYu7n7zkX9oqwJtG2
CigILP/TRt4lbk+Fo/Lwr3ahlofntOJ0AHmuH5XTMEutLfhWc31xrPjkBQHwEicR
EGWfOwHJ17XCgflynjfC90BJRpqQN7TBj/XFMuefZ7WtlHmKPiUMhyN0VnIsuGca
GihBs0Y65T+svZ+hjLMMgI8qaeMnYKOFXtmzVxGb7nYpeEIY36noQtK3zwTTnonv
cHZ+LixGo0XhQptu3LsQaUxmu67gNWs+jQT64u9emMrp72QTmWvbNvjSxs9c1Pls
ixBv2fjs0/ozPEjuA8sr046f//Uy68AuHt3qqF58z0ClqXs8JZpWX1voWT7hGCMS
4atET2cxHeR2R08DpK6SzHMPsPBrh0Q+J4/xqNO60tSUJxaXQWieENVF4UFhcenH
ZkynUZ9B1JZQfMAdKzUp5mqAQQTTYvoSuUkiTC0gkOiih6sZP8tNFPsUxGF1KMm0
VFu9Mr96tQB2TzbeRCPGEH12YlX8RBCQLl1kHKCUWwkSXI0NGPLWvNVDxNp6EdqO
Pq0nDBdzkriMq8Qhfkd2K6SLulefeBKpk6dc9rMx7pZnXmpS3m+8juyLVztT11qp
fUYsTmcBQtT40Hp3LvKJxVU75TYSc5PqcLiZfqDU0dC1YuWTEBD65z30YxLVfYPM
s1se/OXBtVB0rKMxw9F40he68KozhlWuspmI4wi/kel+mpkMhhT2dSmGH9uuk08e
tO39rpwzWwdem+yW3Jlbek6cGalpAT5cZYshjcAkyN3bI586n9kh52g+ig/iJe0A
fMQBIYzjhkqYCzeBPeb11s7sbuCUtr/Fm712fPqYWaDyI/f0zeGV770QdPSqEmtA
5r0NzGg03n6v8hKREhmHQ9OYc81Eg45+Hu0YdOzxoKeGoxPR17Y7gERxFDvXu6qH
PNNdFTBFkp86yPUrjLW0YiMlCHxQyf9iURuGI+muYJYGZy5xw3wMgR1cQvQHl9dQ
KfskJH8qw2jlAUId5i2YGVKR6kmOWaA1XLxZqT6++nTAy67l+2waxMQ3ggC9pZBf
m5XoDBamaAjydcwXEdPaEP+HCA7Ikumvp3VVnOI+cXCCHG1rJ7RbL+aMR9rgUKOE
iZnKfg+23tAuklPNeu81JZjYgY8+iHZPOI0mqvK/60+aDb57kctYljfHInUW+Naa
8plWYgRTNbgRS/OoGpIoV3Vkq6OkK7pS4XejZOAWt4ouTRSNurSpqn34ESx2l2h0
wZkkD/xJYsVZb5u4VfgRhEeKkkWGbjccA9RFW0jbdSK8eSUSw9/p2J+57W2iRgF2
sOV+o+MF/a4QlZfiguRQfYytvrH0iE6N5Wnntp0zlcpLVK9kFDkdCRAr2PIpDmrX
sQ/VL6GJTADvk3jzvX5VglM09QkZXUFWifQWZd5A0IPFdar4vweqSZM9QbYSzEpy
a68XFnbYulLyrwXz16UTHrtFuGdhM17S2ykHkPysDiKGJ0tMKunBKPGk+B3HOxXM
uczBSgdo86ROVe/QNTlEohsBI73LPwin6sGfkZ95tSSKY2dNyLmkaKWABvX5ENFO
iXy2zhDIYYKMQ4crfKCiOdG4AxWcaNeJRCkyudEekoARuzl0cagYx3J0U+w+D/+d
wD9iiMmWyakpxDAytLpVIoJhvtT4KCXM6AxyArLMSoWOBOmJ3V8Ph6cQnTQ59NJ/
CocVFMiVy/OklR4kRORKIDbSHaVG+Tu/nd/49B+0CmbYmhclFJ3vpkh9kx2T7sfk
wq23mCYAR5H/UmyOiJ94WExgWfkqNXfSurh6ohfgaXn9rTo6e8knW6CI7Yme+I94
lIv4JVxKYfpHDdYTvd6OrwXEX/HC0rGtz3zXsGAbs2la0t5H3ywfMX1AffXAr/2A
d0s48EHAg0h1lJeB2gf5FF1NJFiPy6dBtn2Bcsi5zGU=
`protect END_PROTECTED