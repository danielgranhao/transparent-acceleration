-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ntMwkE67LMiEkkyfmHwdBQcl1cJevE8ZfncmqxykwIhHeLqaDbDBv6i3J8aiuyER
n2z4KgwJFn9ynFTslpJ2juxNyrZxL5T/qOddS804BXaTBb7ntVzNgsOkK2MwuQ6N
aZlPpMOuFHmWHIfRtjjnCXWC1WorYSrAqt2OvcPkpx0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 42948)

`protect DATA_BLOCK
BZKi3oyIgk5opobSBi702PUmV4of5Rb+/YqyEl/c6ZvTuv2UeFbxrMAWsCCJ8Aun
TasV7KTSzypZLoU7hDxB4joj9+JwrEtAOdzkfqz9BTdwA+y5cN9gHlEEt64oELKd
nFc2SQN80CO4coGtH5l32BfR+JIDMq1f08u/Frza40c/+00iDM3A+jsaZmBNsuT/
281gBmrNrLE0pY2ycxWKKvHH0/IzD4t/74eN8A7m24axTv31dVXRbDHo9Xy+4MnA
0OWIAIo2VR9AbeQEZeOL418PXcq3bYDeBpXu6KZRMV6dbxfcioj13nHloUDSYc6K
TcMmjUy56BRwW9jpqBFBIqZ+elvHhNBKP/T5npUr72Rez3JrlbyhDXHiVP/U5vLg
e7xRXnWG8pUe+JSwwMkSA6ZbhB+Dx4j8hOH5xqZvc8XwEs7ERhw/arTb0efxTeJ+
l/9Z6J0QlNSn2z4P66rKqMSQ2+RhkaFUcfU2muMEJepWpB5FWkzUNM82utyIfTsX
dFz6p8BSPUDsJVzKtYzDlZjRGshXCJj1O+E5rL/fsuvzaR/s8B7qzwdnTtuznuBc
SliyOXHznD00kHBNdKV8DFWA2TdhyPS3cyRFMxUdXoDyROs3qCL6VtPjjuYkn2OK
zUS5FhKfiquoG7CfePJqy4mrUxqfNDhsWFoOFuuKdpGeOLRXQSV5lQnGnmNbVjmt
RJbQEcZNLDGonLuW3jXDs2PNa861nYoacUuDQkAjjWzZrAiCNAoVpAfJhibjJuIJ
A7rP0UJjJNTS+hsC0jgT8ejXVwjrmJ2pTa2CwUuEH5iBCVUxX2Ez8Zn25XfZCCJt
uE75tTG1kA06YDCDqTr0AtYbM54Hc05YCczew2Wp9QSygobIT6wiuP3Qhj/krsIN
kOX002Jg7Lz4xotyeV+oBKYCFGvJE9U6W8a4/VVAmgxbb6qVCFzS2wF9P0ldFSzD
z3qeSaNnkMPHzCJa5n/jDKkU7sMdJFCrQFq1tOd9OmLBV8PRHFFCyRcT9jql4Lwo
67fEdvfV0pFQudemCYcEnMukZFolViVhJnJ8RgaPWmiT4yqWwwqedqajm+FVWnGO
QY0yb5lAdhpKvfBNBfN+p82AKDZ+xAJvhQibgjVvYugXEbvlf1TH1S3GsbtF2Xb2
0M2JbTvdRJY71eExJZjdYz7isV8HUg7sZFAp3JNfBFaJ3SXw44aTWa7S4phKpLTr
N6dsH2Ux48qxOJO8du8k9TUJPJgUtgZ85IF/JjGG5RxZNPeUcS0R8y66ymXiKydx
vtSsmqFITPDIOSvWsctCMGg6foHOpY2oCDZcs54mQ42YgUkHpMQGrY3ydNhi2Kqu
Ew/MmfvYCHV0McvMY6qPpzo+b7+/ho0GAS6hs6BCZ7v+r/AxtCo6TkF8hBgdYGYB
J6FUbCxbQmRzlQ9vb0d9WFxmW/6rL4vCqtkBCSUbAZHCg37n6beZlWkfxdrBrFU/
481j8k8S/pf6ptUk8CE2ldCjw9nbyWF5Ynz6zNzKXcCvEktjgbOxOtWhIXuWSmEp
0g/JU90nzjKi7ilhtmsBc+I/CjpRz37tt+1PJxhguzP3OBtZmrX3GgqZnTOmSmVS
hgBK99xbduqGwuSOsirTiw0ESE57XnH/MqnHwPRBTI+pulBNP1xfvVdtEvz8BgbK
0xv7sPW3wX6bPQIbCIfJlmIO/huiBKPEoOoDj8YmhUfj3IMJzzYjCQJ04Uo/oVk1
fSaAIrWnL/x2wopLYa4BZh+yt8rofp1D54Zhi9V21ay9iJfDcIFB53zja6Omq1CO
YbgL603k0F1hpT+CX11c5aTkswpZD20R5qrwym21WcglQdcDeVPULwhihmCGCbRe
6H1p+nvhVvuSz6E9R0LwS+umhvp7/3xHvePc7DIEmbCqHMPdVbIMVfgBvhanSfpX
8Z6a3p6F1yKqtlmr4zmmmyFr/3c8Hz3Hp5fzAFn4uOKCHLyoAxr2PgaV+BKQPMgD
l0i2QqFE92wuj62+P4aDvQP4PKSgg7lDvwjfmt8RJ78uy5ysLDjj+/56/SoMhge+
2o7QwB+WimVHvrWT0PGtg3/pTPEiqI7h0ydfZCiwaUTrSUeZ5G+n/sV9QHJ0CWGd
BnWnWuwG10tThMfxc3yYjK3p5D4PDAdXH/FYugfLmaA0cUZtP/oigit1qfruy+yC
wtGIAaj0+mXQIcHfKa3DIy+Meiu2parf/vTpUMsX4uGFy6Da5Fy0ZPNMMR5/LVDR
dlGZnskkRNbIZX2dmyTpjwYcOkOOTzwopA6+78+EjPgTbc3VqZhU9zR3r0r8yPio
26Bs0TRoNszIhwE6Tq1Cq/FbM1TT4vFRdnq6U/NKUNsOAor4d9eRxIupLzYgmRkw
DIC66cWctCwu7liFmX/nPebIyN0xb0T3+HruxZiNQYiMVRLl8t4iJ9iDuBEKnBgr
nvWlbCBw5B/5fzsVBMqWA1kFlSTWxgOBh09z/tWMj8ni2JC6kQ1+J+PdyqFgpZre
dpK5RwUrkQ/BI97vZENRTzC9rfkWEmdnbBfrDQ+Frgzt7kXdYDTrzgN3YDbaSGve
+N55hJi5BeOroG+ZLj+jYVA01NNSrg9kNThdGLeZncJXURJg/7j6JkXQE+FwIIC3
lZ4XNS/0ZgKE5k7hzvFN/K2WXqJGuhMgUbcP0UG+CAQMsRqEd6yw8vkCF9XFYUYZ
oT6Zjv7B7pVxG/xwrskn4AZ2Ywh8r2LKMvtnGzvAI/F1KEJz1HWwgJJZm6x0Y8xt
TpyzIM5kxLvhmLquDwV3Nh7x2UpJJsIUFl0+Xl+paUwLTORmSyWX5+oOKroEIHWO
eDBO4+QsvyxzT3jQciMlQtKgd6CW7gwzlLnpoqRrLxCDqCcBvqGBBmgsAu1fCrV7
hAl5vblQDd7K3narlcvHSLMZmjkrQPF+x3x79vBgRM3bHuLYoIgtd9lRuvfuXNtu
PQEqIcoUSt0yWLCb8AZP92jB7F0tD6ry8gEV1+OwwP4IS3iM/rfMynRc0m35SgV0
NSJWdZcW58QmwnpAM6ZlwMwZQPjlTxPExp8RgBZFCuM4ATFNdyX57DI4WGbQqUOY
hRKuFPKxuJusC0SrtZyPtrgCkK/VNd1C3EeG50K1sUjlfWvmK/wwd/yZOF8u96t9
QhT1KNof74fRIi9C+igbaV7I2fmOmfEanhFtdaj3B5WL9+sfwUDvLm5ePQHV8wlB
N8T0E6b6m4E8tM8/1AkXpbaW45THKyBi9LgsqRGNoBA7uWQMj/eHfA6bHbPp2tEf
G3Pwz2Ec6+Gg4Pdd6VoQaD2zEeU5yCYNl/B2CDybPJU3+eGbRfMBuginJiIKMA54
9XDa9aApVxCCYgIiOURGQsv+iiJTHcmknNAaLOylt+XBjX9+bQQJxaNpPS4TjVzT
AAmfUyBtiGJnfPq/M3lLgf8RqbwbbsbEFI/EUvSjoebcTo8cPac7zK/kHDTC2SAx
xxxDq7xp6w3MdzEM2CcMye56n2LQvnSmRxB6mFiWAoAhnZMUKC/emcDC7mGxu8LK
w5js4KRR7mXvZFDzbut+SJ2SSqZRhBmBL4qQsQDK/s8ucqmhSiYRdhSLMpR/UYMV
OWvFHju9FtDowBYbXKKNnMGtN9eef1sty3FSyjBn0pNtAeJ3iMKzIGsGtXEyjqXt
4Suw+Tx3fA02BwGIArrq0ZsLeiVnPm6BCe20nPnX1NWAvOJpoW9elcTyA+IZBkIc
i3vk13fH8X/FegGbtXpfd80ww1fRGLt58rqdkg7qPFus5rhceSH1C5yqHYPonlhb
Nl9L7SwG443Q5I2w57IEvwzO6wLdSInYjvJ6dufsaX8ySS15ecquoxvI9853Nmwp
0AxS+pjYsvC9mfEj0h29ZKC/WWDGVf0gLgmvG3Hu4G2/ayu65gFCBG5DeprpvsX/
+vEzf1IMbbbmvZ+QAoZ9qNR6q01viX8srI1EmGldhomcq5+8R7fAL+KX6sRx4LZU
GZk7FmsZnyi9B0a+HBwIFx7FHAj/fMWP2qf0z5W2YrZBE27rhWHk4xPzKdk9ra4t
wue0XNKfatTQlhNGEwsIIR5aemwmJ/cvbARWgyRdgNsahOZxmDIlSq17aVwp0Z8D
ueF+0K0jKVSHDY6rzvRlMIDWcJg6/1gzT7We0nOj+Lt3HEGvM0dfIQOXPaw+MJ7f
48inMZVoFTyZMden29qTiAUaBIp0Q3oM2H+XDtSuhfPpDgo1nfY+OtczEzCUKxB4
VjIVNoBsDTHzjdfs9mgWdYn6X77uNpkPfOkRFojpcYgZWy7q11BIdRN+YJOAsZgy
AYlhcQiToNEBGRSB2P0VwfHTS8y+6TisKrV6DAzsJi6PTyXWRLC+xA5QvgOxHsKG
OaNrnM88V8ww+ZQ1LYlLjMrEU7Zrw9inZj6TdxKXjyc78QqxYh3p3BR4J2JY5f29
2KJACLBQ84UV3XhZPuqwU+Z86k9q0nPTKJd07578J+aEf8voEXSldnKLutkb83sa
9AuTN65aYtECS1V+x0wS04NCyuZ7gdRB7hqgaRwqib5u2soRAlG+WJzN7N1Rspiy
X98BpbO4whQyoIXLoXpkpo3qTJL0ABUT6mRaFlajEnBVpdgXnaQcpml2DpBL2KIa
hD8xU1JGnY+BGykNRpMn0GEDiVf1gWREHeqR1adhCyGuv71cZJEWRspF/OIbkoG/
1dmYBJLSMGPeQzH22ADv/1L+FkWuWQZaViV9ayZrexIQZP3I9q5FQDNa/FqyaXJh
3vWDx6LPR4hNNZGHkuCUpJcq9oUx3nLDkyFDb84i3pODHsohVkdgkpUgB5Jg/K7u
eI26/Xrh2WskR0wOqWZ4mAAp5E/gOzSeyz9W3HoGLhrsKAGFM4mcMWafi/sHlhBt
UsbFlT0MJDPxqdA30nFV8NoJ0GPv72KrXlB58i1rQ/wIwH9cB5WvEivlr/Ovwan3
N/kConCwnDVmEKQrnUx585O0aNRfDmp6V+nWbzqY3GnvEEqnOtyuMSEPy96UFwOK
9X72ieDVUSqS3+iKgOgPjrgEuU2V5ds6UgiInnROlKsz3XFv9Zo8JHjdv3Czlc43
x3LlfEA652KlTbBzEj/A0zGjRPnxhhZc8QBLW09PhwN20Nz+5VuuZzimrxHkgJgn
E5hTfBACCLPLqHg9NlQYvIyCV5DKXmI/qQUVyQN+gD/aeAOTdd1u/MRCFYa9ksVd
vWqb83LX5qJbFFeg3j4lW/vweZNeAG2XfpeGCCJoJEZLdFsHKGOJNM6XpTqxoJAH
6MV0iIes1QeLjNp5xY933DhEOf2dbcC6AsXZ6rNbZu1Vy3xklFCIZ72GpiZDxQEl
b8izGhdExWEd8AL2gSDMW3DoxQN0n5guPuJ1fhAOurbkKud3Ey9lZDDP4O7Mgb0o
Rdkpp7FHeEUTpQoN485gSW/BeS+oG5GyssNEH2gsNYyWMUVsKaIE2CmLNQ3XeTZW
huQ0TJZtEM3i7YLZbxi5cj95E4vxB1Az7WrtxtvzjQ36D4mhmMin8eqvX5PBSClt
RagoEBBDvGSAbEvj/efBTLAf7d54r2df/uXCOKJNYOVC64WivoOffF3dSQhT/4xS
5OoiQkQPdn7GU+7Rz4ch+/y8vQpF1RexFwTja1xz8//GOn5TxfPmAXWQmnMPpgHV
5GSojR1Ny7Xw6Ub2gSR4IRQir9VA31tCFxmW0pCo7JR0vEk5UUJeyacvXomLoQhW
cm6KwUAHNhIqb3LGQdXMe103b9XjP034WkpdplLxtWuTDexnorOromhrnKcMNbin
v5eYpgK9aDTFH3hc85VU7TOuypWqds3IkHX4/7smqhIAK2oScOOIJAMA1MWsv+R2
pa0R/8rL19QKyKBCCUhhMYv156HNHNDZS1FoT/Ips0GgjsHBBmrxpUYI7MCJlT1n
fhJGeuBdAic6fRyFgPyfBTh0+tx1J31pHwFYo1iAx6b5hE0YHNsY7ZAMfEgTgW8d
9jsD1UQ928dIOgTwH7WGkQa8+vUcf/OwJvN7Wxy2UaDg6p/UdEOwyhRJOsHUuKcO
OsvGpL8udubkdb2W+IhM5xzMWBtY2eIXK3PEjGZSkfpnOpa3zOgpSt6+4ZdYrbj4
AOUMh6kl2YXzP2mB1yahMnB+EpI0JpvCerMbRytExW2Ar7FlMoCvOdFqmUBsSwYj
/JlEss9Bz755jW0UsQg85Wsuq5gfsVKP8RYiQuEIS5Dv6O5pyFHZrZmXKZMT+Qye
X7+syi1VOmMjFpWQbVyBPpKdCkcniLqo0QWL55pzG0xf9GtVtOlTUEfNGgRNE9E0
9KYZqBdqiDhVJsEMF5c4LIFuID+IjPJex9/ho0RgV05E4tMOdvelhd3VCxNBHXMB
Dq5ebvmAapwg0AQ0+xvy98PduaPq9WTMEwfqRZvBIdfv+n9IDsWpPxGfG0ZxRoL+
K2UXZt58iG7tpMyMXGGcPksxrO+O9YopTInVhthhLh4zBsrJVwJpQC/j+KjbQ10u
fTw2Dq1a2sxYGoC7l9WanQf4FAglzjv2UdZBN9uqmFHbhpVYlNY1stMOGlKu48bi
6U3gxA6Q/zmbhcziMqdw22229JcH63m8jIubEnbRV3I5P0eRgmfeGnipcgmEecgl
EQV8tvPTGj2X5H8rl7XN0LzMjA2htPqFXs8pinodC+MRTEOBotJkhZY4FnEPL83Z
LYH2jBCYOU/aD+rdpcpi5TJ/CM+UTkpWky0W401Pq5F0D9cn6DZtKkJY9KKWK4Jk
Ea9lC93S5wskPqyWWji4Bjx+tFEcfRWHqPReGS8pcpHJOdpx6FPkC56vLWMK+uS4
/4u+V6GthDDfB8GGd41W5kAFLz6ZRfhCjeMelcyUSRGWeHHl3AjtKvAIMoyjm+oU
wG/eqZkT8NhTjwWPC8NJpTpug7Z3JIMUdumYsz2AwuxPD7KG7ouNCbg1fUEA3UWf
4LQde5I81q0+NpgOCPBBBP9Wet2rg+Zhqf1TGjJ+s0iwXumOCCqv8TdxPB5D1BtG
qR4xEGvJ9X1iP4jM3nYngo6WdxpZgOP7deZVbFBjgdKXhPiw/QHjWAsA4gdTZ/Gd
N5B3iWcVeM4pR/odqI83ti8M2fXHwUcUNLSw1U4frfikJjpGhoZ+NfYQsNdxf0i1
ucpWEE5amnoUXQ+MDMip/iOiyFu1nLtgS9KNbNdJMba3pYAVpvnHGNkbYXvCoy7Z
qjE1HuhMdlch67Id/gAgDwUfdKHiR4zk8R9nBF8HjmLxtpwn7zTyPYRd2DAzVFuH
gzBJhVFMoX+WAdMhD2oBMa9aE22sWwAU5uWrVi1V3JHE4HuQ/n1aYqBmlidZEM/Y
n94dLj2NixnLby02XNX6DVziF+sUPIFj3SfJSi7bYPuMGiwx4nBUDo0+wa13brIP
xZWwMTXVib5KHk6XW7Va+E85SApGS+Du5UI9kI9gFftHaSrMnZbKpcbTuDEFl0hv
OmcMeXqA/bHxSffNQiVeLy7/0KSoGQ0mDdjAjExMVgDxFSDXxy+KtEXYMBTIhldk
9byi4c5vwmFm4yMTStJOZTPTkgvDcntGChcYaEJwwIzmZsftFFSFqmOXHykBlnCs
TI4R4B3fPYaJ9Bhwuz6B1wJ2i2HvRmIEJAa6sGs19O3aF1vA1HoXJ6c9xoCVp5M+
JQfGZGpvfjvwsRawbfL7wftjJQBpw/fR3fUFZneic0qzwjlKSdF91GTeHYqrF8kn
0rYJneEnYATZt4I4brGXwLm1+z3qG29CvgmVOPbPvQnvWUM2JdaNKtN+9yKVn0LM
9C/qHZBK34WxajtD7tLyqMJ6/LsuQ2dQkG6j5ahj0qmFDWjJvrelO1MciFgbOBTX
UhlmfxRIrH5yaMWpi7MBTgfEL269fQy5T6iQ1N4T7tH/j6G905rzLPL+7pO0z13D
36qUgPACUxQzykCKLXraRx4dddXARZMT085QwxJIuzSPFn356Xzey30b+GWK4oa0
LSWf+yYLqyPwWw5CUqYrWUwKxkNt0BQmXxTCvaOey117wiw1fkZtke2YnLpyRXwe
gyP1pXvs7x7t7h2Li3lHmWcVVjXNu9wCeehi/S002+dEPnbzHM+W6ibbsTfdpA+7
JjooDOPnXB56wUEDy5eWcyRW9/utsUcs9BVa0WqRuB1prAOGLDBWH6IrGsyboSSS
PpS++2RLabxk0KGrdecLEJ6WPHIwxi0rQH/iZhLl2yBglN69rO2be0gvaGju6Z9i
Bt6vkV7dxlCQ3B0+RnPsRMwmPu8XUK3nIcJ++CLiHclp/CEHjfdteybxlYllEwrU
Oyqj1LIb4DkKUhT+HClTAwoLzAf2mBF2j/B/QzHcpOvueqYuydoDLdZMX5MT2a3Z
Ply/2XVNW44KelhGubtt6JW5J5i2ogk9FNv7gkRoU/MglYkPKZAtHbZweHhJmrCR
JrPjEh0Xzo4MlgEoLtlY+G3exyUNlfQpPvttMbNJMQPhlDgyzW26dPaDWNXQEzW0
f5ZmxArRibyfHATtxwwZeYoVoMoXivTWxOTOulmSAng1gPeY1qImBrY+Bbpl3hC9
3WAio1b64qKjc8Bf2IxmPnipQCfiX4rQZLwZCIC6U7o8BTNAj6I2DCJ4NyG4rSLc
AcgdBxQNhg7sVZRIFLhmvX+qtfeoS5glCdAdUZopm5XC8qvU11VzD9b0U4B/+AAo
2xrnuMNQG9TEcqAodfER0ailbMIZ7V3lNoCfQjKm6Im5rTxZb9IV83XZqpjKizmL
Acsm7Z3e7qzFrHkVfNEZJGPCpiXGEFE3i4xhuU9Yvq9QYSJhEtgzZAgYkCWFKVtE
sJFjnT3CAzEXKgLN9sffpNO7XT07K50xNKfBwEVHzMc/PekfhdSS4eDdOKP647wL
aTkGEUFB4mNoggmcJLGc9wiUjZepZdrRiRuLFkbcDBTLZgkPs7RvDTgBc3xvG9Nh
A1uJmX4S7ojial1JuuUk1W41Xwq9ZpDfBrmKH3Dg1yhqrW0Qb0g3EGOZzOl0mDES
4Ydi0SHVj8vIGJLMA9b2ouxkp9eotWVRZGmK6ZZi4YbEsAO1HEPDfq+4tTteIcxd
C0w+DFecXdrQU88oIgnl5Il5pIadTTDsSR+2npfIU542NomU0IpfXixCGimvdGiv
Peid/Hrrl+6DRo3SfneN5KkR9aFaX253PX8R5PUCJzOLmG46cZ3kBLrSjbS5iRhu
26dseuHKTC350JJKe6vX2WG5J9Y9QrNqkwn9EvzlhPD1+0FQlPSTLQeBc8+vlb55
iGsvjDAUWoO4tluHIzg5yy3H6DAuj5zmRR9FTI73LPXTeCdtpmI7yxSwoT4fNVRZ
P+wqDJGyD2oZpkSBN3l0oxYtdqhqhMbSKyhzkxSun1Fte0+oGvzPFE3kNnQJnZ5R
dF4mo7WNGour4m22dkD8E33Jae8j+7E4Tm25K0EBc65bwYgCouSB9s/ipVs9mJ6n
TFD+RzhbctYzgDWZJHZEIkITSufZYflTkPE7pBrUTnuoZQBDMW6zg2we+Lf0ezSG
O6bQ0jSzFwBvTO2748e3V81/B8+9kOlHU1dnqriq9JzsjC4KeqzaLGEtmqSYbCGR
+1yMVD5uDpQBJh+NeMOrK33RjXoU7LHiW8xI3KwXPo2/wjxKPvtww7sGF4wPmY23
PCXC78Vvh5E+GZTSPeLpbvA3THkbV6Xt5KbTvV0GAn5PY+0ijDYRQYJEdlgCqeRe
76bBIBbZCu9k5T0AN5Eu514OIjwe/aASDhRYv1QJsFCR8x7CFFQ60Dh+/TcbpLPQ
6zk2wDdY5kd8ljNDV9cI2BcffMRDowfyR8VIeIyMhCb3olF9U9TCl7RjYbFT6uHc
g/z6Mt8q8PJRVB3rYW+IgMWrUYpquLG22PMo8Hvz5I2zzUQm32HIBz26IMKe6BBu
3mV416QjBwQmOcxNglhqAlFc1JQoEVipN8SMdQdM5qJtLqBtLg7Qi/8vwbxbJ8/W
CaX0JE1RI3PeRfyee1+lZBtf45SVpO5bAJEaBaKyrolroJ29KSvU/kgij1cs/+nq
jzMSU3ITR0Ke4siy3fJiZtOMa8dwQyCH/zesUhkdgZaaSSPHsDkxN/W2cph0hDZv
AMbEZqyd9K1gnw6jn6Za6wbewom8zPeglcTXFS3L1itP9QLTynOoYTIKrAY/ae1L
SFQOtmKHO2CaJ6UD/qU6sVJ+alQfADlDi0feH8z9fKSSmWMnQXUA5ydoyv3vrF1V
hnzYh2a2E/nIj8IuYzaWH84UFNr4c7yt+sG75oamGctWo8d7luaO8WJitUUz0qh5
z5KF8XTE7EUPKlgoTKaeBo37yTJXRtMz0B+8Jl+JcPMN3aCBmXT+eQW8olyBxuNW
QGOrWAvbf56raY+YAdg5+4i8b32mWo510Ha2U/GKOe6HSpz61Yx7FnVSsrgUZhxw
MELXRLdT5nvE1GwNi4ehLr6j6TMr5A9TUKbfYE1RNteeRswmmkvxqx505v4sDKbj
rKB1bD2Y2i5TtHioP5P3njtJ/g8bjRsAeKL3oAahR3s84vJUuwospuAWAKEdSbvW
sFhWuer1F4c4Yg4EfKff3dOoo5z1WyZc9vV0XD7kiK272S9EiWGLQldiEUH+ZIUB
PJ2xzmWeWQHmUqI4lb1PAI0G6zeIs+tFNQ3YCdAHpZKw5JtAFOhKyYfKIj7RiD2u
OgIo0Jqqi/WRjYbJ7+TcdyMfBJr/SY4YnOSn9hUhCBtXNXK9zSVi5Qd3EhgF0phi
iBQOO2ES9n4Wxo7FYDNiqXQ0p8ERbZjLXJf6ecp4LcD+zweKeeVzLOK/P+SOcOZj
2nC0zAePLF4piDemA7BCjeeGShZtUDEhiYdQGTABVWi/Qdgnka1gwc+Fmlt1TiYT
d390dcjVcbRHkQ4qcCLu73hHWVbfWkl/twiRpWrT7FsHooozKUKDRvIKi5K7iYup
RvsJcuYoVhu9au1b/Ff+2rzifBjw/c5V8Tmv82t9X/AaSzYpcZpHYNylOsWBZ34S
4KwQBH4GeDYMBVPnmTbhVddRr1JFSwYc98XPmNPA7FwXkEWrpiUnXm5BFOj6SSPI
SjxVk9xBZK1cR5kEEYJXn8+UZm0sUSjxEo79arBCTOKFascxFSQ8bYdbogUNvZhb
jzOa9y8vJVSW8aehDr+nI85vJ/9JST9knlPQGbMfDfLvLmXjhq2kCqfMYkmifTlc
rejXSPhJ/d6aC0KRBFOibFRc8YSobKz0+ZxbhBIyym6Kjr7hR1yeCwhUbeGFqNm1
/A4+0A1xrFuMb0jQQRKSgGYDf+XKdc0panNNut6LwBpDCuWK2chpKHvdLmCJPQiv
qpCqvlEn1PKglqV/45dGYPpopwyYZWaxGu1hl4rngnmVeDedc02oIGE14OKjdYB7
x9BTFtfo9bNtW66HP2LGMnXR+6204+GYfbQAcH39HxLiG5O+XF1/EweNBAfZ2b8V
m0p+a60rh/zI8a4C9NrO6EO/+aru95Aen3+iRI+cfvhIGkdfwnF7qpoCzQdEVNwZ
V7jreK9sa0ibBnwH5BWxv4hvF0fNudLx54vEZ7eo5pSdr7mb8kVIjlfNcad52ZlY
ToW6DsNUhqhsXU73PsTOB1b0Vu8bdLSBC6riUaujz3pfq/YJM30PCmwGDq8Km3YC
ObJosGffe2ZUBf1BJJJVfhVCvTsI1vPz7Y1rOT5JtveCzDyXrAEcsX6vzgdCq8Lg
wxYZeRlyDoCfB0PYJytBdqyoDJGhIGz+Tx4zZPxAZF7j1wsM2UXoYeXvmvBbXowL
MgDRLQDnfntmpzLE0ihMhLJOOD+sjvyX5EOtXLShRgaHMBtzlBUNBlkwJmStHYd3
Gsh8h2sseFnYEIWnvaq2zwDlFJIQXNGQpm6atCvYH/HGNK68JuQeH7AlFwIgNOl9
bvOfOk86GiXSwXZrC5aJ+oEuFnlrxdJzSZ3KDbcSzRVdvhXSGuV6q6aU0AEQXl6a
tN2k3bwgFTR1WSCCGDU89G4ndtETfRUIdoheoFRl5IDF+Hki9mcljhSG/mvpsy0l
FRsvMLEoQCLsxhXzCOuO047GKIHtFg2pmioIjIlittoBwjV9rR0LkDu4vViUy/Lx
57grufveDBWG9yRxBdf4XK/zwbmBy9GRmIryraMg/uy5qZg51syfvHR4kIAF7RDM
tqKnCEiHpznBChogwQUB3kpVMOVBNRimmEAPc7qOlfuq6OtbXJ6CLBWXWeLB2gwC
f98O8ss8j7yK/8usoFPNZ0WfRIyNTfDQpXXXvgPhSayeXP/f4qv6h0cRHwuNuoD+
FX83NtcoURLkBWf0Ocfg27IVthbmo53PqYh1r76/ZWF5QcpBmYUBmXzX4CJzUdr3
iQh7zyiVxZ0WKt6jTqiirX1XZx9rM9V1HulAcZ3a3kgOzw1C8+nKtHCSP+g9Vo3d
IT7Czkx1xlyCpN2pdlEmjDXgrydyUZPDHUDHPJ8ygybFb5flClY/CgPjC/JNY/wZ
46CwGkkv1wCGVVSnIuKUvVSQv6pOzza3g6PzE/5xWEzWoctt9q8jqhz30uDtKY1r
q1r+6yf3HwYnZ+WnMDB5tBKZndpHY7+4UNfH5xjg2HnW6BrTxCfZF11cauKjqoEN
PxluZIQAyLgf10PXyeaoVg8E2P85vTEvUMpA+kjL/I9yMAkO3G7amQjF6xIQxsLy
fK92h4BcoN5qPZ0hhsV1819zXmUU+44oiRZ9VqTbAgExC9Q4HtbC+TkIGGu9LPR1
4It8JGrTn97W75fHL5BQcWo2CCDCJam3nl56XRDbjxEuUoOPt54YeHQVDrtk+NXM
jrAz/X2tgsqm6PhnaVOfwdV5h5jmtYsY1JLrHb5Sg6X1Z4R1AwK1mNNmh93RR6+z
spJAAnqm2m0UYUE17zq3+YuzJKLD2B6S9iTreQ47FzJP2GfDvlyzzEFP/81uVIRE
4tK5RMgPKBvKhVUFJVl10dgswYQwdB8rvWz9VR1r2cdTfKALAoA3qz7gtCOegXnU
xYeKmTI1axzGKIkoPXBPzsIdjpYA7C0GNe6zTKK1EvvJA2+MoxtEPu/0Hx1H/N/a
IoLfb8zPFvRqfaWEAdNYD6U+GXNkeCNbqPBTkAVmzUeP7us265zhQ0PgTv3VMgdY
RkRcW2b7f2cJhur45T2mm2UGUIN6Ugr/tAQqg7es9HRoOmpie45x7HfJRu11HmBS
Fm83SL5dn8SrmaURATeJ1CjiBeNr4G+WSZpgznMY0qrW3BcRp5kIwgoqJFct708f
NrKN7Nj4Ei0QHLPYzOhSY7UIpPlULtQUBSx78jhJSnJxw5PwMHoWzG6YfjVV31bi
ZmKi6O4+kVAIf6RL9belFETx22FKtdmuxCR0THLPZMYTD2ozfk4zZox/dADHFU/U
WgaErCrTnVi3FEJWPEkS5R5Ys8B1ZRRr8rxqz7SblhDr5+8v+QPmPuwWPcants//
yWpuxPyvc70ZSmrOWjS1Zafua/T7nHh7dnlwHZVkX8h+KM6M+WOkPWJkCYakCeqr
usvbLIIfhKPcRrts01wNLT+NPYd5CS0r1ReUCV1GSwk11cX4Ka9HbAkWAPwh2Hs8
1D1eVoc6uc6hhL6phzejvLO5f3SpfUUAVdp+J+XzUZZIbJw8V9gf7tcTMHZI0rts
P3gDQdfcZYGcbADSpTB7r4E68c8NY7QEM3IeVStK1Dwxr45vs0Xs5ot0zhjV1UKh
tl1/IVpqL9J9GRB2iAtKfq/M88nvVqmnbHBQX+7kdg+PmVquA9sq/YQipCoWbPGF
gd1rDXd7eDAhiir5Ade/lfPc42+nMnE0U8QoFg8mDFyviqkZPX5XJeJDnLtU8iQK
wr9s5g8qBU/+oZCWYQBjQ3o2rYq+p/otjoZdryPueLNI6+BIcod2xFoEK9Nctowa
4fnM/5XoAzBC/nojgn2kN21D+QYAvU0nLKBJUnHtbmx7V2oe7Y8CEc7wBfbRD2nE
wzBJS0w2qJsOF+5lqR/Nk0FEZkXKQFaNdNmSBTOVSaR7Ecc3UsDq/KVBsgpzKqRt
oE3e9v09y+KArMPmoWGO7xXBj29StyUAUwGKZ+9mmc2+RCn0kpYqnsJytt/8XB95
GY/3jUaO/KB852YnujG1R2FP8uhgRBpqvKYft8LWMDuLSJinvW90UEc2XbFhYz5O
HkIYzmhIejYiji0inl1fCz0maCmkxOND2scC9V7422msRwaN6nKM+HLFAtEDfX0j
GeKczzAI/DMKs2jdEE6F37ORaU4VJgp7a8ZdbcTIEoFyvpBgBzmJjsvrv4vfragg
YVOb6X0tVu/kfd5MSoSDXt4vSCzDuUosnVaJ682p49h9dZ2VFByRBFwRiRdmKCdk
R9iZIEd2NRA2iZh5g115LE6uhq5Js0zsYLLICZQ0h3fWWjByaI3U01T1dsVvSO/1
rD8FuSf6LzI4mZjueOqVAEzpQSMXNScwFKdC/mn57vSl5GZ3BA1YAmzZ6/4bv1Iy
psy3zKwmPJewBV6kCUKphkmIDMUpkjX1YBkGk35Mb0ZYV3iMiC96MnWid4CEJORF
co1EsyuJlSiBBnI+yO1Yui4L+OrknntgxR9W7Ffias8P+FXOjkzL4ydSLLGQUtES
BoG3mjxJsjgLWNdQz9HRXiQmfawUjecr/mqW2IvwpJEbvgAZpd4W4p10tg0q5Pwh
7qI1yGfxLsN4HhDyFn+30Q4N+fHeby5C28zrVaO6wo7CCv2lmsWx5UYmz1NN6ybX
mtcfM0R3vLwCfD6IJG7OS4LalIDypT649FOnKdJGGGdhb/m5+AN1Yj0K4VptKFUH
B3DfEYdJfRbJH+YgzhMtQR9YCpy1jrzihcSy6u4gl0udqK7O2YNMXEUq8sHWGCBK
HjncerrTb3ka+sniPTPoZ6rczqG+UfYBDl4ZBclrsziFF+rpKWhf/Ps+k2s43B2J
vPZx6lp7kja00yWWCx43eBopKa/GIX4J2oNLohptM1tcjGMIX99jgDDyO39jxXo8
yBHvHAc6TiRSYYVEQYJEXqA9P1RJHrqfm40gqHZxKpfPhYgFbsOm5gGb4C5d63KF
ovxLb7bKyM824WFPjJuXhsqfSiTe4Z4k16CyFjkpfoHxHGNjgpybboQUWiaFsMJB
dro76BSPlsoOHjOjSRx7gDoJKeFbRrV326FLOFv3Zxd5g2OS0STwGV9/5Ihd4lSK
T3tHgF8rP01m2MrqEyjVwZD2YnRbVf/3serBCRAdpzlv1QozoDuytJHiifapOh54
cFFprpEgFYJkN8eBJC6+XkyN2pavfVcyhRhtLtzR3NgQqmGZI0St7NFLkay2NI09
si+GECqt5IkwVOaeOb+BbVz1TRu9aaXWy3BMqzm/JTt5rLBemvdDlHk3QMtA1Xvo
b2tOReM1yIZL6Wz1obO64MIWL5pTHFO08QnC1t0Lp7uLqXNeNQmUefp8eOkAvggZ
1rM+w4UE6qOpKJYNzf8yL/QRCsGqMJ/AIMvzQDXZRD4UE23xx7FdOsNSR8cP6Bx/
vlDG9FhjT6Gj4a9Qxycof6B4wffdkpwVlK+Zu6BWwukayUTXQW8vEn2d6OdaVJ/q
Kp19TZGREA/L8sm+4YwH603TmQxccDE6FWhCIwO4HG9aOw72S3LfSpgKE48cZiAH
em3/bklWtLfv5+XzdngnbCDRBgoTh9VonkYZNcQoEBif55eOgqJv5OJ+zSODOoFn
c7wDbHZzfZnCiqrkfHeA8p+GyJQ7JW+87gI1GV1w45mD/C6WHmd8fyTAcytoEGFH
J2HO3b6rnfkbspvFNrhuaIq/5pNLIAhnC+3aUDUjm6PhYpmvwAAQkEmT9t4vt/6u
+LQiByWfKXskzgITkaBo2I0ncVkJJhSX+6ydAK+rWI8kmwitnPxJQn1ZDBDcBHcI
JnvPdkuxiI7EAI0y4bEOlnd0TL0Vsx9SiqHcVeLIzr+XQOrH7LJ+I093slV9rTHl
OQFiYPf8Y7OL23F+rho/FisuQR5E7fUjHDyzoJtyf4dOQgReaNbu6NFKi5W1sY2s
4fSBdtznYAYwJz9eQ+wYGjbIarl1kH+FP/x2zfkGMDcGlTMgktpiyAWUWiJ6Pdhq
mvIkF71ZHqrWqRnjjos2SiUSuBeR4z5EcALfVKiba3Fvvt3cNdJU9J/Hhg09TsGX
I2Wv7DoPTv4uhHoROhvXeYy9y/PcbYMpiBTOucJgDx/thqiIsS5PoZNesERxXpmE
32fAcu8q59gb4l9eF+2u16tZ03R9H4SeCrrG+LtS+8hvzds3DQdw26e8eUXzZrl1
tNyI2uaL2lIk/JUS+TlL9OEfwU2gQCjmtR/Q3AAotzXI1fHVKefkSEnWcGkaS4+U
01K4vGhHCxLyorDM5Hx8qE0h9tKIbwZPoevXdwhHNQvuEuD3LB/j7nLvAm24s6EQ
k7yEDfmhcjMfN3IdH+ODGzLP0nh9ACfhY6wbYF3cCXWMF1XbQd4DiITnIHyHNYW7
WL0kC+vSzK8eRhxBjUeAoBIrqVUSM/jTRmKn3cZjBb5uPTsGgWvtmJH6Kdh7lfgW
/P9iPuS1WggjNcZGldn7C7h3Ti3rnk6jHAGT/S8zitaodBHjC3vDYYZmZ/bGzWUj
Y44ThC+FLjSrJ/16w9Q1e0kqg+vhRqLb50VaSFH3EPfdmbCUX26ACTn+jYjDkvUG
3Ve8798TV4V6wbdsxf/7qGVP3o/t7vsVf21vKEgojCQZbK5tV2HPQ+Rf2OWdfwiP
ETqhuHTVB196WUHfqbD410TFfuDfY9SPucuPLe04QosEuq6ZKuTp24Yfn6k7Lz6i
NafXYG2xY5K+TM1NANaN/2Mho5004MCJU45GTTnoPkF07WW9NTjeMRVG7d8T+nrd
zFXQwFysryCGxazZ48OhnMYL3STysDkQ+nb5URAguyQjxQXXkksjs/DyvSusFQ1i
wqsYs3MonEpPBYZK5Q0TvOgbZpAXH2Z2DIdJRTTpeNlvz04fHd5eQPedabvDvGWN
TTkDkW4IewWtUXlqMkJMnmXLfOaOAziMl941a+lku6LOFgCPFWGjj3oe+Onc47rW
edtTateD2TT8bdhFgZOdY/HXgOx/xE7LQMfFyv6CAKlYNTnXxmGSRL70gdieQWPY
yR/TabFkSDm1xD3eDP87zaO+hJe2YL12aXcG3y3+WjjOEnmvyPMjPpmp5s0sOnNM
/r8rYKOFxQiWu0nMUmsfTQt69TldBGTAxzvMjk/TEKSDcs8VT+0uoVKorOBqONqk
6b3uxUo9ZGZRIXKYK5eiXMDhAA5EmGNYqB2CCMmLXlkXHwpWxC9veUdzIgYiSxDA
5fk/P2+OI1lW9HJS8HzEEapoy4hmkbuJ2M484uxCoZ8IQzONJVWsBx0AnaoKTjyj
RBSL5GE5livRl1Oeu0VGWsFFP4P786oNNEGjP1mFrun1bJuAbrvgy8DXUPWzMKWk
CS0+2EFtyx4suw5vblz7KRRrIlBSiG87oKXKIcQDri/ZBHmckWx6R9HWmKmTHAui
q0w0YFCqFUyk7XtvyhmFhcM4vy86Dn/gx15mpZdBc/8KG+8PflnqVwAYV2v+Pfp2
NtoXX6jrXgAnf7luCOOx5HBZghD793st2De8+haZQq1H5X1BGcsasVPZZnySDiyV
ypvSDTHUXLahakgmkkyGTFDJ+8Jp008oDpoNlx1J4PumfxmjD/baB+8ZTJfdqZKJ
RKacek7DrlHmoFw8bc78OpGLOI7+1+nBHmCU7ue3332xcqAvyxxxdU8buFki5snx
vOQeifoeDEWTryeKn/dY7ni83+YthsLm51+AG8tuQjPpPhgMqwC9tMK67NWKamL9
ie26jWoAQuuEWYG2ATwwoBamnaTrr8JbNSsh0jBxeyKFFUkDHmwPsGVAffarEm1v
a5aLHAjuonXkcYt2qjS7VMHp4gGEnc52PHH8dqBvw0VDqna8SYj5jNpXq79Rc6Ru
9HdIOj+sHRk6hg9ldjNxjdtBwiGRgJuIy2FBCOE3dc/hP5u+EceNx1Y9d79lIlXS
zWKez2zhNClKAFx+xmwhNEtNluL+r+Zk0ZSJ3tRKeslyut5clxyoWDYjVgWwqe9C
3NSngRk7FTWLrRby7rwypsUI1F/5Xqu1XDUDFYo8vHODAW6fs07I3aJqsJuL/fM3
foJrR9FFzj0/dmG2HvNIzbtwgZ93xjo6BNp4yDqNBDCFvmFLqN8fYU45sBoHTR0h
O7hofNiEjs858zXpne+RACdisLPaCES9+9E6wA6fWwwzOCn5ckJSyqBePEBKqpTz
Y52V2uFALiDkevgQYasZOc/MKBYQXajF+G+hFty3XHuWMDVYNPcnn4fNlblMs9Y+
v8yBgtE3VO9/eOJbpCJWwdlfMt4VBWu4pL/70oU0xWIHYAV8KIPb0bkegU9ngaMO
GaIdnUcHshzYHTkPfBT7qmFyaABEwnkcwZIpul1aQLC9xDLxSOPp/HGwxFbBDleD
AKfwsSO+3COktk3FLEj3ImUIY6NdFLUOpc5FCLr0lJsLS/vl04oObfO1K3wtyyWs
ZljLZ8vyPg28H3vl2B2HG8aQmIOb22lo4AbOVW6XkX0KmPX8o3GzRjhoYPo5sQ7B
lWCU1RZy8l/dANXxQ7tuZIuasZ1pQWhTEvcBuGkovDN4PFZlp9q3Dd3NeNj1aZTP
KJzH8/8F0yY1YTNeZrp1amR8s/VOLWCfNLbIo1xxPQHeL6lRq2+Rl9wOQ69BTQBW
nJUtAFbK2+auJU32gROFVrr4e79nZSSliDau/CiUDUsOz5OEW7WMsFhzPr2HNGOU
ChwE1xHNrmY+d5XQ/VvLpS0QWeb/ZO19qkgGNu/LkyvtFB03hcyr+pPta6VrhReN
8ndNRX8ZovmHS2vWAEGiSoK/5gK/YCqppAWZlzKnggJvTpu5ltVkDf4HJrx7S8oL
VgaeLXdwmjDuoaUZGbJqWa4dn5vXuZ3fIcTlhD0ebtELVYDJjR0xcNshH4EpKePR
IuFq3B3Znwte0gO05gtR88RP2RyoiD+VVcqADzgBgK7pCoH+b47aSv9m8ks29j5T
2i9/2WEFHKvnklSFFhd8zP+IWBDiXd+SzCH7LqSHRitNzAe58/v+4+yoNPYyZKYH
35U0afHLn+APqJ+/0CKt+7AxEp+wiR9XmK2+Ytg0gDAqwpHnKsy1AUu/qZv7H4ZW
M+AyCWO2UyThAtTMZxpz2u9uQnxKHkmsrMkbFfOP5bnIMd1TOem1kKexf1Je/GcC
utZGWHwWOZV2bhJ2yJ4AsJGrTZ3EziwACVdbtMiCyoTKYpECCJhEHxJ6Iagb3eXL
63hlQ8GeB2g3UP7xMij+HlYcy/C9w1Exr0GNRoyo6Kmy3UKafpbKX/UzerOwOBM+
eE+H1xndSK+j0MCshZJ3M482+b5j18bXhbswzEwEiDjJnL/DCsJve5B2eYVjqXG5
BRKNgLLwE+BHid201wHUNU1R/r2zp68vayihZPSqcNscD8/qQ9zGXXiIGa6jsnbJ
KdFV/X65RUVu0QaoR1eP1EAdt7KeJ2/MziUdgbIF1T81uJ+/EdeDxYiD8P3Ci73A
hyXN9/mKv9wjOCRkNwA4lQ6FE+azzNWinXs87g2vpEeilll41EpD0n84Lu78rgp2
v4pxhzkkr+mxD/OQiAXYznCBJi44qywv1TScMsby8lKUYxhwjpdFsOKm+S//IpPD
Jvrt8gjxjUM/NnFSPlEXxvqk/s1k/rkHWbYUv6eSI1eCNimdzzjU9BZQHsy3cxAk
ogEiBApZngqa7dAyEyvYeFZy17V5KwJquaCh5RT4y0nPoI7+Vt6P+TWFYMYzggKO
aSiJ88vGu2w4inN9QZDLZKOyDUFfxPXAGnS3n4ga0h3/D6+C5mVQEt6MnpmKJFlg
M/bVnQGywvEhS/Jq+fvYOGiL9iF5M5GqXaPPMMUd7f52fCFLd81VjXe4Gqe0uem3
qEhMTm5x9VrpLhmzfVvu0BHXfMOpWJATmbhgwyd/brLyeh73k6HYt92+wJm3Evxw
yZlkZpDJJmixkuf8ITCzBaFYj/8V5+K4UG+lSvf5HvwsoZibUEJUn6GJFCzQdCtf
K3AGqj2GxADW2ZtXucwy5opyF8093D5cv9W7qHZj8RoGDH9mcrQhTpTGl/UlAK5M
J3mcad4+uDLEywpzofl8D7bmaE+XiwdyN7xZT1Z96W30LY+wTM3b4re8olVlPkCz
WNrTgfkT7XMApWI1TPi0mPlwpVqCWJFiFSvJGabOeSUc5x6DY9k0Br80Syn80xHC
Y5NvWkJtEwux63S8eIHvVGjy9KuRcBLlYFOCN2vrd0p2ueUNXrnqYhSWevZC1+Bn
hvfYtGs4HBXtzY65rffoicB45r9OSY+/voBwQ7M1V7kfkoT/zZd6FzPGL+TyR205
gvpOrnlD8PlwjTZouWGFxxlTxLLYpggDQ1iwBohwSACwSPJg9xpHG2nJT55ZKBHP
2D3bxRsUNn6UB7vpGN1smDgTWyw6KL0boQWwiaNtRBZ+LrDC+91Ydf9zzaPvNNTc
8IePPupr1CPZugrvp8/obo4op+8vuMBCvjJkUERDyf2G2aeluEWM8bcEG2T5Gjei
hk34Qo4G+/7iqdfITJm5BFzcPlfOP1Uv/EjwnSF2+lz2aWzuzTJXw1B6fOZ0aCqg
X9/OYtxF1Fahxko2+RTXBuwCmSX4nMjI4hFP9jZL4EKNiHO0Y8NQCVcT0An/m1q0
7GaJgdp+Rn/G8JPmTvJibsEiwMvyS5LNDayJBytsC4EnqLc2qcQXgU4UQ6LelKJ7
Q1uaAo9g/UADeeHFhWIf41dTZQQoDE2jqGyie8hGpHVo0iTipNeD51strYiyqPWX
JIrPdu3tk7KYNwljVTHjxPWJuaRs+V0XZ+td0ZCdZ9RBawQu6iCcECldpHhIZjrT
EyDGzISEltDoh4Shjow6iMNcaH+h8QDb4d2Q7X8GhYZ2E9qHIxPKVIRRxQE+gqav
TKqrgiumNEyeiu/ISYDAo3jBK++oAhf943mFHSnn/RuKRBwnaDgzcQ6+WP/w2pHR
ac3Z6LOr2RNpJYpYOf6Fg20itcHtgtaPxhoxmX2kNBkazZWp23r0yFVx4IeCJvyU
/KRiCH1xi1iqqq17sq/GXm8gzg/A1SwTRfTnQJY9O+byI5BW1w8mTelPeiWeU5+x
NEAeES7JTkFEIzZ4PJJPOlDcn5qhFNdsIBrih5RcRGDINENUYKl3/4ReZ0J7bSrO
cjOAtxsVJRjB6iO7TU25kBJI9kS3vt6jIMxnC0amZoDF9u8QddU1zROmWvNEh2t3
GH1pvQ2zQcjWgLv/q4Fr9x2OtjIugLO5L6szxR8ZDUkJPaaXAuOReOXdV2CbrmEh
H+wCZKgB8Lw5axbDyyiByvOOurKc098AKbbKzvnSpVkmG55ZHqb+o9MoIS0VL5R/
Hb02YxRrZ0iHl0cmXp8rPZhbYAPWB1ac7YJoI8y7eMBxKjAhJJeCFFvBGBoBZWSW
f6XRrGO/UAhFUwnnvPyfFK5VhQEUdWy6SyKhaAWmZKun/zjMMywq/W8b9BUDITdi
OIjPgQ0/vQBH+UYrWoleCszHoKeYVAlV87ZOttJyOPCYulKhTbFcKEoPFxxOPXjg
r1G7sWGrDfsHGMeMiIufrQZyS6HSjwbJietORWR7MbZlJgqyqlBtyZ6yGqcLBXOI
OAQZG3IgILDjMKBaE5cAeM8xIz/qWVMsrvGiB9r+CxfxbA2bG/E52mVTnGhDvsRe
nDGZAqhwQ1D3gd+WISfcz0t9bO4EkDR0dmFGRtYoAu9TeIXW5OZcV9KcXlEMB8wL
oPY8ycDECGrsNf3LS/5rLprBKcdEvyvbUVHgF6kvFsMy/f/o9o87ChFuPSEhbPmx
JDu85yXgeOxoRLzNTK/fyJltL0X8z4POctVct/xMmxssisZ7Hk9mjLi7qr0AIZyZ
8lQLA3kVdricH5vcQUClZ3LRsoRNDAXI5rYqnxldxFdO5f8FK4jfpjavcbu7L27C
xMEuMGzG9ZX75nXGbLg++PToeZOFRnGIX4rjgG1he5kKQfHx1sPThPFBGJ01Flqd
OB6XCoEP+4XNg81f3Ub/nRRCBZdnOk6jakjJH4MYMgYbbNXybsrKk15QKRqDW9Ua
/sWLhgVtmMuNP7UuUR5IhuGDCE1udKu77P/ig99+rG5e2hxCt+MdYxlJtaZzlk90
x+plRthoXsZ3WJ0nwFRKdGPWU7NMoAchQlG1pdoXN1JV/Ttb4H5KYPiikc2ZZXim
bzmfjGf6oreG0aKlMeDVpK+0IlrNlapUjIMkR0qK0BTi/1KdHI5ki3MvMUrjhZFb
mgfssarNx0PVOx9Yb1bX+U9Rq/T8vtyM1HIUl9mzxATBzMNezEoej4/5YU4wiajX
V1ZlGV9pO4PoxNd+/K99JWDnCn2a+0xM6JFDiyQV6h5RgVNsZ0jIVIJQ3VFzDa73
xtmDArRXG6cYaujkdkpyBNJULDAGlqBmdl8HZ4zxguON4jcHctrcbHc4LIJNn76t
GhZd/6gLuMlSpw+Ji6OGwtarQo9WFrwnMOI4mD4KZIXKkoheK8VJrSGG0T+ELhTJ
wl1e7Gox5c5/KITwU14Ff+hBfrpejtG65Qmce2A/z04iGkG8NaISPyyvu4LFLrSL
4Kj150UF/eoX/CEDdiXk0Lms50kqtDlNN5TN0naufBjx0r45IvhBzYkWXuxOvt/b
NxvDpclxCHXn17HxhoJ1kO7sg8tVrToce9e2gEAgBtFPzB9Z2krBos2ACpxq+C/U
4OzocTFlRMgM9HcKXk/784ZBleKw9EuHlnbg0bO1J5y8Gq2dBu2ozOO5q6axm2nH
crSe2OJkyiJNpqdwm9BI+SNO1NBa5qiA7+EpaChP+Ag0aUxkkvmRSJvRBGBNgpx9
ph5hDLgdAxsUnDT0wICPyb0RI8IU4vXyOh9EJn5GNED4DlygpAKihQA8eebw2WWa
dffX3UJWhfKJcnz5bouIkawwgbgeOjcLQb9M/qDzi7/eckX/vIgahbgg6/smc4YG
0yhrnQ2wTzjG/b1XJIPcScdgQkIfL0b5AK+VXxYsw46A9PqiSqhxp7FZDd12vw0t
CHfEGAk//53chJcTIHbFpLqoEemkJREHqcNkNcgfFh8wbGN4rLthlWgq3gpkoeK9
UoGdTydkjRpvrTINupm1BarWCcWk+ENIfFP3bZ6dZSgF9VZn0wTEI4hmcPY9WJWN
4JlszyHAmAxPkgGaC3AmtlmNPtjO1fsLi5v0zl+oWi4bKM2xAouCbG9z8BTzLoKY
MUoPZ75rU1oc+xZseK1o59v/W4aG5K4YCiWk9RNXd0+YP3phTbZO1YOtnMiHbM1H
vBId3kSHLmiEsFwUag/1afLGhKYUcRot1wYVT1027J7JV2j1w85z1NUt5N0boHph
LFmA0IbCep7oN0Qo7g2OIVY7ji4gl1IkEEPVnguDW4RIkrA9qv2bU86V+2r+d9Vo
9nERdE81hkQ12d2loNmdVsjcwTlRKJtbVzB6wZM8VT2e/mRXijFvi+JRrOoNcvEv
PIPaEDbGpc4L7wi1VmEth9l8TaisH5nfITv+m4pDpMBGPC2nDm5LvqRLf70355yu
s33ZWEN3nvsyd51lgqBAdE5KKUIBdij2Q545tRG6PF+iC7ggTLaa018+BsVNyOK8
00SMqrMCMzPPFfKSfdGz0FtmvPZkkV8/C4xJov3zFfOGsYe+u6Ssv+MaLxRJuieS
wURE1n80dnhLdpZdUH6bZULuuEIGiICeYtHR4NSkJvin0RDvvGBuc2QBVB9++wbU
WUqhH0CiM5GoiLRNJIo/hiCl3a6OZpnbQGzx+DSIJulFWV88uGRTEXSBfZ5wIrnE
AUhldIx2KPMRLH9d/C3ope3qaj7Dko3g36BOO+KG/cJbxZYBlwNkdKMaMrhp9Ix3
bGNnMZUt8nVph4F7g3FqNmIKUYampCg7J3iAN31S4ZmCQwRtCTVsGXMU1y/jA4N6
D6CUvX3Ky8RynVZU2gsL87PmUJ+A9GH3zy7PN6knQw3wLtV9GuMuZr1o8aojJ4zX
s5F/ntXo+JVuOMh3lkOgod9NIUM89mLqha2DBFuyYZJ6tO1KB2XJKBJKV3G83i7P
Z7Jn1XYBWw8nFxvvIK3v23jIqIUP2ueaLMNMHGGf0Mmza3U/s23WRqXSzRCzvNii
pd3XGNyrHqeuVB4hQbfUwXFvRLSxCV1NWlGnD6xdgMwRYE6YmWEeaNeYkKFl5BAQ
650FMI95B29PB6mnYmBKcmi7DaHOdidDC7/gSw6OiwRawoDfo1xPZkfGvrFJSeMk
59iuo/R/gv+uzeJMt3xrRrqpjk4mumLjLY+ZiGCwDlCrPsiKJcZc/RzmZHes3xRn
cGUC/hvzHdjPRDANRTSxO+LK5CUMA06DCVryQkruHwgzBcxMYjZv7JJ60E9znnuk
Fsq+iKW0jiVkDbz2Sd6oJMu3NxQAE2j2yajN1fCR3VYsNI6+1W6rpsBl6GU4Y24z
L985nnaxwBZ8rx0xsFj7vw9ZxadYZFdYHJ2a8ebTzH+0/5ldReyVXm0YQQR/Krwr
7jJ+CMRE1ZJIV087n8resFtZkjeptJfZ8ejw6BNFM63CBHshk/RxD90vj52I6O9n
XgXCDY2iliKZQ4KA0UzGurQJG2KxXknO9aA1+Cv8tqxNtg3f7mbVAyQK3uWJw5Ar
bhG4B+SSz+DpyLyV4mDlTf20VZqDMgV8onjvyqtyEI+9waMRS89LUOe5WSZa2nLo
gkV8d74i2GqbuETVk7v+Yb0OgrG8ja13lbFm4lIeiFYXBsKx+yXzcFqzfbKDW1G/
lrUlNGvOfTc7dYVjgfcsT6qs4FwjUbu0hD41/tDswFD5z6qo8hWDgvxGYPQqXmOQ
ZWdVdOJ2EFFnveMtM8hPVlZoNvZcHw/2Th9b5yj9ykg+rnOpbcwAidPgGLyUx6QE
BtOkZggS7qD7VsbodOEFiGC0Dg2O5f+/ONewJEfwVsOIpI5ZLWTJ0rTK+8Gi+2ka
InGhVJMsptngYYvjzXa/wcnhd2GHA763T+ChXRNwLQikRA1h2iXF1mnPETZsoNYN
Wx5IiwBHe+sgMwssIEWSm++xqOHxgfZvYkXjtt8BH7x2CO8yDxC2668Kjs5pOW8L
YGtuGCw8IOUp8LtqnXMb9OHcgNbrMFHd7s7oQD+d2aVIyh/BU0BU/lr7aSl1jvSS
eqpmcy7vL0S3AzfV4J93M2OXJz058Vtm9qPk1AqQJIrFSZTrkTyLuU3AwidZOXUr
U+9muRQY+LLE3f5+nuYyDeqSKfQnR2C+y2+SnsUAASBFctnQEYU3eAtt9X0sLLh2
gf/BvBG3vfS7f+mbPyd9gMThkEee+FRYEFdkNJijBPijKTxtzfGfhWezIjCHHmml
veRsKR37hFpygbizClSV/kbZY4ts7I1osQfso7wbsnrp3gSxcs6ds49WEa2oMoiR
H1mADkGzPos7OG10NMTO8glaBIX12+Rv4sHINrAnSvl77e7btv781WAF+24srE3h
fFZjTnJ+4AdVX33OtK48Hr7n/K1xWZ9L18X1cGt7RJMi+OhSEVKcu0QLropC5Y/3
XkCG2ZKM9sQ+eRVBzrZ8SRHzMshTsgFx9cWRtldE1RQRDQcI0UgRIYCKiNSb0ph8
TPGnCdjwXn34o/M1GJ5RMPSQzGfVeaa/uXSYXokkr3hGOUFB+S4Yveyd29ZxB6GQ
Zyrgewy+0Ha0qH797V+q3SINuHyOhZI2g3F1juXJyCd0fh6KlE5yaXaLMT2WiviB
WPvU894zkuhibLejKSEfT2QmcyvJJZ9GYAlr6nv4f7fro0Ujc7pGwwuYGTGvC1ue
dbkCeM38ZRGoWr/g2V7P5Rvf716YucngZ1ZXqeJAQJM200fCubKGgaqm6LtPYi6l
eBa3Yf+s7Y3Ar0eRkxkOM4CT3cxrE4bs9S4SVU7znWF+2NcBsmeBb9lWT3yl7U9a
8/le7/6TTfqd40UJ28gPjPl+L/lQvMNlkKgqw6wo1qXvR6eyZc5ywPKufteknoHo
07B+Hm07Rnto0By7AYqNahixbDP+xm4NklijIIu9b1Faw6u0GNckxcaf2vTlOHj6
MryGhenMhHbg7drHKIodNdz3bhbSNRhHGBEGA1LPFg3YReU/SdN1SQryg0uYBFLU
hhqTXdGtdkJgWexiPn9jPsPTxOpCw8DPRC/GOQ7y/XZdC5Bx/A8Gggd4vGfICI2M
kQUGbSsgDmBx2tg0CL0TYQyzbe6jyksznSdAtcjbHdnYkmhl0MeUfS6OzIKce1Oy
GFKmzd5aaE9N7xeYmsOFEtXHdu8GaRNtqG4nKDnFQ0dsePeiqwg2qBsiCvsgi15x
iiLt/z9JIvezN0KfognoUtNLmtJSxxRyk6t3sagtLHNGadey04VZ/mdqRukGrccL
VO7pHreK4Zan5UFsQQVebCsnBtq9z+0viZiwAxt+TPrDjFYj2fdjGWACQsXl9yND
zLDVp4OyZ5gmdxnx+OGvUEBIKofJBN1hH7z+RA5IM6pXc2JwQDxzJX09E0OYV1Jo
M1VNP3nyVgtIwD0jREWsAXiWihn1s4g0HwybThQt+v96e/FCkHsypM6QLOg/tyr1
OEtHE4Qc3EWqhWKSu8fcGzsU2Ptup2bWPPoKrsikZTCWzdkXKYc2C6Wc5s54Scgp
20L/1J18X4UUE64O9rmJopK0dklikUGKuX6ZFRFMac1sKwnsib4aCQXAylVA0rVX
a8BKYE3NADZYeWLj2iDx+aTiQIpRTgDyaHCSqCqGuI++fwvxOX/D0FKuIUZWllEb
IlrQIe4rI4G3vnoFMr1OzGkB2s9Uw6UBX8bkSgiwAcnDCATAT3pjS7DhlxETc2mb
y+Gis3PQqrryOzbLhjz0UnR+ltp2ZEd+9K+WfUJBgI2NGMbUBs740NE5NLM7ecTj
vbdn2h8WNXU9uxfV3biGJBitls7vFos2tPTBLjF2NsSW9vZ9m3xYEjXraOjrgJJz
nBNzFj000lMfFRBmWtBiLVwcgQ+SadpnSGGJM1MRvQLmRQBE8032rR4fhmGN40d9
fK+yju/e8CFhduC8eB86YJQcijUj/kyOt/Va03d8BUHZb9yojNBLICv4xzEei5Fl
mBDjNNouLkPsRK3U/KypcjEeDdaDYTN7WNDg/TmVUdi26/s1Mf6GsfBa1Xc2DKS5
/7m5cnrrTXeFaaecA5mS5ruvdL179T3+3mipaU8DNHA2zUMVg5qoC9VytJkiUl0i
FQoPM8WdKU8msZImAycomvHSYI2Yl5oa5L04TLDrjBY6acYg8nc8NB80HSYznqzr
ADtlJ4vQyjHEIedVG4qOkQ0LuStSOU6Le8Kia9AFaGLUbFnXXpIFSTCDcQiGE/34
SfuQWyNZ+Kvh9YhsKTb0HhlvRdl+3lzH1ePKiWPRjwX/lbQGYVO6/3FfPpuGRJgt
Sn6f5xwCh4LHaKzXAUclTxkGEIDvLmk7mZ0PHC3ukutAckRGExrLEP3TxYOqCp9A
JwwMkBPmBakSZwwTh2kQScARkPWGrvEXHWkflmY+IJxJBRQbM1aVzerx/BIliFD2
VMRIfVLdi/poG8gNVkjzfAeIdcquxMwUY4yJvJtdP+JMHUkcP3keR2E3eoi/RXGh
W2tUBJZR8agzWIF0dHxXiSTYBEXqjlyGq5NAEL8RDdonEF2QgKHAbyaka/We/nr0
Pj/kUUzqOOMewu5bCBvSzHFaBfpbEjbm1EJs/K8lQL61hUoR1La7YEA9EtzKpe3Y
pNYhEjfu4xzse3gY7o3VWSUMMXYXOQoxWtFcwcR5jg2bpmkhAPn4zZeI9KypTMRc
cyqSXsteQmUgwkgAAvut8QwZLSlD2uL0bqbAXzQd+WHdc3r8bWH4+PtnApsW9K97
svP6Nk1FqCzPeriIwmLtJjmvNhdVs8JjQx9yg77rXmMOSNNmNhaM8Gpx0sg1Goxv
78o0j555wQnCQwhUb+uM3Qd5EK471mfkfe6UTGf7fzBZzA5nFufo5wRUM3gRrSi1
MRigGC+0qwitO4vIAQacDuan7rVHz75BqYOcsSfsvgO3i4iiCwP9+wJVCPsUKYql
pw8BVJfMlrd+fqzgapOoL7jbB8asmMbHPsf4XH2Ra2NzO7aL4fbZP1x35iu+qdJL
ViJ8rrkrenl4/fNft1gUbEBtzhJ2SlzBZ8j9c+PYN73Dg3z+kVXzLaAHXvTF/LDG
6A9MOQ9OLvbM4mHZn1iyQxdFlt7Iz7YDGSv5GlVHicbDBwYVfegMbSUJ9KXnu32K
pKqnQgp3oeEVLHguqEJ9PM0oNqgMSpWchNcQ5I+qVRRK+kD7qcxZZ9idLL8XMStE
0RU0W80XxqJOsJGNHUAMGuFWdnxQY2kRw6XuWp0SR600pVgVxcbBviwZ1yJIp9fz
2w6M/NxtKvSygS4eb49YZ+rGA6u3a1/0eJpuGwRg2gdWN15Xbn0XLfitWW2lniV/
iyat0EWuO1Gjw0S3UiV3sQavKsDZVCTVc+FhUz/KAU0WHFtGZGpqonq/mAhIPVMd
mLEZQHVK3fzc3vW0CxfPpEncSpLrS4C6vj3jEh16SHiDH/qsfVI8O+QZfgtJPkGE
knkE9fhhUAc9g/Vkfv0XosHL3AkTDCgs+AX+pa2cF/15Zh70sq9dFNRhT65HCBwn
xZ9FeikJJqWsK9wslDEJXfkc5yDukjW2MEIr1t5X+NvKT4HmfDde/qNmAj6U6Ch9
Gqmmx1YhfHrCLcKlEJl9oR5W2q662aDAPQTzQT1hhoaj5WM0xXCOlppB5DThh5Y2
i+9wtrB0ubBo1OJIz5Z07PhEoXc8OXSy7+4/MAjrKqB5PyiRBsk/Hc1lzU1EhArz
UG41KdJb01O+9fZD04noSVT8Ro8dwdaxYTpCncji7+cFER9hsN5uZoBNl4zI6wW3
Aah/QLDs66Kxqh9N7VydYF3O85t4553ZBi2ElRPUNK/VgKYMgOZ75JKkakJSIUSp
eC0WoixubI/VxbN0sDGhRWZWahmNw3RAwG+x+MFy2hxx4V5WFlbai4Vr8caHnGvl
jdggEpnq641YYcWY+KKxuTkxhYDNUl7Kltx+4q9PJBjY0alJuLibs/v2x3EO1hRY
ho+/xc9K4h7+/MsDr4NNkkXTSsxQ59RptGi2E8FTTI3EZU9mLlDhjyqfmKV7casK
AxTfjn7NFWJKLzYj2/2+1bBm8+PmY6vuJm5hjL3Dtp9BLNzGcHrL3el/GNmj2Ojd
cv6glPuL8y51ANJ1uEZexbY4KgPN7mcTCb4NHrW1ZjBJTCQfdt/Ia1hmfggO7Ym3
D4cLv5iByclD9+Arcv+chxH5/9P1xgXYkzOBQ5cxReohnhoZJTNcu36W5RkQH5DD
HYkfX2R6TI6amGFc301CvqN6EmVTxovgf7CPSnRPZxV596u3gpCZNm3sEkdMbxHS
dF3nckoxLCJP8JenkSzI5OqFsggUkJa1elzqxUKFZ4jN1DgM9VgYR8a08d6SYcSW
aJFY82XS1/YgFZM9Y4VZeCUxpujipAfDe+2MJU5IHAiuves+CGaik6Uwo5hDEAPG
FfweDqjiOi9CZuKOHiqDUbInSnaATcIa96kK9HU2cmXjD9CEH8ZfQUFCXbaGu2/6
0OEjeGsLxsEygImsNww//NpUn1qSdlk9thjIX1Gai7snsLbKmAyK74K+JFtMl7Ez
m4gdjdbJWVtsdMRH+OGUoDJCxZcrpVMW1TX4Q0DhYJxApk6xpa9oYwrehp3VGL2z
GK7OD7C+C7YyCg0dpQG95QaG17NWaZAGR1/+0qcQfmZ/ZCnYSoapLOijHNkqN6/P
bkRk7eN8f5GiEYjrvVa8RRPMk7AZVfJdHzp/EfHO6ojwDWY2oafZzilm3gt1VID7
M52JIAOWpBM9qAlBU6WRXWk7CaTaOcFABZEowNqgNQFrD2PrN6sleMtf9NvVTMEy
58m4ZdEYJIq0l2LJvLbkBRJ6e2yTDJRnZfN9oZFGWi9/kCvSG8l65j8ghw7lPbwG
gZUAuxsQt9DhylSvJd3YnkKm/1+jkzMPFDByZ3LAXQ2SmKEL1xcmWYLaVOaufdQJ
7FZy69r1Nvs0+g6n1KZlmVVui4EQcEQCsh2BRvkEwi0I8kOXMh6dJbr3X45L9Eg+
Ku6c/xGhrFnMeIgHzlVyavFVMHUTlFhYo2pS4QZ61tr/gzRyJnq2NeZmICyw2kHh
7JwiMlsbpDEs97u4htFNIliM/CBs7thjXFxI3IgGKJHT/DI9ybEfb2vXU1nlpr4C
Ls4vhyrmCGlZZVbiuqqnPNKl+NvLPvmzkQICqAbGNJfkHV3BYmWKrGbTIi4eW5j2
qdKHnKYwSeCkQLh63UW1B0vh9gsl6FrglqwCJFibe6bs5ZWfMoSiytjIW6hJrg51
/6oxdpc1Dk8XvvPiqVP5wDOnKkgznONyHYr75C+lBl0hdLBBTAlqjC8NruSPf73A
y9Neu718NWDzGcz7cI6s8vqjlrfnFCn91YVPeM+zGqVvlXv7rKLswNAQD+6l9o/Q
6BeXZc0Qdz5jdtaW6TO0KL6BqwcG6r/b4lAq5Ifv7wPvFyulZTybvORmQLL+n9+R
LxkNxw9GP8ABN37N/Wr6MLVPZXfzsB92Z5FF6waIvoQhoBELA85UFvGbi8LBiHy0
VWjyvSknd4JeID63g7+RC8T64QNJesOB5n+5PcoNIdHQXZ35ECTmijkGO2hzlU7V
gSqlBXHN7icb4R/7XG4CKisUELXnaIRUJFHRS88XPTLEoCE3LP2diR3N/gdFzd62
ZEv+sY3IngfKMatjnQZ5BIW7C1y4q8ILQx8T0xmLkQ8qkpwLkZ71SGZRAhmHjijA
j8oaT0jceE1rZ+wXKw84m4h1MXxfVpd3vxVfOQDIc6wAzIYmUTHJlXc1U/yw7xLL
iePiub7NDtGBdb/tLqnfqrPo3rP+q1ye5ZUUd0CE+zV3LTSVAgkytpd55+R8Q8xO
MWImk2uAmWwAa7km/x+iX/3ppWQgqSpkQaFzJwEu/z7C+b5f1aXOst6+iklX5IgH
r2wiNCY/ycUAoZSbnTg5lLkWx2y1KJznbskUDZ4pEN1oK8xeOzSFUQIrn0NZlmK5
0F11EsNc+pNUyMPq1VK6H1GGMF7zzZcPtzD2fZQ32vFTY+DnV/gk9grSopj+kTPG
Uev1MCG8yY+qVC0YhiwqiOVoq0CBHYzSctfyAbFCsNAAi9btvmsMHQLBbtnduxvz
PGhbf4BJS/s15IPKkgJRrgIDfzIfRZs2w3mSjOFwSRd0gbtiPkry3/U45c6oREaf
hB39cFfr+CFbeD2NXdjMXuc8Cs7j/1Tl6ftij38dmS6uoLsi8mW/k8UlezSRdqcU
Xi4y0kHJGqJMeXVtDc+0f/Z58BFjWwIo5kqCnlmC4AUZNrwVd5vkpFemuLphXRAI
gMEU7cNMsDM3CyTT60mcYInKOX5SSZ7ne0u9LdByNlC6TEGQYc0H+JabxwC8+tAO
qYRevG9c6gLyUG8YgPyJIJAJdp2rfCePlBEU2WxSgLX25a9TsDribaLqZRAxsZlc
6voOjguWvgsW3//ltFYkdO7S/5X5/ErJ6ahAiFVdh8aE65PtYRhNRSacIEMkCdr0
PxY83gkvxEydkym9Qex2tOI7g6Nq6Np/Hm6uO6U7VZq6ShQmaSPP2hSZv1O8Qg7q
zpuTmEOjCUI/WF970Np3In9oYlgqjJ7AJ9bggESgBPwKUbqBoWbdfOoXGgqOIyOJ
2A3yl6iFi0fA6tSMdTI7klfQBTTTeIlkIVWHGAzkydxRIAELZLDAyeQv0OhptnTA
yP4zeC/mMnDYE6oeAqU7m1vEA/jOuAxaUzwiWvYwZozYCJspGOLozzyFKrTwWljy
fPqXDnYOeCXqeyJfyJzW8OHH8VXAsyzUWBY7vpQHnfdVVzVebsPbSUJwJR+FKyLl
0v40e84+8dj8JAyZ0H6z47YWfGrtLlFc4YK/tcPcoa+zrymWcq451IU1xlyKAEEe
di95/9n2mu7i5jh/XKEKwKSoUvWUW/qw7pLZDEYWE+3iiM/tMH0WYz/kkAJL20tl
8scZeVXPrsHt+zYh5K3YA+o1nhS7sgFU5/mS2pLGOqyNUxlKo1fwD0t8EV3oVfJi
imNI2tLVYdswdNTD9GA/dQvDLOdgyc526Z06oqpfvX8T9bHnHlesRgKGGaBmPpNo
urm9wmPhD0zEmnBpBl7pPaDqFVikjhuL1rNjW/iRQbb+FBh5F1+mE6lPsFvAnLWg
SdtUeCgIGwbi+ndj2BAgCzO4Nm7TZ03Sn8LgUhvIphBbyAe9XK9qq2NYbMAxKm8L
Rh6aZzXtH3KU33DZ4GX74K7E5BSp4+k7HDz0c1w4D38TQxU+WcodsQudhLiFXyZz
uav5HEBOXYm0fpd6EHLcLuOwNHhRgPzjdO2KVBvNiQtroN4yLr3/sYe1dw5gNNrm
ygr4IEMCW2m++VHyknI8cO9Kl53Y0TjWhynumt8b7m9DBUDRzblAxzZB69t6BIhd
4awMs19lgzDNEx37Ucrv1xYn489IgWbEW4NR0p0AC2jZ4IIye/jBTsWdhDSqFsji
s7M8ZhuF7YT2f8nZwc2279+akATG8wSzA+VWWV9B7FSCb5p92XJ4WBFhI5lCUUzo
uxyuVHoQPqwFvOUU7tsDkraECpC76RsB84pVNJ1pD7A6b3cHXjTzlRyrUjVCl6Jz
3uBlPXJSy3xLdYcU2nIze6rRyaX2fbB8Jxqy1FrFpnSQirFm9zWkR+j8b6h9jGox
jguHrbZt/fLSCe77yyLEt1agSYKMhLPBXl60F/K4TghwzKWdm3qVrN4kiUFtfDvl
uhSA/Hmtqg3L/WUGQueQsK2F1+uxDHNDgKP7A9vjk4zWIg/F2p1G3bKOT+y1FIas
MSI1Kc14R6DBzdNkMYiNcsYmrzIYCwYZqfeQSuUPqYz4YuztYthK3hQ63ZmFayGP
M7xDSRNjwIb8qgrg5WZb98VLYd0pXL9iu6BDYKbQhtk6iCJ4cRznS0vAkRznj/pa
SleaYcO2bjxBoFT6zWBC5GR+JuN3HCstfi6St0p4IBNTP++vxsd8iaFFvre0HU+o
Jr/j6N0ELxQDcAWSOarzKOAXD/T/y6PSTiSNuP0V+6J2YgVcw0CB975rSgEEdmB5
XcrX13qOIYlsCTykVq5SMNsnus6Ia/cHiSi6GVJ7OJHaK5X1AiuaoQiiVTTEjatI
vRWWkg5xc1Kol/heaNACovS6XwonZ279r5X5nzeJFH8ven4SaaycWSRPoiQV43yZ
aOvNnq++CQUaz4MrpTsYxFciCIgsNeBzeLiRT0Ru2Vkiqufqb28tl3G+YTs+qa0g
KSboAHncoxEoCP9m1uS5tNkD1gGjhctLFsiSsHwpS5D4Ajq0+7MHsmBhpKKq1udR
YQ0/gBHL7NjW6onEER8N5zd9EVo+F2BrDuR4OvmzUyrYcOauKvZyOLnXWs1oAYlB
pleSJX5h2KNs45lFxGWZUdnrLd300bYqwdU3Ohq9oqQInByCIs1GEuG8TFCQ6Vxb
03HoaU0bs6x6P1iKPVflj7qa6dBhWZcAT3L7/vUe87mSUIMHsMkQeXuITnUhFKpg
eBzJ053sD2zoRXUfm7hWv3OQJMrauNGhmAD5LKuoZnbGBELpEiLqGQ02shkWy9uh
9ipO7BIXxkghbrcKEovUD21WU+4JxJ8oK6McaDYCYAf5yYREQqKiyfDUyetNYrg+
O8xoxuYLWMag8qS1k9XL27RDL3/Q/eAt880SmxbEf063jMTP8uenShQQtwpGo3H6
CPji6YiNZ0ExtnWpWGfGAeTWc04q5r3+g6NPSmCPF41xcGKWE2i85fd6E1IWGd5p
xXyUC0Utuc60snaYJrnJNW1n3lMiyQvmyS0O5ZFeuQXMUIHQ4KcW+88UX9D+rzqK
nx3b8kWU74uqopnyGLR6/sjzzFlJQ7nguo7ymSWaGCzSEcNLx/RsvB6zALAhzs8n
xNqREl4kKWXjk8hgEe01ASAB1sxvAj2B83ZswVSyNqaOCsNtex1X7ALafYNEnBuV
+Mj6ARzRyjmzJwadNQ79TyDWF8R2YDNtRr2zqRt0qIqVorkQiQSsFD7e0Mum34pb
2vdT5/zTFQe7xi4dZx+Ui7Vnqeec3hwds+Aa5EH5wNxLdOdysWi5+OKQecTAKzyu
s6VITjbR0KbKX9CuK6O8sQDm6sAi/BLDQ+d58DlT0QSBZ0nzH12NMx4oP7UiWwO7
XaLz0Hgo1PBoyC9+234R4VUYjq7uykn8QnQKK45ELtZup6F/W0EJ0LJ3nMlMW0gQ
caxEDtZmU6p49fJKf+0U4Bi0E09wBPfika4isB95JH1p0KAnHPx/+zKIfYV8vjBO
ZtUG9X+ZrPwkG943uOmdJC5PH8HrT9dAweQdyoDyQCOUiIbXypVLtdoK9WXz/r1c
3jxkgSDGtkR5ZBrSbLgXz2Koc9kMqzmmcOZocdCSCOlnALzhv3qTA68tuNJel87Z
8cq4LqJLYDzg7+AT3xEU0bVgIG6DN6cWAu2DwMyZo34eO5oU/N4epZF1jOIcpMbQ
ZQ1rZ3i0buf/dIKw4pdd8B9P12tCoyxxxT99Wo7s9vj/Wug2oTELNryE2MkFeKlj
v+Vm+8bYkk3L3rErtSYCHZvI9/y23njqK+kAndhiDwIAwqLJs9hdy/fVsSEPNiYK
lcWwqGz4DupEyINV08gon07ZIMuaeYDOCRcud5YK98oqLpH3sCxqb39HIjFclWwa
0tXLIKTa16n8edPISd5Ot1jrUwx65zYQHEPsBn/qyxeMmvCpVcGEAwOJNvih5AxH
wAg/dQckTGPlk84jTwejj99hM3Bb680JKq6NCdgKnfEEcnfkgS6JM6L4K9AMqSkp
3cVElJBDswhXyMp2K0UDv7bmkgZjShDzSrfIgOli5NDchHz+dDPxLywit/IdvmUG
ic0ooIkbx1Muh4fJ9sl4Vd+gemIDCPc8kRHXuSEITmGG9J0iduLgjk0hzYrWAd/f
St3oYLGp2P0yq5+muIYBGUdcilVmXn9FIhr1BFwXkPivO0r6k30BpinPXvX48tkk
WTtGWdiu/w/ITGrB8AmLRTIWH+RCC4y3Pm57RcqR3r9QhBkWTNkZMeC5fswFPhPc
6sErpW44kDKrDuW0oqxf5moboYx+kJ/Q+lzvKf3s0yaPom5kHKKbdQzF8bASSdbd
teAR/nPT1S/an+ahZ+pA22ZKFxl29dGzuKW2pGWulK12AzM4jOUBbev/7p9xtt8X
/edwcw/snD4OIQA2E/acuhaBL9LxViATDUUZMQS6TWgFy02im/4wmKJwv6AzMZXU
unFLD7oJU9ENWIupnixE14r48nWOxq1V2CTaf3eO8884SRz9kCrK2wVW/5TWs29V
x0X4yCusbIh5zfEU4YOQo7VfI1tswGSEnmRrCHybwxhCao4s7HhOvmU25vM6JAGn
Key3fd4El6Gb26HQVSAXQWljCsrt1my7KSyeZD8S1Ka1JYlKg54b7QZyfS0bhJvG
pG12iN+KA52kfKTtRaNwWfrejd6TurZ472lW1Vx3QhFVXpCPYDdkOsbvxalj/LWz
UefpMSBdosfT7uTKwAQFq76+V//4UT9MtglFNWyz0jmuHXG/u8kODN/WJnGfCXDy
dPiNaMEuEnnCNyq9ivC5fqOVXXymZwiXPzYyQ2hyolemiJM5SZxgXX9qYvUEkry+
/IEzuWvx7jW+vaF62wm+CJF67fYAchOvYFYuac+4wMIDkx42jiIVgRBJQvc2+7Tz
Yks0U/3J5IhlT15NVCGO34B0AFErxA5Ois2/jZ+51CFWYtkwryZpUWh9tu/vAb9A
5e4emPFZpaBdXLeBswVIUvO5q7qBV3GMQKf4ZJAUbFg+gSOPsnNi24m9WB5xU4pS
8UdNh+gbHGbsolV9HeePniuo4hQdqKt5CxqAj/xFeoRu2TSNxOK1ojXjjoSIOr7T
YkpJM/aLT5UX/Lwuvoz+tCXPQCdbc/kbCosI+9wR0yTIrG6cplr14zE8v/3zBsf2
IT3zO3t4geIxVACUem+iiE5i2zD4A15zj7m+1l9hmxpium86ERE9edf13+SDD99f
rIx818wXQVqSDynBO4lUw6Pan2x2YYR8x8uuuQ/CJ4vHW8HNplKRQ4GT+bM17kFC
Q2DVVKp2lyX2IagwedouXkjDEKLDJmZLJN7QFQN6oD6YbpZ+qytzHmtIu2U9scmk
s81G1jVXtAjAm+0zyQ68RN7pSiBl/3Sf2/3d6rIpmjnSPl7Iz/Rw0mTCIJJv9BRp
eWbM2PCn1jm67jTgztmJs3Y61eyGXoXmSaw3Cxtw3UC9DGJdAeCdSGnCdex6HrKV
0V5EYjDz7Whui0+kpo+ZdBKGFNzX0EFJ7DmGSSnJYdzn+sWFueeT7k8O2evcG8ln
TpYYiFQQ1HnCiJx6J5F+/MHlFU+Wno2Jw03QMMrOA4XEtRYKvbx77nHDtvqW07R+
H9OOmAg724wWDnnEoDfZBwPKH42NZ4nX/xcnDZMI9yUyKufskE7NGXGl3eNJjp3k
/Xmg70a4pNd/C4ah17G17ynbz72gngBKkXtg/EAVGF432Tah6ThBfdgvm8MLXia7
tYv2PzY8e+dBLGsQpmogV8HXYSxKECK4LK/RIhtFqi7EqEEhbhLMRcUZ5qdoH1bC
6y5WwM1YnKZm/h2IfeX8Xu1z2SYOZJSGQJlZjr8oDE6QuXKr3uTjtKQdtRkcZMRe
NsqcWNvRg5OVjPPJWvVpmIoOvyPNBft3+sVDhA2D/Jn98QIGnwb9aIwZL3SeWYRi
lAJ6TYaHLMKIQ5kxHZ/DmvRvP8nQAT9OqPEKYsMVG8C9z5//4Npe0qJLpqM0/La2
m7kkb9KI24rKC/ZBe2/ej5Ec/m+WEiPxCIRBDbt/x4yB0GSLXpBrT4bi7SwycqMy
s+fAzewj7oj7FGzW5mE/zhWTZ9SjceUQ6jDfD1gc0pVWhuluHZmfAyeqc3YgY1Hq
emgz1S37bPo4o9OLpbgGPQbhc5gPkddtwchE+ODe2rTsG7BEvorCrKi/6J6okWDT
XZOkpCQ2Tx7Y72/npXEtReZUtpYLHo4Os9pVqv2As7ein8LUv7aI4mJ6cUdCa9uE
7Vfoypl1uDg1zMS1G7YeljzOSVqf7KucoeK9+ejRWDuImE4uxgzQNcpygF7CdXw3
aiKlaOr/AY2Wc2eF4xF3t3RSWsGhm/oMvXXwEoaPKViLyz5oc1HQoHxlJ84k4Urc
H2Y31DUtbGGmQiljJouf06ClgGBFKjLP6EArO2cTRomeXhL4K6V03Z8qULMhIHsC
jGorjnuwZMuWspBSDhMbVXCL1kwXwtIUWEM1yYR85tFKivAtdrfBxM7JbNB4YaME
9WY9yYLh3mmDvucKU7YsHMEURJ4UAiM2ahrSXwj4VjsF2ZxjLBLIg9PcflqA0vut
tOf3ESBHj7d9WaG1InowfWUqCm0E0X/8x9nCOdSTeg0yAWwykY9V5BG/rtu0393A
duPo3S/UVsQBjXCYisCbBnkb630W8YSEB/MJxTv0JYZbXhvZn2JRMMRzZ+RJI7Mv
RMyEKrOPYYv3E9TNCzd/fEYaGS5L90ZVPp3uRaxf+395K8k5opQEdvfcXhXj7x8+
Wh4E4YPTdSUDMQvIb4KdJ69ZftTbj+rxIbddjE2ucCHOW4cU0+CkQihACKXbcszn
cQuCekqoCDV/Zdw/WTwKBm3RDD6X6KW3uIF4gANi6opvuZS4TQFnFUyivAQFwqHP
WPogqVRWd9bNjsLB68XVG8BTQ4vrD8AGBHme96UlKR6QGDrEq+xKCcEjZ4gpC38j
34PCtlnN3PTfipS1JZiqVWipeLKenReI7AtsRVqdzzcvC6kCRyh040/lnPsMUoSO
FdZP/QoUSVRN+w7NX01/Cjp9NGK6269gCg6ryDH9qfOH23aTAMN2r3LgBhTX818U
JL18QS9t4Rzwzq98VgV26aVNXF8P2Ylt2kaAOPBbK4GT0hs3r/1OaMsGEhczPsqR
a0u6L7ZF/xTNCFjWMSlPhQI+rQEwwwYxaBvvo1BfqKB2YXhNIGfrHUVkWnz077qg
GinDU4JziWqGc77LnVedxO1GGZr4ihZFmBA09XrzGe7/5YMOMl9D2PYXjSWFwMox
Dg2QRSzJHlRZecxdaipznUNU5qQ3ZyL3Oa6WHpNcwJ+H2z6x4s92jAz2WCiF95tF
uld90EEkFgV+Jbl+qb5RB89UtSGDtl54xNoyGy9dn8GKFswn/ABXrWXtSUFOwMP7
oGT9yBnqEAE7eN+Q5qHhSSXfBQfsEKmH4U67qo1G3eRui2qZv7ZBRxG0dKjFRh8b
Ds4v/xGJBS+EYVEeYTZ11MyYvLqYKJk3yJrWGVEZw1gkEH5jgPmZa0HwDnoR26OE
QhA3golsC6m3VN+K1moX4DnruXMMiwfGNQY4w8ydYXafZxWpCiuAsIn83LPLuPnK
ZMFTm33NI755brQOjMIpJsAikTMO1FndevyjfEW6P4wAE44pZBGf/wqyS+JA/K2u
bVGLsMuwY94SSF85YO0XRuzH5C1bddHigLQynr58HNCenVYk8dR5H9zkOqgBQ1cz
Kp0yXcZaC3IjnSPwiA/zz2XTQ4CH6JAwB+ISQGqxnzYVlnT0jaxr/qzHK1Gu2rWj
Q00fi0+OhV/0DT4a63kbYa0dJRCUgTrpbhNmiXC5Ayi81iqzxBsIb5OlKz0v0vQV
OMYqgvo8YjwkphwpnWvRVVifZTL5Cz1l8xUV/hBb1S1WnPbT0+bIzrR4fnwi3GUq
1aO1IKRqr148Qwgp46dFb9z0XZYkT8/0cqdiUnCcpNtoRdx8Qf4OcBU+xoYFlMAs
F+3e5gBX4qvD3ECp1PfiBprj+H8464QM453xf0M++sHnZG9o1v+YWewBnNl7fvLm
WSDyKcJsJc1rWuhWZzu5uQxvzkT0A7frItltdL35aq6a5XMcVFoivO05tBATxfBk
lGw6TrKxcplv05L01OIb89w4m1OsV9ckhulk24w8wYjyRycqSwbtXrzhp6obUDPQ
lXU4BPOF7NLTaSMwmGiAQkSSKztxdnq3r4IOEeg3dK0gwlidXssYToQ0gfIbKwLB
k6OnQlapeenK74Z9OHNpnKUSpN1t9U8CZsT5EM3PewgoLHuhnNc6x+xL1+pLWMAA
MYSpzWu67+l3oJbK0VjYHrvwyJjqaPsMP7Zbw4tLw4BkzFbUiRJCkvvyUlcqOBSB
DKoS+QeEILiu6TU8jJIL58J9tGlicaoEN+YwiOc+cDf7VNVzFVzO7up00t2WqzjS
CgYicjDlZdcu7XFYWXkQAsUcwqdG+XjOO90R9cTKPZiINkKspRpQYLLiY63IxnGv
bxD95tnqbdk1BWtjcjw9bGDubqSB/phnXx9ol4pzs6pAh+k8qTrf8WbB07fP0Ug8
mYRkhN0N/sT4Kl9DjTSfdHXcNE3MgNn3J4J38oDNecgbHqZ0iDycGPBEHaPISfw2
e9HvR+9INSikA+jPf6zcq+F0iUi7QT3429n3nrmauzYQ9F1BnuG+O9mAeZOWMAj5
0uofBWl1A/8w1DXH6oOSaN+PStmcKqsjKNp14oLbr1eQab0g4/ZyHGFb/udPmFsH
rdjZlYjo2zEOMw+Fs6MyWArBIT5DhkImTWqC6S7RbGO76SUV03MyOdBc2dXvVK2+
R76C0Ac4pGseefFZ9DQs7phM9webXYNGtoNutihpP2RNC63tInENNNDd9ZcltFxW
+PmGRqAkBl/AVzA/+PvMzrXaIFSpP+8kej6SPqIOugSeHgyjwGI2S7G94pFSNScg
W5OzjdCVWxQ6NWYmqNpS/lOz3eAbkOqIi5+fvLXuMcCUlnalecDuAeD5XaK5aYew
R9FMbd1mQGC99QYPWA1ekD9AsjsfccD2JhWBxfw1+x7GAxedA+xtohmDVAlBL6ZQ
BRkAHuRVueBOmkinfd3QkV8phZecG3joQpAbJmqDxb6aUACCzgnkeBtWm+Fsi7h6
5kMUrKLulPPAwcCIGyTf+DqP4I0gmn5g5jqYE0zTLn3trJk6PpvprTHIXkhP/eEb
bOrwYEDUyiHJGNyxPEmYSVa3cQfst+wxHgWN7Ouq599l+481qhbvk/FJUYJCMVxw
vPT/C0i9Fw67esHfJFf1ZYRO0NL8F0AgPDg5jpH04pCmk+sddbrWVoC4b9R46FC4
nubnNmApRrXuCLvvo4RVkqFeHweDRnbc3JJizoafWesX1f4i9WOCtt1ksoBhCW2y
WD1e70XeAfSsKNhMcBqM32BcUh175+5mdpRP7QLR48WhudmGEAvciI/UF3ap0aqf
Z7jIAWYiSmz8pbyFjyuZNgYqD8XUwyqnTuFWIKIokJsfVvyvgTE4NXC/qbGwyhfX
xJ91bosSOK7ALQ905qwVvM05oHZqlp3tkc0dIDwlI1lkcs/SsRlPBgllExsoVitV
xygZhnrcXOV/CAnYp4WeMusAAAh2rakayj6A0P7nwBb/pqJkvtzF/GF8oDrrOX4M
v4zM1EkYyGhlF4EhT5ZTDN6Wfa438F/WMvJkJCIkCulVCEbj4bZTw+thDR5T8BYM
mELK5FPtatamVljluJsygjBpvMGqTYR/+L5c3WxFOfB9m7vOGY9do6rk2tRnpxmZ
dO/6zKP1XGhbIxm8DWa9syx8baNoEcDJcIbm0UXVQOjnunU+3vkSntwUeLjaY5eb
tqCBQXR6cQH6zmAJE7g55eQK8taHA0xOT/txI9I6arY+Z+/05Qy0/SqLZiaOVnOw
rBTyQisU5vfL2ywA4cUPtnfD0SgT8HLShlVinb470C751VcnwKYqKhJwiKtNcF9Y
6Q/ES1Mt67bUqxEldz7fbgSFyyjTB1DFiTPCbpwR9RhUeXnk5N63MizFT9A1d9Y9
+ztMkFPCzqWAiDONgASO7LqzbY2xWu+jBTMkFl7EirpYmq8FQmxeNaJfzISz9T0y
ncTDhSQ48Mj7ZeRZjexRCyZHHYFzjtZx7I72AguoINSEY3rzVMn5FJJ1dXVwpIp2
Hpzo0OCTxVO9NuNd4rBNqCQxvJwR5R1/+RDn8kaPT/dk7FAzeUIDJOOkrHVVKZd7
O8k3VwqDt3dFsc63Aj8B3oqTOUpGltg0P+uwKBY1cAX63mu3PyfvJ3CKB+QjQMT8
Yk6nhrJjl2lXXX1U+EltHC4On9d9dulLBi0fVowVYiYWmJQJEIsHZ13sqoyvNfTQ
xv0yP2UoHzPdxnXgvlC9GvBNsUDP5AplY9RZWFEGXFHT61YZ6xT453E0712d9Os0
DN3mWhG97WDLJyI3XOCvqSY78L2OmF4qeNFMZqKVQzPnrytUyoa1gjeW40X30Pgs
S7Qsa/Z2f2VMDXElW98iJf1jBf0qLKT6vyxelh6NPlYaBnqzpzntewqZPspR4C5W
lLIzablbbk/CqNVzNcmFtSHR2glSc3GWZSlfDD9La7XRh8ia5PyLDCaulw3UvuO8
USrKZJ6rATRC5vJ3evRFIRB54MrRMsgYIiuNeOcogxOMXIz4GOQfPE73WjJsmkOG
GA1Etjz+8FTky44RXHDA4qwigZY7oBy4wqwI3fVCL9MhTGpqd54MWeex9i0axV+j
B/SxWV3UYUZirnuUl1QeYSEqD/99YjNWs0VU2TU+rzqNOmA32VUPmr7y7jQ4hpNb
dO4bFiouhk8iYGxiiu3zyDEcRScAlt3IHNYyy4hsLUe+jLl90d4MA+gLcPBj/NjD
Ua48mszS8NwB4pY0L192GmSIW9Ugbl/sQ0Vulabfl57R+wDPVVtNvfK4nIS6NP/+
TFoQn62lCBD80SzRgDWFI//v7yPnaeK8suqlsYgaeszuH36urO26YJhzIVlIW6ZW
7bI8EE6MA6BAj/wwVqm8q1tApmtT8h2Qy0beLUZrxF0l4T6SnsFrXnVKOSY20dTd
1pdpWQ8xiievIvixsLeGfzHR6a1KQJ05jFZsBvMf0t0dMZsacdNmW0T8rzsOvlIl
MiqEbclTL24lkxj9ONBM3wWdFRrXZ6M3wLSS1dZ+Syn+t43lJvCglS42SXnp8Lxg
CVv6pM0XlMeXjspfzLhSAfOl5hk7gAT5e53zEyAW68B4dDzEKgByJ8YacRIUa9Sf
05CuIoR1Jm7oS61LwxfPwjApVfjYunB/h5P+u2HOWZkvdioQ/RS5wIn5Bkn/F9eH
Mlw0Xs13o+sA6ZBnWQQqGqBpfN4XYg/T6p7F0zbiUK87QREXf7u/zcp12ViCeH0p
cmb+FBjLKbHOWihwu4T2v/kYgFJpbGhghfvq9L4kGCO4a2C3gHP+E9nZT1Abr0VE
OARyYOd5TOBI2qNaDQ31jbG6qyg31MGs7NNqzJfISc5NKJDLXvaOFmBeG2EcBShm
vwNHB+rc/5nSG/yFphjkujqwZ8zI81xv4sbsH3ZqySAp5gNbVuqbSRmdkkvFrz2f
eW5UQuu0rObVrj2XA9onh7MGTTOPml06iBiioZ7pVT2YzWCojw4OQS0Bz+ADKLuQ
hqJKUPjNt6vKZNIeCnjUF9z16gWkITwsXXUGCjn1QBpOnyQ56sYxLXACq5qJ7DgP
bWhfpR1s2AdtmGMOupGxh+F5ZNE086kej7lJ4U6X3SXxia+l9SSjKU2tQ4RvnMCm
U0MjY+tbWYBMbDnXa/7n+LUU/7uFM2FenBfvxcirHTTuS+WqdYpFZsbccGNvESTg
9eSQ4O6DvvOH5nhfRSffX3RLM3YHDkCvuMePyiW0jtzGLobQhEVeGaV3y2sQZcUG
BqYT48HWZM01Ki4C+kwKYrcis+IPQTacsAuFMaMQJthcLypvcc84umuDyEplPsCG
IdedAqcjSx12CIcWwKhFCIDLVeemkY9ZUjh5raE7v8rcOfB0yirJpoALRsRKyu1S
FQuB0Amrrn2lYtLd6Rb+YDnChd7dhOvV8pECy3GZk23ObYIKhTlWyMc2u2YtOHZb
80i1ffiioNPdcOhzkC2V7onpe4BW/rTNquP0VO71EiAW9BIEvp9/6CnMPuuM8V3H
cdKMxXhj3QXhxn0Q3hc+UIam9RQTqlVmhNjtg5j2Mnl9TAzn5XqJHqyOJP18Ro9m
dJNzkYN9lQbBRLhCGeOurqlp8flSxIPISEWTlP/GrHBvOWjaiycNa/7hLcNN544A
B9GggLCrCUIWjSCI/uxzrFeC1OZSuhQGbDv1cvTz7ZzW5loxiHaNUjT2mzPynEh6
a67oTIcDOQL+S21rbLFt3+U+PjouaHG+c2+TGXYHwtbj54FnuOpcSSBF/a9LjUxj
xZEoX8pHtT3KmTfw7LEi8oVQNo4JL7KHWgs7SdcUKtLPa/KGM1sUZbw8GMZOFrNT
NUUgAxp45l+Wk67OfqLzOlGGbtTj7xL4Cg0L3npiq4zBGXA5D+W+613ndMGiS7QT
bdeCdJzlkDxZVlL0Kt/R2vmntJilfrCprhEU6LRAtYz3nZz+upX+1U50WP5RM4x2
KCY9OBREZiA7NQlPzUXPLEIBCD2SpCf50aWEts9sGLZ+aiq1t6IZyKk2JTldhyk9
ywkhAGCgKbeL+mKXJja6clsp6sgPphndNgoH29V/M3nuzhIGpLKIPhC8JXdoSpj1
egzxo2Zn/xfQ2ruV5D3/kFRlRgmm/qXW6+QefMwchlCuOi2ydeLHUXE3o8gdVz1s
vZFqg3vZzmOBX6Y4PFb2/7mbzeuH62j/oY5qKTfYoJ991BSxQlXm3na1wAf6luBA
NPCw/hDNR6XgevrqemD41IpO0mggP9pFVa+jsdLcG7E46nGljJcQ7Hlf7qPCtywY
Hw9RCMqDhCIbtaWRp+MVS5aTJH6RMRlFdZmFJlSBTHXhkh89NvT81ZHyH3bmUOf7
GunHU8hbftXlzAkBkzW19UCjpEkNEIhOM9JR2t+ADzxbteHBt7TsoLZJd1lKSVqt
/vyJx538SLHfF/yh6O0daENAVfWsssbxRumajpMQJT2tVDxye4hlz3+ufPKaFhO9
n6Ye5aLtH78FT0g24JpWUIva3l6cjQJ4r8Xy7LoFC2gNYRcsVSASqn+PHqyVjihf
htHSnzz5W6PMAPYyYlTauhcC3wZS3d3qOU0IkPPENh8+sq/CN6/xeVwy5rDgeTEa
1AgFPfDaV9Fden6GZYijEUc8dTHfBdyRa7TrMHoghxswaPUYWVSwMxyCPUcIcUg9
PE0P/EYZa4A3x7giZjqFVIbhamJeBGa6qv8znKyTYUYZ5MFhr/rgTU3x4Kmrk8mb
qU7z5SilE32NhCoDR3qDkc174yTwtyMfSaXkhM6NO6jJBX2Uq1+uRx0H0U+x3Iw/
krSMctmrEepr6+ZwlmqgSvORr6N32PFg4QSAcDKnIC/3WkztRctkel1br8hJUVcI
xBomcdIeoHUqykN8lZAkRYsWQm8Q5uqAQ/ljhhDjM/cLVxGSgQ1wG7ej9i29fS9i
PUX8a2KdPBf640JCS5rNjBKFjdnhfh7zUTQAR7lziQG1GmVt3NZv0bXkDAKBJhKM
j6Qd6LrJsb3ftOY16r6YH4do28HTPLj4oTKDSwwxlG9mygWcHQstU0O1XdUV+Hme
8skNhPRmfAz68T1ul+/QuAByH2l5G4mhMl21g/2qdgAT5mIpjKYHmteAQVbLRPua
6AU34H9hTa7ix3QoP96h/WqQw/w5OWTcnSjKWkfmhIFkzWhtR8/imjMTzd5xuhpK
Hs7Nw+Bk1ZJp3kCJSEpH0ZxgMCR72yHVPH23XaIrFaEKbRpZWwwXWnJYr6VhKCNu
Wi4wakJXQJtkosjfeu7XiQCRVtm8hDd/ZE8mQlSW1agLcZzAqIhggFLPn5g+8X6T
xvFwihFnDot0jLPw/bDLh7Z0XcPwcMFBO9AbyqOk6qTjQxJqm+CWZ/XU2Ku4KLd+
w1pTHL4ExdJpZspdS0zCmuc3tIPqKVqh+XDv8mEVaRH4mxPXvgPlZgwsioafnEIY
q9rzMMi1hNAW7ChUcWN/BJROo2YVgMHoewS94cesZA8YlxwsH6IE6mlgdP9iWjUM
e70YAlowzEfpkSPxLazrxCKvTuP9XbrTnxD5S4b3iSFLX8LeX4p3xbGrOm9hcwn0
yaHvLSFQvTOAnF20uU4kZj65wGixr3fAqrQpH4Lts48f81sFGrHFHCUQWAa/sbro
dNfeOBJq+GhWlh0yV0y5iP7xHifUKRrodCzJTkIvl2tnr6wO98G8bb6/udQIg0KX
guMObhUsycyq8sZ6UrvfGiYR4zWpjITEbbf9cm39jI0Jt9IeR1qiO2ho6UAMl+OO
YkGmIRdhmfOObY9SOi1Th61Z91DRIfuT6zBUmBM0o/8peWL/cX9CzrtLiLlIkqyB
HdDdAsz8uA2KPgGXSzvdrVaiYtqUIeWjl37xEjDTortdZPKIWi1Jq6Gzw3Sghd1O
3kE1qZoUBS4GOtfIDi2NGh6tpgtWQjq5GfyQBSoY1Ov8ASHIROjY9n9H2TnjAJW+
z4c/dF/SETx8BDzRZg52dKhZv5tP1UQ+SsM+v0DiO88Gy5RvfM+Pjg/pMJQkB4P/
Pqk+sm7qlmvk2yFMqX907omOhYPIRmf6T3NzPqFPnRJ44A3j0zy7RBROPJcc7/oe
+vL8l/clp2MXu9tUrDzHtfxeNY9+Q8p+6ky5a7b2+B60/Z9NxolYWR7jqbERivel
H8UQdL1fG178pPAsy++5KjUsm0mAUHQ6fC0xWFULjVE9KuejR7uGTuh5fL190//e
PGVbkh1k9I/kjqUTuvtmQlpiX1ba/91xtO23VBJg3X3JZLESr1Pe34k3vHrUvyB0
z8mT0PPpsz1Ecnt843KYZJahstPk6Bo76zQpKl2ZVteWNFF2nzQfNFpx5nfSHBS8
rUWSLZu0qhOVTmR+gGjAzoGZrUeSsGSHIFrvKaFfyJ/Z1GYyWy0ytbKOFOJfR557
GAt6BRQ5SwsrP3fpTQORyJ72fpwrGdf1wxz8B6mg04o2GSk+aOc4UdRpwsLasE+G
4q1DxrnL/53qlni2w5cGcA/xf+YKLtlc8b/ylSWXz02M8Mcvnx/sOEVnph/A0mbV
g2zxhRNH803/HHhNOwSC8K3+N+O8UQW9w+ZEeWDo9YxM45jlk+DZk5Q8RalK3DBz
vrFL3CxePRVVnCtjE1kkzEpD5Xm1xbAjGFBy6/X0DgPTOQLitlQeEoVyhJ6U0U5p
KSHDfsVxqoh2/h69ruGxFl6v6xmnDPwUg7rcAdz2Fr+DTkIoXNmUbUlhcjdP7I3u
yO7dI9lgx3f+5i5SSbOrvKiQV6HBxugGQ6av2mXUfyRsFUPxfAP3SvtSNfJQ+isL
EoaVddnzG0MFq5SyEAj/KOk/WfiXu7oxjvHUO/P2nNSU09xorpu+PmuPgnKzcRxe
UsXIgmqsvpNx7t+NCc7JEEQ56M3xKMQijAU0vPk0dpByTku3SoUlKkoOkHR7oI8a
59ie4Dgqetm79NDfMpigiIQS0SkOgXA23oPqLDt1XylJb2FBZXeHhQDOsvBRzBt2
svDglCGgthKIoP1SyU7jurnCkCUg0zH6Qt77KODctrxKUSGuElSZ1ysnlaXe9/ZS
k0Z5tG2AaugCD+wRjycZVqYtA2gqP27/JaY98IfceTFaheP9bx2G0Jp7UjfpdLIQ
62meXuQe0CgJm3duKVECgSpXv9OjMIFttXynn6Meatp7QhJ8G1e/TBUqAr++WhfH
QuCTDJNVkfupRmgvSA0pQpP6HOIgWQhpjEllGOWhps/QtppjHMiCqhy+PPy2RWsS
uQ28ErYZS5pqxBHM4zc65fJwAcTG7Rq+xSKif6hDkIZyUuKJMi7SlDkykqQKbfXA
0OPzLOaCUQXFRkkTnQbwl+6FTc3vbydSkErsxpxlzOq5VMK4+3Bi62JB1uzfOFlN
vSi0rym7gal7QeGtsz5CoOvqXxvU32do+bgdNgV8PAWX33kM1+ZOHbsOX7sBApDE
4hMMQ1HZJ3pVUE1xG9cREDZiSaApYnu5+hUWmtHYpO1bTZM6FGZmfEsT0e+fSoyq
bS8Dw//lFg0AgRVJuwWlOZ8qgnv3HWudQ9kNkzjJsjFQoJOsyq7dJLpHZPaho4wW
yQNvqsF7svjztO9gOhJxcM9rW+0yePzMZrdYwncCRLx1kV1prtizy7rR/AZy3ALv
zaokcJkIrKKLvDzP2IAQRm2Vh3ZVq4pIb2I1BM3npJyktf726glqy2M8LBnxwkg9
6AUaB9N0Eisfg8WdUxs0rrRiMz6p+ZDBzeJrEZAGxdLZXxVtIDAQhErxVB54QKGK
mNDQMvl65yLL2HEyakEDPJP7I6wv2VdsUAcktZr8LQ3f7geamjNoyJY0tS50Ui5k
bhEaCKVt19uWzkBXY12OsbpqlabXUJzKcvB3raNephQGIf6VZ4NaMHBIWLKSF/OW
u/ts7hkJ/fiMNjxYK21LZWSriRQLU2h8fiKsjfDjfqlSxRdwLba8hNj5PSl/ReVA
Kd9Q2wzIWzIGaYp5d4EgeywH93RsUw52qMARd033zy1ZTve6dA97EpBRMj45ClHq
yFOvtFoJ9QjfQXGWxo4RP+t9U0wQx4VdZP1i9jNguXLgusy1rGR0WPSzGG89Ru6X
ulAlsJoj0wTnP1Pxlyvs/loP7sKjRy5vgthtCptbeBuMtmxnu4M7/7s0KE72VeOd
zznRINcUGy4SrUL4tT0dzz39QlCSYhqcVi0FfTU8m3PUfujQdNOuo5Rh/mBq4aj1
JM/lOlkkzp4TJscNDpwcsIgxbhLbJrEVa8unIyeIlRBhTJYfPEM11YlApoWxgWn9
I7wIfyb6oFvrQPT8KMzJOMkG2/zozZNC40MM3UTXNODDwGcvzXCDFlK0kDlkiJmT
OoubWFL3OmbgzmQqYzs6hTS00A/T14K4GRqX0ibzJqg9y/uD3rNBJQTX29wqq5Uo
+RetdAzJZbsR8hC3+vKibtVlx7i1KWKwv4q7wMHPL7ERhWbv4RWAZYqwRz4q6p1q
KwoUe9t5+PLFD+rOPZAm+ZuD0gXEP/9m2Cg+q9x9oePzuMCklzDFr9Seek8v5gwo
R6FBvQn3hMSmAYvuDMUqHb4elCEu13nmOCkh94JGrN2XFnPOJnkFb1ZHGEegui7W
BjRkM9ucDLOsTzt5jRAACcC/uYDuzlWdohTmWCRiAUEdno1MB89jvwpgkBjDtuNx
zcRbR+egRS6TM3rf2nS8STMzWlT4hWqdUTBIAWHBRUUmLBP2hGf4PKANCgwnLBdP
eS/HFTNVxCOz29l/IzNuEnS2FRbM3yAPA8iN9Kk1c0SM0vr41cwNSDQ167eegxMl
52rD+FAlJLVfcdMrCabGLp0lpMJ4WTqXhKYhkqSdO0bK4t6U0Ksd30CRc5yNZqaG
UXM1sshZo9GGmNEbpQhJTfzNLXN9se/G/JpjB0/b9e3PW/0Jk/+ZKBrLr81DOpU2
UgSbw5SDR7G2pb8GIzPa/nB+B73jc1A2LzLV1Rb8iY7NOxxiXDclgWY+0griaoSm
gK5yL09KGeXTajJK3FNQjB9E0v7sNmdGhsTaKAWFfGKMOHjsRM6a+ewnlDJZnPrT
RCSeJEE9OeD1N4zb6/+4wyiMH10CkaACskgJSuoy/4ePbxNYixbgECUbbYpBZ1PB
W0cGC9Ei4PKQobW8kGQNJU3X2rpNdsSOnjg9kBjUdmLy2KlkQhQESfd3OJdqa2/o
aTZykp3LcyHwz87iZ7ipqnGLttB3SlH8/oElPTIDeqbeu1u6jfwt5HdbmhQSQ+4X
V8kZTW+076SBuqIjaoNKMXGYq7Rkl+l10Ntshr7xeoaA228Jj8Cgtcvu/axjPeNK
yh5mA/6wI2JgKm7I7DtEQtLkNcr5Eu26ju3qjaH1tOtOEZd6Wq008LHYmuKQfkXj
93g5wN6oYzA/saPAM2bZoVeazGj8zSjppW7VxVpVnIxmaQz1xZySgQETcWXlpwUI
fUrsw31YCi0MqKROprJfaK/IB8+gXmH0JC0cFXjg7Azd+JSjCQKKfCEB+lQkG0Wf
cKvmWR9/W8M/KyT7JIi5gFrN5uOcIAofT+8uqjl5cKAd0qZq64PXvlYJaZnuzVtM
iJftGCGkaOJk3loKdaWLbCo8jVXLBqQPhE9Sk2U8B7R+sF84A17HMbTsQVSsPmM9
XFyNV+NhmtrzUC59AWGG1XS34tX8lC5/YffB8NbgsLwMDjkXliXFV66D8T7+7nHI
nD7aFlXmj2QvQkhw1E80QdXSzyS2iBA7h9ymNbWBRoeMVZtMsLaaMx0JppVij27/
FbLLKfLbfPo9UCKTNSmwIhQ9JiiF5Xb0UYRrMZiGBkZ8jUoKx6MaX1OCWMnrQhlr
4XDeAB6amtwH1SQq6obsSPVS1tXdXsI1wElklVC3ESCg0+XQZFaiuK0KEISmtTYd
qqf1HNiWLbp4RKcmI+nJD1mg6tvJlCFaeMQcOmylHpsChOTEPFTPnwKmEXljpbDX
3wJNMmkuLhRZlvVVZe9Ncc8TLeIP5IXqHvHLx5I3I8nAk5J5g8FER32Cv/8sI6lj
+pQlOL1SnzRQO0SGR8llzB0pGq6zJGSjBplx2DTHLeeGX4h5RyMQzLQvGvuHLJRz
IkXuU5nZ07aPjMNWVSziREI1b7le8gDSAiKHiAJiU7XQ5NzGwtFh0RLOZXZlHd7g
3OHs4fjh9lD8TdqeCYsIKjOWNqpjkODN+TKiDbAFbzLI44v3SoByi91NedTf+ODn
oEil2MAqi29il0kMMN+p2rMIiZ1TRmtnOyiORE9TIKz7/BMaCATXcxqNwsfvQD46
PMM2ugXO8MxPHDwrhiw/vBBNOzgZNi+si1tT2+aaHVQNThPfAfLSQeNqZ9D25320
rFBXit2S2YZ1NXQSg2zt3qKKg/pObHTpZKC1I0rbqps3iuqL8RkMiEmvUs2ITMAq
qcTr7c7EMAVKcluf8nWsH2yu8aNn8KFuffpTF+Rrc9VyoUSU4kwYCSSOl7860l1B
sc6bx83u6ZO+wDZrmpzGQfbhvw6lT+Q9XjPKMCKX0PXet32KwNbg+O0ZWRJeHJfl
ZrmJM81Km7Gi3UgPe/cH5dzB0dfQJmZHGBhkivC5YqubSN0pjaWdlgBVMLKL4Lpg
RaOSkMZ/mU/LzoVs6hv5PH4xGC6AGKwSOPZoSTPYcMq7oOXlLumXlKZlrmehLQld
YuKr8bAG1C6DX5uiJXaIOseri0dOF9WsfQaWE8w+QVgaDzcF/zVG/nU1Xlx6hXOv
Ca2qIyu/DUNfcUUnIyO3M281UD/XkF8f1w9q8WsIsc39IlM2VOc1iObjZ0D3gaOT
h6i2UHx0P5mGKsJS0TOFm+me5R9Wclbjdln/gTExniIzZSXjk1jPvOcZOrcpss8Y
A0UoZqDkfxGk/gTHg7gW41NKRv2HpqdhLIz3e3YswNZqi7+ZpeEmv+NaRI30CdFg
HAZJCXPUv1JjzhDstYG0NzBXL3I8Zyp3o0NVTjwrp4WeNbM+oSDBxeDNniQONamF
Xpr4W2q1sNaILWwmKf3zHHVvwSSzMTTamliwt7e22pkhy4SiggBpYDAfZcfRyZG+
562McIyQyncYdhMCo30OoRe3e6PBMy9gnumD0WBsoqddrfx0uL1V3W00Ltk07q0b
sdFndjaXFggGHb9qnbVa3izWfb3LQ4uBIUnG5xqP1lKrbS/4pv24omVPQ2ReSnxE
QYRucod7xABg4SdzMZyx+xHnB3tsjmlekROfCWXwscGx8ljjUMI5nVLDEmH2TnvC
BWR8S1SOsmj7I6WQuU++KctyNRcLmPjVOnx0xk2kATL4/yWQ08tZz2gcHt/sKqmV
QKOs/fNLrIoZjmOLMxJydPjdVwWDNseZTVwR0Zb293X0lVpag9pI6Fzt4OsyD1CG
nA1M6slHdfxtBxLcGtalqiHEmevKejzeI4NbRUKea/zEStkXF8nXI2/xOFD3bO0A
ghdF5WUIgrfVY9fsRwFd0YTieNXi3tibGLZroiPmJk5b6FMln3IlSmATOHFkpRnR
97YwZK9hLtcs5inkGhcPY8A95l4tEXhNUYEvF6/74yzENCiX9AYCJhruuXSOOM6U
g6q8m6I3gC9r7tdnbxllg+VzCg4vHQeSbwjGiP3zKj5OmMhnBAbyErjmcONdkZMq
/Tn0xFvbSas+T5f2FqC93BAMBP7+XnjKL2Rkibh4msr5h0cBy0YhVr7r+LMtg/rE
j46OEnCJyuEmIPISpU1UEmsB6c9laMUiUJthkgZk3RxHYLc94GGjQ87Ijh1nyHCm
Fs6f07HFfIIG1E2uMdoXIrkFZrxFu90KFjPhvzI9YieDWsb1EbAzBKKhhMb3nwmJ
f/l4w2sVvRWyHaFu+FouKt2gghtOhUBYPN1lsvTaCgw/hDg/9gkyhwUthi7oDpgE
z11xcvN2a3h9R11LBeEVyjLiHSb+FBSZ2VsHSWfgSFBBq/oHODKOsw7u+aDiYQZV
GuPlYSanv5gAAOYISCiLRmNTO/+0yKeeGZH7e35KqdK1E/dpJ5Q4F4PoEBZyzrDh
aZQOSbmpMfihlJucEEolluchMvI3aKTUS6CAYEbUc0+iGnDrbBgkrnzBxNm8no3e
voaSC7++W+Yk4i3wB/06otbqDs6gI3ARXqkc/jULTp7AAeAPHirkxZ6ggILsg7FW
e49WJvuUwTdrUPjGE8tyUTohQD3stUd41e6zwQXCvXRakyiHQwjaZUMgApALZkHB
euzvCNNVUl3XPaMfzI1xDSqeUWjAtsNs8mabAv7KSBU0Jy7OCs93PO0OKr/mRP1L
vztw829mjDp3ZbdLZ3YGMldoW3TMwkbhJ4rNDfmQH7iZtUaSvcPNWMgJzvJK7JLO
qQNU/hTD9Q+suPqV0KnhjMoJMJPJyilHVoj7qvAHJbiwF9fdGJZ6h/AUWogooItL
SW0Es3dN5vkDX6Zx+WU7cxXD5BQmd9LSomIpxJMX+/6nTH6+TPWTeeKtZBqqFB3S
a8c3zDsnxYyKBIz4amQf7/GF0zV4TZr+APobH/fvG7r31d0LVXjqJDNq3rnsDR2l
LaLRhOv/t9BlPQIA+b+EByNT7mPobKkSPXAvykuGwvhMYwVnE93UGlkl5/Zfnlif
YqQG/ret8T7x3WRzEat0UVVCJCHtKQ7czJQT7DGOTQcnx0Ec5uIpqr4su/DT7zqU
tJDOyqDlAdnSIfT9RgZn6zJUMIfUwg2Xe63ihWXHUhpnbH8VVeb3SUGHwKVOcgHM
RwZamXrvv3tfwW1JJFq81Or1/0O+CGlutFtsDTdKsLHIT+apzn6pRelSkOpbUbJb
91Mv9ftDDIKobRO4I4xCxOTNeDIe3GdA+bx4NFgI0HaF7LoDRZeSuabiZZ2rAcwM
h/9kH9W5fvKKDQFb0kU4hshzXvT+WS2KJCN1DHk0dRfwFIEBTX5l4yBjkjoZ6vRV
PKV48eGbjwDwjrD17NPUpHODJS5yLEQUkPDkT4OC8amnQGYbmNbxcsTDLW0cuwOX
uebo6HyLUbk6ka3IB50hyrdT0yPOwCirAxgzfgcykbRSQRfKSGYCYGVva8Jlwy/J
ZZIf25OeAPxOxF5s91LoI3BEUOhDRhig9teHVVoyR5cMLwVzGs+XGw87xHhMxL9R
DG7Fs1NY2BND1Dzt6B43W4Fp0SZ3mks7JvPKc5qLtTA+NsuX9FJIrn8xuhlMjJ+w
QyUb5JYFxNflWVl1+c1ayZo/6fa9Tu24VB86UgSeDv1znoc0YJMULhicmxax4BS3
tpJ4U2zwpBqhXBD9PR6rwaXge2DQZv3Tkhu9lfl+kNvTKBqdBDoCAgAniDvGif5F
WKeyrx1TpcyMS7iaUuD0mHNxK/qXpeHUKy3wMzfGrxs68tMXqCIjaCJsBuVo8iMk
YFnnyKf1wUT8HV7MUp0vQNpLKEBNpfPdx9EtHbRUeo3CcPvnUIzQzisUeBn7VfcZ
71irYPw3Ig7GLGZouTWGIN1V5NHRMji7jgIHDlJKrk4YxfkRXISZJAXzCZ5RM+xH
iRE6rn1IxE77m5QQMjVnvG8MomnDgoSMxSry0WGPkxo6Nn/em/ZiamDta05jwIRo
/LYh1vCDVMOzSAFMKeP3vs8tQM2ZKXzUktG0wdBETNGK22ci+tIl7BoitLSvJM7p
iYM07r7r6aN3EKE7Jj4mOffSADvdAFL0XHgCXFY1xrOv+9M/HTLL9Qq5ua0ayvyE
cIeyjpHu9TR7TAtfL2DMBL4tuENMpW52/EwxxpfHdzsrrzpjeYEotW9SgJeqqMUj
n9EOntftcXfpHuKK5E/0JKG+E689novPEwY31vNu/5D10hVMN9Gd4xbHM+m+wzxD
lVrmzeYDDbweEw7P5U8KDPcwt1/LArGKB21E9jwMyj5s4I+8CHfJP7yXdbz9eyPV
JZz6jeWGuKxfIP7VF5JzRYK8ftnTF85UJfri8K1uTlP+XuQsf7rzshVeiLB0kDwL
OL8min61+BaH4BsKng91VH9wuEfcxNPF653xvyDX9KE7+Qmn/ivIYvS4YHAC3xf+
1zPH6svcDwXcdxp+Betbws3zMY3zSg80zcf1r4jKxIk2sT2KOVU9DiqSCo6Q52tL
+RoXc+SGvcB2x/NUAs7GqSShut7tIdMyHksSrSzATtmX4PMo6in/xM+6FsV3GMol
QRGps6IhtfHHziYRWUlekMDtPFls1xbYMhcACNpPh9GDiuApf9GfKpFdEcisgsXe
x0emEx6kcl/1/lmI7HKi1FhqiMFvaRkG2gXLOzqY4vbJp/Ot5OTYM/KbbtUGuMZ0
TG7Ss83WBPzcoqpgO3mzKmj7W1FPkujsQDCos/aqbfvMcsBWt2EHclp9uVYXs8lT
5NlOELE/ZndLsRJ0GJZ4xh/lQXBcAF6UttJRroS4DRxA0R+NzQPKgU4w5VryqbHz
96r977yl1MqK42Gc3wZ47jUloROfBmG2c+P/vqflqC0bij8cNG6ZJXWZvVAzBVvC
PXIzhXz/nRo+bYQX4fKhTc8rM41exx3vfJKKbp/LIm1ZbNosQcTuebzXEim9Lsht
GWwlqnfqtz913iwtKJgq4m8WdGNL4j1HpNmqOt1r/Iazo5NQj3pR8IIKeGCMeRdh
Qk74CGe8LDIOob9htOn4H0TdOzoDDHdI7fNrDTEBQMvGh9FYv8JUr3DH2+LizMce
jdvm2mY/iQoF+Jz6titgkc3ZmpWPiRJpndTo2Wgjbf/+Z95UVWX6MC8Fp8RT4HUS
ov1fV3QzCNUY8NH1ZhNKKnmyv0xH1MAVr0/PPMyjctJvTFyKkU0FEayW6VcRZvp9
bCqQctwKn3ChTu/ZoI4oE8/GDr9teaU8LephcpxOkEy2pG6JUY9bZbf2Nd/aag9k
KHq6K3IWen7bNCso1VF6IjW5pufoF6dBBbaDBSKtfkMUW0PRbMtxGWnWdDeR4cYl
P12rLyYkfPeH93NwuiiBKzWlObEU1t4Rw0x9+u4RNwZlPQjgjmKi5cR82x5XFOcX
WRDxNxa4RYpQcQSoOyzMTXjKvJenijOxYXxWGSCchtaeuC3oV+eu+kIE1MrJ0X8r
9KJyzm1OR/n6oFK8tgO6SqkQaXnMCg2imuTaaq9fudl3FR7VK9iWNKr96o7Ma/tf
nv17pgy82PAl+c/pcMR8qTgMFPlsDVsT+OcV+pUdGD53iXHJ5GRm3kdDnhYZhCPH
wZQTnGKsvDNYg6zONyW0NBqFFj8U1eXNLsS2/GwmawV5d7tZYdQKPSRput1BqRcy
S/ZY+ia7PsKpeWfTVxxk8QUMK5jvPGQECDaSwXPSiQtbWwbz7arv9R9jl9Rl8zyS
D0Noe7VhARojVHzQIreRXX9mtsLEy6Kc4AnNeIRkCHI2qpUwlIq+tiBqSyA1+Ktc
+/a7HZ9M8+z5ln5gIJc5S497U8VsfZG9ktAHrV5gfpmwHgZPC/wvAxWtq6xNyvKs
u+mKeE+q2O3hqCOa5GQaCiNWowkPwqVwrwVKuOSYEoL2mfxNdUMAM1Cnihvcm30G
ela98D2TubQ+81ghg2wybTSqt3YmxEHU6BTl0AA40lw4sjUGe6fF/9cXQy1CYMjs
OYkimqezu3pBno22f8uQ+TL0jAXZm84KUtM2CoPY0/RNvDNdHTFXnNNsrxbV686b
uj9hOA9ZVdmJlC9FswINqoMY7lkzexeK1nnVS5214kchHuoB0LidTkApBw9dZbr5
DL3fauCzB22EnFbcB/lAL/R+k/wxSeYgCYknR7GgnzjjSfgavVLBPvzSQ26Sl4/5
+OOEu/BMkb5HDA1F/lyLd+FjjlNjVsykRpM4cGTH37Ncxjbjf2IdPaMUkAXbLmMI
b0sYjhZXEglo+tPUacDZgsaFhsct3rFB8J0FMJ9ytEn9tDskyOHD0uQuejp7xJ6X
lu5j5AuEc9vkHbdWqSZWOvT2Up4Oa+jYZBk4IyijiG97Xsr9bI4oScLjJNgvsC12
L0/TNdLF3XGrcO9HS95MtbIJ+o8WTV9pCHHsD5nTCbaCMqDZ1UMpWye/mAd5wrLi
t9Voc1JkpjUjWy6B0gaYhYumkT0AS1pjrU+Cy/fU88XAZmxsoLIdyTXmL6LU4CXM
sZGDsDn+n3fxHyafemTeKlNxal97+zOlg8+1M/TrSgOsq3BuBxZW4VM8xa52PHVo
/MWrPRfNf9t3/T7YYHLTqVeMKZIvCRzXNiYDDo+cLdrMg97P8RKRzSkPBj2V0pNn
NqYbK+grjz4VGrve7bdHJfRib1JpdUTDb45+Atv5yY2Ayc8l2gXPBg0RybpNE/Uc
sXtOwQfA8UcoLHixn4dwhxlTDQ0tOitllMbXh/yuqph10VBd0bT8UA31XoO5S8I4
Ff13/Fa4Il3bD280hEWGnN0GleD6LTv3g6dywcTAtCfp9plKl/+xsjkUXhLStBkz
L/uywxksBG2ToQ7ulfFGSg53kVhRIZrLX0jNpciDUYg76H7R/2GFEiBg6iBigy5v
afG1jAUg+l7WDZwm6vkpeTz3FxVMyM1VnG7jWX5e9E2GyJGbjWHeM9PnmoxhTZWp
6Knz9dEsTXkY+/370d8F6F0N3Dj8wMenFPk1B09jFW8gjeVaQwbd14atCMBqnmCL
osR9kYHu7BDEWZHLyYyKyKEMIpoTF5xb1kBvmP7Nv43SBLMMO9AOgkeh1vYCZfVM
hFNOpBj+QFZShfLW9AwIGZw9+8JWaHZYfguywFKeTomobZP3ShSECT2E0teGuctl
kSZLn4ND2p+xTULC7lHlpbHvHEyML8npp2qmuOpN3oNPfTbW3R0Gx2f8DpzMcItK
zSSTmVFDxdMfWV0YwFHyoP6XaW62oY9//mpn1SjVwBCaN91+I9tC9b5+VY2747Wo
M80/924cuhd3TyBHmz4n2ibLJJu/Ltbyv546N1ItyOrXGGkogPiI64xx72TU0Sv9
+OOJUSBMlZb6Xc6SwSwDNk1GVuSYg7NWE0/J5mNKx11cmz/wB22DUshv7zk5HuR0
nawaCyARvFbH/aCcybqkyaZbzVDAqct81C3wh40QZv0T5MxxqzBkAO1jSS/1oRUF
lYV5iTF629cepFE4O6Nu8VKZE21oEz9TnW0Iqu3+OfuuWIf+oyF9mwp1Bsl5KcCi
tev4rbWwZwEl84l0LPPlJ6UpoGNdi4DHLHwIcgJbtLhvsUNRI2MgNrf+Z2yLm92q
Um6ik//mLlX+JpNRmqa3IEoTTE7R8otGohKVS9FwzjLB7OexvZ4MX/ctWb3Kwf1j
0RPp5f0nJ8Ia4BpaMpmLRfOU/F+W71B8FGuopLZvhgDFaOrEKL4pvBtkRLE5bn47
1uDNDMAp3MNzbK9BuGp8dRF1WSQBV7Gojs6uWE60mOliesig5a9Nn4krhn1h7BIR
GCHalHlHJCaLZ4deTMHqNgsUzXy8GOpxE0pRMdCOjntWvUJFyYNMikIXkdczu6ua
XrA4KFCOrYARY1+vzSiFaak0AbtURjX22ALv8MnJjSzvYnREAfPRKJ4OW9IVoolp
o+MsoIuFLS+y4JRJU6s+JYj0TvfhpU/k+Y6ozg4XZF60ZTvNz/3amtZP/P0V+9YK
EVm+6uzF4AJz1wV8vjdyaDAqb2e+efTNKYF78n47zN7o/FJ9sjZR/cOREowYRM/v
3D/2cSy7iLeEh/BQplTXUSLVCl7sKpRnhj4PtU+lg/pamSc0lcW9kXMRqkElgxOt
x+HWRUZoh+WUubK0n/ynLZ6+e5qFgmL8nQPbblr1/b6jNPPR1tJxtD5EHSTkw4yu
7xdElMsbczW9CT/4hUKjsCVac9dr+LAxHhY8nq5fRJsZreVs5YWiYPwLwhnkjqoV
YVWIiXWps3Rn025radbBu7JAOZFcoqlYWNHAZnI34YjMCuCBCsZV/vbgjTKvTvx2
MU5GCjY5xNSqOgjw3wnqJ1yvIyP3lqYxEeaBegCw2F6RQj+PJFTuDUpd7WIkurOH
vJlMMkIsPnY9qbCuuywXTyf6rZ6OxEo4cG0yTfnlt7KNHWYUbmjaSCEMF4lwtrH3
xu7K5AfR8BRyjHE0PBiofQ==
`protect END_PROTECTED