-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Ggi/AeZTDdHfpbqdCK6FrLvt3FlqwPSkNHjIsBWVvTXKCXramFQSJ2fywUibKfHRnhPvBncPX86x
ksr7sMybdQUYWSheJ2VTl7kmBIbaZ7gDVqgLosZHOox5q3TObPYIPC+/626bjrPe7KtTaW2b6cle
efRgrDqJoJIq/d/nFfQCNiDq51L5LOMxPacmX8qtTyEjoetS6oSmyEHH0PLkOTz8BzCKK/3QTVok
ASooTTYpyW2KgJskmBvdZYeXktQyAeXaPLY6U+gMS7SKOD9CKGFArgxQI6KwouGP4chWu808JDiW
vjYEq3klg2yZEAYdDdxt26ZBUQ0qiOqV4StvRQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6000)
`protect data_block
ECjOL0rsQGx/deYOl/FqPWVeBn1w/5zGi1bz3rbfqWDy2u7fpqsgU5Y2OTWj95GO1Ob0Y2ogkVWR
1echp3Ky2BlQbLZ3vlcQ3gJ4QJydeBVdLRPW466mOK46Hgwshxgs2orTvoR8JEPKRJgDCTZWYyIv
6ue8Jht+2Nyd/P9TeX7fgdYg9YHxOVAMnKXvX2aSVljBx+mOUnO8QECR4Abf3aHZU4chhl2osjCd
QjWQV908BxLHFi6upgE/GYxw53w4Nl6zQ/BZIZR9MhbuvL3koGLnB5EBV25yS1lIeDOXRNHE4X7+
iZxemiUg8FcSv8wHVF5qj+siDM7RJZOxhute6Xp5DOXm/16GS36sxIfXbYUw4Vz6BEBfD0smP4Fv
WzhsaqIwOswE68a9drMPRWfyWRDzWXUNKtF77pn6R9an0mHC4igJcH95NjzDLGkAxF2fr6Xe5DQZ
3ovesCd4Jl93eovMG6jJPa5nzksJ6VQ01Ulw0SYEXu5yzg3mGzcgwiSHbXNR5LGDJUhGgrMC6A9C
tWCqhBNcBlyJnIMU1mSABzHyCt9HvQVMec9duF7CvyEDtXX/NFRAciYV2pfzlh8VerE64kHxvWxe
hakNwh3dxWv93gIQhtTnnPWw8xTaAJwEn0V2OIJelfTk3U1EFAMUQYm+PkzgWa3SQY230lcz1+NI
dG8JMfRPs6VropShtR3vsF8JQ/AGhJ9ggfi1KCT0/SiE/tSKCSUZ7ksqP+Zpk4A8r5QN9bmFkqFZ
BuQwyZJI6cfi4RsezogRXYdintvFrPGfYPXYdesdOzkjyKrmpV5B1dZvJtG2gbJC8v26xTUIy7C6
pS8h8j2wad1crIt5oaDUj+zC0YTtVEIoWggonhYAlExIViYfP7rKOnMq6J/VCcpRaT6IkBDQDL4i
mMJMZnpQMoRdsPBNmqPWUjR+0o3P/fufXH4+Jbeknzam09ZxW0XJDf8yGsPeMI5uFVKInBh26oEg
+ozUraVrdinQogqKwJqka7zKtDyZPlWoxGogohOu+t5Iunsw/BLfuHSBMXf5V4oTaAUteFQEbZiW
V+tSsFewOMOJfbFBDwL3Xgi7Q91kWTiMVDbzpCl5tg0en2K5sS9n2Pkl4/SPGpRD6jAPCB6fUbDI
iRgj1EL1vo1ddvt9yvWCu9drbFrHr7RQiyMD2nUmsHinSsXYBrowdkM7wl/GqlT/Tz3edZjBtHE4
gPtIE9aQS4qhywTT8DcMnn//Gf82NW+jcXmq95abmpz+kdlwB4Fs2/SrR7VaOh7CvmdA852vrQFU
P6UWXp+qTJWkq84+zgLWD9tpX9J1VR5cKc9QSy4PbgCdAYVA7zOHuHPW/9LT2GiYfMx4f3go7M29
tpAU68CCuBDrhzAdQT7/wytmQQQlRnwDbn1YUI9OOk/wlCSHVMPBTVOfRq++G3u+UomutW9vmL/b
CLgLLMYHeRhgtWb/rp5BQ4Fw6TSbiYCUY1zi/ijAn/4lWTpWWIZh6ONwN+J6ms5Nkb/K6/17p64J
Q6MuP3mxzjHDBRrYxTwRkSSYeL6KjEx/T6iZ3IrQDx/U38u11dvju4ePFpLKHLmtVkp/+1/C/mQQ
3jeEZOWj2lAB1EqTqpGz+Mu1dOD+G8fNO/KfaIDc69/ybWhIQjYtBEnDvZI2eLo4w68ekq9XNZLF
h1FbiiPf5I3v8v078ZsOoTFE6FsKVZM8PjnXR8SfvMJlXiaJvlw6+ExRCjhqz3C5h1nvogxr6LS0
cNCaVW7ThhUEwJh2iqDRqVUChWCe5e11X++0SOan5QCSMyOt6jpUAqduqBSBc3ijgxp1wGKhFQxA
Zl3++EMK300PoQuvLR+AsDYr265a8Rp11sFolsnRz68fVt8zaDOyL3gWsrP/RjEmObyB1uThoVNr
J/CUdPVjfxzbJhvcCOueXXrvidhSL1qo1W8w7FaPexT3rUzLNYUxcW/d02EPXh0YQgxH7LrO31hK
b/FsWqCGo8Np5P18ONVeF4NUwQYgYeflWWQrHGfUcnsulU6rLakKr7jL8UzpGEJsye+v//2GVI2w
16KUjcR1kXpM1Pg6SrDMdPM+MnZ5DflWAY0OxQAFyOZ7SHLT3dd20EYhbm10yApoIKQvgdsdiPuO
QdhOlUqVHXVqpMuyhY+HrTIyYxL6q3vct/K2bLDQrHMVmMHjzSSj0F8qlxduiuq7N02DvDq6vmmI
CIXoq1UM5nsXSTjVAbd1IQqH7zjFquxBMF/J4/21DH8MQD7HhWPbkAS4Ssz8VJPJvHhj2Wgg2iZF
u5bZ+aby0LkqS9EsfPavjQwZ2AX2Ld4cPVGiTvq6xK8TPqMxW/UIvGavs582P08KM6D1futiP05D
uvTbGw3fYE+svZl5lHFo8mCkthGsHZ5ikP3eH5piaB5yOWxfr7aV8VxNeeqEvnQuV71Bb01hVck6
ZXpG7jGFd8hs46DfznmUSZDrsPBbgsy2CfRkk1XvQbrvanr24pUzWrbVBxlfFgopFOh0tgUMZ586
q7Wrne/Rc23jbI/9Bok9t7PGDOQFx2tCajeQFL1FWFzQloAM4uhThqosy4H/8oZE3Jf1SSJ5/tsu
eNPT50qQW9eKbZefG48ztTT8Qcl4Nhq5Sm5RcFWEu+hBvBU//oN5aIwvVl+r6u0fLu1tojocp+dv
BYR3FHMmxkFp3M1GFmZeEW8dEYFJhSbvNDkjQKIcSnF2DQ1eLva9a9owt9RHcNsf4fD6nctzpUc+
1MmVvU76/I5BgyeIPrxlph1Ico7kMlnSRaaPbRmBx5lmU0QRdPLeus9M/XrE/cYZGN64x8nKtRzn
lKOiQ0MTx4cH4ecKe5m6E31dBN2SlkACMzlwC6zRJ+izIEY/GWjRsaK/BY8cpQ5uFpnKn4WzDra+
ptEIl9VsXvCPXE8eIc6QBikT5t3AnyO3XeljAu0IKR4bcgyPflnZpnl74FRkJKSggFKZRCZwKwKy
olTKe14h2/biZkViQFmB897dqi4knvkE+aeZhJQD+om3Ui7O6bw2/Xot7dW+MZ0449PTbFr8/8Ts
EGI72CUNLhTbXzNd+quaiOsD/2/LU55BTTXmAOSEgvfn6NqdgPPEt2z2/xBECUa3i6pKfoEw+XUq
PczY7WhSkNTKlAw+cmwhhDgPw0fPG2X1PxazyGFndIe3R5kDVTAFKEtLwZPEg8LNDY7yopGZf8/W
SMkip4GMIumQHhtiRZLuPzZWVxbcjGwof0pCDnd98B5WdqKU99I2mzRP3XNPkbqQQxqeLzL2ry3/
D1pRUUgQYW/MXyyhTlRAbC/JYG84UB8aFEMeqVD7z5xIHtVXM8oX6XNmrGkeZYZbwmIUwNToaJoQ
cElUPQh9W7EPSz/o4TnAd25znwANGC3rQKsPsZfztItil4bQJmwtlhhA2oTp6orseXdRyyajYWzQ
AZbYasGw7axwZTb4xFBS9iDoD3U0S4JbF/ktfn2c+h3Eho2PnR6qNhvxypgRZsOlia49Il3ZByGy
eZMUfhGyY6mKvgE2Z+nCSbGhNU9U62hVydlRzX1ZRgrjQm93KNi41Kw1KoqNNHd1ymyruQcSJQof
GotJBP74VfjkVVeLMdEKUyDqVlgYZjLUOlGESGTMIcxCrLEJmwLozsaVhOcfB2C/c2UV3CypauDg
oA4w9+mNbOVYsbZRUz3m0mUo/OibGzmTjbtrDNkkuod3pzOaUTGx1T8+antVsJfgbUy8xfpdZEgg
5XTVId9pdftiFHOP7lphs8aYtBeufxnsLalTOPm4y9dpFtIiAgN2o4Dd3LdNbi6S1uThd91Toxeo
aKJOhdZA6AghwlpnT038IZs9rZ/OfIG/qx59oO2Q5VLWA/1+FHBcHpJwxpBXcDmQEQBz1q8rBVt1
SHMvxkw6X+7aysMze6hRKAEcJr3VbL5B57mSWacAKtmLQEcfLND/Wz9biTkcr5+3h3ZQv0eoaKDs
UdatOWG3YCFbCrMWQIJ67JB3F49Kqfb/Q89ZTOBZGC18ybxuo1xgxf5unAxQ63rQvJYls38rkp/a
GDgqYSXeH4Xn1Caxeq6HpHeqsOwd+kBBuqVuMEh4ziwk4hln311OclTqhbbVbTU+X0lEcjJbK4XG
lsKo9eJ5evXejDPc+BQxNRUbUqapzbvuMetXViYQ2CYvlE/nF95oRU7VhF7Whdlw07TUeBG3KJiv
DPwkFIYfpFOB7BTBneBXZQyZ/jXWQbjditD25Ic8sds9qI7TuA0tTJJ/KTaLl6Rr8IQHvPyGBc63
vXqhcR5sLYjgxpjNkJi9nm3FjClUKgcIKBOEMRRGeIIml8obFTsQL04CEGsCyTUt/Ifbq28o8Mjs
Hw7cG2MtAQjSZxEnbsyaoahF9+Flk3fx9F4nvL44bdrmbK32J877VEUecmJk26EnAeaQfspP3da5
goeIS1SC+UKzwmt41LAcboRrhBiB77UWQd4BuWWfxKWsSkkS9T3nq1gxLTm92Z+fiMMIeb5R25zq
6NdRAtZD8avpq2skHIh0EFHAIANo/CtI8yxFWMFUXZNUe3dZa5bbwDj1SMT80H75HSBZDMTx2970
BxsgJJB7X1QbPnerZSJYDxvnbeRTo/Y+YEhTRwGZwHlZ8hYscLV9REyyeWgKlEAbGrDgxYIIiEMa
RMZ5mQQ4KumhKlPX2m+J6LZaOjEJMk6Jxpa8OJfsedYTuiSycX+CWHGoIEPCjqgywG81p6ymUgj1
KqnUVF8WYkTYF/Ysl4Qnn7HAnOEXtdc6AuEHQLv+/5tovJQVAWKsn9MIXNU5aqW0d9bQBBKTnGdy
Vx9pmjVwjBJQ2W4hPUfHWO2V6+YBNaaRyHqYQMq6+C9m/Wm1Kww5BvQWwAjtWSP4PZOMzba/NIAO
B3lGRqzPsUsob/W15Qn565/tms9UWMUQLa/ZPjIsLG/pcWYZCdMvySm3F9NDQolhpUh65XnhiMBw
jygR1xDL+9QQk77GGbHLBItZNnileipmo77mFn/f+au85UQapcdL4tj/gwsSW3bNahpw0k0cMUOs
iT0mjnCfEtp9ssc/2tnZsPopKsW25GkPe2d8+ezXRem5PW1OV4wL0sm08ocyj4upVvq2gKp8KJv6
mgo0WshSbDqIN43Ylwt5uXp4dSWxYwVm26MYOJa4X1eIMgYpS5/7n9M6T3/q1BRIe5NXua/CLWgF
GoOVcN7XL3pAJBn5+qFIHepm41kzSbu4CNUE4yovHzp7AhQIvZ/76iBb/dtqoEePWCSdNlamOnBL
8kfGeBtl6s/Quc6E1mL1TeLGCgpWeYACZ2ixZQbOEXGf6Q9ctMzLGVuGD9+T89ATK+hfpMmMmeIf
W03inzZyGGru8smMSuXCXvCTKLHjBCb64+iD6qhPMTXLzt6fzaldqVxfthpgb3pcbR3uQ0BZ/Kpc
kDvRmY2pSZiEnwjdK13Jy869IcPRwHbzNEQxmwyj10E8ESNJq3aSFEeEfW6r0uZWl7Z7QRRsYcwo
I31WcqCD02DGobt/lT9xt9U+3DqRn8wvMmnq5CytskjOflNS5C4NlXG0FI8A3mOMc8KGKkKv5u7W
ZRarhOgGrS5+E7ww5VJsysJqwDy4uU+YcQ7z22evtzI/SuU7khTCgbJHMb1FPc5SKzTfDLn0IYr/
CanQIGXA/h+mK8j0skYj/rMQd4nmdUZT8+dxEWL7+H+MZHG6FSohtdCiC+jMmlbXLoBUpPr0CaFR
oUsNIHKXaLDqBT4kvnLSFQ5kgqvWzkw+u29vltkkldtpr7hU+TMGVXfhDICVWQioHBZunsjMw0ZI
tsntlM7dGQlmKAF9WPgQ+oaY2U3Z06TQhAc9xnHCGVK/F4f7Vo2U9QDbJF7HeDQpbog8H/H1Ew6s
Ap0ohP7nFQfZdXuHAoK+O3EMx/ixeDv7HKvCBuGLTTlFQI36WfCC/z6pHb2w9VVRxknWxiTS1mZ7
Cd0E48f+9IKjmk0HLIdjXIApoo+zT8WPNkBgrNZn5KEschkh9RFnSRtUjfQV8XoKfR05g71wdThx
DnkDWNd4Tyd1Pb2zOwx6cuPlAIJyxbS0rfnfmka9bI6aNhGsjqFAOrwHlADAyrSaibo4Ejv5GQ43
b6XBSr6sHXdkd1PUrkFvtOlpkU4f/qcBhLVC1Y7vs0KYgXNtYrq+MYOQCBTuMQUJ9n25V/wmOfK9
t8TSIt6ztbsDbxyfMWnjJHhf3FzK/0xCSUnLjRY2FXUpJhivljVWDT213YzLx3ZdPV2O33stst5z
o1aZ9sSG2UPE4O6pYahN0HUUrjRuDDyctwmB8iSbQC6TeUPCWMb4U7juU3J+xyleVo+kxx/iGvJt
s06s1Ftj7VX9zdTtBQkKIjCLndH+poPYQilHHi6qFzVEIrYkBgZajy/FTaHdyorxAsfHBZ6tg3jH
+SgOH7T/zdRvwENk9frlWsKb+wBwdVAaapyifylqD5Cnal5MUbaq/yuDmq+W4wUMZdtoThxwVJSU
squVsPDlG+LZHhlnjytS6+sbUMEZJCHLIV7S7NrqLSYXAs5Wkkebuf7ixESTgkeZWeS6FxWc6cso
hBKm6bjt7r8JFNhySY1WXnBIuo9hXRCFQqAUUoz0XC5XCBXNOQuyMqgorGNEFKT0x/NK7Hr0kmaQ
heMOaP8FuqgaEHGD1dVqZZf5k8rnsiR+EHjhWXr3a6rvkPvKgQ19RF+FZ5voZLbIYGevYBqjhgFT
EQK3M6Tz4n/AQzjXKDCSsp1DB2+yl4gpduEq7nHEI/Mhl96HK8Z8R2cIgV84Qiyu5AAKPDCcMVOa
IWHCC+Yvgk+YaQja7v1Y/WzSG6SisDfa1+gyV7eCjN0ff9ScYmTT+R6ykcA6EKRYHNr9/N8VTEhN
VSaNZk61LObspTfnG/WNreJ8B9tPVPkFojClNsZLHZtbcU7SadflxBQzWufn1LPkVf2hix+ZA+26
lSYg5auGSIAkoVPwQ7EdJVjY7N5RvMbXa6MZu5Audw/YUShuWLzUx4MedziJmSI3pK2Rvg94p0ta
04MDbgNpodVuadQ8Piq+ZBN1XCU1uh7qXc3XG6aJDiSvI2y4oZCF9J+19cyp8cXZpIfl/hLlgiXy
r4hOudo7hLHiRoAJoUWiDRPIJlcW8wJilGYFH0QSeTZdujHLlV8DlI10VWn1ZEZ6Spp+JDcDpMAo
KUMZoZUcKsixbF9d/drjGhrvIs0YIUTnUAKRTnGzslidSVZavAyJRx4rd/BO/gBf0dC0V9yBDyDp
yQvOQ5m5j0y4spbrylRD8/xcrCsZNebuKvOQe9wy9dKZGhW7S0gZDizwvAeC+lm0Mwt+rj2ABRkg
IZIdI9j69n1ub8p6FE71VAkTvtmS4dYzuCH8Gc8TqUMGAZYkrlILAcWBKDxkbkUHVdyJvlZ2OI9R
hOrfAUOfXa6mUAxxaVAOlrgVfg/A8HgdJCdWP32OYeGVSQsvhk3F2zdmm33GMRiuYNnNExrJkMH7
WnAztQxHbMOYKPX5o/zn7q4fwS3De6fBxyOxubz25nj4oR3xG/qd167wv8viZ1ECjb7qY30zaSjv
d4BW3ZIFPkLsIy7/WJo3S6QDnvCOWdIc30WF2u8bH4RhE67F3y8w6WnoePo6JGKtI2VLbVFkEf+u
zoBZmbHKvG60MO09gX8XBiaa/PCLkiHhYQeQ958fO+Um9tTtbeouaF/KYgJQT6MtjNS3Ys/ghD08
+X2aX1MAYfr4uQbbd9JXmxTVcnQblhHgzAstMDca4en4Rr+JummRjxjAhlqwy15NQfwcud+d0J9e
9CAI/r7pHpEEi+r04I6FibErJQAR2U8hHmG+EFa216bluf5KaK+bHuwYmEvHum672aUFJfhNJZlY
Sifqkstc8tIRJzUeWvWOx1+1L0MsExTY9bDVUTo6gFkQBpK86Agmas5td+BFnnGIRpHyonCKKL4c
HpWeLKXvvsvyo3EsAv0yUdAQHZe+U5ZvmxE9kdSXTok9OxueMLarfjN7MiJONiJVagLK8gt9+EfY
GBDkr4xoD1p8FPBSnvZF
`protect end_protected
