-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
YZEzi9uUlokqAXwT/4lVwfJbDShsQ9xCIlcE5zs7t1z/DwRAb3WcjeeW6hnLbjDy
+DHebWS1H4MsZslHw+6b9dibSEUoouqxq58YRsrhb/Eq6AjjhPHu8MCrz0sDJTVj
vx91dWVkd46Tr9Jhgn8b9mHjPG6CwabrNJMgn2Typ4E=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5991)

`protect DATA_BLOCK
NKi6M2NyrvQ9aYwLDcOLByhsoLcPxNGAGcTjE+Mbv5Gt5EfPlIQJBIocpfhVgSiK
xF1EOZ9FcvUih4Pu8kAwRawNHHvKylYJvBaq6GLtSedAvAdgK3HafF5VXkOoHN0Y
Vo+nzOuDoqFNVStFpLNilKvrdoKBmTDXdyi+3aGGXk1aONjhB9+EWhBJ4MCMA5L6
wR9CxuGdXCQgJij2jP2nZkQLbH3UuJYf7TWRXONiBrwA33YSzP6b0Y7Wd2lX7UHk
lRlTBrNNNbECK327kHN9B2snwmfij8IoexsxzBZOEAlUyhd/MuM9ErpGgpaHa5Qy
AJNfYvJSME1WSRGt8ohWSs6VOBIUUvIOe35JUiae28r/Me8ny6pn+O5JIKOhDMBt
6mzaxoQgKcO1z/dEL/vdc0nuIbCqAyewUzppByGgvALbaoS5AW2bLlpMHyr4/Vyl
1ecK8Tmjr1i+E521hCsIp28pluRKpsng7ZkEHUB5BWM7WsJwyj2spp2BSNw4XZg8
+Hj/t3ckCXcEYUi67vYx5tDopBbXutgPJIbrzCPCmiwX/QNCGV91AdTx40FwXNc1
gEpORHt/RZ6ZgtmGdGlrOu0NK6+ecLjGeiH/9DwlijZrFuqzMQihbITgyzaPGtGi
F+TMQC5/TwHyEYccOwEs/I9iG1x1/thnJK6dUVU5XfjEEZChRFck43ZZ0OecTvUF
rT+7MYCkWp40RALDgWOsEjvVq0uvvHv5QxCCCRmU6w7Jj7vtbxuZ0g9BDQlnBpkn
N2yPovMZ0k6yr8cT8Dv0UlBVgcnOb9hIUisMWkKmsaqHG3hEc7Dj6o2R7CqtfGwN
dLEd/sdXvLkfkhms88v5kKqrJanzDHHJ+A6obyWgF7eVdrDf9+hpQONNc42P6V1p
Tkv+t8kdsYXlHpXPaHT8zgUMDmo2BxzKJe4o/PmgFIaLeMN0NcLBEqkgUOuUmn2b
nSj40rY7sIi4P9KdaxdE5qU9dZNC2dBpUDHT+OwLBI73XhngRDcSuEmzE9R6CiMC
Laa97x6VLauLD+DV1+DifiPp9k4+y/EN0yNywNwf6CvtaGVuQDoHWMWUFksZZFIb
rRnYdG6BLP2hkX48Tm7T1Wt37HfNQqw5wFYcloy0MW52FEYr0Aw0DZS+7SJH2HjX
pq4ovpJtKUIsqUCE5rt4oDpAUgIq9jEdsbDn2g4oEYlrCzof2kOje1KdBlJxVFL4
gnupEPcaORWFrzxLGPnRUoArKr9FfTzn5jbWmdG6rcNbVSxEHKCUEi7QBLNAQoWh
129o97w+zCbt2LzG0YVuWLaik3N98EszHTmYx0pp1f8cnKv7xEOt0r+VRwBtYKCc
u5ecAqkML7VQTTjnDUYCKqs5PFRaOO1y2usa6E0nA2kjUbJWXGTEcG4fHDdRkCnB
mB3GXbJc4zVPacxlqLjtcbU7s2AOt1D3z9JaBCh0Ze2sanIUqzPsasOlDLww6AkW
Pjwq9Szp8zv2tg+vS7zIW7LFGYSrXfuDOCbHBe/dgmfDorJi1Vnf7kB4D+zsv3YC
afR2RAZ9R5Kg6GAEpwSZ/ycrjc7jbP3s6i6S/2zxpvoPGvEB32QN4ivGQ7NrfHcB
KFxT+JQp49skwWwOLrLVUr3adwSIO/Q/QAmtZoFHiaoL9eWVLm4jYzrar5FcdamA
Z8xji7kXV7YXHY2V2NQwezZsyGHuAkvkXMUwJGTldeM69FOvYz3yzjA85MYsb88N
m8bL3v6FGZXPjsn/xPj2jF3KsOI0ZizPkGVkiAxHB0zodJVPyznidE8R/5IBwBAx
cCQrbXAQPN7xW+ZnHw5gWgFfdOmRIV7NFze6AOIgsVJZIq/BYiYFYTCniP+c4B2F
hpAfhYiCowSU/JtIPv3VN1a649fGCmcgZf99oVdY/QqYW45B0/ZB/725wHRDuca8
nfKrLz4oMgQ3ThWRA9DAb1FC/tPMYAaHq5fRlmSXMv5sXecbenVkowP5FFUm+TLG
jRcaVpHjc0XpJoduGwrzvCf719k5IQ8hDNe3UYL53u/7t++YujRtBqg+WzczwVxH
NQ2RdrVDVi2rXT8Yxz+/77b2hbF8JsbCc2fPPKhYfXIiYpM2QeZsuWsnqqRmcNx0
shp4rz9AefTY5I3KmrEoC1yfnSuj+POmz7p91pJJlgMuju2nvPDq7j+DjdiMLMCL
omDILLME1Ch2nY6Y06xwdVZ5IdwOJ8i4nyD/LU4CaC2ollG4pT0HWR2kc8C4SBTp
vCwowN9NO23yFGn+m3wjgFgLoemwFV3mgH6507KVTD+pEq2xhNXDG2F1jn2vYluX
7MVmP35aWsf4/2aggcpJaX3DxwGOUbyYZ7wB50mH90+k8s+mgrAaUZ44S65OsW7d
uFlUyT5SFIpPX6g2FyPHfU9yuaTecmBqchQl8AEeIqQUxdVuL9WFCtbeAhb3dZvu
YjafK+B5lzghkbld1/22akMEbXuEsuurfFfMCvfjs+r7zkFFsh3cHclmxTxpkCBm
O82PFz6+EpDJ7+nlD+KQwXwdIH+j5xW3/m7/qk6CMq0XvdQ+AxsST4Q5T0jBrvdz
+C0G6IpyJTRtf1ET2MIHIQ0Pew37Di+S5zNc8cpRP4FysizJ/l76Tj24znFRb3BK
1YujifzDLiiBwePpmYNh86TdUCXy3bGaSPdS8pROF7Hanitth/2lLQHjO7V89abK
9agG2weOLRrdg3Ys2c7oqCQiVEF7o8SCyVnKXaaaajsFXXm55C1BNUg6sMAJYwTt
q5pHrxsuVwc147OM18rUcDOaQib2jAWh6Ryk5t2vkxGRbeZJCoyJQJ0BdXDYDa5K
VMZEV7LvKJcPSyjV7E58eC3Q8H8c6EC/RiMHTer/+x+73OMGpLGz4JZxc+U/k1+f
+BrPfspzH0740oCpSqHtWcDoGM19iXe5P2LDPkK0p5O+JkfzTUYXakNUhjv2hS2u
tgwojBZqJZbq2XRFMgbRLf2X3xPV3DEothoSsLcttU6bYKzGq7yv/HOmWkTmKSgB
giIaBHq+3qfXeN4npbMbxlg7WqNlZCe3k9RF1zE4nc6/+94fHoI1Cn/dyLLXEiVP
EvFJD6czPrEnHkSdo+ihQlny48Takx/6lviJA+bovTsPi6bMzA56D6+IlmKJUlKs
5iBhpYZVt9eS5nYkhKiwGTjkKtpAFDR1m/vRRlRRCsaC5k+yoMgAiGIGC9El4FKx
Hu6xRboUCZcSYBGNexgjuMhE5R9Zz2v6ruWPaq/5n35RlqTPO2MK5GV+BqurCR8I
djGlYZuHKHJNrTPrMGffJx6lZGK/vLmJDOg0IIfm9ecDRjmJEkeoQ74rY1r0PEKh
Pwei8Nbt8dxrQA8+Z29U8UnEIzFRgAyl8Lu03mCqtuMgdrmpRk/zMM8TJME29/7q
oIRUpBfkt6jzYZR73Ffq7YM3qhI3/0DeGez2D7Qk3F6ancMRVodmA/kZeAxw11SE
n9m8XgNr2NGLSvPCodcv/LLFnxpi/FLInRGtOVPo0ZWEiGoq0uQB3aknu8rlUBGd
sQvLkn0oHHbn7LmI6ef9YS8s5NWG/SdJzZOP67Q6JEihOXG9Nc6zsudpZXkwukdO
XD4mmAbovfRHR7QAknJpXYd17Gr0XI3bKHqB/h0tuppC/R0IQQHg5c//BQdjBv8c
36eVt1vKM/7q91Xjf81TPG+6XaKlTn135zxnJPvEp+BLi6GSf6hLUHY1oDhujvmi
JVgYjNs5uPraVvo8RGG74v/tagE/Em6CTERHr0//9WLtVneO0d8r+NPcjFIDAtN+
mAvBEy1lVvL73/tEPg0lN8DIYfXOZL+pMTtSxpFBh3SO5bzNf+zpQDS2BQxDEuZe
PLRrfEp6In6io1jPMg9lpjCIkvll440o5+n3NjeicXuTJrb1YBrXOf+CltFeEBtM
8iq3hZIAvpMF1skYAm1CPo95IlPt474mbIYyIgIzWCOK4rMhUsbvU6E5ShzxAXL6
0UWiBL5quBJsMbaFQUf2+492fJdR59+apHO7soxZIH+zjxzcDZ9acthUCanL6yTs
//iBXu5uUQFDJUjI7v5riqPnLOgl8zJnANGBZJfFUTDPn23zuDWjmnvuqya3rXyD
KvIV5gCZxsWl7toWbt103pN/Dw8BbMU1rIubF9dr2T9gqrGk77b6iIBkLmgCfXCs
/zfeVrdcWsyFmCaJ+ohCwP/KRHRbwMiveDt9bYbVwKbKP1lvmwi0tSeyJqZC2i+B
nTt90cee6LeWlKNY9Zd/V3fh2fubSsBIwjnwfOdclwgP5NNgb9juW6BRWGLf8Muz
fZgFtfuwgxqnDP10rT+9HXMyTHGIYeVhv7HZZAFngxdGWUhh7HvuuMy1Muvuc2nk
ka1+zlgxKJIgny7toHc8e5Lqh9AIDMDOsR5KDeLSwB6HYZMrlkqt3TEZviJ/GNER
0zdm3G6XhVMlh3GNEl6uuVif3/WlHZkdv2mF7baa2TOKxSFhZNDg1B4wZK5RE3Qe
QdVaR+8LovRukfRl6FhAsJU2fQp10fQG3wtJm1otEvacT6OsCoumo6pBGeq48WiE
nYdTnOLVMJB9JAGqzhRV3PkAICzccGwY8d+KSX/uuTYhTFV5FhceLq5maOHlyzoA
OjI8xVl2YVSAhKUoQRFk9QGau9cUDxt1aRGkJcE9S1ebC7BKSJUzVQ34EKDE+f/H
JxzGLERcJqSyJH9LoWNyg0PzLBC8MTT1QCK7T62TV5fHwbeyf2o3cvFQ8pJVvB55
CJHkbrm8D6FqO4UA8n4wP5zomIw5IAjh0/U2bXzfrfnKRpaFIybJ0GiD3DS3vsYT
x2rT/Tc5HSDfiWwsOMmqGsHsPFqqd/xMarhtANx7mcY9PuttKPXyKiwvdgqnNqy4
izTA3e0MhAcRV5Mw1MpZkyDv4sdpRHvpOlsJD6I5P/vaA4PhJALD8lTLOiCr3Ks5
+NMl89DqD/yJ+QiVr4eSdK6J7Etf9rAUa7i4s12t64ChNJO2US5afSgcK5xOdUsG
H7P33DZ38FpFzCZtFVxa4Ljy8WZNksG0Cp6Ek/NSH7st31dP0P9zTeNeguaRlR2j
V2rcwWvBcm0ZjA9X2ixjLnS61GacfSOyGYZS/AZVGXPzTliaS6oU5M6MPqy79ucl
I7vrjJ6vzOhzLl2IWtaCtrjTAZ0Z+6UycM2xs4mgwbdYxwbo7+BwPVktKGH9MBD5
7rphc4T8vVkJb5IhlIjbRk2gS7a+romLO+9FnNstSGQqWQqBMSDYHd4rIhoN6EvQ
h7JP/f70o+pysDgSO7k1npyj3BXQoy1f/XnrFamgY6Dy6vSfcdN/4vf1itQPUQyK
X1aOImwRb0HX3szT+VHpuQ8QoagDqoNW4x9QBZF7x3TZALHbIsOnx9EQff2oasLw
aNPoipVkY1tu11cLwu7CBOB1Yk72PfYd/xil3ecslihlhOYD+VvOnnfCjYLyJTwl
VuZ3vOo1udIAQlzfGb9I/riQxykRcYEvEun+4zy1b42QDzYQnbw2BjisbV7zaYVm
FtPViGkYbl7fXFazYm5kIN4YqUEEW7rITzGyR0pwM8B0yR/e2dPpZGFukNksEvub
4BPa+BPfVQ8FQDjeifeAhy+7kX8QAKqTZgC8fsbQ54eVh++xCTim8OvLRkOQrDWp
SQCdXvVlLJVJyfuwzZVqPVkRQhrbbmIddEjbIljLUMotWZSdHmf80kfZ1ZQiR9F9
KEorxVcpWV9OqtNNJPpXHOgYMH/qLSuSJ4PMbRhKRgURlyIb//1NstmsgnETcF65
he0CuVz270PVjuLheMeuHQry3/jrU+j0wbBmgX2N4lGsmg310MoR9F41sVAo2YVt
rY94LeIiGhKmODVeLu1+jzyxIj5FbSEdnxBu/9ivf0tY75aXDS0kJdTvqst6w92u
pljFtyaUAzAxaNN7XiJY8h7BSfO1pFwGTSHe+YUoZ/OAxaykJfPNp74s+wByMvS6
RtaIzN4t3h2/wEtD+hvrC7amhk2RMeRumnDrbEpgRrq4ClGT9wI0rbk7nuD4e+Nu
UpYb0AJGRPl95zmZdLRDszShNeUnwjBKX8Gx0ipP01G/ByLJxiFxKxVg4Zod5DrL
FqDSiZJHyY+7UQNgWXtZvGqwApm3l4lDMtZePnPbBA18TP2jRHKMBwyKPvikTyNb
MsTbf4laVjfeTohMs9yJxxqRNXbeggdT7XbnubF/qezvOZn35dnj7a/4SEgnbpI7
CSH5gn7aHxXX+Ts5DTAFvmwiw2NiXPri/Dyh8QWOm2WLHcNjd93ADFKhwvk7d4s8
GNU2O+xaDHBPBXsUUojAMML9BiSwxde9ftTvQeqknXIQDqJ+TlVivt1cu7iDtB4C
JZYKsMhopUs35hZv/XEWxJMCitwM8GqPnCcUxuhIubDL067qMxkguLwxP7XKYuJG
7bAk7dSpUME3cm+llP1706MKcMPIeDrT0/+41yCKGZMi0t+cIjNnXxCmD4cPtYx1
BCn17WX7vK7SeXHyQtVIFPpRKqZE31rqaKlWNyunmFdm1VYZBrBsGfLA8xqCd0CA
yyJZEUfYTy0xsCnfPjVge7/2gNwaTkYFn/qQLN1vB6LlXogaFfDBY1paKWsbaErP
VemPH4hJ1oWxMm76Zu8BqlVwUKKTBenhoNzz4HD0tuN+7HXwCLBQiQKFHYTYyzVg
dWqOsl9zPjO3DhX1GpL1CCogSYZg+eE+Rmc3GgSCH++5v0tQjdrOy0gS12t7nuun
Ee9x/j7aNHCylZ0AQ9CL5KmQhDKvpgEMwM4W4WoL0ZL4fsDJvMhz4UGo02Y5YQLG
tu5z0s3tMeZTNwuJ9vs0ApfpVDs3crPZ2wkGVRw79aGWYdDgP3lqDQvXDPWi0VfT
DDGZtLT7e4WnMVS2OHzkCrFLFLnV8VUg3tYlGllWPToAgXrXhsSWQc22AzHPjhRj
Et7fr6PpScJuDwj7dkiE6hgsaMBjxeT3KmNEJXzOXPanAJIUCBtQzT0gOdHbg3Uo
stNdDdbowLDPbmif1JYyvV07nmMQfp9DyBREjKtKQZau0U9cGURTSKcE0ZVAlXr9
y5E1f6/yDUQsmPyV/tQWDS7MWkodlWY7pW9aUyjxETyYM40DzX/b1bvmTHQwRFJZ
gKxzb5gZObIe4DoXdmQrE1axaSQjn7Bq+sZmIHxx9l4mP6CGFj0EYGSYCYTYNjbj
oYMXiWEjtP8sLzg9izHRTt6IE5fbEtLv37X5IkBot4AamaIX51mE23ikFBux39eu
WKqvqxnjQCHV0Os89hS/s3QtNFqIYdqpMRF1DewJE5v6ON22OJ9/MxEqr6yJq87V
ohOWIH9rf+uCEfLhztoENqzQZTOkh3ANKseONqPAOLQNRgW2JiumyxL8bNk1V4Zx
Gn6R1z7wY8cigCSE8e3kaoh9HxfsmhgTe0ZSDVvhS9Sd3llxWawMTqpzqJgD1naJ
CWVw28oL07USj+xKrbxO5WVRTeevHf6LFIRNuzo2KK45d4Gu3EpSU4FjqVU9Mylt
qU3v8rSGE3lMbu+IW2LU4dSyCSYELXCnxbU56oRXw4s4Kof9YGezTk4eF7HjeiWn
M/Li6zvpeVCGew0PT7C5EliF4ifr51JLNVq6eM9OyO2ib4fdLz/3brP7YLR/iv8Y
C38nUY2fLx5xHdOa9zOzFmEml0tvBeRlQhwap/7JB/bRPPlPTJZgp9v/ZTUMYw3s
F5+L3sWM0tqOIzRzn0NxgKcsIxFyH/GdvXOSEWPNgWcoV8UMg7agowSgq34omUnm
Sc7GYENyU1Td/213Q6QzR/A476T31Odo3EMZlRSFzC00zk7Lkk9iGUjg45IBHImJ
F2BRDlvziAf2/zAOfG36beMfUnQWXlyt9cRkFyLMCq4ekcSLGdjN2OOYoErEcbZF
mRIoHAY2PoCLOmE31t49hqZjxpxAuB3kCHim+XczPtYY+Eiwv+OPX8ldtJveZq92
XTpv8wa/In9G5elxkhumba76o5WVh3yW1oF3DGmO9u8GBkjJKW2ZDRR8tsIPSVhq
WQwAu0VT6ao8Lh3EIk828w==
`protect END_PROTECTED