-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
bwrmD8m4vuivcbZa3F1eqdw5A2mz2hNY7Az2v8FHEKCngca2NI6qVlV/ZoAPY/oy
7+xgUUQgLCVaVqWwMcDxdw/pJv0uSmGXvjWkjKFKF/Sc6skAe0y8gn/6Nw5zhX+t
1+u8TlcLTJpIgj1D0HjxLfIVtomgR6sfRSoB1B5UHmk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13560)

`protect DATA_BLOCK
e+9QfYgotHYIsYZz24IvmoAlq4RrX1dgVPprticEvdazbkV0a85JPPfQYxFfrGQW
9E+YqPLLhRwxJlD73LKCl+aEm9RJMJicGXh/gIIB+xSKhqH8WT4tj+V95D63wEwp
nl1rncZljtmZLJWVz8T17tu6pH5Dd1TOCmPFGk/zaUqSkOUj/vwZy7flK80D/bK+
026/1ARDCNJJCJTDU5qH4LrdBhNs0Oj+6Ae/Vs8lPneVlXMUD8GvJLCKEmICdYQh
6h3tlHvAcoKyvMnRqX97+RuQ7YvECaV1DHFDLTjp56OKZ0cvqv4S5tN4iUx4h7Yk
7/z/UqR82PHCarRH5tlRFSeOt26GlAIz93074CyfJMHNBv6HbUjKyjftw/l0JrZ5
emp4N7UJmMh/VforiozgL+vsfQfT6lcxHbbFX3mGkBhjJBTz6w+AiPA5CkzRoE87
8Qz0Jhuvwkh2mz0daicGdE6brSsRjMcpWqViLa07fTiwiuv+Et+C9G3rHSRDlbgi
W+R0ApSaUIw50/hI6k75nvpu3coJ/46E8N/4qZEhcNuZssnT+lcyOhqT5JxsqwdP
EeionxaWToNOT1v8+6ufXXMxI/HdlWQ43/mPjkzD1GND4kwpThsLdSTk8tPhsXQs
JMnQoRjqvjB5XjRUGDVqzshrHcNg9PU8VNnZwC5nkvwHWJTTeqUnV4Lxxn9VlxGv
4hc5KjK2Sere0vSqhqJQDe1V00maf3eC63cVGZNWtYUlgRXEDi9Gq6kMT/DyKLc1
RBbKmq/krPvHMM0ZY5kr6hQ/SKKzS85mSPDh5ukG3z87Rw8pEAdnyFpBCMbJnC7x
s3OuCz4NNWP/K2wC+zZblFC/XG5QzfOkMf+u/HOsRuseZt+hR8x7/HAx6ihZ7UhN
/zLQKEKjzcRtNYX4/JfF0UVw8Yqdt6qzzGeQOEg/TI+Nx0z4YY4Wx2TMXg2bUj09
NBcIbk/6LH0rrTSyVqKBFS7ycocf9lezB9df1VhGCjxHvX1tC6TX86a/FQtTN/iv
iY709nVQ+yTA4iXcnu6+OqQVppNKBbsBAi4qERPHDACw7BmG2Bkt2Q4sgUz5G+NJ
3J7HYkhQt4S3QUWchsKdG6+KwMwDRqgxg0OkTU3RywiCUWDQmLgrXy0Gfg5hYN94
hMlCiRUgdBP8DoVwyZOvd02iojxDm9Yl36MEV3J6f2h7INpcdH0rG9LAVw2BePmP
RNl621Ry42Uny/54I1W4N0LRnt4Ng7cqy1XnMdy4DTy1UAMcS60t9+5u/B+dJtk8
XJ6PgFpVXqvGcIHKmrJOekaTfbxkhccCGv3HqRE1K6QbMI1eUBgTG/8JwUroilaC
VPtyGzV8j1ERt+SmXAyTuauEZIPgHMMjCIG1GkR6EKEqnub8VnJLKWdo6xXAzzCO
A5aNphd4u6GwpEcNmBb39etpZ8xGFs1EA/mNJLscuxrStt8pMr1bWK0POuHH+GsE
78ytLmL7JKWMpzWkJbLUWqr4EC0H0w7/7L35BcVkt/Eb7xxsbw6zM+begnumQ59e
Dify1S2lyvkWTxRXAxpp+SAnCvHaHmm6RpJQtYcN+M985YD6uO6jijXrsc/VNI2S
UdN72u9MfSny3a008WKGldkSJf8xGrUGNA0+0dX6dA8Va6D7QDfoKkUF1rxUwLOh
Z2lVbytM3TMgHTS9N0o232c9ZQ+t2WsaO99wmgDal1cE1dCSEhd6L8VEwAql3T3F
wfWKgUI90Rh6HdnMd12mg2cwlT0Og4Ty+SQiJC9dscwjBEM37v5BOXaQHZmZQ23o
TKc4BhQuSTnihnyAFxFVjsywW5bEeW+3hIFwTRX2CgDTkEXxJ61lDnKOzhApMWUT
gPFoH2g7gvnO0v0HQsftwHRYSl/AzR+zFjoRiRXG2AOuI5scgdok++Ii9IbBrirC
RKpVgn85iBa1qgNAKN4nPnfh8/3MQK3OghB9V61SOwB5oBSUHJznU7EnFrVL33nD
ia3dCyjNGCQtVbpUzD5rulccTH/psfUcFouXsuaVRqFKelVU599cNUXqSEQvWnMZ
ntmVVja1fyU1FboUJxqvnQN7tQ4HPBQ2pa8WeO9wgVojK6s1z/zWRXKryONul6GU
IWepYLIkDg5TLra8N35hlctiUskUf+CpMant4eA62kMP1Exe3Zfa/b4niUJf1Kgo
qguFHTF1ZCWP5GzN1hF6caeiX24KjVD99+9wgjr2WxGfvGJkstessOf4EV5MEPuX
53cCEMKGXacB0UjzbW5q3NO/cJYBcouz9za9CVSxW9buPCqTEI1JYDfCJLcaoPjs
m//xH6iofbqy8A+t84tcF3DS+ioCenNo3ohSy64rGdv+n8eRoErxr1LW/b4gVMGT
w8C1DEWY1CoCLL3WGmJ8cuUz4Py5dUshv0eEv1wM7WeqLzYsUyBC+Z8fhMbIwrQD
ET/MEYloVLFJB38vlEhegMWv51ZB4tgJfnq/l2B3uwaXkX+VIf9q0pnkCdowLcDl
/1pKeC/tEYsICm+QpczzrFxafW7CXghqEZ7wShaWVv7YmJdisViIlAVE1tRKfVd9
NEt15+EDz1TQWn18UYFQBWZZx5nEXE/LcmoknWLSXCImskQP11fDJjOPiay8r7Zd
QRtJjCuxS+B9+6JhzE5keW8YxPvQltyYtMb63BWXE/wqcLgFwdQqHyyycdpkfwME
OhmXhYjvNBQJLm2hIYRVIRWC0sRnycKS0Yg2mMKu+FnFhpRRSDENtehrckaTulCP
KjlleJkgbha7TJ0zLV6ZPU1bh8L7D5xdH6Mg7IaS49SffTzFRqPGz04U1vtsXEF5
LcVsLEOKsNMZppo3dvXyF9tqYAuamaGYp5L2X4Xkhz95Qmubm58rM8QOTYa6S/EB
boRyUoDA7aZBCHULY2kOBxUbhjIgzcowZmMD87Ios0yKEhLgzVFPOFZIs7K52mrB
kg9cFoEy04Bai8xyvxX9Yh+lruvwpn2YJMhSNo/7RWZA+Sj0zvkvgQnowxTG0l52
oVOVc5ublqaRKUi/6GezjsLy+/XTHEA8GZ+jq//uK5dBvNzCYsftjDJid5tstYrG
nlgoBMoRmwZXfkSejMeBwO2rweQrUjC2tcJ4FI+wBYuAIm+qLn950WsxL1JjMS9f
ZOu7MiBf8P1zYw8aIaw4rKPgJuddaAefvQrds6ASUuruhU+AbJrCzWrSlVml4kde
7E9yoV/MayIwyqryMrQ0msUNDICrRl1I52aSfcXOWuc1p0PvRsYXlyqfET+hwd1s
p/RDuxtCvHscTVrGBPyGLRtkVStYNKJzzm2FPuG0Yp5S1BqprCzWU1vwmXfcSQsk
YfoI+5rbyNa0fYqDpXUw+Vq0NL8emSQLXjOm5HJWeYCiYx5KeJiEVy+K8yWCZg4a
KeL1uNa99GR6gsCBkJsmZlLD9umIsfUS1SMgQ5edOp2tTFQdfiRAxWeBnYJ0L9tc
PIco6uqjoDr92vp4LMyXiJe2Cv+ciaqYuT4vox/JjgM1kMUT1aKtK/hoYmC9fif6
qgy0NUyCGr5GRJxNvIiHrURIeUM9rCyTjguL58ZdW/uo2j2+UKnRhFsqE346tVqX
nlop6LJstrc091AK2gTvcGCJQZRHr3xAUt1W/Qz0Cn5eQjQLPmLzi31fl2f4ieoP
kN2Z22anlFoRnwNNPqBlCQrstCv3aRJEe9gTobrIQHQiy0o9Em73yn8B6wamyhn9
mo6W2gFNXDsKiCh7yrTa3yMdc/rI5d3bs1+VbFYqDOAgZcFhKOg3jLcBruT1zXbK
sVUU19xPvJUozaJRmq3BCqRfF6XLIckNeA2UwKBoT6P6wKQYPqXFjCBTqOKZtfVL
hnN+iE3liUd1HGh/6gbiqgZ/vSgHFMrLAh+uypO2ZZAUUu/aUxYF3lF1tnOV2VMb
QjZA5pin51zd6IipgVprcgzhnxJFXA8Tq0+AK3eINtMtXr3Yj+4Uhggydna8D4ST
C4R0HXt19ViyPLBW6T9iQHHZ9QKWgub2jcG0a5T1sxuVfUfWsn6wgJS+GJOTIDkv
zdplOIYNgwesOYF3usTnpGN2JYFGKLmHUl6UgiLbGMJt7Q7HpXpeB8VjI1Kil3/H
lnc2YauOO5vwZi59GhMnuXF5l4oBTXHAKKKqdymBguRAWuoru/674dKkhp7jB/yk
XWTD2yDxNCicAyxtN+JBQ9QQ8pceu7vbuJUUPql9I4KrPm+ItrMR1lklZ6MN6LH4
HAID5xXiXwvDeDgDsVwUHlhWz/MnjWQt3Wtg1w6a8W4imx4E/Sa3zcqUQ+vYSEgT
qjJu4nH1t6SvN8Y+0dIV3z7e68Ktv9rBGj6QK7xwwK97hYcwIg5B5QGKyq4zPTCW
SJhFovk0fGWbvOOkP8q/LrU6hJHQzZIMsoP1hWvu7A95x7p2yQgYU0BXcFzmKIzW
QwQsHXPtVBc9ZXahzZyGNrOR0mqAXYGZeeAPmpELA73hd524CEfH5drm7j9Y+9tq
/AFe3NKGOf71xNaZWnoYySICmE3SAx18RIrSr7XLvRvfONr3Dk79MR6J62z5laa7
iMurByUOGBNzeU62f6uSiJ/Klf+jEMuIlNHAqKWK25EJMThZ+wbwVEQYeYG0YMXn
np95epgXC+4hq4kX34+gagYtbmhQVGyGuzAn2PmCwsrfydwE89CZT2TjctVl9nOm
rfVeELu2uL6mVKzYGVjqJZGhFd3urAKVawU6H4ee/3zWUaaptRS16p6KwT6YJXvh
KGNVIiH1GM0ajkANBcl0Rt7oSpnFSzgF6js9QxXCOWDhg60DZ+2wwwkC+Qhz7AvL
ib+fcyH7ILvW3qhncGf6KY2psS5sD0jn5vGeDvP8MY9HN+trcAvpQWgFz5NnaCG0
BoXyAE3hBBONGD5WjQVtzfMpon5DURKckaZOxZTxw7W8ULdICc/2RlkTogcC+EnR
39IWhUJcF2VcB+nYlnzofRe/Czpi0eU3BXp3l+5H4lilC/t1CcCJ6ZPOqAArc2nO
gmTzdTERX1uvTsuSV7czIUA0mOz2RlGfMCGkkWFtMso/P2Vh2/WJ2U9mFbelucXC
L6478nwVziiiNdWtYzzx96baK+kn0ojwQrOC6hMPFIwVvWVRNtLewW0BeRGQ/R+z
TK20sI8Y7t/hQZydbQDvuZ5qOG0kEH2Kw974O4xSg+rVYEvW1dVnm3m6EhLxmIir
+uQP244hpYnK5/F1yjeHwZMZ1qlzmUbAenr6jIRurhGuWTW1l7A2gztdH/VLJjCi
5AEaCzYxlSqFgJhj7A7+Tsc1VEVj5Gw68FolWNDOncONXzwEd2hQJChSsxOW3ZvP
Y9GmI2F+cs3DVQiLNvRIpqO2uxin1B/8vxtvdHTjCgHvkvc8NkScJt8aF+yBZm5n
HI9rkHxk5ABYIw8l8DHnCk+pNw2hHCYnbxjylP/hz6ZJb9kyI+td3NannELaQmAV
05AgrzKNIXm4QVQRPxwukRY4BPqo87vvMnqkf7bzucX4AmAIUDyBHwWpEX1Nz8Dh
GRLdusIIhD5sXA72/hN3u2BoMvp24i8NXhk5O8aCJkfkfSHl23m7dQEhjnHr5nWG
6kaf9uUPpNwKa1Y7sMLYhqfn4/VXCr6bHYbF7N8lWV7zPY95uYPQt9dTAxu3BMy2
EG6j+lWXa69cIEXAm0HngRRTnFmvJ3PEGsauwJvDOkfhHKq/7bWZJya+EypO64za
Sn7BTpNZJxGFhfEeroMIdjfIvp/2FUmkBLdWZwsXm56sZ0CqEncGYo2WK/GsO9qj
zb1xwTFeRt5EliWyx8dKtr+3QZ/C5s+Sz+ITbJId8M2uvsf9ebXqhISmAvShQDtX
FcsEmZMPq0hRtgrCa521EanoGR8U1ctYiT0VorJhgst2GT7Bbpm0Bs/mDCJ/ibnI
S4dOVx88HVhDtuDW9Liqqvhz+NkYGYf4NMKIVstHiJPURLHiMF9d7NlXW3GhBXso
psT/laN7yWgTIYPXyhHTmnd70djou1P1lhDPvEGiCFS0NvXZBKwIVaDFW8S0M6Gc
QNgbXQgHP4gUMk8TGGYuQ3oq7ztu7Z0al2QNEERLX6nImII6lUU6QunA1aa7077A
LAptIDm4/5hx0YMs/tHxhYgHxBnnschIAIKjua2GtY02VfeOROLK8NXIO2wd278Q
Ysj63qWPlfTqlCQ8kqpSZFs58wiFU0EF4CNCdq32veKXxf5dqOe3WfCCLE1aIfaC
KqDtdQwWN+nEVbx8Z2RflOK9g+vGnlRYHBS1+aF9gLlxj8YOKetJUkglq+vEYWBv
wHXxkgbWu5khn0/kc6EtNRio9+K5GkHpgfo4nTfb0m1HrzMVffDt+ErDK4lVoZAc
YfnjEpyRqO4tbuNX2z6Y3gIWZJG7RnrJMOLtzpyvJ9OsCVZsh4pY4UTLRyjP2KcV
KSAaVdG2XPo06zO6cPBIEpjDuw1v9knrN70V63tP+cFboOOpWJS3ixFVyA7ITQB/
U7YD8lPFThqYehW/E9IgGK0SZvx6z8lfHHff+XX31dsjOP02FHgSmwIKYxxn9Wp6
Asd4RqAq/oSq/Dp89Ee3R7RkNidFUN9CUp0KEYeYVsHnrV0wt7ZauLLhqr3WkA9W
yCFFID3/GNYgw7jnFp/gTN4iAoEUvNgyZv7p36N57ekZAemayjHPG4/fMuH6NpOT
uiYL4kFC6xvDCF+HCNbv4PLDIpr2ujE7N468NwTyie/Cj6ASmGOI0vv8jjGzGlCF
C0nny1cHrun3x5+kbu/wBDEvptbHynTSLgOnBta4djXw2/mwqqqVaziCCvlikAIl
NsRo+M22jnzlZyfqLbHNAUz50v2UKvRS0hHTFtLb//b6K6yh5AZd4d9VHDNFX+y2
+N7FCa0V+wfSnlbM3JFxl/yxN2bgAtZETzqrYB/EdY6cR9NdHoh1VZPa1ZOAZJGD
eCoRVRDZgxb93rnLcZKL675/FGOU0x914yflghAvz8FIojeJDsL4x8eB4t7ilYNH
IPbqlHPTYTC5HijzYiwi0VyXaR7GS7lP+cJIqJow2PAkduKCVm/IzkhEqMEH85d6
4ZKekj+lL3mHhxFhUQLMcwAGP5nz4czzVUDuNW4bKN5eMge4SizoZjM0Xarn36jF
8RBPz6La08Cuwc1Tp8B2FBYN6iaSx15NQXaZ6YQLWg2f24VziLsvJKpCKSWv28kw
lFN8ik6Ai/gjkOOHsbkIsLbqao0f2uRlusRKK2RlDZp+WfQPcm7HBxnt/PSPTtyy
/kDS7N0dNA+as1PiGXGeCPDRNgtcteveRUIF1SC1FIAjYUSK+hTXfoFirlaUfFQ1
6xkLB9+3/rzO1n2DUa5f7tqE4WqpWHQutBrbAJUPBsA1eOwkrWYTONcDPcP78KB5
z/LbYyrncbby51eYJorKGUVcMNjjKZCVLD58lt45FEdHitXPXOKkBAorgymHC/HX
ti+z/keEEVotStgOy0WiK3YFu1LU4QAi4cBiEd7EeedDxio8VP4XmFCwfn3gnvx1
usOtYOx1DhRSSU+TS+PDci3g3aZz0VHZ+Q294cfbNJUEP4A6PCS5V6wT6QGpb/yX
BcbsJvKSedOnr6ayF06BgvO791CJ0XiJlhM2uwErNHp8aIeMKOtJjf0+3NvxUNyM
vCliive3tzhO8JDf9nLxsuygNzJLHGiemd6FAXaRbafmmytF4X2WlB5bG6gf1Koz
uKe8xqt9GLVWVBIphvg2BXFFLrmvNZ1JKIQjy9tr8V0/JGenlXQ5E86gJzZG3DAe
ChhNPCcv1w9BWZv3A+vMFjUVzs3MQg9Y977IhmGwULPZoYeIMNiZENOppm5j1KTd
JFcKbcSCNQGNybTOpXgnaB8Zq5qCMICRDbVXG6JDuDqhDstaDkRzC2nzPT3TnJv0
cR4lNlg7e+xiARFaF0dcZPa3x1iVS1lvrmSfxlWX3Xbdt2NHaLFWZyVBglfEIZyJ
ZwCHgyjIcGlqpA8xeRtgOd+svme7HDdiyYcPsdApwYVJXan3j8ja3MGhQhVRAaCG
ZGuSLK7X9STI6ZnxYfS8c2R18qsXR9Sh4OgWqj6uiGBQelsARDVwjPZxqtG8t6e/
GRAtvg66i02wXZDBWOnTq5bMNeiXMGU3hx1x/fUALwh5CXn8dD7v1THBIracCfDL
ooJY3ZzRuRe2MoHBacNxk9jB9KPelT1xNxFVwlNpus8nfUsaKj3NIzEmUDHf753D
awA+aLQzGaFq5p0xTuvOUKf60MZqKQaC2UBtsD8t7m0v4WnFqMrJiQtqGnIzahTG
7ct9GZuKtM4Diy8WasuYhd6o8IqQEoCM7wwJCaC7P3XKnuLhGTzmQgSlV6xssuWf
QrVWT2ACpG5omgaVuII08oMOXI0Q6glwG4nA8ID17Uc9ArwswUGZ7FCelw/Oc2FB
lwRyXaspzSGa9FfXDbq9hx1O9WXS13B7rMkhOMQ8U7XqUPqhzFmxbqZN+5KYgV41
QvTu7Ev0V3YfX3g7nEvAxkb7hTa6nHYdU9swYz75kxwv/LarQKfjCVlIp+gUv8pb
SJ6vJjSDR0yuENOah+BR4Oxlt8GqakrusvgDwKXeONN8DhvvgI6n1tJK8AfJDLp0
HJLoZ/QeXfsyy+WznT+IJdwz1TvSApKiTgz1e86ou+ubpzVADtT2W898fQXqkFYu
K3BrkTan96deMVmVduWh40/9h4VaqLqymmWMZ97Tj9xxKX6U7g4rON6gUigJLAIe
GuOKSbF54dbAHwNIiuoVI6vtUS+8PEGOtpKIFVgDxi4wVGJrHr7sMDPF7c4x+l6m
JehhENPZynKy2RaLHW77qhVu+r4GB0omEjHTMt57qaYSNqBk+zHMUsDoUR5zXjMU
TzJDG/01epbslO93N49S+CV2dAtgqgmNgF5ltD5DlDjbBFdtoCbAiglnm7byO4py
oUGOZtasd9sdaddusrzgx+BZbemMY1mOd6AvV2ZPOvG5kEjaY40s1GoiR14Xea4e
XFi8C9bhx5fvDpg/SsJ09eCAGc1mN2f+i1KgVp1UGNYVaDWqJvSDnyP4CfPsUF1W
T9hESRfq1aBaqjb4vP1W9xQ4BUt20BkJh3xi2droszTRDOGW+xXKl67UvfNlKZYA
ieGJOuP64sgCKOA2Ix6BLVrUrkKjkbzeF2naVLejgZBprA5ksdkE572BORMr6ET6
M4e9ApSF5d9mN0fx3qw4WH3HQcrQWfp9gw4TcVpUlqXjPxJ+l8goWEVbk1oYCkMC
n1BalLd8JoQfqZ9VZk1vAwZYQAlsbgsoG7zbLlVACl4I4cbAvYzln1lfTg6aocaT
DmxyLW3JRKptk9Rqvt19XJaROnwh5FmyVHgRK4jTdHR3bhD3qTGmavGJVin9VI1v
mIQXJkV/XMQdGXvxFhonzGQTPdev09pswukOnq0E2KW9fHTOpguQc6jBwvk5u57U
WKGsS4e6HGvsVH5ZdXes0qO2XyEa19V/MnRRgY1RxGkt+IT1AbXnR1TLeOBJRvjv
OIkjE1kJ57daM4NR1ktxtUF9qTG5vC1vVd6aFZ8Jt7pxHFK2FMSORxUHuvkqeR8s
tDkvJLXBqjv7hBK7Ug53v4riTDvNlRVJDqRT5MbAKdiQkGm30XL3LegU4wehWIZg
lzUMM8mOsvhIjKzidncgfjDnSOTCR4BGPrCVg9Tvpp9H7qtVRjw53zLj01y4s0bO
toAXFodi5rfZ409Kz5WviCnFmuXDTPzRxTAQdQ9o2eASAR94AkBcGAinDR72kkGu
9pEU5uRZWIklHSgpjXtGEI54H44VwwSAr4BlaVVCIhyeK9FZbXEa3hrBSZpX7cqN
LP10F7lvG0isFIlV1Dvfj0HehFzDNfH9wvlC6xkPvcz+cTeMXLg57WXdNkh+5/g7
GGVtaASdIGTm7zIM7dOUSTQ2P0Ox3B7J1QoY9Mym399TCjUfUkqXdFBIJG7mpptU
H4Dxijs3Z1nwKCoXovQVltodgEm7CUAT/626cnzpHg5xt7VbODPuED3usIPBul+B
lIZO3OIgDwykn91UWxYPspLMur1PkRgngj8szN5wOd4sQu24v2D98NG4Oc4vUNcu
GRjqOFQAfISVzKek7/q6mqEJMrELCk38eF9X+/OYzwiEep5d6V/CC2SU33Ib9G1Y
gm37JlFl9yL60W9fCGKqAMEaetqNgEvvkpHGlteJzhkFblEzriFUbwxnKXf5yJU7
fSdcQVAtOJO0n57adML48Z7e3QEzidTHwplMVFMdDNMoeD/d6Zc1R5imcLwHbOkf
YPhH4kn7ATGKU6oyd0QfT2AeIsVHnCBMb9STiCVg8LqhAk7Hy+eUyTJDjzxbW94c
3e/HO2qh5eYyPdpeH7VDQ2Rifn7w7usURyAPEPUAM/ECLgSPNdvUYIpX8jOl1g6l
kVUHuw8/ZJBkLilR0V7exwPKzQMZRBeQyOE+actrm3qO9asoIHEvJ9fny9VI/8T4
35PNwXBuP1/DVKZ93UJA34nBU5JDn38sl6IAMGYu0/veZiPZnIDYNPI/VdEE3Ej9
oWL/UE61nI+QOF6NZNPDePJT0Wh0IS/4D9Q1fJ9lNp00D5GqDmeeE1gXQfBIGXRl
ZQucE+yELDLz7/haHnzxQEYV2BzN8vmRfTQzpxvwXQY60peeTB6CzuqdPDStzTse
E4EPmjRpzVlKn2kNnkn6H/eAOM18vBOm8Vu3MGVUbwbMUST0o6FjEli8kieSeMMV
3Y7O/U1/YQ2kB4Jv+PlgOnMJdZjnhvZQWsf7qfivySAZhif8uXpbbF/2CGFCrOuq
I8/vkuh+6t6UWfzrOE4UW0Y3lf8Sd8SZhuYi51cbC8uL6yJdtMJGXpQZkWQKpOxT
xjXfvJJcoO31qzYaFmcdAceNu/nghxrNTEQ4COOfS8c2JpQWXYyKnXSw4LrHlFWy
eDpw/pf9Dexb/52J0VCZsjimvicdaUi4+5wrcBobH4mS02haDPvKG7021bmzBvJJ
EmMq7Twpsp7lmri153HupwURIjVJRuVgBDtFRUAsPnMLaKMIHcYQdqc9rJYWICSV
WmioL85p3miq9Pc29yb98Laf0WKW0PhRcdD37WMxROZw20hYBzxjRU4UaxlsPx7P
/qAHEOMRrxMsSrxbPQlBnVTq3tt7CpT/5k0EPucci/7sLbBt6vRfu8aXRaZsybND
7h4Va08oRGUnYfJ7DbGZNaGucIYiII76gV/e8/JSDcBViI+kvD4JF2wh9KsXOE5E
0pBijtJnpATyJFdw/RJCZwcznZM1VoBkhXaryDFaEC3QcKwN65aztHoOXBD1kA9k
0itPLLdmhkCorFkxcudf6TKzLa74SO1q6mKNW1GV940ITO+DfYLp/ENb9T1k+pI0
BMQDJOGUj/DSvwz9NLIZa3QQarKDW60vWPapT9dIj8ROuN+wo0zrhNZJ7DWHPnsM
aXWiVuvgZvcrOYUZ2dSfyAoDcQO/cMhcQuUYjsxFJllRBycHRrTOXsdGFn87/zQu
US9zwz0o6+XhLe0rwWWk5ZOCjgNtwaILaJUE1cd+qslRTRck6J4qdPj9LGoh/LZX
cmGNWWl9bw+2scVo/XcHjNl3rKPbfTtUMIPa9HxIJ5XuAYf2aQ5ycaplYc6Xvz1b
jQB96LN0SG48aajZRZojqA2Yr9AJcYEjFlE2AbrEaQi/fiIGhI55bGKT33AdVkJG
ROfGqyHQx4Hw9oCqMXw9f+4klctdu6VylhY57H//MVfS21oublg4Jj2bO8ggO1XO
KBYkIVP4WwTQqyUimqPvYoaSnDUfxRqnBuZAqXKod8+du2BnWdvrpUYP6Pu6IPmd
3iJ5d8gXd9pZZ6ZiNEzS8sgBdlGtAxz5zFiNESIOQcfFLqWlZ7FODUcjy7oPespI
dsJ6PQWrKlBQE0KiHUBijyd3t6ewFm+1xpTY0CkpxGWLI1LobXWsqHhqfmJNN8K9
yMMsZrkl7vmZej7r442WEWPGlOifoG9qhOIIcG+4DCQHXVjZUkJ6a4YVdkYjk2Iv
QERdzTue8LlqTflDSBRwiXCarXTDH+pzX/thTjDoQIoTHDjq08cvQFEAVOcvEu/K
JHUUJlRE0KoEjt1Bm2z9F/HLHUBiBxh+WHER2n3oIgEfAlGIaNENyjrgo3GlPndI
6S3kscoHLNqgUszMlwOuGIkW52p8QQAkBnR5tcorQmOTHgKrMaTBulZENjS5bk25
Pp16/A/+OkxdQoVe4DH7TGrXj/DQZuz+kIdpu/orG4rvtH7OW5r+qRfkyfiHFeHr
Ff8M5GZcPTWqdLB+YyPUcdrzS3KYMIcqFyE4wFJsSZ4cBJ3k/d5re2WlAc66xkhQ
1t7uhpMJ+vbYQN/FYjoaWQgivztxd/jIT/jfpzD8cxNGGs1/1tgJyjaumAh1CP2l
xcK79SF+Nk2ETrL52/YikYDmChY5WW3pYE8tLXK1P4U6FUFURMVA7nMVbXM19Jgy
YmmmmL02aRoEUE8OFz68Gz6s7Pg2Xb746fNcYrGVBnCUGYRLyk8NVQt0NhxovkYK
INPI+YFRFhcgeDeoeE1QJA5D+akTjewFK0UMDOd0MHunFtM7u1rakg27sl2uUiAW
R1GZw/aoUZ8zJWgzl6uJrVGZwKRRlDzFxigcnc+1yD9avPmrIplkTAtQVJ5Cl638
G6HvbwH4amd6vyUegzIKZH9iYtaUgkyvsbRXNLcduB8D51ag2XWKkmLgYgQGn01T
deS0eGdFWdIefp6aeN3X8N0FpEuhPyWgJBzdCoBtyRzs5YxDpwnr2uMi5RFUk0zt
SYwkSzhr/jlVhrB186ep8t8V8/+CW761EUFq22bm4bEPkD4zpd3fMyleD6adz6qx
Ic+hFFnT7W7ybR0wL/byM8W3+QsjDlfhBV+JJFFg+UitXTf2h13m8ikt0//zyZaF
k6w+i4JEoGBSmKAJD4VJCMth6Hc0eqU/37kut7qWvz6n+g1IqIO6ysZFtLhnd3F1
u9EY2PdinIszWUGdHpNPz72beoTb4qKVudI21yqGMCkZCr4Coe4oRXTBOf76v/9p
Cyk6oA4kBg2S9L9pwwZPefZUNmLzG2+V2bjytdDRlwP08FJqEepC/5Ieuql14oMb
e/Tf3xIwxeCi4rDNvr/TlbUKhRAWLLYMTpKf6zwanfW7TYZoNchzhvgfsWa/T/hp
9qKjXq5xitAeOaMygwgId7rZUwIOnsoLBkDhdQldcztlqns9KJdiYH1QaQQwNAtu
IgaqVtsTNGWvDvMXn9vWcysZdNMpDC5raM1qNZsaEY21lgvd6EPYByoX8APomtnU
QHB1LGcwoQKDdCW6sRNHpo1qooW3IaawCHOu8cFVhOV4BRW8SuEZxdvtCbshNfjk
onwNJjzQlEUAMdZylmRSq9Ti+CSq/r/2Ar0EVnYFCMJYttGHG1R2KGlLQM2Mcy3f
M+hE/bufIDBHrQ3l5RmvNIhzo7L3DIkVrD2pk3F8OXpsgFbwbbJmjBH601YzZ2C0
apGfq9ToKGdXeXje9MOCJ7oy/MXNX26k4oYXd8yy1/siEShmX3KI5/eXGFuH89LR
7Q0QTsHmjILQKDJ37ahSd/XFGnWpxCP548r6WzlqCNScMFecFxZVGvs3arcEg9Un
pkQpizYev2RHrK/Qtta/9mQNFfMg9Tqdec/d8g7Xt9oHFYXs72FDzAEIpV5WRgtA
i+ZEA6xWPX3RTOuaRtzkUMQM+9S1gLmJWNSewg27OYfHjF6HDPw7ELBpgE+gj6LU
oL1RXunb/OAB3isgaonbrMPRhtJ6SYDKBC1I9iuaHIMJGxnnpGqjTYjzB1rM720W
GyPBhtrhvFyVhZJBxsKLoN/lVMKAMEYr9Fie3HUaZyKO5Z0Ns9c8Biy4r+mD1Q6A
YIVt2FPOlSSze8AS0Fmpzbqmn/NcilGvNJD+SeJ2zlNFqzD65vRfbh+KE6z5R09J
aWcrLVY755rBr/S80/I5CseAUIki7QUgq8XlmAr56Z0FzT4bWTZ2bcfmDoaS1XgK
uGgB/03LJBzYdLf+CD2baymK+XJPsyj3afqRnehvbhEikCPXCOs/GXKXNzRvgSzI
lXe2wKcoafwHrt1VC0JzzVqBXWFkLBA65jpdDHFxJ13b2919ijebsFlXKKbZ7lMm
rdxHxXrdSQFBVVNtVRaon/K2efonhtWI0mxJT5sLtjS+RwmJKgcfHGoJaZsF9677
RebGNfS6z8oC5xB5vGwWmKggYDWuMmcSfehxOFsuZQHSo55EGvnBVuB77zQFlITF
RamaiFkTUoRIcVpqpMQoKU4f0Z+OIyf2BpZ/cQp23op0S3GO8CFf0q51p5nF/RNJ
WNyAkQ+b86ejlF09J1SmesX2EPggRWzQdvyPKNWx1a4AOchaRAlQ1dIEtIQn5/fj
/BW6qEn/hVKrQr60/o5/qEwmx00GlYVopJOjl00bz4o34RxZqgL+rtlbuQybfSkT
Gg5wDAwQyIhD3DFh+cXgwyfWBX4XQPgDKwX3EB91V73xncVpO6MWkATjMbAMUleE
juqxgNzwnn+NpaaZXZaPspjdLzcc3ELJQvYASCBeTs62S90TUVP2k92cNcl4KGDl
P0REeCwCmlXvJkxXrvLS9NChE0mzfGpCl9jf84a28AkhAeLIbrg2e6qdvZmARSdV
Sib0T+yy/FmbDyB0P5ugmoWQS2JEK3KRT1FjLxLOBOtYkjGksUvnZ+C5yPXGKK4W
B7fNRHrl6zzhGYG3Mu1s32jazLlaajr4Ad2AOd+mIqFZztJDCbmNcc9cbc/ojtyo
iJpCqSO8fRbKZ6mIp3bEvFVZho9I0R/oAAt0hhMVKhqifxroBhvaAgpjKEmNn+NG
m6lklAj8OBDReUjtJNkvEnSR4LUHXMy2A1uG76LVXbtfQzliKzgF2W4+vk5Xih4w
jy/fK82UsBz8NRne8anp2ZW51M/HW741IutB4np+E0roi8uK6b7Tngr3/O713+OB
pBNN8fJreWwUt5kpkQAhMIMIyEvCTqtRAb9sdM/VV/Hk5mpSmKLZTDK92ZZrWtuR
CwiLyAe5iIsBtG2e2S9tELRHaxelNOvD4f94T5JzkQ7g6xcx3uOvfSYvjmNsAhlm
UCIoYw8Gp8qMsNU6IWsM0zzg3+gEj6OvViu8WxF0KAk20krSPVN/sVu0GAtUsB99
lp3Jb6AYdLmCSn1WoVjllS3DpAZcF0poBcYXPUKTeaAfbH/da9LMlqr0P2uAPbLv
Ryc7GHp8V9kUou4EwNecGL7U10Loayl6Oh12HG49ZG7WMJ0/RHwnMWQaWpQrWBWO
Nmst56QzvLbsRXYV+lxkTactKfEhFvEIpDAxctWf+aEWRVaMwsGqoL5UBpmKO4kk
l41BF4n+28Y952TXROtICqKoZWIHOdEneQuOiOr0Z2m6LG3PKlMXJlEChL30iQRC
tQ6st8zeql/EMdrRXnd/X/8SaQtglzdFPl5GnEvMmLKMDgupI6Cvi1rA/DDll1e2
BjS43QP2FRItKXbraYZ6XuLgsGbsZVhiY2GQbltUPACmVJjl1RW6jIr/sB0aBxFw
oF8OetOLWp2Oa1J5nHjGl0yI4lHvAuWUucMdO5RSCXbpaH/FgFlJTihXa+PUVq0q
krbzdInlHHO0V1Y0oDcohZyltpv4GqfMU4gzQLJ49Gyp6+hkvv7hejAgboXA29+o
gZDiHRCJ0ciY2Bwiw4HuJv64bDS8MPLSKU8YWvUhrOaJzU8qtsVp8LmfnGAZrfbK
HbGRwhKzqHL5PC01ZFdCNmwEs6AWSOfW7Y+TOmJX6cN9tD0At7xpJ+dUHwnkUepH
1urctI6vibPAFddtcjcdl2Jb0RlORoDyEakXUc9LsrIKO6+FvJ9x1g2raWjJ1XQv
fJZSVZfVbDaxpbpyAx26efTC1IwWwsd5mhv+Yk7CJvnQbhHYb5fUUDnZFRyOEak3
EgKz+jid4mtrqUUPw7G1enhe2LsiwvrxftLflHIqt27zxqRb6dDfu5XsdOgZKg6H
nlIoXjViaZG7zVQOceDaMhUitgticvTxWiXFCS3V3qtO6DG2jypp0pNrBwajN6cn
2qM5YcRlWjKC8JgW21DMis72gt1qhKY9oWARcVkPq56DAb7S7tM034+ewEu3G0dr
fxHWJfAm6QGNbqhM/lKQPLcEOHh75lH3d/iXHITTyfFpczYm66DhddDetN5oYbY2
6eusoHAFJ7fHR3x3ozg/TqB6zT5UgEb4sKtKHXlYaLuYKbLqysEKUZq2Dt1rJ511
92BDLvRGmxnti1dpWfitEK448P41+wLXvKNB/aYNS1dRk0ODXuzy/V8itzeI27xF
SfZ1i0GNhKpG415P1bvU8ovpnsYPUJ/Bc3yOkeUsPzQWAKLzV+xLShDhUaZxAPRB
pwnSXOLAuyOMimczrCu7kK5edPaYUzECVTJ70iLb+vGIjTQyuo9QKIgasZyQgNJ9
fGSN+/sY2fsAoNF5C9o5MdXn73pB7L/xYt/Rz5bMRSVxOz+WxU97XTz6/oWXCSrh
/3FiVbqYRWob8ZSfsBNweOkFj/aptj1J1uh0nDZyFPYOppxQAxbVqon8jZSmNZH4
Uws4QONkxpivpgkZv4fjZwlV0bOP9nin3rkI0Szcs0aAX0gO4/sEfu2h9kJnaUaM
U+aviRpbWmseNw05FCe3JDqJVdS4Qe9EkYY8KWabDr22ovlBeBRGP/fVlHNZk8r3
wGq8MO1MRpfFYG9SiuqT7wN1xmaYWI7B/iQXOoT7wu/ERlxd3QsDQ4TaJt9W0WGv
YRja0vnd7bFVNyRwJ54UEh7p4BqjquVDdwRsc/GdoMdmxvHvklQddV4lm8MxsWrK
DBgjGyi2ruMvqYwpNnhkXeDsjVVhXo0Z/CwxqqThFtEcKohgUlC/SDo0eyZw3nWh
yiEFht/Dj/qUSiRQXbnn9cDzGSFfVxTVNv93AuQoaE+ihVuJLyG8HiYSTpTZlbGY
PVtMGTYJrQ7jbSCRpRd1bLPC8NYIuTaEruiDOXezEMt/mBrlYYzM5AnQjAq6Ggvq
plESJFdv8v+8zqDE9X+mwiHsYl7J+CWrjvnYAG09cXugenv9nd7ARN51/TmCTjNq
CnthhOa7WJys8p/pTSeMDlMiL3YuUY7G/oLotEsQF8ogkhXoVQ1pXs+63WGGZeiH
qZDhW9UmhramQIHGSmsWobwmmv6I6bPuNuYNSyOFVH7oEQIL3j5F8u1nmz1StxOX
s/k3T7u1tmAkIdhgae5qXnUoZaURw5qOLYxpiZSs9hFRkAlsMpOv5EetVufRiWWy
mk79KD39lB7+b9z/z0AjuOSafWVQGY5+0bmZKKk//tHv6M+8HkicaCsIyWMpBV3e
nI4F4Lx0p7KzmcWKPlKoQi9Q4qGU9Ggb263tWaQZ76Fh5vYHb9HpX1ngBXbJPfm1
Qp642DqPVg9FTDv3Si6MnanggQLagj+3ONm0fnjRwPElIlgk4bJ32pXCX4fjzBwT
A7UnLgez5Z2MLHvtyqXviehdyWJqULbp6MJqd9aG4UV6NPrdHauMQ8nEnQO+Pd+g
IV1mM8zo8IdghH1zehN8C1yMI8gKyYMd+oVakbkqcDm6eV1V3MbaS+mwBTjm4sWc
Oh4cBukLVWz12v04La6LZwFS1xGN5S6ksgtpnzH1sqP2fm8PXwCR5xqluA14iQqh
aXoDRAJF1c55tKa2IQAcW1H7IuEk1ZUYHg7BHc1ChENw9OxMWyIwo2ly3qG57TW/
ZA/yuhjcnhTm3eknyNi5ycxLgiBjN882xMAfuhg3uydZ23KVlLsL/XgYyhQnIU/d
UY71pKeq26U8L9fXssjpr+LA3UGoKRq0IFyEdqGU1SzbaRLYok1tUF0SX0T7xCm+
5zfjPPU1DfsZjx9tZRXXn8lckmZTfHD6nS5xjxg5FG6hC6jQEuGrcG+36hiFGDXP
RPBAIbMQcEQNb3vwP2x1CgcT7nSRMK8gGyujbggbR+oPwi6eoH8FypggHELLO3sU
pjYl3ybaE98u+n4y54EtojYNiL9Lt47LRil36oS7PHjy8v/TUz39OPVZ6/60wnva
1FX4xH03ExY2E3TJhSKi9+g+rEEV8MA0cFA+nCqYQUz+4Jqkwd6H1TX7uOXde+kk
87cZTQhasDTWEKnVBwwDgWUURwXYr0gN53ig3HLW/jzaAbudvnDzr/g+QISsqOk1
`protect END_PROTECTED