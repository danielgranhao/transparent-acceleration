-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
v1ffsN5HVC8qmtIiJsgKaJEv7Xb5n12XcWa4VTAWMI/XTFPZRkDa6ZntEWf++3ww
7cZTlGglmYhLDMFyGu6FuxfY6rWdiu5aLU8hVKEAKSyCJ7CQLf6Lyy4cF9CS3OEz
uHHbNV7GHP6j9egs7jEJ9u0LWgCa/nj7izdK1WFnloQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6896)
`protect data_block
owaWV8l4KRqtoVYHekOsiJOdaPLJR2P4R88HiU3rKqrZf7HgU6w+KpL5bWbOQowq
vdjs46pd5bJinrV+hOGlQ++68W2oP6ZERlRO1V6Wmv5yoNZPBPSat5THmFoq6luL
w+oQr/IfHksartTbX8uToVuGpMb7gSPr82Wfu2qSWcMmXSm767w0OmBvhPsJ5H2i
PUsDE2uMJ4Xlg6SBGUq0ZSFj9TB0762sFm+iyWUyLqQwKoV7Q2MwtPrtL02a5aed
iDoPOAEmInqXJoCkFnQJvT5NJIFCikaWinmfbLHoKG8IMmQemxNtbR+xAKG2a9nU
JCGyjiWubbFxOg+9YJWLojsJdi/L6/7eKTPESwhJali/gZbd/PmNiiL94cKPuO2x
ZeBjXtb5Qh6LUBbaUJWY/R5FvhONhxwrVYAVVU6TPsuIgUHXo7xA/2FKMPYCNc6w
xjU7JHnYVjSS5hik34J/tzzGtB5E56ukuQUFyQGP5sf64CJgxFqMGba7Sm9QVeA5
eO//vcjCEaEIl9k9Rqp0/MyisjXskpQltQZ+AqCU4LleWd7j3AURwVsKyqDkMg1a
qJZ7wcYKbc+TSjFLKeFp4uwhg5/m7+N3gdmoSngNtE90krR00a6vTHfPhbZFz4dR
zs4lYg05a2fuTUWgLJIh8Wxo7EfeLoq1mdn+S099f9tgzqEaAY/iZFXUj06ChVXH
K2rCLHk/vakfpM73jY/EFYui686kHmg07xvqS/cA+7mKHCsbhPvIfLrLXVMLdsnJ
qlv0dq8x/QopK2fT+hFkIGil5z8nzgTxGWHfC95w69NORDbZO5OhUff5GWRVJ2sc
mSPezJUeb3cpxMNM3IMp5wwm8j5ceiuJrRYwUuRl51VBAm6fJzTFfmpWX7l5ms2d
dBjnnL9ObVnQ6Lns+Pxpcsw08lIzfT041qSZItM2afKyHYkmV492xyY72HE24uOt
rg1N045678n+N+V1hlAmz5u8ewNk92dmLrmOVBRcZcg6SCty5UCR6WwQbiBjHYgl
UYXZK7wLtm/7HHhbq0dSlitKRZuteoaNU2criSGtPQJpgSDx188C26ApIdl23oEs
5wbBobGr5PKu+x+ApYahY3EG5TPGJtgj966N5PYXGfmdLh+opgUyHxzSwWFa1ZJR
TKZLe2AqINHN1iLni9rYnG40UkfIZxI4YG7xq5JULkkyXer9Oorj+uaeh4sg6RvB
APYkr7rrLr/+8cmC7DCj4Mv1Oc2KrKCBTktd9NPoy/Y8oytHfRpRv+Ug9vZtbX3y
kxTLl70wg6h/iJCFxyHIdBrb2qB8c4AqFUM0WZ7dKt+qGYA/g2Mbds36LKllFSMr
huqSnpoIUlQYaTcja4oFyGN+ACpad6JVQjPyEzOn0keZtWDg3cLu1p1tu0NvAC7P
AO8v0xHRGsxNL0J4itkvKtLiGp03FGscW1nYxMtqeNzBB6rFL+cfVtW+DtHvW0l7
TmlRiEFEU2Tj99ZwynE8LUaMOh35cqav77tdEvy/a2RUIJPpLFfDsb/Gu57xO+h1
aNslwtnhl6z18PproV4RHPqsRCnmXrBXIByzPnawm8AE8AUdmZxld/Jmi+j14vM0
ZZTwLtDAZMar4l4ORXjyl45C1786Cy7p9VNJPpvcleNFikbI5X7J3t2CcS2JKHSc
kOl8tawPSn8pYG4vueATi2ljG+jrsvZSrphOy2iqDDKZj17K7JT7jBqJtjBZFJTX
YjsiEp6hxkVfjvJ/rhuraqfwbZzCNqde76Tib0v0tKfrvK0NV1msgLO2mS8dHQfn
uezTKRQOrJw0yagDxqdtFK5hGZ+wjqfTEMzVFP0xUyakQuzL1NIA7Z0abIlEHwh7
Og49b8rE4Ph/Z2ts7S54toUFr8XxdVlmmfJScO/kWc79+SAOs4FWf16U6YISJ0Zm
zcKu68+VbOf/S70n+vbxX/ag1rWNN3Z55HdLiN86FJdqoN5Ik/Bq/lLk4ShlUabQ
AaYBofD7mQ/HT4Day08q6v+3Pms7dLzU+LUXBWjX6bdiL1Sm/2MR70hsPb9ovaXY
MNCvQLvUhwqzr0e47DafpW1Vsi9ViWfCNpqkCvBlPz3f9EdQrIEUfmsZkFYDPs3Q
GVFmxcsrVSQGm/EfXytHOTz1Rmgj25an3+eqtR2A0GAeQgkSfN0+HJH2RsHtx29q
W3iW/cqxykuzOiXjfm9kEn3iH75lHvNYuo25ewlh2venuKkTJGrvtFKCyNnPYCgE
35W9AXBA+o7aCZechZ2XzwqkSV5WZqqtJb5ihlqBJhtfG3cZUtXb2bmB8vRM5IZY
2wNcHxC3iMHpXNZnLIY3FvAVKTeqpw3VpnGTIDznJfmpiT+vueLf20GrM9p7YHJa
AEJcDP1HP4Q2GS02T+p78BeRfnMootZoNhwHyz26qjOSBzgOlsiOQyYkcCF+26Zr
9K3RbhDvbvWBRhp/VoD+kkZsbdu98GBfFawQp0kH/OP6EHUiEOEh0/LM5Mgrdism
zf7vPYmbyJdih7vJ1Hkx4HAVXF05sy8AlrAM3dGJo+ppjSpmwmBbrSy87YUWgvQk
0fZOg11sSNOdKbOM18trXYg8Vi0MKeSrbFikeC9G0ruZ8gdZMme3lmJMM9kja4H5
idzWlLXga1ZjGaHYcwF3bgT27MEWWV/wfEFy9aAPYMS2uypvHPimdT75AfVjVHpo
t2Et1/2Esiedm91hKIroGSzkeaDWPbwnsShIeP2950h1MphBB9LFWy9mf1Qw4CgP
6WEq8V+u+JUldtqYds5gWOB77xHJqZ9i23YOG51NLClnk+TXHqmiL1PSp/T02I0X
18Fs+Umw96h+4CmRmV/sXlKWWQuqfq/qqAOOP+6RhQQ1OU8Tk8TgAAPJy3MgkRjg
ZtiOAC4m6IQu4OAW24AAPRmZqyvLc5h+cRJR8jgZNvWoSfshMCEcpN8+kndNC5jR
3XgbCL4hMKRZCoZurjCaik38UX4XAwPTyMDQB+SYk9ewAUbWXjGgmqNelcxuvOZE
qlqiHpv+PPpKdbs/CiMmfQeL62HyNNed5O2iN9SLfvVdfZ4521hnJMgas60o/EOt
XfNNnxCgyucHmcGGeDaShsOlNMYPLQiKiXycohIx6emKgZwHrXB+nR6V8lIXgVid
8B8tteGQ6YtkuMPWYMn8WfVHlASTQSoxvrXvLB8q7LJHUOEc2bKwWrrtJOm3zwDi
6RniFoCvm+gfOIFmjF/xzjEez5mLdeGZ5T8JZutxKHqk6NMiqAr/kn1/KoFK+KRc
K2PhLP3X5NWUhX4U8J0QVKhvDjx5kDBBCbGlHC5hWnCRD7MOpdp7Y6kr3EfIeCgf
wfOY9IEyhIWPLv6ZYXv7XXH9TYZmmpwxBIDXUh+9sai7AnNT3PD/eIuXX1t/kLmv
ZVBf+hIZmnz3s0p0iB8EHlyulMiGYvets4vMLVVpY0w2NhkHbasu4hYrjF4bNTve
5hRJDQ5asQXM0jmoEjehnR38UBsUNG5LMOo90Qvvdjgn3WbeNBjLPqIUQ4Xq2OHZ
orboQ+lDcTFktcDti1/8VeF+h+Il8pRfqbmJ8u4Grr7sEKdx5nyujo/PrSMTajVP
NtMUmmanTh1tf4MZ6COrdGu6uOp4+nVoblwHVn0qbxv/F1flw3pyT85xGAzL/c5x
YyQCvB4NPiv7ZN/1Y0Cvp4Tmtn38xnTG/oPLfuge1GB35sv4ImZLJHCbHWSkub0I
YieQbc912pB385cyOvubcWanvOZyUpbcbLCLWLk4FmXyqkIjKy9FaXl1BqZXaewI
syef8SfJ3fxnl+hYrnmL4enMbyEyLjLE0+fTdysGLktgWiMERx8Z3MPhQv56HBcG
BLznER8TarfSVSSmHtOT3PzToBKRHlRESUcoQBeHQE6p0rRKi8xF7bwGu7Xy4qOh
EqGwIQuFsCy22x7k+kmYAF38tx0Bs1A3VuJGqE62oI8xB9r1gujiYeZLeqSJwGqz
uo2gy2BonGJmTv4i1f+C4nSTLq4Reo3K4n5fhXvYNEMdVo34ZHX0WjMnxPAaJaui
tVwKnUiKGoEKS1rzhUJkBqvqYKFn2IFirE56MX/H1FJOa28xTiIXbF426+koXZ4S
EG4KHGhBYZhIzN+O6qGPSJM49TYrUOGxaR/g13Eq6OXVohe/42hITzg9m1B6geIX
zFXzFneRjhZcTV39ZN0v+cLJ/424Ggabz3eZaDiLUQXR9dLcHBw+p4dIZYo5IicW
jwMwFzbTAugrvVocWBf2VyneakqylCfZjS+YNIh7L4Du6kRVbWCZwQbLCeNDc7aG
+4UalzDeYfUMKSd7Tuav2Oh0xCDh6vO0qei9xUVJ/CRV/mVQsBXeiGFUUGIXa23P
p7ftpM4CNGnVFNYKuGAUdqGHz6gpj6nqEsh/Mf9tPTymx9HE/GdlD+uBHi+HHZGV
tNNdEhxEdM/SFtJIkNxtVz/KMKCSLrTPVEoabZKQ8gN2KUunme5NKzKBHob4ACe/
cugdw5QigTq7q3OJXjgkddK5ePamVxgpJFYkjWkuc2HKfEy9YMjSJfEMKRBLMDgQ
6KuITVFHDRgZaW5pg1Y96n3B8cH0cN8FaM8BXKSeJCUgTIuzR4gdLQoZ+R7sukfN
AeSm3Pb9nsHiNOXni3XpSjtVnFfnSwC62NraXYqamuQWvRBl2CTDTetAWVrYK9f7
y1BnscOkHyT9zPaaWWVHVeDuBpYTHKvZWCgTQGKgpP5gnItbclMt69ou9I9uWbVO
Fff02mpp8JaqWFDzY7bHrlZwcv+k/E6SzZNxvt8VpQauMUMl83IaHIx7iICrXUz8
QRwoeaG3roMO8lh/YFngxJeOv8G6YHEK3dZz7v4uMKGDRu6oGQxeiLOxwwlvNVDI
Sl8SMIhYOr20R2rpf41bNlMwmSa2yqXDAacfQRGJYLEBGc10rFg08kxlIVNl/P9o
k2sUEZ45qs6Gj/cAPXuJFDN9krmleT5n+iLiQ+RxOGU4d07TCJGdOlD8mmePAcqJ
IXvbncwswBBB8i4puHhCtIq5C2t6dNPvpeON/tic2xq3bVRA4eEh1qKEygru5+CZ
IZ8Fd7hPcscl46O0kFdMAR58buEPZVUrceJW/ihZUEwQw1tOjExVsfb+pTUwUerv
8YIkCw7HgRGBTlnuaneu6taQgI+FaZUvyHlR5+XVLF6kND7ujcP5q6ZJ4CtN1fL+
o6zy7XnPtFtVzrHUKsp+0jPmn+IsBTPmMV7/94EewrcvL3uChiXlnSFsS1i9Zqqc
2ZCExbD4HqueNj5lBJNZxxMy6MlRf51uJ02LZc0qaeTbaW/6BwACJ1pG6yYcblWW
R8zVnCXKuZM/X+f3HlnwHVGFXVJ4fzmbMDQlZt4wa4lxTYCgM1I/b7VWrCeFZGuL
5Hqc8/t/Zrtj7rVhdvLCkLOPc+blX8H5F944zjlQ48fDq77L3s79Md1xLIXVULP+
LIuqQ0mB5Nen5ssZJVgBiai1sJu00OFfqh1AkA2tvx/BpLQx52/3n0OrMbFAsr8/
BDcv08AyRHCunC4zMWRisRMZPZW41ewgAoULTwy5CfZZPVO7wr2Ii5uHEOMXJ/Ak
CPyg/TJjkY0XyEfUlir4ZYUYdT7Ktn0U8TKwldo01wl1HzMRVu5UjenX8OOR1tCE
qdQOf67gl+bIrH8Hmtj9FWq6fIUTI48klss+CFTecbRqOX7Lc3B9OyoWP7MbAIZP
voKMsBX+MY0gzZkr2YD6IGTyBlandtewgViezrOGaupHcHlmSTK6JvdQeqlgeDOB
19GVhF15wKPmfldNrRc67DOxvzrFqbzJne+WeBE3dOSdDb5d32LspnWLxG2cacga
1xktdOmThghvivkMaONu2MeDgd1DXKihfx2BQUGcmdKG/nDf/rVb9hOj7ADkdXFU
MBZe6sviTFIewbeqidFsL3bbrcFkBQuj/G809vrNe24hqPn2V5qECM0+nHhzJluO
CekUyj8vpd12RcygYzMCMnYuChmukRZsO3SVGle/cGmfRJRA1pEf0n+SeQZAKkdS
6FS0YJUnjyXov6cmH20z1NRux5VASFsHCFRyTmeo8ehBHP68So2KdRUf7WNiBlsu
ETzSkevp7XBbdeydVUxUzBPrMsmNjA1CD6kw2iPRhbFD+8efs7tK5DQnu6nd38q2
mZ52uFUDg88VMUyy/ackiPE8Fuc3MGJhRmeb8eQxL3hgGnkz2RoEABmLz6drySvl
6X+6EKcnPBsWF5Zo0OHFoc9kfA7UXNkDI7YeCQLNZwhph/aAKjNIBhFEn3swfwZI
qSTRGjCyu6bQ/YyRyhst+BKJgWCFV/lS8lbyRnqzlXnrrrUN7sJlm+eiotOCOUn4
DisrpKGRyURqyVDyTwnfE+TRE/IIBF0OO3YGALebitP/ERY0n2wnO700Byjt6JNT
USMwPaSTUa8Virx+KA+Hgvd5juGVmUhhW6Z8ilviVpJ1Hto2z48jnPoFJzMfGiaR
GT10Zs+XoKEWf673sp+26b4ioDCOcJzUlROsF81RGYcj3a5J0IdXqWhQ6WmoUTen
GYffPsi5tMGL1wEaJlJfcFm8Ge9gaK30hS+0ibzggVdp74h1/XxuB2htNLAygtMy
HdFlyunfsBjVOt3eDnLr3h3u2P26cAwPLxdR+kqsmFpNccEX8ab2rrMFLc4JqZ2f
ysT/Cz9xSeWtv6CCgTXGmcJx+kIyZM+iBwh575zvtsDiiJy1YSCoapTusmx9kyxG
dlYHEyf3l7b3rJwg4K+TFYGEAwoLMwTTFEzQhdNsphHFgLE059LghlieN7FUXM/L
WZXW0GRr9/kZKWh3/OwHQTz7RMf34PLhZP4vgPSSm+iXyLeyiQ7JHAOqnnWSMOvA
ao5xaThUVot9PwXcBRcF4oi8aNyFXDe8+x4xqsYoRv/9WOnHCbzfX/IwuhHNt0WU
9bCLzWavJsAb+qjAmWda15Qed084TbNlX7F9YCg2Y3Ie/EsXy+G4QmkKSj710xsR
MoPwJzeYpTg9rBFEnDLBSMaXDqPTq6ufOQ5z8hWsl0sQq5C0epvbqpRfZK/g2jAV
Eyq6ldlZtNmp2Q0+NWIs2mZ33PJufKsHDMP4jnWKNU1OYO0tWUji+T1We9bX41Fb
rRlTcV+7PvpAPrpvscWDeLDE4geq2OdMAN3bso2soOk2Rssob6JiS59iVPihePKl
UN9/1HghK+v0bfixsFE3odoILP43VwuY+O8JosOJHhV6Brtoo29DSKP0N3HoMi9Q
AfVMkzG2rfNNh+GlUGU6aHPaxaAMPLBB5vWAqAs5Rrw0gASrN5RY5Pd9Cxo5GZHo
ApInn+ytST6fdXutvN20ap80blhp0LTJ/XUYvOKCprZOvKbI91LRWt921cSulbD9
p8OFa1SgVbxA1j7oucqUNTr6Lb+/O5iqRUBR8jdMSd/TeEIjMFFZKWZ16/tqHuCN
1C3vs4EmVd8BoCjaamNOxBUYc4e25MvU+40VFA1+COKenVHv04TNOBxhF3jIdtv9
M10H/XBf16aooXPLHt5UsVC74u729kmD56PQs0SfOrXQa1vuqqop0h4cyNNiDidx
akv87yrTaD7iVhGUpaoEuN1aq9R4mF6rzykTXfDPX41AcX7sXltsHlaqqBj8/DZS
9/vTYM0EDZUML5bCNwCfydmyFCMasbWLsFbZvzfDqvVTOu8zfRUoN/7ImfPpIki3
1FS5TyN7f3GM1s+R8iX9Dz6ME4Xw4pZu9ypUIEDeDEvz/0F0/zezCGQr2wN5Dfng
ko4Q45r9zeNeBnECzjcccYEURbIhkM1W0Xjl2rwc/dMgkWoMBUV0kuN191DVeld2
cFPCzjb09eyigx4L2wXxceOZua4oF2ZE5FWBoz19fXOeQMYRwAxib06N9NfYH/f+
sDAb5pOiSFq4lkaRM/6f3+o5o+s9K33Z9IaWQgxFAod1dPcrNuiVLXtgvByMgcxN
Hh0lAY+WWMAPYlxPzUCWHmLQkKy+ptgKGtkv5vV2+avCAY8MMv1KHgqP9USoZNCV
mp80WyJTmC1L7rWxUu2Xna11tLNNdbWC1uV5oOWbQl1C8cbknav6bqFWtTeMFPI/
eobaS5fZtOwz5tyX7x4WjyI9LEz76mB68L0TxPararjsYP9r+rWa2fyJyZrMrE2e
M/TCfKK73yw0BkbaFF91KtF4QxJwGzovpqqFO4ZeNHB0hJYtgpd/zGRUozeNrR/l
c9Ws9Syb0iSl0TWmh+G+UTm8apMueoDLhd+pDFNlAWGabxWIeqfr6c1ENp+ZC44f
DRH0S3koVHo2fIiUUYW8f9PuN6DLLtaEmGxzZ0sveuByAJunpQiI43bN2NS3hXp9
Y5R2f66ZbJZpbfE+7h0W76YAmb5DPihDtQoWUPywcdnzdFJlEyOTPYt0K3x4G/2b
bFKj6xnw078L+j6M6kD4Q+WTCZsl400o3GsJHA82jexIRmCql9VJ1oZIK7yTNFq6
snXfgMwOsBsrFGyY8IrFNfees5wSFyD25kZDzfTFWnPOhvCnjZg+cPMxB2PZtmah
+mp5UUhtNggvaeTDFY2toRrty8RCQ3FhWWqFTwQjCOvAGWF6Gw9wKF8XomZhbOx1
D2TYzGHo4l6okQDQolv0GLZRwTX4gPr3E2kqt/vdTihu8u9h/hwv9BnaOJONoaoh
+TZmCNRlzcXp999SKqhbkFuinUnmoO61E3BhwYTVfM4wsYUOnMe9bZz6yMJkxIcW
SgGfgclgbZmZdF4BlqDIHKPZxW/yG0bjhR5Rz/S3GArNrJWnIBS1dqlGC4BpMrcN
5fWVKBVbzrrsmk3InDfQjN3omr5yLXa9XoJJsPWrXxbWNZSWulG2sG1yPSyk6zoO
K8+qu1b8NQK3PsgS2s9uHBIoHopj1PjR3UsaRjENvp+wW2a73GSuQ4xeaowoqcQl
xSGdoVdAoDE6H0V44mCUsGY38CPw5iIHiV4gRbbrCXHIbSd5OPunOus/5ubVKLcW
xS2scoz6FYR/6KsUgwHG5CJz3VXNYsN9QshPwhEsroRAgNl29mdoj4hCMt4zRjhd
j/KbSngI4J8rwHrfyvmguEZxOxk0rNRSsmcvMBMlQQqE/09KKiYfU9P9BK0Irrn4
naJ87eR06CelB9a0mTfFatpipLTycHtaVfXBrOPndkJnUN7jV2p58jZAyz7IsSc0
fM76U/rWea8hswZ3kRpljfuLbkNCfhI/Y/atwhfHhbw=
`protect end_protected
