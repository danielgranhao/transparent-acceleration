-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ZgQO9Qpz0w0POD8yvG7k7advLKdLLpq+cM6h0dGNE29QhIconNt91AEBD2SHlA65
vs2nHLldSc5sngeyE/3GPACNZEQ+6IxiwAK4kSy0zkNQ7brM0U43bPW6wg5skg7V
7f/1JsooVfwDf8/S+zDacYGdLPyuMy0cnVSroOaGxqE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5458)

`protect DATA_BLOCK
ioAeuZfVt6Y6EKeJbEiub7vk0Y3yKCOW7CAaAOwdM7/DwEgNGUjbv2BUAzVer39y
eOldvsF3vG/6gMpBbcQTxiWhFBAVCWpMgNiyxOqu2uIQM50rZYt0WODJhMfqS818
10T5DctSH4GBYhtqqUcZIQCovbi3eMU4LZ989ua9htO/M5nYa/VTGzPKD9eBPu8r
fyEMffX1i9KSV0Azhh1+T70jyaKGWTmITN2CVVTtgFMJJ99Rh1MCNF8zs1+H/C6v
RTBdUO84LRAXnJOXK3YvUSrllBZyu2hUFJ2IlFVh3iQnIV1z7tmKDf389uO8AZ/w
cH5FI6f/4l0pWiGgXjt/2P/4+1BoK2tOyp4zihD9pFAfBFhGO5v8UjMqD0vgjZkg
uSEXFqPuBa9VyBiEz85QhU931X10mUwAZHYSi0GiyQDNCjcPZ34Sou6FEyn3S4ko
1d7BKiG6ySfSrFk7VZo98MRnbSzmYs/BVWyWtFFVdbssGargKw+ZsjD4oaNMf+4a
up20YGm1ySdBZny2D8aNzH6NfbWVxQESallJfMP1SYMbHhVGJdxs9lfYx0aRkbBC
sR96lmBon9nfm9ImRfktxqr7JNIm7+DHy3iNL2ZwGYUpirw7wFF5Bv2RUwdV/YrK
aKuMF+IkEd0P3vbR+SYpBRkFNCh8HNptb3GXtNXfa02lY4GxUhFaWuW4312Mz2Bz
MFVXHZkJHJqzbJSYhHriAOUZLwSu+lD4qooWZTJyAAmuYB98zz0kRaZBUvdCMg7c
9I2ibuoEXaLsofzGKOHv4zcPRht30NMLdl+CJoHMRfKZmu+wgYe8m8c7E4h39E3o
IPOzySOJWMrOCOMDiTeO1GYb+FD7QBgb+jkkMHnul0RahU9mtNCoQH7riYx11pnz
AOXfF7hQXaj1SrKlKd45o9HwwEVWOKc2OpWh1Lvb6LPnI37EuLTYhdSbNuEtimYR
zIC9pizh9HXuL9VSlPcP944wqg5dXaYlnykP5fg9mi05kw9NvHJO9opVuV9pwEjT
pUFvIl8WZvDnjR2S1tnIsFY2XUbwJt+JrOAKppIrrWjy2VgT2XgQy/OuroOkr5mm
WhFRKwY5Gm5JdsF1QG0dYeX8XjbN7jCXvYkmpmOZXZhKqgWXUm0HGh90pEs1r0Mk
NBENBDq2eIOnLoXwk+AeRkEfdjmZeitKlqd1SYeDQOwQHIq+JZb+SfDlSPpCo16J
DcjTo8R/UPA+BnlGDBALwV27zsANj/R45lWEjKoWogSeEcSKGz41o2fSeqxYWfU1
uoK9iOdKTqVROeq1vRJbGGQpD5ZOcoYEgxjW55tjRQwnBln/Na61LkZ88BeJKnDR
sMw+wRc0J2MHBPEMf1NN/1+MZHF7v1HUpQLkteDzH9ldn+hSfWfYoDSi7JGFVPaZ
vMO1UEvsKo1qoCu+kOTyFrSfuDdRX/23O9oJZHckLhmrvGG1GZzxoMLgwhdwxw8v
BMirNRG+A4HG93ecBmwppAKMhn5VEUDL3Zn5ZJ8eYKV9PGPLbA+GkVwAnzfFxm9z
kYyIEpHDzFNHBGu5ATmiLoYMSTnyDGDMlX7qWmWEwsYxzSH3UMvDahcLqwpi0bCv
Rk2+pEaSYRK/kUXG0J3c2znVUqu8AocC+NWbGxNqr1A1WKBOXnGfm+tuuGgOocBa
CcPqBQdhUVcxdZV+qE09vTlfSkdcJNCQfJgwNoBclN+my6D1qITSRZ5nj1kHes2f
gYY9cP1D3+1TkK6tR+0XeMffaSXy6rIrpUCyHk7ETJawnGlYHXrq+PWmlzG3uwwu
ntlF1cp6UUxWDbFMJ4MgCdRmzKPq91rvWzOUJKouP5lBCvAulnqQ+XAnJNxUxJNY
1FbD8eXIM2qUKZsRavFqryN1h8sxPoGus6KIJdKvWZeTN6phHR8/VQSvf2YHHzId
MWfwjbgvzcK7DEi2ryxz4too68hlXmk1Xb0rk3+hsdnrYHICRDMC2KVOF/0BqpPS
EFZZ762MFgIQodU/QM9u5c5g56GiPCOGfdJ+oSuFQy69eVbtxTFvDWJKkC9LrSNo
AcPaPFLnBuS3lDrpkFztvKJ6JfA66dBJL/d8lQhhSDvccfGLn7tVoAMtzScpUB0U
JirMNgz/s/EimaLll8h47NpmwhHhq4CnHQ1vy4r8ursPd5DPOnRg/LiKc7XHkkSc
JFFEVLtve84Hp0Lg40+Jl0B06JkIwQpz7BusY0DbQ7XeV9kqSRNx27PvXw6XQnEd
uWIUWBf3xpQ8jYrmSqNccVn5D2ygIp5a2BHo4N/7Br8dwnasXwAF9bA9yyqy1+/N
CtnKN72r1R3mtLVUBJiYbZEsBdpaGLyxziXHVcoAcFg8i8vLErAr/JjCEE9WucJj
pZ60B6AR4Fp9a6gJRtGqRCCkssTEGzA0FEUqgftdJHAhgE/V6izAJEgJBlil4l0o
cIogX/84Czud//06F5bxhSqiJZDjlU+H2/HJfeeY9uMh3O/ZpD1a4UrH609KiJXF
ujK4Xjl9aKyHYWkHlEMYug8xxfM+zpQN/sC5t0zuMyuLDeUn6LPi0d0TSd/Jvsxh
pSfjmhHUvgASSno1GrGYoYawqy79Tf0XWmmHesmoIDxinCWv+FREPL9Z04F0hp0j
O8O76cDfyh4WBA6XH8m0zIu1uwQ0qThM1mM0zXaWzspSFnrbJhMVZ6zZX4IHs3yu
IyeUAG/Hlxy7+hMAQDRBRj//IEHayzw/neGVj0bxsxaQu8vefI1y6uL6q+TaX++K
YsNZSrVDR92AwU6yjMFQ9QFyZrFeh0PFEmMPmlQ9nqezLL/yl8E4bNExmPn7bOrA
kvRQgT7V6eG6XKPWyqiqfsvaLF9hWiohat86BLJKVj8m+1tlr80r0S9UWMteOaXB
lL4mX0EW8LIUGYJnttzCqa/NrE4XyIDNkHCl+pPqbzGKg1TGlEgoXcO6IcfDZ5ZL
3LzPVVfCk1lJXs3JDLkjSerwUcavzgQ1+sx35U8o/xtpIoc2sXMgZstsFPGZSiCH
sqDpwQwzWp4nG9SdA0sVuX9SGGs6ntYln4F0tjh1D/9iXGOOOiReNqZcOKmvHU2b
fiu2D9Y6CbY6RPA7KW19PvK6q3wgndli8vB/yUi+6jKFDILO8/mKtVnqkFYOr0we
N0qsSUC5KMwkCbc44otHedq9+vEcIwmXABvmBwzSM60x+mKjv/VnjNCT3/2j7MkZ
K05kDJRTnNYSl4GHTIHH+z61vgRHaBBCqGcN0uQEBdCpwTGaGf65JAaWXZinie4R
ri9/gcjFCdRu8q1TSvo6X8wH4ZUhGoOPG895eMzPL9niVSi55mgWOUIdRfzTLL04
wqKMVyLHTM0dPkgKsBPM7Tqy7N1xjFmWHNby288eqP+6OfiTM1Zkp9Rd7bHs6rP0
u9D731eYBKCsvODjmmLC6G3tZfXyF+Z8eWxSuWBgdCIQK6cx3eF2rf8xg944wgQ3
qIzHlXPTYcWd2p3tDvFopzU9mXVUSXZz6pbQ6ODB7Zdgi/mulb8dcIkMDE2tA/Ln
S46tvHH72d742pYjCub+E3JwNfVq7WBc001+17p2xkedbsBvvZte2YA5r6fP6wO1
CPOkGhk5iH4nFU037yFu+xhM0Ih4AhLFt5IKFzCA8K5tkzydNZnCDW/FQP+lbhyu
vgUUZvbsHqNfSavXPRlbz5QguN08YBEaPFaF6LkvNHJUwS0VPzE9kGVIM5XOdIVF
oX5uszUJMZb8pY5FLC1LxAAQsShFucKK6b2fVxPKDaW49P5j9AmnuZ9YE1BZzzOF
bSp2t5UoDp91uIsLbDmwCZ5zjwMgvXmMrnVYMn9/4DwTsKGcwjMO2YNlT+wJloTN
5eVUGK7VI2d6BYa9+x6NqZwm++apnzdp3UPFyOovasQFEv9qgrbnudpB4n5X0/Ec
Km0TMSLji4u+9r1xoaJeH6g6ZImKH2fep0Qab9MGp5LMP3nOu5UtWPRxLYZYC2NK
7Qj/cHZU6qM5KruzNFkU38i6sYWxfSN2O+xWdlr+PELGJSE47/AP/gWpeXHGU5yj
aci+8uAxK51qMQtEafPjCAed+n60Vdt5axDcf01TGBcXAMFSNyui3B7hPGBSKU4u
7DmCehX6luIhtGbCSq/6/oE21Q7Un7MG+bsLZo1dFA6f/ER4O4o51FOASI2S22pJ
ulwN+nHvu0YS1sE2Xlffq/qIzR/kpTYS7ep4rgnPPGBweRc0T/Ab4WVtDfthcO5Q
BsCpm8B7CoAyCfQolxewZ952oNs5tV0Wu2E1JNHtVJ4ifvEOZHXvgpK6GRZauPiZ
XAkZVwP0+thZloKecMlelkngS3YCzFRCOCBjF2472p6sNlc+EbuzWPuxpCSGtVnV
eK+VoreiKN/gRuLB5ZiI86dCy7qjCl5h6kenFHVA5jH9uIFufQr9Se3BUoYz3IAz
frbChFpnA1RYo6xfO7Yj8DyGfGfa/ojXZJIKb32HfI9fI6RzlGPbmCSERxzj8+Ar
jdoaNPUTks1hghfw2JLNiWYYGTMuziVOUXcHiH34zIZQl0aFCHWev2Syo4TNV6xv
BGMBNBAFAy0Ycx1ehvKiSAnpUTlqQhBTOw1/T2ksFqS09hUlD5JcvhdwIqzyTQ9v
zfBNCQjR8HajyBL5cx8FfaOn8R8Gid5OnVGqZcF1GRyg3FmVSNIxQkvo1lGo6yal
SIsC5vvGZnsV+ZigAi7+q8JGdZNWKetLfjWm6XUH75Uds1DYTA/o2Xb9xH56wntO
s3e2Qzn3yynT2d/6sObeaFA1v5+whpg3gdksS4C22HxOmOSSDzs0LSbyXhTqLCil
1BQsUOfPwiDty9YFdLldW5uFllYeTp7wvFIGKIJA+Vt0Ad2DPmF9D7IbXW1kVzxq
bfakM2xe22/th0cOpvZWae89WZ7hcxkcm/2yEqggEtyer4K1M0N1GJmBWqBzpbpu
rmfvDV7NouJNMtfRFnJG8XEHwewzk9ocsJwgRYhHK2O8O6FseHYg8RgpDAynDSBW
PPaf/WM1HOjy+k+ZnS4O0eTgRVFfoega3YZRBTIQMTZjB/igsYDQjGz4gg91eGWR
u9drffDDHG1cG22euC0yXQraR+oW3xwe2Lkomi4BqD0GPNWetj4nMdcWuT4QCj12
G3KRjjQJd9dKdYrI1HiOOMBXK1c6z/54m/XcCVQc6y2YqHf0t6R7txgHZbm7Kw0Z
kNMhmaVxbIR6rvQuBvrPsHFNf68y8SAzDFL/icmZIkF1+bXh8OdYMN/9IHOvZ6fJ
+Ndc2Sep9G5wrVs1p93TkkU9we0az0ZbRE4Ai5Q6arWed6JeexSR8nPgG1JrnQkZ
DSRX+poIMyrhYynov5fST4x66ycMIqyhgGPdYCubUIVAuw1dYdFjHdRONbEsWkee
JhK5m2nZnJy/KPCAQHp9brNHPRDjO2CwBeO3IzMM1CYBrxpmU003Q3XcsHn03Akl
MYi6hSwZ+SRahQpu5KbTCLWwMT1GEKQkTAwLVYLwGRs7TUzoRZVCgRXEiaiTGSoU
yfyli3HiYj7vINhOle28UajmsuIOWODlWka4Mnf3IINtPF6JScDnMeAv4AwJFD+k
LXPijcK5v4JYzJDJiKVc8fRbQbuUyA6J8cDlQBDWjnFbX9VNPbngvYMDJg9HeV8z
tc0XwF9LVEB8EkraBHDT9Kqj+UOhTqLuNpGM0IEC1RRim2Wr7bauUzljX8q9uVZU
NMzB1oYbZsVwxya2ShdTp4jFUGyupH0n5LJBSMTPx9QA47JPr53/kPO43dQv2pw5
M2qs/iMyZarRil0k2tIkMBNj1N9BbxSpJ2k3/mKWiP0e8UwXTD2/dlROl0f1iYiK
PSdua7ml9etpXus5XwqCeZS2W4ECQTNQ+hRrJTfL6KCRsKmv3BIVzM4Q3mpo+PO3
cyXX7ZrlZBXuLEpsujqz6SEboEukgRK69UxdqrE2uObA/xGuCaJFrz+fWBl7pq3/
Md1lR6UKMKf10pMszSef+BQFhBrKhC7Ov6C1W0uxhu7Mr8EkoXCQbpvvUburTkDv
dtAcIXkZohR3s+BY26e96bcI7LtGv1HGAagbF1n3Ii2TVSuiCGkMEgDoxFRbNqjs
katiqK1XErRLCuUz6kYtKn7LemrFdEJrIfqXjsDZSlxQccm8gzbn8NObYYMtxDnH
ct4ZSGdaDqvBY58St5zW302cGM3IxWpHPtLolVA2WP46RExvyVUpf20N1qlDKMTt
Qj0asCuL0P34cXfs3U2SfLCzES/m5Nho5zgoadMRyA+tV0PdSh3Df/9HvrKjY1B+
QMe5hNV2kGv03V3AeMKhgn8eZAiA+p+QlWvf0il5xCqZbeFgw0gwutF1/08cY5ne
kgIDYO9/Plza0wmCqh+1/EG8y0VpERu2H8R242odKkktpewxbnfNgxuMMLufJrDf
Wle41+4eRElepN1Q7ur9CeHzKCNB11CjH1TOBZTXi+rFV3uDxkjQdrnk45/6ym8e
srGPjbbEw3XlnWwgBCNaD32Kf8IfL7MxwcYvvH/e/CsZERII/cniNF7uiA1D83Og
j6tksqUMak9V+Ep/Rz3UUcgH7lwF7JJ9S+qFDwtGiK7s/Caw7Z/NmqHRrp02Ptmr
x9YhriJLl8qTv5Y6rUk/aDz8+WeetMpr5rBLLLtYUDrQqw+yHocqq4rQiecmBkRd
H7/E9YQB4PpDW6Bc0tE4rYuXqVW6wDb23K5qngJHIjuMiebsim8FTh7pVxGzeQQB
oanjQRaW74Mo2TLwak/7+wei26Sn0f3u+BNkvchqZ68HsHjBHmthQ9VkMbdjM7gA
3xpOrXZRqdlbh3Duav68bwaXesYlFLk248y0xGgVE/perP28kQn2Ketb8Ivpvazo
t8QIAQqxVHJhRyZ/V8oFwHASiu+ctFRquvxQXFWJwWwkGhmZCZb7BXq1VQfuqOKv
aKMsRB1ZFM4KPK0vpzV2mNHBaTMTg9Q/MUYG3fv06QS/IEiIafDYT+w7vtF4q+ZY
Y3zsdKdy4xM6jvj15Z0O8Igdea0KAvpVeC6GWd49L2ITHfiKQfU6W/uNP6zF9txU
LhHcL4/NiuGhmf7QoHknt9gsAfYgOIBN7/SwlYTzgrZ4p5dQ3oGreiejUSiAP41k
diagJUdadGEuFbfyiWHXerVKhsgS21msTOsnRTLtGIXMbk1KIroOYVDm/8ONjeuX
RQTPHNvQzWlBgbJQcKqX7F0BPd5nJmHnu8oRl3XLJNu2L8WZ0/rnDTkkfD4/oXrF
/RLLpoA9dcxx1iS/RCMpV72dUb4Vd7h8jBITUj1bo1SOZVfVrj3DCrDVBu7syxXN
GKMwHNHF4lzEx3kDZ1Xjrw==
`protect END_PROTECTED