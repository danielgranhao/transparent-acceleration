-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fcqFEdw3+NHq3thzDpWUDhydTZrPDdb/npYT3slZq50a9FiriK2iAfFBseI5C/Tg
EZe6J1O3BUg+Jr80zbJ9jn6CfkpPHE+WWRhmzUOy4I48jJPYfVhD34LBpXnb108f
IL7LHYufZDBFGvcRVJveJasKWarytxiUCv5FeiFbLdo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 11530)

`protect DATA_BLOCK
xOkR1+JLU4opuVF7rVSSwSgzndoHz/3dpNYiV4TCqqtYqYy29bANMD87tYm1xcQA
Z3v+GM4P7O+EdhlStEoXqvIyv6nX715e/6ppf9irLq0Rmhl3IHtAZsvC0jrOaeSW
Gd37WQJMCdHXq3wBuym7qfg4oN0enpAull4S/MWr+E8KIxz3KlvL1dtm3fd5mcPj
mvEkRV6sxSqRO7Ni11Zju0rnDePBBQ0+EvVtCBheLKSOQFpRd8yG5vkDRf+sM4OW
kgt0BJ+uBx4K7hoDJZfDSSOlzf0pvSbYY33W6eVspa7xpaWK7gJZESryG9IbnJxE
sbN5gDb3yXV2Fcz6rl+I6YCuRh1Tu8ylvfhUsx3ywjrPtWXuQJuIiGt5L+lxFMYN
tz6L2eQbzi2moyWhuS94BPMqIx8IvJCGIvLCRIlGGTjO8+osuBJfmNTjuVerHgFE
4Jqtw5UQL5I2RrldIwq0FBR01vQKFG9HAcuuR2EIG9m4ZFsalO9j4k+i2RPRN9IH
GOnu4Ogm/CF8THsvrukqyottfzYn7GiztHq+57HhR+luml+T2+FvLRfJrEGb1MgO
9Xb3e/hnSn/u09eeiH8KOTWJARz0iWoNBROpS9J8EnmbriO7Miy0a/oon/rQoja5
4oawBFrH/v0+8F4DCrgejY4HNpW2GtEUQNYnKELfGZT4XqssBDcKu/CdmVXLi52n
rSjuWTVCL0l7YpBFhnP+nGB1whEGUTpH6B9mCpf2HvX3gPQdx5cDQzqV7kUl1d3D
RRrE+y4zbJrMomq8zTWJE0JvGMHjPbepGZuTdIq1PPzb0PcWYLKHzwKQEwwP5PgT
Z6lxwT64A0VQ30SRMoLa/MBoGlVGuncOdvBsbcJMNZe1gll5YuatiuUpGqRvLTrw
M8+/KT8cA+clWQTNwA9GnxWijZFzdrCFZ/DC5N0ZaGaGR2cimqFVny7D5onkhzh6
wGFcTSu4rSzz9nHe2qawubGO7hoFgXpgOwhz7ju9yrszWkakdzn+tldjWrRVVjSM
EW+wZHIv4mavFL1b8WL0h/9T+Bmmq2YNBqe31UNV7oNYgwbTNymMmh5pPJPyQdQs
WfTHLs9M57FzEZGAcrbdWPXrjwSuO9M5AWoFemrYRgypVN9mGqhs7/JZn2j6Ynwx
ziqwEZcvMvVsxaRGGqsx1Re1k9k+NIv285a348hhYTkcOlpbntrL5hIUEFMLJ0Pf
dotc/jH9pCVI4GyWKaXJ1Zp3jtEZPgE3OwNVwqFgxEH3k8CSUMzoIvam1twpV8y4
1ZC8cgYI4E+q1JLbNd6XN386pIWor9+vTLYVoppcW5jxpgbRv41okLYkEUHRM+dm
vvfh978XexYWpuEY+feT5LnlM4z5tVQkKPb096jCRLBUdyYMZoUtLICbKw47ufe6
nP0rTGZdGa4RR4pTzZnRNXHzIwD/VVwjO5h+zE8ggLzIuJIqANHpfGkeYUaabOIi
Spw5zAVumzUYXr9/rURswIvyvpGlxhJYy2zZ9MrPRJ5PmqhC/jMFO9mEgyDy1vMQ
G46+2ZAF/DgwQ7EKis5BzP0/NVckOH4tCLO98c4B+TBKU/d2vt4J85pg8hD9Oj6p
ZsRUY5bOYjgqCYEI6dWI8jh4SHY2IiU8I9hztWZc4jALI/4HOhRYHFVWtHgYR4av
1raCIuOu4/3Odk8OMpd10IGbCmbcLGNmOkNKwZ/OGc5mYpNBKFr7gThJMTDCBUGw
T6aLrhtW+WryhVfGBP3W6q26bpj6qr6rb1eAmvqCiY2rxmxIS3NuJbJbhc8yRZGI
dG+HkiISYYTn8ijIW8HRJCulva1Dl/vyiXZ7hl14xbZXFPhX2F49cCc38uB0HynT
/WQRTZ71KB+U0Y/ZWu84mRyBf2D5jCgI/f5fEGr6inGpKLoVEOdt4L+wqM/neaBq
Odzet5QkkcGe/ujZ7cAb3ckTiGHS31XZxzgmUegeywtg4c2EjEr3W8CaoKESOz0t
qBHKwPtpTZ6eRtD1UX4Giga0MStbmAm15dhWSfLH8oUs65B/S9tBuaCCvCpBsaum
l1fNT7cBLkJzvvGgGDwS40QHqeRQ6y2j5ZktSLKKjaFsNsIwmHrN71SkLI4FQakZ
xwFEiSgCulKlexMRoJNlskEIX1b+0MpCS/4mfC/WDB9ll65sKcvsQ0uqxY2iHMrN
3sVLsrWDMitI7EGYqFvtL8zxQyXO6Y+wa0SgstBLGeyt1RBdem5csd3KBeyp6mc5
E0oVrEnZE3TeYroB9AJ72KY/TpgVUyUHHy11U2ciX8cIN3pZu8dJ0Br8V4h7yljh
x2Z9b+/BGScwvW4dAyb03dOgv3w0ddsmaxIQ4GnSK6QYdvlqBtOhtKyNjEqALnvu
nq4nX1SC3+lrd+1amY0gX25juwaciXNluKyIHAsbvUkFjOQPEiroqVzA5rYKTtQB
ByRUM0FLiUfHav43JaCB2plbguSZFhTVx2iqZKuwUCbftACiHoark5/2EGbp/Rtw
vV/FU7a49/O9jzfrYROEtPNneXQ9ceABygf5BH2Sflrzl2+eJhGJNvZBROVENLPq
QY7k9tIQb0rGFIiakMpRBGswfPSLZM+Yzqxc333DTHCgvuuMI+tFLDHPyO4y8X6i
grO+tn2Ojb6j69MVm4QAnbjEjLozywt15JdNjxmGkZaONDaS0oDefdy8WG4AE+2t
EUCZBTgLFE1QqM0OpHh5sdtZRI+18lCWE/Au7cvc/5atia0Pt4CXJ5uU3m+Vtr+u
Y7ZUzcg0i62BYia2gkRrFWQWd3MGYudT9lm+ETSmcH8Z7s42W2PCQSTCe2ZilZAI
joog9gH4mY+LnzFo5150KBnMV4lRNjAYJVl4Kq54t6BxXrJCIMbaYj8ARlJwwN0C
Ba9+db8dQfRQ4bQVnPjmaSD9RB+hf2WnVo+MHmE3owF4/CsHHPmE8aB6lWTTpsYp
61ptSq8dFqQoNuDTmVKp53BAv+paesnObJFCpSad4DzElJaJZE1pHm4KU60aT1TW
lgaBnBpUmx8p2NrxOLK4VtXrM+6XQrNUyWna8RM9I+wEkftVNqw6J6P8eBZBESrK
VKbV6z5mPqqQ2Wwonjs27TgHH6yzHHwD3yXSipyPNZwr5xS9PJAZ6gVzzs2lykA9
e21SPcw1OEchOSuC2qzTLI1lzVGSY4qiqYKf8kDpMApMOMXkia5UCgk/CMD81DJ2
KvGT9kPXhQbyi40jlYk06qbS5UP+oGrcSyf4dMrsVwnI5k6fHDLHeW7QVwWLsm6D
tH9GJxzr8sNYc30LhmN6j7tXOMMa8PO3SwenYJ9kDl7xEzfDkq9jNpGAs0HcqOr9
ftr9BIWlxWWx/5PBESYFibMQ+WbSAwcNzwjvJZnqtsf+EiaavONMSfJsYIDaFBcN
FvcFe/ahNrl4hbO+CTdNuqXc/aAYy1Mbhk5TjxXtuQEGAi7qCyLc7kR9J/mkTzGx
jBel6BgY2q+AGo1o6Gf+Vrd5Pf4zJmgXMnzgBIR3wYNy7ZbJ1klA+vrPLIpqcbWr
OnIyTL0Dp802tfKpe/67sRyylrZCSkIy+ArfcCZIzK7W7e/y2S3Nefo6tH9XB+wa
g3Fl1//EBvR/23F8AQanEpd6ayhutrY7VmRjAN/TLsr5MV+rgherM2Joiip0Fhie
3zSVnBE4HoAs22jYGm6ny9oVBtstzlNcNCp2pIyEwq90sifFBWn1W8SdtaUFMVTL
hEvs7MgeeJJ0GMT6VHvEQyeX+JXZFhI+ned9mU/xTJpDTiepOAqlzJKS+qtDEZ36
tdMJpeHOk8m2k4OAzRRtmmt3i8nwl/RxdGhDnbz1zqQGA7vbendVqnWzB0nBzeXz
5YX+q5gyI1W2sHRhdow+GC+Il1ArG4wt5G3sc4uZqSOXlanLRzLEINKD3e7+IaPR
bjpkoxvOnJ5y89Mhw6M+mUPr0CYYBU3OXWJKA1T8Vl0igIAR0T57clJbdEk14eqA
A3qq5pzv4fcURc9WxBsIhmx+QvlLYw/QQF4ITdRVsf1gbAN5htfYNq/aKFbZd4ZC
xxuCiqOhQC8cUpYiETYZVokm3C0dfeonzIF6C5cRa36zUnuHRMVNuCpAxyyelX9S
0q0KkAFhx3uI4833SpmC8PbwH492ubahnEZq8b05NPbfG2etyWyCUCEnWgEKaEgb
TYxUAGA99ykgj1u+nw8gIFOo/3UKY0uGryrWrekgRLMWE/09qdVBr4NR7A6EYzl5
SpaquehM39eX5rkd/wRCMZGcwuLKQMu32d3C/hcDHqNSEQuno1zHP+X7kIGDwiOi
F7YV67W/uQpSuoHVvjM3HhZMZmg2r733P/1XR+PURcWgiuRFE9lts7YWXAN1Blia
9c9CnGmtd7M7EJrn/MzyZTcps24wcf1sUER0OEvHGmjURJ+nRLXz1xBzePg5+DFr
UFNsn/C3FaFifOVEDarNlJpuj6+XHRQMH4Z8xVs35mI9SkDKSLXPBf0JPk5n9UV+
uIUsE/aQjUWDdb0VXbrWQ33QpnJmrsxpBbgztHIT33TUgMIBEWvk0Namsn2Icvii
eU8evsrONdO3BZqq+JHlHozHvI9QqZUkuyXpeEUlmff5GEnM7DBCXPnlIiNvOdTw
p2Eys43IoZ25ItGgHoF/ef4EROakVAtr6JklbWNfh4BLzJF4WQvnGvrXqLlx9cYM
1Sf2Rb2yjlpnCMrN5Yikdgcj3KY30Gxe7b3bIsp+jiag8yU4FmjWx3K5CvBCXst5
Ch3hKSdYlPK0W5C5rAORPMjTXTI8QsNl1Yx0LK7xgQeuejBwY4B2wgaBeMx5/ZdY
qcyMeUDYBW6m26XCl+1e59lxUfQboSIzoSHJEg5ZeTUq8n5Lwws/4d7/xTBKp2TT
jzGu85IDSAUwd0g/8bqOQLmHns7X4vxz8KtxkXx5eFZxbPH0OvKD3jpNMiB+R01s
3hRmiBO148pH9pb5eyePKCtEV/EX5Cv/7+mGMDmMjvgIyCHqB7u2V32ZkYyTx55h
sC9OVZpMGzAc/bO9V5fr/PtIg7I7LzioYM+EOMX16EUwrTMQWkhz1MCkDvtdzAqT
+mgZSWxXsDEvun/FmQ+KsDrbHUqkssYZ53fNs15M954gHqVKyggsB1XmIUSUPLLd
oHGfghecllbs/vY3gSRseWlXIj8M0jOt+oAI4jleVIRLHxR0mWoWJoAP17QgVT5X
4d2XJsiaXVf7pnlRkjFQROVsQjRIOFcdKUXfsq6Q2fouv9yR/cuUsxzU95TpytF7
WYfcM5gG8LLgCLszJFFUUfIxt+7+hchJGp7AwfC3ZocVYj+8C+KxVIQWKiSNuZVW
L7CR8Qk5ySkbUTxZHAg1f4uudmsQuPUZOH1Oh2DBCs2DHa1D5N/Lb8HH5cOAktuW
tZDq2WWQMwmNghPSdyvzFT9K8e33rYUIK9x2fXOwPO37JGMY+4NF+oQW3DTRRVXb
44BgvEAZ6UbrmbqHvCRTHo90vSJb6hlUwWHpYpVgChd3JhdD1Ro44lkO5AUU1yQ3
xJ8SNRovV4ul8bvTDlYuZ7pDJ6AZSS200Z5BzYiwkkcjz6C/LN5Moe3fkKAihBkX
6JmbwCpATVXaETGZroLF7vTCgzIYGR2PcSQ6kP5uTqNVs1ddMaUb2w0mHdTusZb2
LRgBu/CNgZeYbBiKnblTzkH97lehkPE67E33jVcmil2mxPDlj8BI4K/93jDiQZLR
SJ1FyXrQXjVA/maCmW/MtQFfCrWZDCFHT9IMnzPGy45EzAJN57eNY+1n7V2kvZMh
WBIT3LD9t9uo+/mq6QGOcxwaXpOegLIuG75IuKIpzuNnEj/lGli27EwCy3hyCzby
XO+lISxkRE5Nfa7dSIKvMcxFOLIlnJOHHIhjfcWT39Lj+NMhj06LJ1EjoYrsu2W3
nm9CQ2jMVqoWccRA6lzcjQpdzw1d8r2uOpK3PIq/+E2EKZsJ4t2/ij/SO+pcWm48
cfDeGpvey3NWyBsHSrFuOCDR4A/ea5DlNmQkCTzbbkKI8bhfhUMN4j62V/rwTZo8
90MAEUAY01QaX8GrYEOT/uKilxUk6UCn8bMxeqkc6H4BDqjlDdZTpLyU4gYmZ++H
FAUZauIm38UcOesA1+Cf5JZvQWfJlN7t2CnPKZiRR1/3hN8WHsJyo5D1YfiWVm/R
YPxRU74lt/+BDkoQUMdaoHoix2qu/4aJOHbGUo+ODsal2cOScn2qnaW3NBMXoDMq
HAbNeHiFEEZivX1/K2C9YUKbVu5g5Gp4qjCdOrhJI+MP5I2uGtXV/rlb1WvcEPOd
qzvrUC3UzZ4dd00/niorbLry+ZALqD+ALkyfxZDbEJ2AAtac/0QexgxUtgZPssLI
7QMsrqOFiVatuIhZ60LkAE6SObcGGRZTO/qKtsCAqQEYbA6PskZCzoXeg962IwVL
JvAP0oLjbNNB8QWmIPt8HTsZNoOn2J0aF5+PBdMrV0GYQ7LBh/45NQG7A7g57G1T
9t7N5s6o0n0pise+ybC22HWW9qOro52yjOAdpKo1n93UoHJoyGn9oQ+u0zh+8OL7
rpdOevPMEZdcQdpPxYZVdGwetL+iLIKu9fPTGuXXOC1K35OXeI7PObkwXyBS0VCD
q+8x1Ub2em/HikQFMIl4BnH/uxo5/fsQTshkj3zWO8wOE1sXqdjo0GmMdntkyLay
FVdYF5W/jysKM73JjL4XNkoMiUAKN3eSmDltUzntAvh8u6Hq3i5bVd28a4Hp/bvC
WqyDhfKJk6dg6dfDfL8bDreKjufS+2V0W2C9NVmnnisPKUqVVCmXYcZfpTCIh6DX
sx0+YB4L8UZ1yCj7i8uvsKZ5R2fmL6utYqSc7Ba6KwjDuQd3ObKa3jm9hbU+3Ng3
iI0cMlxmzWcAeZ79g+Xh/Zwi/6hA63ySal2yjm8em/CbC+c/j8zG5xCxgzfwzCfr
J2Fu5kv9XX5PcsPPhx55yrZoN35X66+VBWX18Mgfu9H1sGN5xcUZd/1VRVLC75Ot
Lanl5n8Cfth47zCOlVNVtgQ97mXQ5T6+f4452lO2xnbYwUtQvMs6kf/pQhMXZWjp
/zHQ3l5GMz/TWGydgwJbt3d0NbnqCxRb0iPH9TFTVTFvOxz2+A3bJ60WDfqF2mAv
GZ0wKecmCU1/db1iXY+vPMgrbyxh9df4A4KvZUWuh9uvu6ZBWqePD+6rjmaKmib6
ZX71b6qQUlp6uo2eSGIsOr3DJiN4jk3oXLwdy6mt+PqSSSHojpvRjsgklr0Q2hyl
bHXE3lHzYUwGJKPI4bDGsQUhJZfV1h9oYHD318TbaovP0PlQHTKONLX7yGTya83d
azPG50KH4uSXAGgG8dJV1WsVEpmVuAELgoQ4JpJjcBVBznhyK3Z1ab9koiLFM3Li
nBP+NbRUHHZLQen6zjUJDmqEJPoZZscAhkvkdT7JqUhTOweABC0KJnpaRZv6Gaqc
jfzqp5cz8bG0hlvtt6yEabYURLo6Vt2sgpo+IVuZQ45r6peh/HoxS4o7CaBAEZWo
mB44SxGuXkgf8Qa1IoGqVA+ohDxRsH7ws3g1sutDEalraPekWpKpokRl9Bbruw5m
jqBjcrDID/vC3hL25QBQTbW0DHctvtOwsuYNGRdO9v2WmQKE8JNBhmGiXwSESeZ3
nzktGYy+8KXT0IMwNWB7E1kDwqIoyNqf6B3+FPdYGDHwI8K6NRf3PiNNAMJJdULM
CbYH6hPQ2vHYChInFSVSApyyUCU5FutA3YxKRTD0/gGfHdvvUIAdqvG2nh8C/OY/
HoouNVLYpG//xXz5ZDyvqLVXFw/llaoBF+WoFeCNVahhyQAyek7/BneTNtkPBI/a
tzKNgCzke/Xk2ZZra7V2NmjANad1SRbG/dQu1mmkOK9O9UzGeHCVMKi/ypVjrDFN
VGHMNewAKK9P3r3f4Dh3p5qTyiT2fL2tmrIVur4c0G2jom/1GvUtNpVMWHDd2YW4
PhQbuKsPhSKpdfExQUxDG78FL1gZB4EkfO5k2AIxiRYtSr7Wv5ly7Rgu+IUgM0ut
ZkPL7Y6eraKFGVgptvQF1U+BmK935B3iK7gUzav8YKMrHNNfcEkKm4JcLal8NJmA
9RCfOShk10lODnMRNhkjN4G9MIGclmMyMg+j/fMIRL0NQkM+1UDh7DxfB2jB8AyD
jld3m4tzs0poJ+AP0blkKiKNkBUKZgHSLmu1wr9a0n1zcqtw3Wyz4JdxEr0B5dIR
9a3cH0cOUJcwIYIpxJ0/Dd2x+TfcbhzLCd9es8QsxuP8uziN5q7I0b8CQNdHAZ5e
iRyEQsf6OgGiCw1jIEbZQJKdBZ7sjKNfnfUX/XpK6KtbJRJaujkEM7o9snkFF084
0mPgMLbjChukbkoEwIgtMN3Z1KxJnciYFHeDfcwDWgVI1qwA8Zr8uUiPmVWYD36i
Fc1GsTcxcaBNS7tqm9HdJexjy2yZ8Vr0Zu2XxlHf9PIw0EN11CoBnh4rOA8EBR+U
U3RrPz623LWwTEAmFPCXpA+9vUNLfymLLKHDGA0CFudinai5wenNgexumDq9IO0E
G8ZXixr7xuUal3f4e1mHpQZvhw2gyBpcXtYxbhJC2d+EVwN4Y8Slku2U9AYbJS9c
sgnGHYKqv2XWA/kFEXu2JUApe6k1ZyfXyKhyeAib9JFVVaH1GSXBH7wClq9+Qx+n
QVuOG5otGoN4l4vdEeYtIaqRJDtNnhaIze3SnYMwucR4OF4Xl5qJYViTnCNDqaR2
2E6brAYGPuwPX6rHoZ0vr7Cjt9svZcNLmlo0PQDk1tbGAcuVsicKoYbWDN1TwVEm
SypaJecyBGRe28VHNR2IPAtFftaE1RGyDhuEwkZrktcf3iYwG4Xnt1t2Ojm90Dvp
3tUv7U39+02GNavxHL1A3uw+mPghQFlGV6+KXdtXGz+ALcWpC6Zap7027V6/dlyK
9Je2x7oyCpmzrK4fPYNYuM04A0Lkn8X+a5q2I9m/FdpxYWRvWGhD2s/wjSNfHwCr
8kc/5q9VMZ2bwtK5I0wMxBh0UVEkPmjPVlkBLDCrV+KdusFZaH08kzoD5WkMrmav
mk56yBUKzjkNPp9nsQ3OensKDLqYI8TjDfpgyglaZ52Ua1GTv+VxxZHYJK6y1bU1
nkdKgdgNow8GPQnH0YTspBHAoz4vuoS8f6/wUq8z5/z/qM11GMiQZOcJWs3/LYWk
L8uao5sPfmhfIeZM7Zh9rD5oHXA6ZfmLVK5BwDQf4JkHzft/A0bffN4t/4F/gmO0
7c6+DiczRVXuc894X7Zf4UIirfQ5rD1+Y0unh3CN+USwnSNT2Vhh9/oDKLMDwQjH
Yv0z6kNIfGwpryIpBE1eJjcJgGxQLVOKUpTldz+C4e43lhw86ahaiQAn5QluPIs2
38RNtoAEZxCMFLOJDfR/j8knMaswZz54EkxcXVVXVuDStdcYwBNQ5A9oLYfNazUL
YcFVTkZkwCqGv/Wd8Uyg/5s5zsp8ro8eiGhTHP38SLVfuPzVVqVKxjSm7xSBf6xD
cseXhurIZzvnayGMWhUFvq+A4EdwkKRsib20y4zWIA7T7TynCqDvi0MDnRF8fcjN
D82skIlvZb3T136Z2IUtnCs3SsOOUsctUQQJfXH1V4YiFhQk0XIZiHsIJ76EHmwY
q7saoIUvHD0eZOpanKJYHpDmduYaYoaisy4vgBNmfanmabO3n3zC8GwDdrarIMIS
TQaL7CcDHQV/ZR9qnH1iq9gkVwRZcnYUM1SUAOYCve0nQqcW7oEf/jb4ByZNmlH6
BOlPvkC/uNsLjEGuGn8o3Mz4zYbyVc6zX+q89LedbihKKJTdVq31vtnWKudGOWqe
jL4lBHf1J09cynxpzIySd9hMco5W4iQ/kkETupgeE9d3wkYTrDQE2A3FU3W2oW0d
AeJ1WCAOHJJ17n8QI+ekQ6sfNgwWaXa3tk32ARJKsKMZ0JmmaPpQyg2lH0PAHSyb
Ktz7PHG//uCuA5O2DFSs+1csdyy+si/fFvnPUAz1LJBA3ED0FdLPw3Uac8rx6kE3
0+hinxth8rtVrJL2t8tQ2TB9u1cyVF/iQqgb4T0dm9DdQMesfEDm7Pq2LIm8aE4g
pXB4/BVi/iXgVvD8sgmE3LFCoknxGYX6jScLmfFONcaAWlvGoUbf8Ie4keCdfbb1
Xk9wQMOYvZ/mJ+OkVBmdX3Q+H+W7rEAH5rOUwyVfVXdJXSWNuu1gYWONNnof4Lqi
v0sl01CujsyovlBYvsyCgutVNKKFV48rdOmb/b214R6lkyxVeEXfYojZh9ESN08u
7y9Jbvp0EBGPvTxP+CmIo05dCgsldu0jMi4KyUiqFspI9RgfNBYPeCCxXSANHK8c
BetgGGB3xVO5AQdtkdD3K8ok6/VeVkxQQ+mQwlupOY2JW9gidedsxonAYqOhqUmI
iM8wKH9CUZiCoyqiUTYl6bCTHWoerTeXEFiYjDcuxEMYHZsquSV5eYORkuee4X2f
4RD8PJnDuQEGQjyPNAKhI/NS7uvX4aqunfVeqjN/kWbvp25FmX5qXck47ICC3zfw
/clTpiJ7rzTSw1AcY6/JA8JwUyNNoKQxcdT7oUdHP044MV6PoqfiV5To4/uJ+Ypl
UtoFiMosbuTXEOe8JKeiGxFfPOibt7Se6gngrGMhb4Y5qk8aD5tONSP3MaqjY+cR
voIgnaXsFOaWClbDY8lI9U9WIfd7h9K7Eji/WRfNKW2CUOw4yl34Sfum1fyo60Sb
bB44KQbO30uMLTqrmdFbuAKu2p8t8WRqJrVaY9r2hYaWZc61NkHLllEoKCmMZS4v
MqxFwZYgcEirvziXOs7tefeXUume2mThKUiOA2oayllEAw8dNljQm/5UnqUWK24z
rSKud72IbPsXHYj1cn37G3yjgFmudtlByFj4ikDD6iOiF4UkimVZEyoKRHlJ4zCG
dQHO10vafvnp5ddkvqc5IJKripiIojDLbC9tkYTcGMbupB4XxyrCo70X3h8jbM32
zi5xcCPEa2aJ+0VhS4hKmQiMD2PudvV6Rkft/SlafMCjmolzB6V/Pfx/RveGrOfl
YdMb2SJvu5pmKLHSk0W2gntcGgl0Sz7P0whhnSbrjhCGAdQ+6Krj/hUY5LEHPAKM
obIYDgUFsaJkQbAwW7NvnVQNFYRs5a2Scs4CaAd4t+f68wLDkQno8yBSoCbPlz9Z
y73F0Ly5W0mi6ZeI6T701mP59wdKYZnmZ417pdoGJRyvSYzkUpU1DJLEGX72f3J1
B3ieNfZLd4C870n77DncxwmT78VZ7J6YDeviGLzJQtdCDFr5P9tG6ad0ofeh19x4
BM8mBRfsXSFXBIlwkDEJodh2kpJ/kpEOw+gOV1ed8uUXUqVmt8S9ku/5MKk/uexs
DB+5s/VsOHd3hnzkUm/DetZOOLxj8QjfrMKMXamdxB7ODmXiLSClXTISTuFHaFxN
anJQ1dISUzUqVlivNtUqFm77EEClJeF/Oj543f/fjP+uhl/CgxZDU0L9WZ/sDQDL
caBD6dPdSReXimp2tpL0JMEuzVkGCmrLR+mFvkQaCTmwgV86tKj3ySfM0xxTdSSt
DbnJtOUVPg7rKprbzqng57ULzn+z4hs2I3zlqA0a0eXgJk3EJJ9HCzsoZ/AY+kFW
TO7DK+/3xvLN0k56/aiBH8+1JucyXaGTG1uwh5qCEf0v5KeHxGQTIjTAqFN/7313
qLVNsCKsoH+c4nGWzz89Gqj1wbADJ/pKQ3WodUilJYEcThF/OKmg9JwVScD2EXZg
gihTQt3BF9ZkX7oaWq1Ys7dyfQqMmnyhqsVCTN4GoG57N6qRXrMXvyXD3Ry9h5EK
PKXykO5vZE2j9kQ9mX6XH2g2y7RZbmjBKJtPMmsflCA0Jx2fJZ9y9kqSgmbzW+rU
WMHGKaZdZ/UhTWPbA2ZgfFh+MmuIjWzEsb9NBV0uP0H9XGLwsYpUVyLKI/FznZO1
QTFoh1OtpzOfCi7AhrZU56IdNYeguXBQfBxZlAQ45TYJInyrot3knRAf3jBAE9Mn
LzrnCiiwR43wBPG4MRpjae4AhGWLDVyo/s9Lh0VPr22cgAR6KOzcVb7UUG9dCpYg
UTi1XC64HAYUF7/7Tw66pmGpV+tp+o4JWdQDakF+07+hSST1lpnBdTevhEaDLnnB
FAgRuHkHkcW+OKPh/gpPjVp0GGv/up1mn6W/gzi2Rwv8WVDMd/U7WFBerX6oUBg7
HAlxdwBKz0z+HXTFkJsMb479wFzl8LPRF/2Pqa2oAzpTqne5vtP7XcKJssQ6+SkE
1jVwfDDHpmt0o4VY7dwBAzu7fddxYv4bBr4hfOg9c6hmBqVgEt8uzYWv95IFndS4
5+Py11UdDedonOfGky/ws0DpFPnHVc6pRBQNJcGqas9c5pPq3L0NwGphn6vU9Il1
1Ebxek64dJiX5P3CJlhX/Atm5TsM+gEGjRNXst/Ml68ZPs3x8TqF5nCDe2rDFwVG
TuqYsM9tP+YVQEFgzTiIIoYgpq+b/VcrjBFX78OdE/94BjEkN5DftvEPDEYCAM97
UVEwHW/rXoYBcYwAYNLoYZW2mTYsb9EcWsk03ZiTkRia7lmKElQnsqMxrqw6Shko
qbzhleEyU1IKnbQkXNqOg8OQwC3dMUDJ3MHn2VnDF3Q2fRSuoF+5BUISXzJi8mDb
Yc+x3w5OjFmUwLjihyhztA8PuwOrjBCeLZYgvXjqjcxgrnKtkrPjaD882lqmFRvS
1vx6WgphjOnEufFoz6tRFAkNopDIpr/xQA2pV/yemJILVsnqaSILV0eGQ7WmO6UE
CSzm18cs/sK0se0qfgiMS7rBuGIk5GpDp+hWG6JKGvBAyK2857xCkW41RQdSr1Jy
QZBAu/LE68l9U5DC0D883BEHdcSoMbNzwlwkQ7Y/lOg2l8imLmpSVpPWR+YjyxBU
20IHeVUBJ6qyCbvVVcFD/SIYaQ40jv56YNGMBXHuMoLyViYFrKfj+VydKIUHreio
UzoTFQeXojLFfhwxMuqwSIKb5/L7ja+Wlokaz+MH6XqWhkr67c7PCgytDMyaHUUC
HisjQQ/XDJsn/wZLPMKZsZAdvyTQf4rWzK2KDHMDGvfz+Rks/5sRGe9EbtOqs6AD
DZjHZBZn2iACbGNXzZx+TZpq4ESlHsfbdii0sgFqmRyAfiJqNuuOE4uQ9pLcXn9I
GzLlKyIexlHlpyF3dC1MT2/ZBDdQauC1Yffrn+s+qKl5cZ6VdIAi3ADL5QPsW09Q
MLkDbPAgFZnQKPVbOUc3/Yl1uvAfM1YRFPMZSQmIjI5nt9wXHRBOwYqGVsy4q6cD
5UzT5C1zK8Z5nyudHx92wvOnRPkfZQ+29+PNRL5FW7jo4ZE68UzNjmIJR7fYeIrl
I4k1Er1MeeJ7eVly2O79rcPZp315sL1vdfJSmCzU9bdQfA/mvZvNqvjw2iN3svCw
kyie+ZHB/xeIx/sBcSyDYv+AXogogeTHPjtuGkTAg6ntqRETRyWDMO3gEnXkHv6H
fW16/piIVBE/adatq9X/YDfh0jVCJt1G47c7gzEpz3cq0um0A8k26yAxNX8cLLTC
DsdPFUOC57xgyCPiOdnJkHuon7PjRJYK3nre7bA8sFO+ky7lYYv9iljYVb+gD8cM
hw/67EVAk+gr5ptfNTIoCvCBatUyffzBE5cVC0X1ya2fvzwYyjYU23C7JDWIX0/k
z0aQPg6k3yEoJkJzmMYC+edy2xsZ0WCdbyYtHWz60JVDAdiZCMSCvyeAjZPT6CLH
pkG46CUlwpiYfcDydMyWck69VW6kSB9Q5hP3vLEEHeJMcRizd+5ApIFXJhDrgxzc
XlRkeJewrWmlPhQ6yOr5jfIIIi/ifylThG8KDYe6xIMmksfHShO0N7N188mtt9Js
6YSP7Vw/phKznOfoPOY/MflNpAq+wCwgHA1lVnVLuQaE6mR3K0NkZavwpYP4/arv
b2jaGVJwgtLx4OYXCIpZmNTJairv7DKCdAKCxbqnPu8C/WelLYCOiviT6FjoyLn0
hs9LHe2t2+Xn1WP5fI73DyvEsikKoH9KgiZK0uBEJ0T47wIpdmRkPTxOPzthhQyq
KdsVRhicqQLv7vJkJB3JGFCXqCbJkIYLAQBlfcp4YYWsOOI8eYa/i9zbpvX/VIEu
zVQqRLO7K3dEB5PfHiBbp1vKms2+Y95XLuZcFHwhkXGG9+1fW6Cpdm3Bt8gGfoE5
aqESHeOkD6muEM1LrV0kfkqx7D5zcokbDWf8gJcLpowZ/aPXmFZXNnocz0WbhoOE
evCb58QsaffXRMcjPX0bU+1Lk5/ZSXqlb0+rx6pKHU4pE7/CPz+LF+L5Iv1htMNX
4DFM1yUlhKTZ220prX0gPpO0YZpU25zVAo5qc1VYwNAMkmYsMehaxHoYsXvyIZzu
emSypC/qbRpHJhdVlowistY3TQNZR8Jss35/oglqfIUZS9hFYNSN66X7ZWpX9CeM
2SS1O3GO/tVm1+XyzBjtDMqpC22Ii7XWoMbBoUNRM8nnFxDcDBGruhlTpeQk+qMi
2QcS4W2x8P0xkSfGeZx9IEcLth9Ny9CjXtXR54k3lqm4p+DsqzNgHjd86WUTODE7
xj33QEYqu2U78TVakMLO6AsgkKahoucAVC8+WEHphwWhyAQeUhgnwMloSdY7igvH
N/xx0WvRvOFrbPloplEL9/d664WI9nG+Dx0cTlmXp/m8be+Bs8FGq24QTFudFSVf
fCs6uypAATLGDYoSsExMPovU1EQlhq3a1oZBAXlyl+sALPST3n859/To+7bHA8oN
Jkl11UXelVet2zQZ74pVhIU+5CEmnDVcARqQS2OqefLq8gIal3I9obLxYTyiEWUo
pmOxkHuwAtK812YbFmQxQFkreHDDsnNlAqb3mzXdowO7DlapRZ6DYKMfGDPt45Yq
s6QdHwVfHsqua0BwU9qso/24ef0z7pDoKHuFk5MBYTvdDLkaRr41bOY2D7Bbk8KX
hkXO30jYz12lH5KsIQMlrEb1sZU2fcICENY2qYpnn8z2y9Y+61rm78LZMdWhhPDK
+EM1kGM5uF3NrZnTEveqGYX0dK5+Q+AiyxL39bcb99GzSWa4bqJop4wc9C7bd2tn
5GkkDUChavYLnzwihzj37lPNpDNCdIuseqIPRY36e9qoEx0f2hb0LyPI8kZiRmnY
JvgMl5xA+id4hPMpoRuhyL3KhSL/onnCoMZprRg5nsu0Oy0D8DneBp3sm4b1X82F
RucPnxG2idtrE7iCY5yyjK8PNPA2CgaqP20AVrIzVDaoI5JpcwCqNwV1nz+bbpDW
pE+NnGkvr9KxlDbdHCxVZooP2Kcan0ziGoULHtSTo786WUjOTXj9JIqYVaxfM2yt
zbc7rOuS7m/OpjH4WHGOmv6WLZnZwrR0jS7p7voEVWO1xktVTZQqhX07ZloceI4R
YhHxzSARDZZ0xnCm8BFOT1wAf0/CBxoVlmB7M+cEJNs=
`protect END_PROTECTED