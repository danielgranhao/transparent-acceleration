-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bTYVcY9CAle1hlsp5kcejgxftoXVHPig/gVOSMWojQwfoI1c5+nhuezBbdZkxQ03iZXCPZn6ZMuX
Nqt+ZG/TvSFOENvp9zXKk+qZqYG7TwuUTTor+0CdjXS1HFVJfdesg61Mk2UEGBUzPWPw/PSn2el9
hKoSZmo9tSI/lpKZzsMInH2funrZfYf3+v3cITmUIum8ncEQ8bYoLc14LlEwdb5hnAGfHXw+V1K6
QQd6FKHaIobEnPpxSfOhWbqhYx1MQsyeNhRWmGuGq7LtTMfmD/gdy5KKGNZLmCMsEOUSWpofRXWQ
1U1nmdEasLPJrzgPBuwe/x4gTyV6B16fpOOVzw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1680)
`protect data_block
RljqJn7euU4tP/gNNrfwD30zKQZpODTnwHP529BQGy+Fdt0frSnt/pdGuqSN5CSjMgVtS+Hg4A16
yqQR1IWQ8r/48YIcIkcrPy3rd74gQa2vQsZvv8QmfjWAxxhLLQJvWh8+R3LvoJ3kOZRAnroy3aJt
e8rzTpZIVtb6Z+URoGa93Jggn8V5jTq3PlXJaPZ1QIUcbz5ZIAOfaLsPePH/mCBM6xdU+YxU+70+
qrrWJMVirrZfM8vd3wFpeZZjUXaG71DYtsrUMeesM078NwlTsDbGxWw0+WpsXgNECSKhnZ/gbgzQ
ew/2gQ//RIdNBB3d/4lNZUtvyNluGf/XJ53tSUDinugfWVjTzM01qzsqMA7mhqduBSl/Lyhx/zCU
dyRIQZ9KsS+PLQZZMHcn/OafwY0UhpJ/Bh/3rs9SgKoReY2M+Z2yQdN+IpBwYYI7zamOGQUhmQh4
M8/Ee5TR/6fG8bH48c9kSnZXrBftVvnQaf+KQtj7Ria7+R3E+9zmm4KBkuN+51hViHdqWpJOSuME
imIdvZ/InVljOj2E3iAJFqC6Xa76XUTMQ/IHjC5BXPwkReyt9BNh16BfeaDu1zEXdvygDxp52t1a
9xrWLMIPcDH47fNoXkc8JHlF3eWH6YMR6fX8WdrVFM7X14/YRzOLVj1U0V+CQw5rIAhgA/cHEKcO
U8T0B0fCTrqveoVqQsNqaNOaBK7xWqy0HALkhvW8hSoCr/CIgKAJjbs9KTjU+winC+NTL/atbpnX
RpmU2CWKM05JRDcc89ReSly0/QJxMWZxAmZAoPZp5F7Mbg+gqCzvJT0nX9yIrL0iFU0O7JWjgrLO
9QdzaFGoT4OhXaSl8pg2+EPpWsIqanxA/ioWZ4PkBUDx2GQXEcw1CyFOO/4Wq7VMhEGfZIetboCK
6xawvwrpYGB7zKiAogxiuBGWjJ5KkqiPXge7QB9ysy/hKguFi6Qr3NUao5V0BvEOD7ms3egkUKgX
dNoUsrjHuWJCvrvZ96XVKu8ada1y5fBqjzGq4t3Dvt52IVUtDtSQwKdVgtu/EWpvl+sANGu6YxWb
jhG5pEOwXQIS53ZSO2LE6NmQV2M4y/BLiE7TOAhV/ejnBowU40GstXO7yL8pogEVHTdbIPOk0oM9
FE0ZmKgcm2j51fHnLkCcghurW0XdjWnH+lFqltTGd+dQ6F7Tgt3T2iYqtNI4HAYQ08mj188Kp4Eo
0QRzV0gmMiJyBt0PGc007ApFlnRZAaUUYqHyb7PAjOjMuZijVuT+3zEgfd1ZB3JzcQeM/BM8nY1O
Cr9qmAbW+XPJebn+tcmhwAKg9gg7hFr2mnftknWk97gbtik8HsS0tnAaF/Rd82wcH8a/gcuu4F1a
kkTTF+AxwrEp7UWzqGBd/LJ+H8CA+lZJDvHjKwixFCQN3qRTqgVABGGOk0IEnQ+Eu28n2ybX0HPD
akxEc9bLs+P1gE4GnkH+b8+TmzU2WtVTlXrJ/Fy86mA7W60zHjfb/WACsUFfH4x2/kiJTGev1lQF
0LBvkVDGAh/x43S1V8dDM0XhT9hQ2YXYIIlsuvUoQaC828+8JNUZc5d7mAeSWbk9RDkmHwQ27ZrT
ZUrnlrtP/O/EjjvNwAxlE445aWw3tD0uibUvCK3Q4N7mjfbW3oY7JS38wHYwiICfEB3nRU5dpqZU
0VbuTYE8HFZ/Gsrvj7FrTHSr/wiXCInlzRmSnjd5wd1l8Bizdqahy9dJzF+/ffziilg9piYJQNBT
iIMmj1CCoNbOi6Eoc/V4Br5VkJgsO3aIKVugzujeWHh2HVJey7MdhcuyVzqK8p+cxRUSuLziqXRA
jLpV6HezxiPlLM8Gj+z4bEGxG7jyj3HT8IJeFy9GgSowFUQmFDGu4PerpUCpNOLktxm0LHuhGC81
3/WiwECEbswCOtvTK0y4+yLlX9eeRaqhDN8B2XVBb2GCYCJzo2BAXTN14UAjQutBTC2Vi2Mm4xnD
yN0aiUIl8wchL4q6LMdGuooo8yjul4mpfqZNz/HDpCKuGGxoTy5c+aRqJrtXUePTu5qGviR5jw/F
r5Bm46PcqOFFcdvCcVJzXIxWrl5JY2i7cyqZtRkPqW94RJEv1lks3zuUO8t85N7eqaSeUf+Remf/
JSOB5mQSo1YfwIGpum68TMKynhkoEfHVK3D8nlz6ayR2jCnuiZjrawV7x6VKO//1okpOLE/fcMrx
M8BkSXRmHTpAzc5SjdddMd9b+R7uTED7QEnr
`protect end_protected
