-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qjCYUJd7XVov3DXp8BeBnbk34D66kYpSup1WNKLHMeOOL85j0RCycSqBV0MFX/93qXe0BL9YIZQY
7NrNd/kA4MrROo+kof05LM5k3PMCwqSmOvA3wWW+bOI5DNRZsdsgbIYGRjvnu2ug/BlHkzLGMkke
oHVvV7lfe2RiIegyw79nWBXmiyjllK7NzKHPpvktabY8mGA9Shd3DdNZnCzxPFrnX9bIS0ouS8iw
1l/0mO2cS+rp8sFBMoNOMPZblrYU69iLQmImxBw9JeYFd0DlBU7thMid/rAuq3Qj46NuEMqXHzIH
vL6bdy/3kmGPbFob+mfh5Xq2Q4DIdrYeE53v2w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 36320)
`protect data_block
pyLncTM/grFsPqL6XW1LhMkNqL8wAyVZHInAl5vRvlc5aW0o7CZ8WPUjniAY8Gm9h7UEr9Dtei9p
mC2Th3qFkSqzKdbbplStfxUrusL9FB9UWXiz6wXxTSuZSK6M5U/R4lIH7gv8Ewadq/RTu/0G3u41
YwFoXk5zDl0F4YFVPzL1CqtYO8TfkjLkU7DN0BbTXBajqVsrLssEtyRdxAV1RUs25dOnAsvXEzlk
p7/pzY8OnKw1lmj8/fhz0HXHE6/IN325gQd3yQUoE6kCrZsf+ialeEogYEKobDAcuF1ZvHphk2jT
fXVcnJ8PltCGRmjsI57/dgh4WkA1OOqu1GkXGyoGr29m5GdtP6ndZQ+jxBQfaWIFGHXPd4Nyj0VK
CmX7c5Atf868oQczzeZVEhAlfnV75BGOhf6RqeBiTvFreDi8pXbofbXRf+Ke78n2nCil+xIbMd1O
paMt96MYqVBpbyYZNoyY1KwoOfaZk/LUBHnBI1rWPFxKJm7NCPxR5z5kfPKsgSii9gfI0q5naADr
MddKggfDRW4cZgu2HtP/KLQHlKnUKvmUftADoQ3pBKhSiPZgR841EVHJhU3KOcVWIRrQzBsmensK
9CD6b0K4KgKg4iFhyWjyGOq+xRBEKlo86I4EyAw1mxsdYrYff/fYmX5LuLArIX8pQCd9DNzeOdxg
vIBZwA7xaeEtyBijVFR0uBJ0UqjMKPp/aZxg7RMDdpr1EZ0DTS8Oko/zOg/cTTBiM2X+mIYHRhk4
9uNJ7+j4hy880RkY8asaS+1sLK/OVW5u0mefOzVVFD2r1P72xE8r02CZk9CkVdMHoNaoRUSf25OD
mrNacgE2lG8YLI6bZlDKKq7uMNVM8KUJjcrKY7oKdRkg5MNHf6GXCQQiTUzZqGjHPzee/3MqPCAl
iZRQ7zWwJIDEa7yxELUmyeh40sSgTU5wh418FUBd8zHjHa3/dGbWhNfE3CcH0z6zW5y41VQAR39y
t/3XrDAU1wNm3mFMAIbOdNDAe5eNACzg+OneQu85XRKHgemvujpziZKYYaDTp1Q7CmphsozYoyVd
UuFri1+evGlZT4r6JNgez9p3p8A7+blOYxufOeJsFtwPPQAxJN5oLQT+xVIk4yrEQpxKoWGK/uDQ
ocrpZoAvkDJb717cxHVO+AqCdOguniDVGgLWVN2fmO2MV95IcmDJFTDVkqez7oP1dz2TK1FMugJX
N+xjO5RzlVbnJyF4TIvNbefsfxeT9/o7Vqoiey6+hzQiZz1WX9AuEL+EtupKszeT7N1JproxLgfJ
dXTdj6AqgXxpnPCn53Wd0W9zMNNGa9FTMAkXMk0/4F0oXGoazYzX1U+ARG73POYEl51qsdKd81dk
fFUNJna7TEiNWiX3Ya9toQCRDhdtrq0YVclJK4FT4KamX4Xg2QkSTTaXajCniKRC+mJWTLkv9gIg
loanlQkGpmtI+8pkwzgOd/6flFrX54buDtGjfo6L911qpBluD0weNO+TV4oP4fHHD4CDtZkBy8lf
q/HmiqL5oJ14Gp6v6euj9aHx+SCWHG0w3vRb6BZaMUeVPz+tVEGeOla9tK4GRzBo4hTs4MkRqSWV
OYCJvSW4e1DQJjRUbeorBpfwrT3+PXRLFhs4MnyTzYvSH7d+ma0EHoy+6no6Wis/641cDLY/HBlT
Dmk6OIwYAIqM2cxFRBedN6fdY9AcPbpBxLP6GSmtGosePvvn6d/hImYJxjzywjC/pzZ0uwf/sJcX
EedU1z1BafROzhjOsU4QZwiX/yx97DBqp72zioxyLN9CWic6UDBYgHRXII8lTrbTa6hd19VccXsc
NTkSVmBICsSF3yiFFAHazYXQEfqMUJCz8vobvFpB2jKkWKWb5czdA5vwqeW93jYXvzosZTrVvOQU
HfjjDN3Bi2+bMQWnKK33Z1J17xjMBQMwDy3tpdpSvqkgDsvnrEpBeC7L+xD6wRmC01xFPzmw+R7x
NGx2tUnG0LlwvowbcnKoPpf8UVY6Cg4imEuZQI5fsZjEaGzlQuIALWSFnGtuQykXUSgFR2CWL1MS
2It7o5ER6B8h1+RFsqeHomqZ7wD9YSPV4yws8caoHIm1FJQvHpRo8AIzf8bJcCdkrIwJ50vxXhIa
2tlXh+uMwSbhX7iCjEH9WqkdqoBtFk0AF8ZhfaAlUJmx53F7TEEDHnA+C0bWGc9i3IniNIXkbcLy
gM5syW1/oURteNMCy9Jbucxkx2a3uesUH3FRGkWOz86D7E6yjXaONED+ng123HeP7dehA/vf8z7X
ae85WEeImCqk/6BZvfglEa96cy4xKUquEN8L0UC9CCKwrqZ6ccNEWVsQj1F7vWHmjFYMMfQqOq7W
ntyESOqhUnODIJNCxzVtz0WP0lXUL4vVpogkCTSG0ltjrGrODNGKf59XW30b1HaF6DvUljwbt7iO
wMgbw/Vcg0PlqVbrUsqBOGxZvohpqgGBrUlMiuS3Y4NoJiSQuy9d3i5NW5Zx5Z23MbI07QPXJIN9
4BQLPZYqaxGpD1vBGFpcx+FBbIFkRHIF91hQ1M9sdmCJ+m7Xj3VlGGibzVoLD/XT/CCj66t5kA4j
L5+GXqFOn5meTm6MPwXZcx2yeTKRWvjMdkKxsEA1kaw9/0PQ4LbsxNecUShhZVXECb2mulY92fj5
ee9xH1CIX0E53qZjya/JMObUP3lOGLhePprMoQrxyR7/kNjHZjfZceYgHAp8Ac5wuKDJmdne0yRU
cWm3rP3oCIa2HprPRttHkXg+iz4o1l06Y6kXIGq1AoSreug7l9rdPmhGagdQa7ABmPEodpPBRc0P
qRmmNQ8U+eRUpt3XlVPEWAcjh8ILOuN+rF7S7agmnI6I0AuNxVrLEkFbQD/9EKJ42Lp4mCnqC3jx
wn6YFAp5Lpxb6Cs8Pao2Jph25brqcfKd/PhEepxBRuqQiZiXyF3oWbyVCKhQTNeSDToaeGlMdHs7
Y/eXQ9NRucZCnoVjkZN+C7v9iImnS1izzXt45+AQoMGIF/48anRqamXK5wjtjJAFX15q6QTCAnu8
O+Lyc7YCQSjTqnkOhQYXF6AjNF+baZuOyU5UpN5R+TjgzRCbe+HTBoxlekUlz84W7UQauY3DMy5x
4dGCsYSyc1tCqjOWiCQKDRwvKbr4xaG5Z7+k/gaul0LUBT9iC7/T/H+/ktqc8kW+cxnXBj1ASA0w
tdDsMWZbptnIlHj4STWztq9Iwk/JhIWCLDQxAmS96Gq2Xpr6DI/1xm7OM5B0M263OSjaimJVysAX
XzhQIJzQIgzhQqpZb9/oAbsI49G/8Q/cn0AwYM6pHdsmO58QxEVRv+LKZJyoGz2GTKtSE5bouQ3Z
chUbBJsSAARvFBypx6Nra+OWQoi/JxCVmjLRZkkWBJfWJwoJf+DOHj4wyP6yocyR3XFPnNco5KaL
4VDnATMPASiJTdSbbQkqN9J5rRa/ewxx/kV4rfYjwpTYUphAMQ9Pg8z9qaDatDqTh+Jj7pXw5Uf/
NLuDuOcnYwmjVdCtS+fSyl4sem/sKYuDlnwgAmm1LRjh1vGMwAqbgm3wVOsjXh5Z9BuTv1N837JE
QPWZ3Bo7lFogivV4PdEWwsdkOnDSkoDgaYSO8HHNiNaGcCZReRdhXfZibMYIRQ8Nt90AI35l0Cb6
cbapZwbFVISPlRaaoJXKcgves3rehIqmH3IDL2rflEgnG8ANsRrUmKnRCKpfj5NzCX7reY0AAoZI
0wNM5n4HNLj8/1+LSEFasG1ewg3XaJeGwqi6kP7zGxxBM26j4YXCpwwgmr9pSQuaqLXMVx4HuyzO
TLhh7slB0ae9ddHg16mY5KImzfN83xqpYAFajp3b5ZQB/5RLKvBAfxRPdrJdR6YfHO3ZxxeGixKe
qWr6pkq/UqGNIKOnksqNCPJ3FqG97czoc9gKg/WePPwFPLa6iJYx7LZ1aYnUIKms8/zW4OgfkZgC
37actUUY/9xC2BiWwcjKW1Gah2PCfVNvml+jqgKA0SoClzWSdHLSwoyNV9e/0Vh2EX6xWsVJa2JJ
/Elcj5eMcO/T9pYswOrdRN2K33WkUuavSjr4amn1qNRDTWuBCTTT5EjgXmYfnW+Ne5zMQjiuvcKq
pRerM21lmCC4N3P/LWGWOFsjvdd58BtpE72fb1uamvuPj+cpam4j6ZZ5lq+6I4zSTayI2MFkVmfK
p0CzQQ3ivr8l/5uuXr1SAgNPGT00xJ5VOtehgaQbkO77zBHOvCD1dVQ7Ru+s5fy+5hWWSPiBMW7K
ojZdyqNENugSUf/t/zGEZvBkTTP0A1ZFR+zqkbeg2fHb1Jl8mxXEBwg00/REWo+HQ4uMEyncUWdp
CSXcBmiyhEGc8wUKSNQ7qpqnl0zETH28k+jgbZNtEZeQKrG8maJ1x89QsK2vJSvYT1+FgxzG2PGh
KiUdB7xenOtOKeLiUJGCxIIzMO3R1mMRFppM0nb1i2rdZx0mf89Du6Qe+eIquUymJYEvmygw5Vio
woKXqP3v2SlAUGucIxvzCmQdh/mKShOU3FaITIynO/HytM/UyHuGSYgIYXHlsmkPeMzCyesWTYW6
aqisqyrQyEfoA/U0k2d8afI8wVVUdSkwB1EmNsZbVCBx7NkhaN3SbPqtdn7Lu91ZEd+csfSzJN/m
rNR+P4y1ui+P69JSm/EOXzc84dWaPErlvXVaRf5FK4nFy3krNMKP3mEh0lWuJyJir9uEQ+YqyyuY
1/zLWrC6CIj/k9tqyyU52viJ75DPc7Uj6JhPeBBPteA4YvEE7BqZXexOYuE1e8iB7uefvJMaEEM7
drson0ru5Fazb3cVqupwu835j0rGha8qDb7cTjKGuSDM4JZctkcrbWRwGKmaG3Q6BwB6+4Tlch7d
NOiVSYCt71R0u1shAzyeeyLvc/Sq/ikYDZTxBUoCtxt6edX7VyepmquUD4U/HioJRhlsS2fs0yhG
nrZqmH3BIm3w2aA6wfjm2liQcYOQq45NCI3N1yeK/bSiq5pO2wn0B3hkhQ2OqOgj9uB09DCJOkiJ
/fIzexakZbhVu6/8Eko0IBJky1Zp8R4cnVBhRz8aS+SaqI+wje1buVTs7DmWIvmc9BND0RVKQQAG
BsI8cNBaBkibedZufe0t3x5mBRtLWIAPK0Jx/RyLbzickM+ZyBZ0GGcOE/4ABTN7Xap3J3GaJni6
fnqW0cAsrD36lxtYcMIWHO6GKjl+A/cdi9Pi4xKtlBnDFyF8eocTBqrnNNv6nw0HXLt1p/0gDP5W
AhtJ8K0Zm01W4mwbA+vlvClbVhVhNI37CcCUrwpa2UywQw0ohyIhg39e+K96v3HZsMGpV/iBCNMw
5ioc7t1QpyYCH979ygb6NHGGk7Npxv8GFwj+s9jE26macm+uwHmDu+WjGgNE27y/yVOUrC1XG72a
+gVtcJcrRdKUm1yXRlwl6M81w/ctH5rK7xV4iak5aLGFWSMCSnGybiwq59ZblGNpiFQYhjq7kzM0
5p202/9eW9IdabMOETw5Vz9owjeajfFtVWsclR4vh/UsqQjQ1wg2hnsSDMbnWozxaYayVVjkvhiJ
Gvf1A/ceSN2mzbLnqZ0JszJAG3dh6au8zXJN/HKqeBQjzOucytO9flhNoWc8uGWZL/6w88k7E3QL
8YkdFwo4tqLDVIsbTzgY12+fGPqyN348ZLc+SGsq6/+/ggPDzdpERylMEiiUzYp+IQzHqhS31bdE
13bsMOkz9trMOKaiDu1zzU7soJX2U8KqKrby9BX/TaeM83pOcMePWJyEuC2neov+JIg47hHOfSyz
M3U2iNFs9fcB5ddFa40o7PMvlwt8NPK5qyc7a+U/LHxxAx1zkuQ0t3Pl0AX/gA3f9e2JLloZtI09
1vdvFzjNZkFNOgvuq+aGad2ONSlcRUspb29gmD4/drIG8pLztVq/fybyXEtnBXTw2F7+k2Gfkerj
Q7EUHTyCD6il4Jh0Z0oDQmIW09mJ+n9Zd0bGZDNLJ8IW81j3CvCMw5Fp+Uh+/Vox9s+pAg2nPehQ
bW0oBUFeODBHrBpJk2sPUscxIJiKVGtADOjqd9HWujim7566o7m8y8vqET/xDRh9DdAqT3E5uidi
djFrkw9Kn7+Dn3TA240kIftZItzPo89dng3nYKTvdxqTH5BtTD/z2kyZdO3zD/UYueTO2JvoUBCD
IFGZIoz/Qp9e+/Vwo3rCj50efRutyQdud3fUl1nXY1CcVF5fPpHn6KwkZ1FTxNRCS3c9OcYlnGh9
jvAnA4g8WeSDWpTh9K2UD3F4TshzdabGakruNL3S0ZW7Jog9gIhaMRh27vu/OTi1eJZIAb8OzKbT
FKpi6Dm40bpg7b6WcdmlISaWqka1B2fxlNDGAN9zXhcv5394/3uIFMoFHj7KBYgzopxrrlK+F5pN
/72KWh6mB2VzWChb6NGi0749NrjCDVGzv1WlPOuNcwY1sAg8LS1hD2uIj1AIF+UhKwJraIYVSfkX
tfaQAkCwCLGOnTPRV/YuKcIBEy7MwYbmw73yVt0oB1ev14RQB7sIMRmwhmBorl90q2ryFhfR6chB
mMTkVT5tvWq53RLOgriK1iPN7RTFSbv9SB8FgMKOw33KPdFz1mtO2HhHkAAalFh5Qj2lEvRKOWPv
lzv96FUfABoMgCufc5tog011kQuARR0sfBU1d53S/jkoF1mOWoN6VXlTNNJQdf/QQpw0KT3uv438
kH5rpT+bZbVMrzusm16WhBGYOEEYI6FQQ3OfeEJEOK4IDP513w8DoFbzU9t02QyA/N7oD4ccPAm2
AZ+B6A6Z3tIEGqGNJ4ZV836+210I++wkzRFeK9rUJm5RDFH9LiseVx6cw2mnfQ2oJL3SzxFWQVRa
eZvQJJM8n0RO9EDD/+P/5EkYXje67dSkiRd0afUnjuYeQkkvspwIF6dTeh2sAZvbw00ar9GtU2G2
PhOzUjaYN5ayqeTckoOhC/S/zFlDHOwWsQ1DZ+jFEhJUZB3tko3Q+641GJ88/VkeCmg6vWPHznOf
rSgY4Q8KuoWyWI15AjvrTkdUVD2lqPttV0BDelzTS30VnYw5FlEv4ws35/nwXRxUni9/FpvHlgEI
OsWOyGqOWusI1+bYglVoQAJENozBUnqPvgyXfA1RDqwiNOA4fsQeXkcPPqTeXHPIcU3MgjYCvF8L
FWbaYpuHJGZvefI8x7rSo4Gxi3j6EoliTL4/8FGTt3Di+FfFKPGPRsC8MKFwdO77do4yUvy+GLrh
sP9PvSWEk+bYMOjrsfTYiAwWED/7VTf3hOtSenXT8Deqi8vZd7LfvlymK5FX/r2HOAq2POqjqufr
lr9ZHZFtGEoztAJ6nxGFXvV8Ie59WT5EL81oqmPJzWT5r4kFt9kvo8Z4QbgmuRZgilj5kK57fNsh
kmycHiT7ShB8UrTM4Q7nHr3ynbZq5azEp3B0ZKJMz+ssa07phOc9mCxS3Zy8fQ16HjEWmPXPs9NN
yCyzFgOfzpsfMkDQRZVmWMWUdhq8CDiYIS1YnOXcSga6UDLmlXos/2hxS85rnCuTilKFGV7edwsM
zamW/S5JdOJC8QJrFMYBwkfQNEGoE0COEYBGa5fiUwynurF3WfTyfRnQUFlsgbMUFyodw2ljmCga
zo14fFZ0x5g1Min+ChlnKPmdfTVz4/yi4lMXoe7L1ATYEbb0LUafsX5SlHj55yPFA2mJq+HWt091
lLXD+0yp9nb+ljH/7rCTccZ/wXB1ZtOBRW7ZJ9qmHpf0YdkHASYEwqWMtiSGYrSe971mQCIdnvzQ
YzX/wvzzd8kYf/WcQWMbJMwLiQOoTuj/Njm/jJzxJcVMkQcKBEWxcQll30sSYtkYm2n2G6gkca7w
k9TecLbGHcwJJN5igz6sL2b5Pq6AmRV9SyZr1K7IkQFUafJX1agmv//KDZyJafmkcBfzxvZn3nO3
RYZNXmCkGX7WXvnUO4eJrvTfRbl/x5/sbgFXzPf8nhGXkoPOoAYcLDxlvt6lv0IanUyvlczfuKF+
6AQ80dGGxUZHKx708lYmSsQZTeA9N6xs5bBNXZMI3Wkqh1Qga6BFPJ5ybgud+ODw9KvGkdDlS5bR
A+RJ9ioa+8HaQifjmB+eBLnpnKkLmSepyZGog2vynN0WrpggnNoM/bJY+OI4Onza2/0UENl9Iq0B
kXNsfrd2cA5Ade6nJx2L3DqkAyZHHgBvJOqJPfxSE3BwW5UDNQJ4ihlKZaDI1790P15C+xbq1fzR
hamlHna5uiLTsfojZBMZ/fjH0W3k8P+HA7CJ+kX/b3HUKVWIuUVSsCXrKKR/gCWWTVX7uYrkoAVp
1I7yobv60eJGe7oameftJ9wKGGp7Ggqq7qoOtZaxHZjwQJI0d+DFLEIwHqp1e5UVcOh53M1Aw7tW
PpCRq4Hf6lTSBPKmp2cmdLsrA2V0nsh5SBPfR/nADXpyz6PokEKpQKrmgNuX3n3MBxOQRmR339mb
fNxqHcWj0GgwW84tqdSrQBCtd3wVwazXE1sVAEJ+WFSjosgNGVPd+AU2uvC3SzTf5otE3Z1YwOIp
p4jqonSheOe5oMvqTfNKD7zBm3qBS8BUhYEh6Q1SASJer7jnIdI3WKh7f4J9DhnUT5Qwz/117Jvw
/PBMyWW+GnLnmp4cEH/ve1f8mx4kX2wUQQBmuWX/gJACsItl+O1YG1Kc4vbORYRHSTpNBCBG+O6u
qCQBX8sD0zxK6XPW1ka0nOQG1n3HDosv4c5JCMNPQFhzKRfcFw1iWo2GPO3TZufXIwbCYgC+erot
MKKH8wnp7D4mUSAlq7+Em8QMLBTtMCccAMoCg+anyWep+gsUtI4hgV3QfJ4BgkxuZRPGvnN4DH+c
kDeHf/mbI9F+tfeh5lFxqizrfRZRKYfZ8twQh8hqMenfwbP0rmaqQY8gpwduRoOGvHkc4V5DA0sG
WcTfdqm2SZ+9vpZuraqsK9fbEn4pGvNBW3TpOwPg0RMpJb3M1dMlAud4NKBH0Loftl6ejzPsWfKp
mWVK7oS3sAHfkre2GXT80Sq6r3rYW1I5PXQlJe93xfkkuvSpCZHlQ1gkMf7dY+a9cTZjEXCj+I8Z
ti/5i4RsC7A56NKOrd2BvjyaFEULnX5fUvv4G97PD6gPadRCuJChoNUMpphTh9deLU/37JtOQPa1
GDWFcdzYIvGMMYU+G4VNWktclasFAv7Gy0YeJxb5aEu+TRO8TtdNfXncd84TeUK14smZsNGCCdIO
VT6BueLKmFJCcpqc6lg0lZ/KGmxYpb7oBcqfIxYw7SHWrRv5Z8cXKfRy8bQ1dhrDI5yZNlJra2JP
Iqt+B11Wr/xS/M7DZNTCm8No6ofinwfNZjmtjbq+vv+LWJpbOAU2uThg5oA7gXvT5sN45zdBk2+a
jZ+nTtRoUhlx29Y5kSOEcyJva7o67Cj2HWFPBbdLJOj/7nh7MJt3sk+L2DYzUc7F4e39I1ngsiAW
UizIM4ajO0yvuYUd1GemgV+KmVaBLg/8WrgLnZ2mCXMv0zEagQIvMTZWi+RYLxNWhP2DxAFr5OwR
VgBhGd1/JrNDwBYKkasxarC84TXVNN2xOYqA/7fvnO8oGjswBJ5jtsTw2RFRKMAP/foGxXOV8qsg
9/Y1+nY+bLnP6Z5aAYZrhoO2P+eMx2+2KWxwWaiGvstZ+CDPIsOQU62AbTEeQqzz5H/HKiIjEnMz
X5XI4Zy+jsqHtyg7nH52vvPYqIR/vNMZ/S/0ENeD7f257Coj6TXWSQyofVehORzHNFgQfNyhFMTz
YKoykZ9Td3SF/XJxNEtdpNG+ov0pDj+db0aZsdQ2nvyJyD2teIhY9G6EAMFtSvzo1nxnfthINpgN
CNlLHJef9UUIm17t/d0LKrRnluuDdb1cFUzEqzoVR8AYHlvrl/0t2JQc7hAcshnw7ggw6j3AUbHi
Shb64h2cg0LylvQ4OCjzpcrwQr7UaAJ0SwHEABChndsXQXCMeGcvbXPpUAwmKJZ5inz0HicD7cp2
IGUtAylB/yDWnOngLYoMG9w+hQ8HF+Pj213+QhMpUVi/VN0O7zLotC0QU0NhiscgV6YSTFCeW3hr
/v0sE5b16L0/jkEmv4L+CRpFML2ovE9NMqUbnfoNtiNO8y/47w1XUYmUMFzTUtHLz6Yj58CZKkmc
DJE1L9DmUzTMldC3dt0/dkcjngfFmZXFRx+FOGgY1VRjwzT55rUC9u2bKDdoFzsaSHNb4UfDwltT
gAr0zB864EOJJlXrWP8jNQM6EZTrwtXDzIO2MSBXF/Ih+EQyRnHPMygiyWh5jUybXk+gLuWE0bZu
3O1in9r9FSKqbyrHqY8UFb4s+r/p6R/Ly3T2Uf4sWbYjCechC1O5482qtXpLRMyc68ncCUM4hXrO
f8gtZPfz7UJep6x+rRHt9igZUxvmb0sVLEn5E+dOX8tC3fFuRr3Zp8M1K3n4SB/sGACud+BPO6hH
DrJ43P76b7pVZBp4j00EyZVBUITuT84nckjgY/AzxeL7pubWMpCKvfFvj4Is2nKrJ44cvD59YDfA
QKrUm5yhahoEyCBBvkEY/Z5np/vpPwqgzQYohcRGEyZm6ZOcpCWaKMqWwwY+H5NwiSwS8xOdhXIQ
/rpJtgr5DmR/b30JobDTrQYwBDscse99Za4Aty44iyUnzgX1yWl05sVxzZl3wtTX0ND6/1E4mXmV
DBKz13fS+TcNz5TmKh6ZFQ0tJEKuqMYQzAsc194rBkHOBlkAu2AWuk5u0pQKTVHqbGMn6/zdmIar
0tEK/xF4rJWcsE8VpdvTAMWbTD5eH2USM7PpnDLSN9eRuFH3+NiDroFyv/py3WT0kkmCudNm6bfb
8W5FZmoeTkpEmBOEP2T3CL75kjEQsU2v2muziqlFjnysCAaljaAqOZK9XCqTGeiaitBgl9KmPmoa
rI9ij87lv7eDsmR5/IBmF5z/W4DGwQBkC+2WkLCjjXZCaEHk5/Ga9DZByDLt1SX/WA/bTYAiJ4cj
QU60Tl0whOG1JN346J3k6NeF/+tqTVg4zuilacc3qoGaHdyCZ/gWnDtjLAM+RN6aqDXD+ApvHGrq
NKjvbMhdGSpfx2At8KVGv6jvsBOXlklxSYeCBE1NlDL6c0gHJLJbBJSaM7wnGHw2L5mQxR40kdPa
422tddZv0NemhZv6qSQAGsFQXEWQkLy3fezRq/PrImKeNe9Y8HOyhWoxG7DRaN3rLmxcE2bkR8Qo
Yj+3TQXdiZrGxtI28qQfuv2VyGk1YczInzy5rDKq3djlkCC2U1gGDTNBuF/hCqcdYNSbqVUxQy6k
tQVPl+O4DHfz97EkvmjNaHnEpVZX4Zs5PnUjlqDm8G4Ar4ow5Rc1awijePeeEDT/Weck8v+6bUNu
qU9UCEeNnZ7Ig8PpXN1f5T8W1KRmEq9H2LpsT0+T3ZpW8UQDe6x6RuHfgQts0ox18vyfyyiLmP7U
88U4sEtY81xrEM8yq3k5Rz4dgeIu7rU34kG0JEmOmNpNQBB+svPZ/ryDIVBzubZIHFicFO3MMMue
OWGMjqD9VhcdI5/SF/seZUx1Z4NwYJ8yRWmRQPd8sR8RyBQ3+XPPE0jkZ7rZb6bxQRqh0FoavqWY
PLCekwYysev8+ENRgPa1MX7FhJecw/22g9HqBd1znFd2wNnNSv1+YIUpyDRhmUXfkl3pTOGP5M37
JHH94EO+nyHnWeiLmqSwZjqGZ443+YhvqYWPITvpPeAm5mCApniFDhPIna4D/Vnj2VWYzd/lJmNt
Wqfw835A8lDQRSr4zCQupuK8l6iX73J7yLM3VqYsg3qeXw01fBSzOJE9KhjEvaJjmZiWU4QstXe5
17KnsbDfuPfETJ0+rz/frUo1J7BKDTwU+/t4R6s6TQmUnCJlB/Xmmm55hey/qzyIej6NB8doHe+w
QTmLMQBOavZ1aVCD9+qUwclBITd/GgcYidrVQYbqm0LfWX+k6fOoQgPYLg/xo000v+8xR3jGs71g
bpadSru6XkXO0N9+MDuSqqufXN8c+6Jy8u5uXmGlY/9rN+1RC2diTwFKXto5/Q4ZrsOz6kYsgZ0H
DE7MP3hOlytQY9EPUBkwpD0tvTtRylfQWnngmgLPfctd3UZj5S/Y3Xxc7K/+rV7VoV75MITo8Zow
Qvu/H3zfQivRc6Giyjq3wZuo5n0mv106QQCA0DGOqDS/SNtcn5WqzQucyAEtbQDjaBLkPfNYIG8O
hN/1Ev1JVOeV47G4M3x5DtiD+hNnJjTj6iPLHINCcG5g0GBzhZKjju8ImhPIomz7GLP/CISur8Sy
AKoDbiKng3mNR2Nkwv2fvQh69S/fjJierGAwa7RMYknggWWe0d3dDAyuytta9iHhNg37rLI2fO4W
/0zigotHIE99g0Ajq2QjHNT+tX0Csm1CTggShEhPu0qmdmDJ2AV9rSU31zSzWVvGq34zm+4reiHc
t9krD6hV3aFfRwQVsuL5k1+z3eWBXlMRYLDGoW8dcYgVjMGwTUKocsmyTamlieMAbeStw8DVu4Js
lGbjllq+LiGdJ1vKqMFYXpgI0D5litfcqDPDXuIBEBSqi/7J/a+13yDMipLOTWbkFu2QWLNzXJO8
wgvfWVklwcd/8hOM7TRoVY8H1nHY4YRikeD/AJtrpaIGwK+qyBcplC6063AZ+nM3X18DnT2nD/HI
EY5jjdRPOx6u1zQ+02JhK2X9vanpwJicfzwkfs42qEpph3gr9LmmgSwtIeB/G2aM1LeVUczf4Jot
Lf1f3JjGRCaBIbL+0vTK2hMPyWDePohf5qUz2kGlev142hI3gwx99Ocr5Z7WIbx2b1+fumClmxRz
bK/IG4ChngJRPShTd/382iIokOzaQ/luiOs9rP92En8bOxpKWokI4fPV56wvVEgsdDP+qKHpt/wI
ObJQWPg/CKOLzBw1g9pzch7WUSxbdtATF6JXspgkAVoDi9HCuYva+ulePDlOi7l1lGn2BU0tK5sR
eIdCLiqs74ty1iwHZf6X1p5mYv+qpLJDHL8xg/16HhuWRIfGoFse5KDjAFjvheqRzpvAzRHDkytM
6SuxgyIZq9MMx0yfvLNgJVfHAgdhRwTQqv9Uqi7W0xRouZmlafxqKa2g7k0qGU3xudWaogJ5mUoH
X5NQHrf8kSqV737efr2T5ZDvmV5nMKuEaL/PlghFuE056XW1qi7vtp4EYCT9PkpJrAYOkSm/7AWC
oTzKF8OPD9j+npYz4WcqzCb1KgFVF/q8OE7NwueadqHYycU66Afz1w2vppCvxGN4FNnm79vNW1tA
ea1+XA33qa4vchTQr8hVsuTXGCws4Pih92wjEzW607XJ1q3wQW87/i7XYzv15ZynLxfrcKbrvk+C
mowyt8R7CCrIP06l66Qu7S/NZG/3VjvcafgbNVdJUSkNBsXkBftRJRYgFp1eZZwHuoub+u+OtFrx
cDvbIvwwvcQF8SGppo4DsWYCDVYDe3FizTAEbQID+NDNK2L5ByirVz8j5CdpJ5DS5Kza0U8yLn81
SNWIPs7tyj59C+XmdG7YzQpdKcB/GdZtw2OoY7sYWmx0jrJl8U4h7v9RB/Kmc1PIqZCx2uKy0OKM
ZBSnmKx6kiXe7ylFSNLuzju8Pmv5i5wlNAeXNmvi/IzDECD4CjZ2o/hi0yx8MUfCxWmB70AA7isU
lybkoEh4S67ljR9CUKV/K0r+PboY8+86aqyLZn5UqiKUYZ1RSlhK4Du6NeEMF1hEUSwM5nRyxhmS
6Z4fWK9qQjRVAoCVNHC3OFpkas+vqJ/OooWwsQTN1PA+vqo0WKFEGaQGT+KPMU1GWN5oSBx2A8My
K3GkHM70xZp0WgKdWTTrxVyve0hBiFlBl9wPEy8qbxmeA7LSek6GWlQwHHmUhcMfmbtjgcKyc7KS
odz3vH3LuaI5cKvd/vTOBDCpbZMR2Y/2rBL/rNCapGEQ8s3Vr3Noqje8T+XJxKwzPLx2OAut7XRE
7/evY9ch/k1kExgQ1lTK/s4qXJyKtA/fplzDOsZ8gvEhTK3bNy5i4KNZMXzL6Xe17VQ2I/ef0DII
mv398Ikg1Dz5X4+ZPVr2yYXy585+q8FKMMVdM10CAQ8ItnT0W6ec7xqM23HPoCwx6/wvgmdf+Q/p
8C1b/iMO88I8hlOEeflGV7OqBXwXyn6Om1HfxK36ZwPHcj30VVRXCmLG94f6qKcLrMUvBGEXsrj0
Mp1q/h2UTeH99RCw6oaL9QOjH4xQVYprceR/E/EwBTmOJwajtHmdRLKRHFAyoZH43JToeC8zIesT
EnnmkvE5b/QKW3ga/lBslbzlOa+KUCTh/F6mfmWqWhZfaxGoPn4uxEnc9Hzrh29kV3+Ibxt11/LX
7x0MJYFJzBoLE1e5YaqoPMquyuX46/7lCBuT4JJu9gFuWa7MYX7R6iTUfmG+bEiZSFn8J+2de3aH
oHrD8XJ4T9HAmtaVXLzaQfiOXZAuUCrKuvugJUSneHLWXBgnZ2iMH4gd7kSOgfOdsGE5b8TvKwb9
Zk2mlHsIWsp2/cex/1fhMirIu/hqnP61XH8tPBlKoQ4FLUqDup+gU3KsVy1+7p6XfZJBd/Wfc3az
wSjStlsNAyAhf8t/GLshOq7mdjQuMZGVNQZpsdtiVBSHpjOc145o3iYEsytXDyI002h872R1rVDe
NS812SdoQUb1l1jpSFC4Pd7engR2YLnnTy8W4LdA0PVWMSDFioEmX6/2GtC52Sia03C0kSzZU1Vv
Y6EJt/Xf6QYtZQlZqrBSxnSSd1UfZbHbWX7Favfrk5fO+zChhDCOzgKZzSpwM9CC6crp22fdsOHZ
Gki9OgNYLCzFc6mIilx25Gy3a+B7AZfBqalffNp/WqP3bHgaBcQwaMH41kFXjXlYVVFTfJIeRs0v
k/bgw0VrBjEkdPVQ7K/xIGEtv1PhDrc7TDO1ifYndLgObpkx/bgAbfLQYLAtH6spU3M5VrxIE5QS
IY5wII2Y36v+RWPhaDFs8teYD13CPzqbvZ7p4Yips2vbUJI27NfTS6GrJAVxee4dHeIapoPC4k13
kdmifiWXsZb3FGyMy00TcvOMfElKAMuWOtFZ2cQAC6wpK743tPkm4EnOIY2/A14DakTbcjZCnW+N
9/zNdHDYd7waubU9rRA4MsunPfMPl/CxAhbrz+VMwt9b+2bpsNaCtqKtNhDOoHKoV6iluj6k0QW3
NRKTB4YCb5m7ZOuoC2h5gqWD7/6v8qa0O8yYXLt2QNe72SYawiRo2KFJyLPtVb70oUHmXQJ7JhXq
Cn3fDg9Q9w0Gj5Y7YxJjw/0So9OLcIrPzhL2DUJmV5QhF+kTCqZgQ+Z4KyiuwzK0uua7bNGKDxjo
Jjtk6vbAIlmCc40Sst/NWPL5DrgsybKExSEQN/il4tDMib18TSWxENQrcK0OXgO6dm7YbMF8QivH
LPsLUMq107dJAb353RHfr6DDnNKNRpVr+vanGYfNBdrb/lbv7+IisDIbX6y1zx2JPLOKUVYqyA4q
+MP9rsBhMtgp8pgeCXuTAG9auVMivqyb2inwWcGlKgiVKFhtXcsKsVhzBNrzpXg0DTZ10VwHJ9bi
+lfttVsEHR3XQTS7FpaI/wV1MWtjxDoaHw+ICd8dgEVWA8fMCmlewXhMOEZQh7l8OdGzKX+/goqv
YJIVqd0ttmBL+Xe4kGXADdGSJqdJw3bBIrcl3EeZjIw1XaS/w4uMNeK0EmMWmNbuB8x42/63ruxH
POlkahyzGbEElcVrSufv6ZBlDxEVyMI21QTD70FMhjc261OJoopmem3AJl1B0QM6PmwiusRtWN8c
q9t2gIqHowTFO9tXhgj90sYE5vn3ynxPZH5a8OX1Yalwas/46tRmmOTW2hqFvI3F7G3nYuu+URyH
mV1gLq4hr5YixFrikRlmWNA2Kd5EXJQD7CSe9hH+yu865J231SmXIIlqKFQyFtCCIyW9iYCNFpYB
uNYo+kYCYktV6PqAYH688axW/NIuYGK6KRyJtWe3GIjfh6sNoj6llGnSB4xqwRvQ/SajsvQjY+y+
ZD3C6qw4v9gyBgx+4MRi9qKtsUhr/QtkZ5PGKCe1xwXQJ7mEW1Cf9xdLXYJbU0xxhR7t/Tw00tew
6QlfJpbWvSSG/eMcV71//NrvuguYra85J6kmwB1J5hgmOgVp/ITxhzq4xmoWJqTWR0S/MFiothn5
jWjxd5c4C8dTC5EXyvfG7sn9fZCiEx7WdfrMAVNDggtV4qpKpIEf1tBxHMvfIYXA57+oXEjCYO7C
EceDMgJ9Eun0zQjq6Co9b2RIXeMBZ2LL6zCXOdPc3IP9g/N64j+9ec+8KabH3OaUw9E6kZAMVgiX
MY4lBCluSs50TbasGKIiOu6ihkG4na+xjcn5GgyWpQRP6pz2EJ668R/UrxPlclpC8fbi1Cr0Uwno
ZOZ1xzmmEWaeyPtAf9UMGi8YmAvP5r1+s8MQnqLDgBC9JcFqw95hVv4O5TkFbL870jCyk6K72Tgi
5d9r2Wfa9j14fz2Lg3shjuUxvwEMFBZLYYJJJfDs4bl2zD8b+b8nCN6mlvjvXuO7YnUU9bAtP8Ub
KkzeERX5r/U7btaPI/Sn4cujQ9S6g3W9bcbYyckxNcUPcE4NkH1mTOEcayaeYPFiYY2fCEMsxEof
6opxwVT7AVb9l9XrNlZE2JIj1W7zg4ckeJWct1n3Szh4KjgF1niv/PJxVKz65ZYsV7nkja1HH4HJ
39G8WPn5+fZ1XhujO1uJrtr7LHj5pwIqbcKqadudHhTG7Mx5v7x2cSLjg9x3ghfm5grKavRHHsqm
Oud9/eDqdeTI14HnMMhXwiDm4TAgWiN9ZDuTqi+PNK3PIeJoPNLcRGzDIZUQxP7f8tDCi6KOh+O5
JAKsTG6ehH24lIL4xQRMUodMdq4mD2Mvk5+zjq6fP/ikkfJ2r61HuJfnFu7fXso0QM3Y5AxNhhcb
2GzZZckHLDPBVEWwkOjFgbGGBzMrClv7jYIg2tqThUDRjwwHxJ2VxcBAp4oui9/su04Y9nPD67rX
/d5m+xxyDI7N3lbLoUHXNr7MI3PJv9yb5cBH9fWJKVHrIfT/vmsYSlVwkU8r2X4xYXapzd+kimT2
W8cUmNqx/BiVL6PYolplYpLRfFqH7JBxadVHX/Pxx3CtZQY1VUFdwB9DEXZs73WpjCFeyl2NQvAV
KyANwHGAHKGWlVlJEw8oJdCWRuWpMBkGvUpc/d+jZSlSvyp6NqYVag9O7xzdG+yktuHSt68AYd0c
0OiQqJHEO3LZbFbKZdGpRFlsVMg/3Lr2EmgJtlO1foK71X7TKpSPAI5QoH0IF84VgZlaI265Ktsg
/CcDUvzaRwdFj/8XJGhH5/Lma3eDEOAUHmwuNmnRgzVzP6LUoB2bcygKviITf3+6Bfw9dDrzz9Ja
iFEgyW2BcxkqT25f6B2lAmDcBT1vArVEwkWEu0HVyzFl3WNHIv1Q6QVLK/Oq++RoO11FAg4O/RV6
YP5Swze23YFSkHe4aHs1VO/aRHQP3fRfh/oH14HyH+EEe7WfgQfl/IR0w6TlVBFCXnZG/qY0CYqb
FzO8m6/y+DYtNuJtVh44sHt0XwJoIj6v1jJqgA4NtXcGbk8Vsj390nBZncfUZxLscEehAxiFSJbt
EdfN++lrZuKGnFgT10F4pl+naTlfiQ6VhOAMYqLcazyHe4Vs0nY6BIZ0attgjoEnhu+7mX9v15BE
OK8B9zhfFgpxxekMxtUWUSD0mBp+klp78r9SO+7+ZSv20CfOUnPsr2tc6p5/FEh1iluWD2aC+EXC
01GvW4hE6z2V/cPWsanA8nl68IJDug7iutP5lJr5kHDwfxdjbjYEUyG9cxG0qXN5x2h2cVZ3w1j4
AldFp0Tg8u89isMCY2YWzScO/LDnVbcvHpQFaitAgieB6fVWEcKOAT8iUodn8MhR/bg+4j/MYgfI
Fp30wNLA0dU27miul6LxSlCvGCuM8CZWrceNKvU3ZGM02zP4w6DSVFC67TlX64SUyZs29fycBgdQ
e2067ZZXMWWsp0ytMMZXVx8q1wdKKVSYqEDNibpYVUmQEh3pAKLht5pSxht+YltrojqjX3ZC6Zrf
vb3yezezD2OvNszafJBuHgfST124r5DGQ3cWIdNp/suWwxD2BHXtGcCuOJ5S70w949VnkVU3Gddm
kAjr1HGMvO57p5xLBiKY5x99KnKB2XLPQu8tQO9RnY8NCgIXbBi24B57Kjsy1AA/XD+O+jQhMFXz
Qbi/YSARVeBFxPkmrgD9T2L8nN/zWMY35bmkk8TdJTNZ+snTLUD9YJ7mAdtZopP1WeAGVFoCZrvy
iU4p/p5nV4U+B25QipI2fpCSRNLYTBwapYXTTTLvetu1srSI9z0nVPMJSuLeNCvEytu6em6SEMiL
ltb0Pek3STYXZjmuaziV9j/YRR4ZYbOFj1cU3T6LP4ve/2Hg2eBLJmpbtElJsLphGqktHGnh9wi8
MyGZDX5lzrflBh5M7WJ6YVsdOa/FhcLPZiw3fUYhLPc+/Ug45oVk+9Qijaz9xvSR7t1685TMgY1S
85yC5mIfiEpC2lJ5u7FfF6HSHevfOT61Flh5DE5iFTRhX6AwxUFax1dmYWgII5HYCSM7O8mJL5k/
BEG0s6YvexzhodLs98PGFqBGrRO88aybOdzX0TN0gP/6GC+ZR6B7nt8TSE0GfPLM5/OAYxsCaQy+
R1Ur1eHjgqsyVck3Ip14tCkqFZBtwn+eLdoKVdsmEaeGiSoANxvFaGTYhF9O6Uz8wgX9vi5WBkIr
6hM4PlT7ngBJBPL9Mh1M1SzSrjWqegsskMTxvSWkFWB58xgNVPZ8qJzc9NDC55JiNLNuz/SNGes3
saF5uzTuso3sf4IMwjXJ4bIOaMy93ZYJky1QBTdoL3VJ5JIlTpVSNzqwoqw3SWfdDbjMqQxEOn6r
GhQADBM3skUXUuaz5TGhs5QFOyLeEJSu+Yxx4ShDELn/nGAL+4Zdj8BYqklWZzQ/sT0zDCUGnxQp
UCNU1UmfZz8Z4GWVvP4BVIP5Y2rYQADPbWv3H2eQgg4sqYwHq4fDXSPeC4kQ3rigxeFT1jWzCFSb
/itCzG4iVE3fILDYenClbXAs5CeX3sY617CHpi5Bx65MEUyBSCdoaMSUmnY6BTCJosq/velhGkSB
+R1aZpyJFDw1fXLNWQ9+8mMk8M2ohI81ZpUATbGizpJEbk/SsMvLRANmUWyN3Q6iifIRPjmuHzZJ
ze8aZHZOBlGwlVxy9v+Oz/M9dYTnoH1u9DsFsfDdI47oPS/YKQSxVCR3l1mJhR1CTrYEskzYZSfM
+KZcjegBUgiHGwS+iUZSEGfchc7q26grEEHnkR9tqWhI8dMLCWAp7aSdZlpCOlcrrdoaJqLQxY8M
wUIO4LKTXnRJJF5eVwdvkWugEz8h5UD+ySBwdV7V9Og4pyKKmYibgl/4tfgAxW2NrSYROetWZUEQ
euEwSeaDfGeBHhYW5bYME6YzT8q0JhRBY5ON2+qIKwLHOgU2EQpwnIJckdvqur4e3pi5NpR+V5y5
1s9LYEyxZmvnf3CupqQOLamy8lKpD5AOBpeMElPtDtS6xm95Yt1vCdPNndlMhbrc4lyB/gfnwxf6
RCkPZ27tCB3y4G/9OcpHxPs3g/zeuxfz0ATeuTt6O5nTkZZPRAdodv8Q/Y9OwtqGJJOPMwFKupCz
S71FzfCEW6gQFOBTwWeMPw+Y/vZ/z79fbmxdas250ZqgMx1bzU6xCaKBXihIcGRYTS8Af38/t9Vs
5EXdv2/noA2qLeF+N8i1jilHFj1ACBMGRViUi2Pc6q6H2fCCKkyYmdyMyRW8TVlRwfk+0fS+UIZK
1SLz5BKtZwOBZ2TZ28/IVpEcTbH9kO3zBH9jj+ledgmNQ1+NyexAog6uBqjaelLB2P3GKhava8kL
T7LJiIuDZURhCDveVC8/756OBMKRx0YwSG+pJ7zwO15fmkEIibC89L2xM6euW2suPmJDgNgf7SSL
eAkGX/YPXPNBxn9C5KQLcUdWHpqPFF2d+kFchCmL7X9ZupD609cZnC3Yek/Zv2u49ZUCKVNpv8NU
a0V/yOPal7TdvIcCS8dRK3EbnV5F0BfmSItGfS3u3I6RYhxfZjJlOvdgO9fpk0/q64dNTiqYstUK
Ctyz3TH0eyEfPRWEuiyOTD1EebqF7OAQjq8ItTsHZWn46Coqa+I28iDN0PQvqxLgibMbHaDTEXbI
CZQSeSauzycCogtq1rRoDhfqYMqbObBvtHb1Kf4ieC7R3/DtO10q+tzdB6roDLoHHY450es11SP3
DZxMIryZb364UTrbgG55615GcWbb9YBi7z8U5mxjOTzOkkVzgZsB9BMpuBkfQBmzcFfgw7qnn/eq
l+UoxpIknoCHAGlzKASdqCuzd0kN+Hp+6NxafT0jGgx/Kpq9pv6AONgKNCV8YOHn192C84TBbIpi
HGkUbTxhO+F9XzRP+IkGdUez2IBaTrGu6XzGTSNbj32x5/V5Gm/msjd68h2qwqk9YEWyh91Ci0jh
NNRpEpIyw6cozPIKuZAr5USxOlxXFHlC9hQ6a4p4X1l0TfZ3WUSlrPWg6DuT76ZhGn2orSVjg7XP
rcS/CPnSaiV3DOVZ67hIkkbYA9A2kGdRxOS+DjdjH8RyLK2P4IAi1F1/M9mqGzOLFo08B80uG4mC
pvdkrLeRdo4zwvuWw+VwpNCpy0xfWVrmtWzyVpBdMvbslg0RiOTPJyVc+7ilaiKEBv7KMnfNzigl
LrbCZp/Nu22EqWnyP7ka3viJtCO8ObiK83SJsTN6+DKz3ii0s56Wxjbn/Kd9HoIWL5o32zvCwKqU
qzI+iYxgdWVtULmh1SWecrWRinAPvkEulr1U+n/vh0w4lKTyuyKQehOZ0Vp8+HlmULXW95PPhujO
z0XYmnRVSbQFfLiJWyVy1S2TYlj5nFBxICx7xAe0F0C3ZNDg34OnC5WjS1ivr9LQQz2KMDeiR4+4
0KADQsIGAKAwq6xL+RCAUabY4FZO1J9sxSoqH7zMWgbkq0jpMZXwF107oMpqFE0hGgv47ZPIyhYf
f1IG2OV3c0hhaWZyzM4rBdTyd5L8h5n9RPq3R7l8JSFRX53z2vsKPE3vC5HKoJu15OogCFMSSy/8
xE8f+DHfHcKPrARbje/+ZodXMrhUtF1EiMcYtm0eF4VSdfFPCMEb5D6ULGqDssGBCNSAlC7s9bs6
MfmNKRFeyP8DJ3Zdbh+ifP3QseqbEbPoXSDAal/KhmX3IYSmaZL5mZnW78xOW18yCg/HbADIdnwt
poF3UBK6WyrC6ZV541XFX8QzPZdA//YYVfnXts/57bQ+QySWly0/bm92h4lFwkTdxVCTgE0HWqOj
XiD7yZvsFETn+l9dL4vxkEMhSCwFtzmrFkMzpzF5N/hyNOLqHIp3pPDEe945oLDMTtTtMnS1+msc
TTDAWj9GiCekw7BeKk+TAmSdAdlChdNwMA+cqw/TQ0mi8gVaiSzOfCM2zKF05ooK14o+cKCeD3tT
p3VtQPziVZoeWOtbrVZS2UHc2zxH0PiRWUV9Vat3TA37owsB9YBq2X40w/n1+ZnT3eWdePWM9qWw
wRYQa5e9OkqaBWPYEtKZym8tCyTmvcOTgcyTkwYxHbgivdo+W6rdQAHloOBg4pUzsIPPwum797x9
Jq/ZD6691n4oq5LEVm9pEMdu8g0XaaBWUwRVI07zY5fCmazMBkvGHu2MKvlNgv2ZWTt+EHE+CpHl
nmNmq93D+j6L+pcDAeVPEUeYnqlpXE2wJiMHhy9DFMLTV26z3EqgjNDEIaUqq+ZU+Zrev6zhBGIh
ZN+Wx+R6B/oheDwp2qmYA1HEj2yyin5IfdRlek2sE9ubmTiGIPtal+ssM686oFPh7zILLZ09Goey
VsSI8/v0PQ7aWw3m3jon1hIiqFoSxRuXYjZdIm1Yq4G8FvASYPdb+ZCN9EdT4wm9OrsLgT2Ks+BB
m9EL3/w0gHzA8KxNHsX3bvdK+fqkDY+n5HuwTeqsOusfcZ7TMDNKWz+GvQUJvLyFnk8oLOF2Dc4P
338G7IHlR4CYqNtpNxWJXS0GkFO519/Mg2yxtqk97nlttolGmOEXle7E9aYhZMoOMO+c0n1A30Rv
9mlx5TNGIyh29rfLC/BOTRS69tk+zUBV4OI0wKhaZOD3A+yx6+16hk9gSomz/o/bljYaP4l7gLA2
MceqKojYS6rjjIhrc1sS63slthqA3EBowNRpzdWk7wIM4qtlG9vxkD/wOWg+8LkIz/SRDA27nq+X
opd23hGuaSamB3AQlDxafr0CIbCkGxBKzGV3nLzxpQ/AtBo9u8Wf7yMg50barCaOrp0dndx5rs5x
Xpn3gSRt6YnvdTULfPviuTNUrEVCmszmr0rej9eD9XCug3jnH0ObAdj3BTKx5uexAk68ikvK9m3x
Gji6zVhpBGWTMy/E+cwfdVereN73e7MUKbmdijxgcE2Kw8KX6HNVfb96orVvyBQHMwqSiaI4Rf38
2CNin/9HV7PK1DTHD2yjz7Z9cLZCdECEm7bCMSBGR91ysPc5pU3f0dA9RiBQPFWNLAIdsPI9oQ74
cMPRCyLqUTvehQ3mfwXbsdYtwPRrRU0VSbUQooFQJpkpcrHOt0JbUpleCPHNfhGDOwZkFpxyv+a1
EEly15gn/1qMoXaTh2f5T6kRIp5W9ohP/818toLPoFA53ywFJYSzBoA4KWerzaUUovHdodKoKi4H
6XYuvHwogoDb7ZZqYtwoE460mNaBqNXFhnOSV0aiEhhk2RVUXG3JWMsnsnwtlvqJlxuV9wZ8IPph
SeTjwMFAxfGc7B9+FH3ZRLLuNcZkDXALmbSGusp5BmYgAfMz0Fk4QoZcqd685r3zqc7nDaVDIvv8
BDDD0N3TpiBz1BQLpDInVC/32lLRBVemCFAoMGPdeHb82RWCWYl1ot49gEBKS24jPD4xCA6QMsgE
R/+TRW+vd0ItB3aE51fZgl9qxL3ww6zYcQ4Y+H/vxLGELSqKk/qoGjyR8V/FeV9zkf0NOgG6Zd2R
tAJ8wz1xha5I4v4JeRzOKoHRdxBcNgMK0YIaLX5ure8gWm1GPybrbc2lry+EJ0ptjhpOPGCH5GOn
+bFCdATTbUPLwG1zpmfIhWhsT+fA7HzXgu0ykPa8MV6WsQb7Y/1TFhkQ2fqiKlG77qDxmI6CvgYD
pzcpm2021JtzRpdOJyvoiImHYw9jorJJsf/xuJm232YewyarsP6hSSzM+9yYpLPsSut4bSwSqZDl
UzmjrFg+KrMb/MRFfIDrdCo+lAelqyspXlUm6RYHE8vU8WZYDlP4lY7Q3NkMM3yWzbN8mw3HKT8V
lD7wI1+i917EfvTwVhKHYxs8tDiwggLP5dY1WDL08ZvewF+kWQpcD7OoZFxitSHcchLA+C8mzGRc
9ssKSVXkib6EfqhSXO6GHAPEts3s7IXUmhJoI0EPtvOIVdBKP2ME0+itWFZetxHJRWfTEpd+qN3y
+QP0TJ+VaS8GRnknN1kDZDA5X5VIIPlTMejukXLiS374tzER+C8h5SJr5U8hXKykOP5jyE+IxOZp
Mxe1KMI/mBIJUkhNyoWtSmndVdLMRj4mGtru8CWZO+HAhKXzEGsrw9GUGev1d/UW3gxW1lJlxVDs
EssLqoiotA9HOyjs3cNsOEbh5W/qw1QoBfWMRHUtbczdZQ1NqFXnxFZbUDMDK7n4cCEuPm+i8c7M
mR0yEcMPF7EAry7s88utt21FXBuRm30SLuMPfYrCu03T9SUkFTQ0LnLjLr4aH/1QlCYZFltJhsoL
q9CjiB8Ox+cTxlgwuFdtEn6OMhbPFVnxuFF8OXMq1i3OrnYQV3GxYw3htRX2hFHRcAqBnCLxk0uw
GB+OgCA4R1PAjFVhRvpmNXbsWPqHycQsJapiV1QyvgGaQHovNKFdv4QEBLJvwER4uOZEN1g07z8u
ES+P4sCFjdQbTezV1/6mG/jL+CG45Mv0JSmnUk9pRVT4jBek8ue97rDF2h2QN4igoacKdSWPNaQd
/uBqtfcsx/LMOKz9n0enWG3V/SX37wo3XWaDBxSq4LEb6KHyyYnYefEURLicqsItz8o4Pae1YZk7
hpI7Brk/VtocObyxxVlGlVNdtWzYJDqpVni6srg25EOC07JyOpPENE/zTXSz12t69ZfgpGs/w6ax
l48ebvyBINHRTDXp4qOt3x45lQ35wftKTYJYJtUa45hZQiih2jTBK4XoOG63qSFHSwhbivh+n80f
u6nMh6T1+fCMYpk/vzwPPo23HlX5rK/vwvVr27OsNJvCNVxs2uDspoofThWkI7d//sAqvdCOhxeQ
G4sepe8MVDfOnRH31tPAp4n0hFkzDAnz/Z35zc11nH6oy+XiCpOwuYuSKlVuabgfr+I/NAwphAbZ
tXqjNgZsR7rUV9mhojKDscvlpMDYtHxWUhLMFHWIsuampv87LxmVu3aGObJJSMiVkTFwUHwaBF0Z
DHvkMiIvj69cBOQjj+mp66ulWg/AxIBcN664chVMR7TV3VhnHjUsv95RA22ZO9onPzFsaPtcV+p+
/wcqDLZ0+fS241hdK12KGGVH2yTXz/VJZWWigEApSaTTZlBocYzqq3yAkpCZlqP7/6ZmsUZF6bNM
FkjD88z6SywlyNsfFS4AGQe3evL+lj9lBNaS7dBoIYNg663FuGDlHXDkdH9uVd83FjeABxRbUZpD
BxVZ/MJDTkkz/wfSwa6YtKUSftdEf+OvR0ABKYQdXdZk7GX5NX5eWshdE9IjOEYxnvX5vElUvWHd
r1MZWn/YDTRKFNNtPnIf0akwlOrcqYGdVkYQ1VWJztj7qnzS/NQzW6U545i5phKNXsCyPrtYWcDV
ZiZuK4ZDLzgiOYY7Bjz3oo/Bo5V0GnxhZT5nTA/TZEV/EAS7+8jrEc7XJGuPHCkIZXW/JB510DIE
3nq2hmqBlW4nYPMc9IMXpRb9kydOBLpHnAXWBSImlMBW09SD/Ngmdtx4JhfR1aXfBzPjCQ0pUAsw
JvHfIZYJdEpmkreJnGL/c4E3czrNhXr8mTc95WbCsBM4AR/nQ5NO3STztWnKYsVRdp58BvatEtgE
oVKAQ+XBWjJAh4jNaB/LKH9stg3hqisgdA4sQGvvA0PfPrkg2gUpsYQQozP9VYjITJROrV8bzJtW
tFS8JflzsSgfaVcVPYJ6ricYgVF17aEATktm/1LYiIVEeDZ+k0+yRtdnOmzv6iVHjsxmk36mQvpL
WXWs49D1/GMEG6BYdKhZpJtUV20PrHu/TjoIrdFBfZQR+v5555lLm+Ahu9eBo5gy/vODQ6mZBIZn
5zjUZR/HhgXen9h0JWMXBPlEYQRyv2H6oujt5F65Soc9DRpcWunIQBXSmlty7d+fwgRndYlVaCvs
TZFgSqjk4NfnmWSgC9YPfkNqD5nJQR66zpEYVXnCn9ViOZNJNQTmWS3qu3Yd7m+MYtQ6fMTTjirA
NH4KfinTVayer0+QqXiHhy+EBMMj6ThJrJzXhE5M7zCTDD/9EEMMa7KmiOx7xIs6RnWqG7HEH01n
i/WpUKB7lTxFVwE5WCQlszLKvjJxX2Xajmi1wJoknlzzS6Nookqc5ju4idQs1cR/xCVQgKeDONUO
lHlquEDQUpqF/9IzLVhqgF+njcNKT7birRoRWaMovgTU0jeR30zFDvqaCbE8d0VuyhYMiAA+ShQy
Dz/+M6AUjQ5nd/SyctbRPmE8WucDRlN5G8NAHIJKN4dNSih5tgtq3KAQCS/FJQx+3aaRmykKjdvK
yTbnrJE3BSD4JnKS/NDOJcejoG169fh8ep4WPI+Wvqi6nZn2g8OSvJ1cgJf4pDPBDaZNeTumiBsb
CryKd8yNgyXTn5jQB2p+2cqiPkTIW9Gm5+sEIlrzzdP2l/0tTdbeiAJ+Prkh+kLD1h4f9yl3CMZo
Bgw1xEleGhVlJ41rM6JWL/atq1R7fqyXy0j2xB9741x34wwHrmQs1IuRZrcYrevhIv7xVjXMsNmz
vI3CtsAuFTigGelgHTTMPUtmuCt2unHcxjqdtTBjw97EJq1bH7YsRPE0el2AS1qeR+lNvXIRYMmR
3oDb+SRMTG/hGex3xkZvlzNVo+xAGNynQ9huCHMsKBHd0XVbCq3ZvLbmCrlih1y2FUiVwWEgQKwj
JH6C6LW6I9Q4VLjs7k+5OAqEjZABCSzbUcMH3cn0eApLUJ0t47JycdSHBGHPzg+mkQOieeT8x4mn
wuhML+rrxoQqii8XzmfoNvHlsiqqOOS/IKBNYHJrLWhk3l8u2tWzMBNlyyaAwclanhOYyaJsAXQ9
i1YfyxHpvsYxLIVpauB7+81zmUaz0/boC7A6Zzj0LU2F+zqySbOkm0slsGyFrK1DKk2ZAXVhUqHu
l4hSqBtCyYb9IHRWVpPg2jHOFhsmCemknzT1U8lsN9scP9h4GjTdN+bNX4p9sKRu0tPb5De/8fsM
q4SHWb5Ew+qCprqO109WG3sGscmlnENSyG4yig/H+wyow0+FNPrMMMXWF3KJWPj/bFeJejGJ7Teu
TPupJ6aU+qgsErrNvSkjo62eFF0tyUdsk+rTpbVl0vqTOJh4zcXs7x8QQWgHQ6MLyFUt2ayCY61P
ynyFqlJqU4pAgkNP9qFYpY0ZUOF2fOEcBz0xvlYKM+RIudEn4F+N/Hawop6Lnax0ZpA53RYSTctq
28Iuv4qxtrxuCvmVQ/qAxetKiwlHjFHkBBVdzCIb/cmmEh1GDE84tNWSFLBBSqT7vXFnp9RrRAwE
NQ9zBP6c42dkXKfOLbcEHogbOBz7fsCK1J9umNCwuDS0RtOWgPvLJXvByPCTso3J3sdolOSt0VyR
8avrdPbbsnYonvSHBOoJxuf0dxXSwABAfkxuIqAp/Mm+xZOTCunH0C9xnTsvPVasfzJpd7u590Jc
YJEAKceFHOj4S+d8Zm3LNvAWW0hUfy91sLBB4Va/iaoSTZg6jm4Uyv4OD217+vZdM0Wcnnz1VejG
u3q2bZGN1nmiB0+8OCPQU2BOIZAW/7SAMNWOm59s1xVm2pt24koVACQ8Yya5B/Q+U1cxSodufZ8v
gWU52haeFTUN8eEUZj8NB9xxxhiZRC2MhkVSC2xaktjoq5BM/dd+2xgpQhi9FQ8L7MLm6fsi7C+c
+EuO/i7+tJ9up4wIsFq547fF9Mi/ESvYbg0jHwsSn0mUAOxJ4uc6OhA5+TKcFU/YHcsKORvufM1K
wLG6ECOC2ZqOw/AcxSFsVLfDPApJXSlh8yXiJn9qLDTJQAtVWcnonjE7cq5H2X9EubT/pw95KfG6
+F8sWLiv9kLdAImVsyQSA32GAxYJEPF5hBv/3ZOAWdCFD+urPnBydMBM5rwSCp64o30NGeK5ZJ8B
gXVrf8zT55oBKEQYtatlLrQbg4FQbRdAQ+UWYTc+E24fzF40e3eCFS6YqYoG7+zaoi7Xv4+W2HzB
H4BvB0f2Q9al0W8SPf6r/k8F2VE/LT0NXkVBRZEjUEWiU+23mh2foG3oit3sP8j6g6KvyG8Gp6b2
2EKZICQyFgldw3fmUKQlYfcV/jSZMgi3rcsrAxuwWFPPE1uoUS1XPfa4pWZKd+L147sayvpy58wH
5YTZNFyBsL4f55yy/q5AWJBiaN67r0EYwcVHZeqj1o1FVSoGcyOEkJEOVmFRGLkchAGyisXAlwmd
CV4LTvnMLyGNZpqf+TaoTq5Joc7Xz+QnV+4Q92bs9zqE1ZOhIwZNMGq4+lyahG4umijz10vX8GpR
gUVQMy5ylmQXp6bjOWPTYC98IfYPtEjnLTF6lVmfkdvfP5PPkG51B4M/PfIZrXqug0cSQfpVOWm0
1RZ1oFd/VtnvBsi0fCRZFYQRXCC5uDWNbp+8fkoqy1oIoONYc62Be568p33QG7WyFLT7MSAu1oxy
GylmoaI+/qkuuRdxLKey/xoBHlCzcErPqGXAOuV/puoHwc8narOunDhRtXXWEYLxcHxXAGwV8VlA
P/gcgZVE8ukKLnH0UmuBKYnsXmS750zGP6/PMiiCMiVT5AveLJqf/f1W8RfRrqG6/GF/6drbWlkV
57+oUlP4oM9FK2XQzJNEm/srZHqeR2UtEGANMjAvPG8+/LLA0yTZ/acWeRIG8B7keJOr39u17q1x
pWut30MJIoY//93hn9s9ATxEQ59R6qTsCCu7ChYvJ4/lt7mJv/ir0TY88gd2ZxzEjt1l60BFJ/lD
VWVPxLbbN+AN0/gJOIFdwuqYljPQ6VrsMNN16WTy7uq1XsSqocb5gr/IijL9bYJmG8ArkqPjYG0Y
8q+1odU31e/gFOC3O2Yaf+n34/MKxa8dZtsLf9l5iEXPb6V6hhPIhKWONOMlbNq6Ko5/YG0OuS9+
XihKC1J/EFCzAj6kLF8Ugs9VpxpMG8sNS6PPAUZX8vcFuI+shyZd8mE8601iEw1RFc25wq3Q4/Fq
QH+sxgmDsN3bNyhregeLQ/VcZJNKLmK1GTxG0Wb4sHBEEWUJ/WG17VzEN6bUhjfdD6D0ljhzycAs
TqgSYNcEtT15FFBDyajzm4BsC7kx2bXzlPg4HlLdgGrzDSTYNBgJZgNaZ3m/ZWpUXBwuIIxzpfJJ
bCUz6gw1uhpBPA9B7vqNLKqO2OE4kJj0I3wI/qr5blXOBAbeRqSPZWsD4ToDM/mELx5jXeHLduvr
CT58Leg/7tGWj+mwKW22fRo2HDxY3pA8RVUPUhNfR+8z47GPQNP9sclNMNEGI/LdWjvetTrroZZU
pyB4xwukQC3bP0KmxzFPeU8uFg/ggwbQRaAOlEt6gj5fwBRXf7mXX95OlQ1JodaHbbcIK6WVdwTU
/1QpnXJHNDpBIgmBa9vffAqO8xA+iVa2Hq/n4mgpWLd7hzhezAT/wFSp6jClOZztblGFn+7Ja3JA
2sA8RC85kFIQCPkXLvxwDY+VtcRS26ErDQNSYdKkmM+IbxNlKX3/l7McaxAyD69eo8zYFHadOzOD
CjX8TxwKPCFUoWPeHGjuROMp6Dd1uYjI80SQLPlgfBrS3ZiOSB2ujBdSMZIXSxLwvZ9lLFDNLuFz
OXeEi89dHq0FRYA5GUADQ1ZmW6ZY5Je/mguwaRWGX91JE67fFIsoCI9YrZgqd3KJhZpE9g8LIQ3L
1YectPR0QdY5ebpGrx3ACzrFNT4riUwFQd9AGi9CZUp0nBBa55/2Ag5CHX0XBMtSrEof5lVMm6PF
rRX5kLTwMdcjdtVMdR1dWx6HaKT1qyugTHAQf2zOshfPWGM4A5WhypaGzl0OJnvXV1f23m/tLFyh
q34Oex7hKVE4NfaVLZh58ouKY5KD22rAPkBOqACXu5aET3n4j7PBgaKeQGfVr/Ux8xBfhOI394a/
LZZJ5C/uCpxlAAFwKEqH6b2e+KeLGGOQVLS4xv2Zul9uko8QFM38G08/GAn9PRkljtJsjDXUH3Ud
1bvsUTYicQtBqyOLyoTI755ks8oi4lKK1yvZDZnf23zT3MqFUgKkWshLCNVEMMb+vaoDej9kqXcw
QmpOc/mlTeXN0O033MTtJpLi4hEVZMFnTt2DzRSOLfNL4DQRkl0X9LCax9cKPFI73qhQ+F4GE3Ii
jnBjC1cPSZqJD+GQcZJY6rveG5WtiHIuB2nJTJAjktWv4EEJpBfcKb2xUiQqlab0SOly1Rh6ci0c
rU3OZosoVCl5dVHSZH5wYhDYd3QY+d3FBn4RLcNp+Ns9XotKra7SDvkqiWfW1+bzOGH+ffVkCtdt
zrY52YZIGsmWsrcLERefxR/PzI9NOMyz5MgoQttI51/lYU8ordWi5BCXW1LuKF/lEyuKj6APin7o
MY2zMgw2bJsXM1urr35UrgjyS1roDvmzsyvdK+kBkFcd+rqm5Y7wvmXzVlSmbCzT3jFtrJMuVvIZ
g7O5EMVozmOFbfaeALMEzQKhXx/ThySVS3DAZ2VXdrKntjNkvV5aAUbZLiktnd2dPdqQ0qVORFjO
R9OKcOxZoA8fbP+/B3UUd0W+td0zqCEMValPa1ukKtauTG5PXapESWYkskMGjL+Z2X1+xAw7TdFQ
0ml46qv0XcDuVzsUlMSrr9yxN8xw8OdQeg4BJ6yMSxDlmPnwxh+R8R2nGyIKIr75+AscywWeTDTJ
tYjDMGMvgPqS/AitC9nl4FLu/etNasMKMmEeImzjVPwSrQmEwPK316nKeRejtBTfFKnjDomP5xkI
o7u+R1c6XWhyyEUpMlAqkRjhKdDekxci2h00spRZHJB3ypJgEz/Icj0J1ALv9zThe1w1pbPP5N6J
fy7sF2Qzwp7B+oDrVzugC6dop6sLTKvtNGXkgZRyHcXG8FkWoMkIlQAOkZ+gJEV/i2gstbD9jTyj
VSsAUrU/Pzp5DJDQF2xo4Zg5O8zYf4JUhveRlDdGJ4GDfnW3jZl7yIPfscZRLLfDH0cOIEsi0tZN
AA1I0zySMHOypfDEq+Oqy/Vc9ZIi6bGKHzdCSCVfwdZOfk+Bf2Prsa4JUD2IuVph7gBt0R24/dfj
SFbaefObDdEo/yI9W1CU7hfBg8/E84Cps1z4JfI+8NMSPsJAeai5f1AfNB3+sJkmt20cSlzKqb7s
ng38pndH/d64+B4iYLM/Hu/OHWqvAoW4fAz8FMFPVQWsIU3yVmRjtu1L1imF6oTTLizyN259dRjq
8+23wDd3uJBuODemUy5zC6RnjGkPNpjrGXpQqsji2/dnuEjKtprqS6vYCfU1nGTWhO36sUU6Vgly
czctWQRQ7Wo6UhMXeyQ6/txZk+hglESystsmc9ffzUwYMQgl7HlEaiGvnHjAL3Re6gImA4IrT3G1
QtIEx7A5BqOiOW4Ney9t8xRDTKTAewiN8zNUgwiMOW3OrMu0ukoTIUudvLfuUjMptvjXBnP3ov0r
KDv4uYrWJVKk77kqUzHk7z84FXnICwKS5jye0hIj1ANF0q4xwkcigLMFOhwb78RgUtJ8cj8TvEFk
nzTUEoi+sTnwB0RVjOuJSyRJIcIJ1zwzP+mzaYtX1nA28/zqFxb6HT5L0iz6ZcevUpVESxhPxTKx
bR3J04tuhxHr46nOKJDd9FMHPdNvhIVZwjJelrt3ywyfZ9bZjpHm6y3+hZX8kv17i8rlFceTb7Bj
2Ht9uv8l2G2NkyPe01JVEsIs9wNzCF6tMJjIlTueWOjEtTcebDLykAxPX4TXmbIOpYbT7eDGlSvZ
NhKLr6o6b3xmzvx+a/rT4UpTf5RhaErKz8VBeH5WylkgCEVEpei1FOnAQw2vFkKQCmD900yGx2UK
d9iR9buLn7ZXcxZJioTTx7KkTc4a9A84WPzzZV8w9xLmtg0uPPwD5fJpTsxZB//t8BNerPOlSvcr
VifBf/7jyQ4c7Mb0ulsuRrqrp8hrAwlsPbu1+M+s0QPzVKF3+1dxCFfg4nccUN0ZKjcINTUUY8h6
Ky5UyXpPjYodgZAVRN6U823jOIjqhSylPB56gNmgCfcP04iYQncGrfC6UZF4JEC40Db2+++Fkmv9
SATxQyKgLTFBagvxtJUBb4Za3R4jg/e4NkLo0J6ekmQ1/ov0ouLLpJRVVbPoZ4C2VS6s3e93XRqi
owj061a/32VoCMJ6E2EfKlXew6gaFjiq3mYwmslZBiMoKmsxMq+2/mo+1iSm3oJ544cu3H+snLkr
rsppIfAhFQ78TeDj3gXqL7cFyaeYmlop3jZJ8Ks7fdQLyesl2qS9d7FzitGfehibVKmKPrvWEBX2
hH13pv3BEmF0NUxubAK4Qa4EkddZjk8KnKHTDuAZ+hHUTPrbLS51syC0gmHlY5z9UPuKfR+Kh5v8
s9AKhRNjEqDstN0FM8R7QUCf/sEBYq+bnEdNn9H8Yy/EpOQCljOSj6XC4muY5eljJZiBkIxE9kkB
4sPR3e/zCErcVe4VSfrMrxTaAsHQyCi/wYNMBTP5UBS4EfGQBrQ+9BjhzUkbSnaGwPEuRCupQWt3
0haAJa8siZpgqL6AFLsVKLIy47J5b/IPK1PPZAhJefh0qhCn9cvQ7L8cOVU0gkwT47B1jMeHZvgu
ypqbmdZm0iaemuXzfqnKh23A97XrfnGoNRwtgw4RKkRYGsR9HNWKRhYTkzzPt6ddhHOK+CBmufGE
Hiem97oNkDzw63SIHXN6H4nesiO1RDIH9y0WQZRmFK6Sm5CS9KkxMO1YHFcg3syeLqouE1/Xxy6b
uSdxfJlD5ZR6L8O+1/UrXTrctIbOYChSivNylAhgOd6u9dVH+rY5AQrlfCd2b23RjVFbW0NFtva+
JVIozhEnV8Aka/fa+qkViVPl/4To6MNBrNReX+F8uVarU/yyA1tGQ+8Nuu1DkpnsY0iBk/EGEKTh
hE4F5AKmttFYpSf96DKQaq/F8yHGjYpE9Mro4mcLwI3NPZ/b+u9udtqkFyJnky5goajIX/fei9xS
Fsa/XTf0lVsbnvh3HGjQo3zPVGYSUOnRBZ0txcLcca/HcsAWSz8c+oUBFED6iJ6MTOolae+2J1eR
KePNNYQqJwTMkBhKpivdOL+gzC+/P9PKY6bNGqeILrqBsMoUA27MdXuNz0pFj40QoFDIWKlNtB1M
RurFgAzqCAeWGXX3PbOeBl8Cn/J8cFU7CnSXzRZWdG7ZlivNmCtnI0TrH5BIigosbMNsMMjsN+7K
AUX9fh4bTWe+bjbpKjSvQm01BXoIk0cCxZdioad+BsT99UescaeA7G1oyuNFqJMXhLl323VIIMwW
AKU7etqfcTLTxKmdogPjKhBnrauTUjuRRUCSoMw2bCa4EPFMaPtFGvurj2K/rrS+H0HCDwAxQxcb
n6pYhrAhPQYmgKyDna608OG5uoOeuDmNRj0PFxHfwAA95uE/lAivHEZOjwCCuobDtE49o69spoN7
7y0e2H2+H5dquHduJ9VDY6RzczZaViFM/Oa9DlwnZLdjAj02G9D/RrhAeQFe6qEHWqJRkeQjMtHX
r4to3ED7pySvGtOGdagDfR47Y6apgAxRJIEmTQXdb3GZ6o3b3JqCR+25EqzRabeQGloh0VfOtRBm
vwRgsfKf7A8I1RmlmrZF4V6JOQ2DwmH4/o+LV9lzyHiwsxx9IBbd6eUWxKW90gofqIhwbFeFcth6
sCyab1h+NsfT3F17w6j4AHcQK7d+zAHG/ZYLpR/Alrgkwky55aDU2p7w3L4UrQBrt4wqa/cU2rX2
xE0tRTRcLFl+65M3dBtHzoYGAzct9ca6r6QsShsLsREDTC8m+OtpUnBjzR/2N0/g/z8ZZSPd4s+6
0mKpFdkLkB8v/x3aSV+LyOrWEzcx+F64F99VLCD6/O+NtnIfU2nMuN5w2y9lfVFr0PUdDFtskIvd
HZEgj8yP5Xs8CNe9Wj/ZE9WRjYu82P/JvqxzxcoksPG6YSTMzMZ1oZquOFrBdcus0a4IeU6LL3E4
ur6S5PW2tc+gmvPsVScPO4mGP+s3stdsO9F2QTr2pjTyQqxsyqEaSUhN4GTNQDGcUelq/9fMxtLU
mGZt6CiOTsZ4eBDE94TNkqq7iuFmiUKtPh6+jiwhtM8Aw31QrRXo0de5L/FiGHrMIL/T352iRuU8
Qd6neFYV1gSlgdSSCNmCSfCBxF81rD9k3bwbFUmLP96btPrZui2FUMxu/X7Vw+XLFdfThAbbB+hU
x2ovwJWSVDgm86jsE+0PBCMVQyOIE6AzNWFXyTcY2vxus7BQJ12iE2c9iYaLsSRU5HwefwG7L0y0
2Fustq5N0GYxkUnFBGzFeISRbxxoB2RmgT2AVdTzJxaMgAEAVkr3Flxe95wLfsxOHtDIhNDv7RAA
jdCCeBq/vxoM6iiZxfFwqxPI8yQS5Ajfy/P6qUZT3St5Fj3lXwYDlUh5ZCc0uiaC1R3cQLblndHV
N1kUFP1BuCB/KTrCeKh8uzviAteBK+Wo7Q0R+WSnSHxyQwB3Yo+XvZvXGazJyegxGsv7l23hHUp0
QTTyzt4wankz0VhRvXiQXZZRkpD/swi89YZq/0vihUKF4VRjXp4nkbaD27l6fRNk6C/5VhM5RyX2
PkJ2xprB/Ul8IEjkZxZxVToQe71L/1qRkK3fa8PHviYIJvNCnda1FsOSbDAJYUCrnaQy9vAak6Z4
80AkhrYSPuyNcj3gFkBNOUooHd2IXtxnC9HIYkveslRCQQbGSqZL3Jo8S5ba26L/Vf5s3XlnAezL
rrMySCK77FN1j0ZH0ClF2QJwqqJ5Vl1ULpV2tbDJoltIigLvlGgh0HvUGMQ7D/loPJuuJ5MRcPrf
x7IYCP2orx+A8UStVoM+IrLScYTfuEGSNUNpmHuGZd+Z9bPY3WU5e/keBepZ8k1BPxqE9mtTSL8i
07DXJTNNTywW1pWL5wMUa4Qa6Z911eANVdT5ZCI2WyQz+9PlAbTSiOyZtaEmVIe1P7jd3POQVzuX
PLa9cgV2jeW/pSivXq3LiCfGcRo2nVi1CxJy1qcNPz69yUWdQIaRZwGfh4o5W1A7VpM7LuqieZVc
iOC8APvirRIA459j/FlrQqSpqOGIitfZFvldrxKm0cK79rNyye87hcct75yW2wPKaNEwXRXj+y//
8IAU7Sc4z1dqOiPOTkG2hkELA83AOtCkUQfIlLtQV9zoingBoAhJ3/eg2osBKSb2sO189AqYV3/L
Rz92u1LsN6p/lxsB0082ao2YnpdoVFGF/IA/rY1l7k4KSyRlwdY6zIOIBUXPfsgbTqwu2Hgf66Cd
HxZiarA+5KmRdch0JFGwrGGutl09+uNgVfsP35Rwl2oLn9CejuX83lbC8h0a6X7sxV7IYIavCj1v
CdJsDUqWbM6UaVEDGCFoq4ywGlQdQYNw5zGb55lht1L9vZdPpHRbItJ7QwldqZaUwT7m8y1eC06J
IuUuUqbgUbRpIiFRWpwQvaKAmhKsVBLPeJFEXDeshCmF//B1m9RqCqJf21nbhjFkdJrV1hm0VQbh
NIyiyfzlmE4rwyohNeeRENF9cHNsr3pbwUrkQZM8LnVl2tsU2UfyGZR9ShqqDHDWNdxebATo06AQ
07+KCPm9xWGpMFRqVO/qIb7kg7JCdgxSzX3FMJ5tsRwUzQNcnFhZfrogtmNSzBAh4EZKD09LVJaM
drAt2YxsmYXyAe+b4lD7wOM3leMuo512ZvBxX5YSYDuCZFCvzBu8VgNEeShjUTYpm6SbcOTRcXqq
4IgTUAyhMAgZuDeP3wXmbo56yvjFRf2KSUjLKu2YNTLhK8Eq91+D4HrR7u2WfRKVz3MK7JTQsnkX
sKTtjYqG4jbaewA9Z8rXgd328r+IeAbv0wN6rW+ma4fM1LbVBdTj/93GxdvlX+2eCzBGv9Up/w2J
XN7BdbtDorGo6hUyw1OkfVL7z0lR6+VmvXPSJ5qqDLclkdzEtLd+SzvElue694+AB5QmNG1MhfTz
MR7nneIryEoMhjad7Wc3aMxTvJ6Xm2KqylGmiagw4QOxLQX5ToSrhSg67+bk6FvUgK94uyTQVhUy
Xtr5pkDV9yjQDIh3OUUDB7bVHu6WDJ/JgwlcIKM7ZN/cl6Gw9heH8L17+1bmL9Z3Bbkq8YBv+7dm
IsXFM0w5I4g9kD4q7mljmn9u9g5lIQYi9tVIV5jvsJGDXOO5kUyvVtvrlsZAW7zeXO94odjAjQHu
Mi0gbDUSDJHFFSatQ4/iXNubMbmC0sP3TOwUEW9xpOpGuVlysGXOPGeGkhH+e/yg+Gg+WAiDHiJ2
5h6SuSC+5y6fmgzaWVvbj4UrT6bpJ8XB9Iy/k1IdNQRFEH5oFxyIH1TZybbTdrE7eLsX4M/NrWk+
cTVK8jIvVQp3EgSnsNjsdlt2dGkQCuq3k7JnmQ/UO/Sgm8zYvc7CvmNCOo2woKlQt8kiczdTd7KI
Rzwq2M+cXfkksmCpJ0omQhpER7krKUJBWuBUbWkrxgT7ivUCTO2urhaUhvou9zP989KSISKYhH+n
idMLDyeclzP+37mXQNuzX8sbSr1FvzVtu6H0CJ/5EzH2jlXGDZHSQXrZGyo50m+PHdImc8FCMH3j
absO4Baif5wa/b2uFGcjtz8IXrGUchnFs/Ti3gbruBHh+AN8VGJStjC5tWxN/W8fkX5AG0B9hsDx
7Ki6qasuJgzKL0Mqm/gTa1dAPqCVoEZb/iuCT1f+f4yz9zIw52dMBGhx2gMNcOJBI4W9Fru0Z/5Y
fjZ8xkhQZADeZ49mDQLnWoFuQ5fdh4hEWznhSMYZGV2JsyoY+1rF9in0wLwoIeJxrNjicAURVMhW
lAinMYyDLsVzqKBXYg/tlD+fwMCLP2WZdxsuOU9OcAb3Mt4/ifo2ayQpKuEnyfHwIEx7VnyHrvfV
DaIJaJNx1hnVdV7T282vY1TtjrExsEuQWt5TzDBv8Keb/zSqStoBXNvPBJtFBvrmXUIqUPR9yT+F
hlesYe0WylL9r3MLKrKUvTL+SjJYqH0vwEKOjPBvbEqO60tGF9yDcCbvBR0/6yYlU/D/BSFCpH5k
N4bytr+7kkM9qe/cBobrrhA939y89o191NJOggrGCQrjJa3jqPVPiWp9+JiDunyKneyT8VIcuT/t
JsHR1O+zJ9Wf1qdK/bxwiIqZ7B7PCvBrSRsn9OQzL/Yr+Nj02cfF9ccO85x4isCl1mJ+hf+vsELo
W+ez91obkhHh7nA7XbOizYhO9lt2w+az4XEGf3ykpIfZLiDAzR1HqX1dhyNOBVlgf5/GKrq261je
cHDKJs0EH2mF7IPUmNEqI9Tk9GSZu9BEyAshyL6uh1wkZur9Md7X4g2zTLMP2/WweDRQbFYk3dov
7bFcFm5l7jpg2q/CGs7kX0dEPqR+Lerb6z6upcG8z/cXBGfkWpVYGdQ+wwQraNF67Yynevm8/P0C
5knep768o4Iu1oXs4qBr3Fx2YG2dW5BO5TcIbVReYY4C46Wikv4Qf9luTuzyngvtsaARABWSJyOH
sDOQIRyN8N84Tm7oliuo8jKR2rAidCzYM6JMiuDFth2QI1ApP8JPLl8wch+n+klP56RhFFDkTa5X
cb7uPAOTBUzcbJegu1ug131PSJ2T632OLyOz18CbFyXV4J/0gJjgrIanNYcvLXou6pCEOGv49+E1
ILzIUz28a4xV9r0xgAWGJ98kbMQpvcIY15L3csEPIzY4vCUMkBoErqRQrJyCj3hPKB3S2x0pN+ne
UrQ9errj8nu+KBQxJYul+yMdJp4JYKwAqmUxucRzDl55bh0z4nstyNAbomOfQ8tHtYRypcUK0UDo
nPTGh9L5nS00xJLzXPIL+ba8aIsAdyWIxypoXlAX85HY3yArIxkUzr+f/6qHPNUnHXqDJxJJcldo
bm9bgC+/I6UDom5zr8tO4VzsQIbzGs/3KgcGPo25YJmi2Cp9s2fFFGWCBndryJigr7y/hUP5sXXB
wPzU2RH7SBmdvg1rfFE6HLnYBmwbYTJbZFcTkETl7bykao+bRInbUDEkx+BjvJiaLRBHsJWMF0O2
sGQgRRP8+p3u7xqYLhI1AT5qLSwHUOsezZ7an3d0yX4jS6K3f0tpKdamv8SVqtEDjwJAWsUBXDFK
1ndGJpJoeFOFFCGpwBNZJ21awqw/HnLiItP5M8OCUpj503YLGjqv+gwQV2Q9FGW4QcpkCXfg4P+1
dH/hzkNUqC619vyJLuVmf/Au8dkf/kjKHe5Ixivr3a38epex3btMJkwJbHcvFaXEhG6v6lC7XEq8
DIqyzt99IHeUyWdsxm+4PveVOe9pWLfjATKfO0RHDovdxPQodG1xsr/WAg75/gGt3cgHg1fkIs7y
p6FCZ8FZEY5zxAIroQ+bLtFFk5Necza1UVMUV3zjbXxQonkRpGbVnBMMtP8WCmAh9+S/BrlbUF72
8rtMOqxRMB3DOuAP0A+AAblqIoc6vwwSQgX5BPstmt55dvAvXgs14UJgnVilh46gXeKjiws2Uobu
GJLUdUOPyiZhb/bHWfImwItGLU1IFF/xXRyImxEeGiXALSBfG6Adkjc8dM13c/4iT6sLLhca/LL/
DaI5eR/weVIiGVXlHkUNSYvsHl7obqTIX/sB3exQtjb0fOsSaZ434g1rC4WTjSuXg/eT0HaDAgdI
gKK/z+qHBEkANy0d9E7/SYtP1fQWtIWelqbbw9JG5MM8PRckzPwQ+sxdAEjJuwUz5Sur0lbq8+tx
nvyy5GteZJDzp2908D28n9mFIqAPo9yDyKaYpy+DMtbxqcSwiyEmFmnnbhXwaud15pvzVEy4H/qW
tMqGhTIRynI7ZYg3E7QxHTjZ8n6Aowh3kilLm6ycG7rbtTr3jDvcd6CD75Tmml3PZ5/ZwgGAms+w
KxX4LpmV0fpSStcBYT4cPA+4CgL+WFzM5Xu4QWhSLjaksFXAEG/ItA13x35NThhOa7pZgdmtlmAF
GYOMaambCu6SlDAEcFHFffUkTGnhvm4LRcIUgtaHMohubVul54HsYEBeWJIZl4lspZ1MoSzI+aQA
5LPtmqKg0Q7JOENvMkYQ/4HcZMsfN4MX9gzY5es40Msb9CpQSxE+EPtRYzRI+cGHgOMVqfp1AHxa
yjf0avkrkuir/eDDuA4p7PaaQnKCSiklmKLsExwEPW2Qoi7OZRiqFeqGJ1nyb+sH+fIjnN+ixIg4
NhsOzZG2XCnvRytMwH5ycLOiFvhStX7dYw0nhh0QaAnbuWlylw8yHHkowCwMD5myo59QNSvO3JIU
PrHufiOEZMKXw+jt9CDQQBG96JTBbeZq8bohMIg5QDz/8xEdS9HlJX9sTnQVqq67/25QdN+li7Z/
b3/F4ms7gm5FQGpHsdTUtdKn9elYoEdpen6aP1UHPhTQgDzVEjXIQgGbLVG4IhScNaL0HJe9EBIf
raUrFNUDfW7ftmQAOUgqIN53Af4tw44rWKCO1LQxfC8VazduKBLDFWIwYDsp+o2i7/iHyjQiYd5v
YzBS/+96TCOr8jE+AQJim7/j06Fmo6auCeB5VCCsqG4vWjsedVHhFZWiIPCYGUFnTsjEURqNlnAa
fOqb7BYRRRNe/9ahbvgVNOW//QUzMlATE3hQ7XtXn63rnA+/eoJAZ+71evuBViehmeHItcJ4igsu
0ZDLfDZIRDQFQv67XxAuEPyNlusLkz4Wra8M4+GKsKjFqkoCCXHii4tmw/4aPSXPhxFgiw2TLlmt
v12yqBZyThRc6WTZG1QvdSgp8H5HqZZYlJWHsSPpu/io0XOqieEZZNs0ZGX9NKhTXqRLu2SyAjmr
FKbYb2lPwzj8k09tXxOEacTDrw8ZlVSYgvGblV52XNcm6yb/PMNAmm1HJvYckWmpCGwuizkNsmsW
rWsFizo38x/4x2qbYQM8fb1r7xQ8AzemjgpCpmmTY/xjRtV2h//PUSuYEGBpS/oLI1+Ei9lwpeba
LLfi87PyeyDePjKQGD1BbtFZbkdgcVCkAmTBxsd5fGnVIJQwLVAcXpg1Y7MH3BpnWoFl3OiYQ6/8
1rQr+vZZ6YLdQ7g685qu9PEiuiQoUlDiVyvKUQ3ohvB2/zN8v4tadUVenhV2fTGgSgFldR0j+pnL
ESn3YFcvAaElL7afIpkhpgjxW75Dvg5sOAS90fVzqm5IElq3wESf5vr9NZQvMBstn0ueMgLxh771
bU/boXYIS5ryVzvNSHrDmawPMDAhj4LjGlKIEcAZkqG8t/f3S0qZDYt3LewbJUAClCnJ15bDCdcZ
oXVCCFOACml2IdcENtHwj5v5umj6Ly6DCk4OFks5F3H75PQqu1+jCq67P7XPBnktPlOLo0titpwO
9ym3po6aHHBpPWlNK4EY1mQjpGD3WQLvARdP5eLljlUFOUai6NfkvboKR3F/n9MmjaNuKEswgpli
AnXz1w4QVUvFsqX4K9NCk2nDnQO31Zy9sSxGydqh4zXmrsuol+hjpM6BEZrtXqd2YYzxgcZvfLsn
+brcXe36o1F73wSupgqNKaBV3EwFwGmZE2JV65vYgc5gWcVKct3aFWTqwaz037PLipRMfi/0y9TQ
+PhIDRtICxVf50uM9Nq7ZyaYfOzmsjH+D22WtfpOi43Q9ar49+3vtGYrPAj5VNFf9Jf2f53f+ya4
RzsScDDkfuhYF7bSVxJ2nYKLNvplcTTWkm8EeG6+SWi75rOARWirlLr1B2NPLSJE72atfkQ6w1vJ
hVSuamp7+Yyz+UDsDR24Sf+MP+5YfZ1Y/iywE6/fx5PU5yyWScEnIZJQTkKIorn79LZYbAxMa/n3
Yh198fBRz1tBp/OJiuFCxlTgPK3smJIcXaff5j4Xja9+nvZJLygGqe4XHvQIULLX6oORFiYWogDb
LDSGcAPbqMsP65VieK7xoRIE1dABRLkPZczFjtHBCht7Ad7iMYZBRbN6r7I7IHAOzHdwSfBEw6o3
4/T59NytAuiE5Hxee2syv/7aGinggTaFAFV9VHi/WDAr8hWoNp0BLVBjvj5mhgYl/Oriz1w0Ithp
zwEbJ69IdBhidT52kLAf0Uh6FQsg53LopMp1HvYll9PyR0WbHemCdY5WIFOvh5p0ZnnDZ/kAnnmD
o1j51HDIrwy+pPMP7FyeZKIQ5COPurKeHkzxWrIRjvPbo0thIWmJqDVPGn7/9QJBoA+x+9ShH3TM
fvKWP+7fCoVrlvBWYJRKOy997dwypNlFwSBbCiAq4iDL+c6UfJU6HC2K6rU9i6KiGHgpGT560cJZ
ClG+lOPXkOSCcPN8LjheBeB5Vd01J+BcUTDollbAkQDWqE0eDw/Xnz5qFmQKc8IzO+l2l363LGHp
3RQxcFkl2h7EkJmCJvOmshe84bAgi0S0HndpZVQm1Lb+IGwJ8X1UlBVr8Y/2aTv1d+ODNt7c7mKf
sx9ffY/ywhwkM5vfy2XoyeAeez2AnEXcu0P5N0U9RM9iLVIQumUwOtrS4kn9qBCMkptHZnjmbOQs
ChhaNA3aYSJacoAJGUi/R2cy4SnIKYDcaz5Li4YePOOpYiGYvp3JZy1hyFw3k68Yk3qfqS1Q4DRn
iczBdt3vC0Z8A5yAfbaTdugKXalgdvZSSp53IYpRAFiHO1+QFFSvXuYu45fti8DfPdvFVx43ESef
m43ryAxED0HQSaWx9oBNziChKGxrKo0c3djgC5oaicPbUXG8sSrDaBB8sMrir4GAYgOP27r1Qlwm
fEcTMPeqJP9yHESKCAIiVFXxYI1TlHrU9zCcUapwJ7jP4WO94dWIIN1opGw1hDjMR+2NwAkHb0NP
rWuhm2JabY3zQNvut6kLMXs3I+/RVavPdZVW/xPm4/TXq9PXCo3MIjzXDvbXYDKSDeI1/iYP1uK7
J1HZBgokzXFUhgV/YSG/phTIf2TGUOE1r38DD6WoQuILGeagRgWRLBVo1XYK98LRwclko1QQIppp
Os1PCtFGZ9R9iWDiOw0MeV68GQVOCdSXPKqydD0oHJUyv3fwEhX68cFvfSSdetzVQm1Og8g0hJmd
JFQXH+s1gTo6z53KaZHcBhDAtuDNEwM/JNTz0PD5LM+qv9394PhlQQctKDfJCGzo6p9b62bt5FXa
rPSMrpqotHbOt1DjyNXU/l0lb0U+zQBWIcQkZERENesMvWuRoq7/C4TjtfQtgPsDXnM7JcZrl4GB
a4O8edcz/Ve/p3KzDcSXTLh+mmCan8n+HPCPaWavsGwM6b8C6p5PBk/G6eYpsWBgBb9XkGHG/Bem
k2O2gkiuK6NsUe8i3O7Tb8nq/y0u0gkWyeLim0iWzgg1mTneJbZwLOVmHICbrzXttFr8ZjanfHMB
BfAU9r/IGPTeKygf3xrjwGvrDYFdtZo6Q841l6Eiwss/JCpdxBKgPH2suqBmKU+5gnPnCFwtf+ZB
BNUdxl9f+F/IjrNqurRQhQhLuGIV8MODAUwo5VAJWPAEkmSIeRDS1C6x48vTVz7oeuHcpJinwZpM
Rjde2TAKwbtnGjw6Z4qLVi6IkChBCoQmKXkQy+IPRtQhnER3btzmrOrExtYWI9BfiS7wN1q8rh05
poB7KJtqhDUEiFqoCnXDbzOJbb+YGJKqjksnjsHJ6vogzqQgwxUY0Pd3Kd5Ec/9wiG+swOzYjHKn
iLXM7zIUGAlgVzkIYMb3wy6Mps8WZl3ERZxLgiEoLVeAknNUvVaqmMtCKTQnAz0jflDwQ0zeVZ5w
ZyIlHe+bSXTiPPWkAC13DAEljnraVi3LHiPtkq1tP7DvzSOvHdENYLOZQ+jbnC5VNQt7KkKK8ftR
GmKHM/YRtx3G13O9E+7RWeH7jz5KFCvTpzQm1kuy0+ZRwagz+8sETi5P4cpfy9B8hQz4Hy4KlIHP
ImB7mOjfsEZYOP1y/HIQSZGcL+pVCv3jn4u+Hiun7PGk84IlRSAfmneV28a0Ij2Vj0SWdTAJazB/
tTquGDCTNO+nP8d4vQ7tGiXQDDyfcNmDZxa9/Om0R3LtsNUSkmBOHUts/GrA3qwliH1dDK9Ytqss
s68nJsV9M9svBPa34veZC89yvMyLBpjDk3NX526rY52yHlDrdVypNPtrA7BjEFm+PBBfWNcA9gyM
isFfUJcN2wgEKMebXitQVupyn04OB/tpK0tsPVp0OmeobHL+PCPCjVcVx4fsVJKLlQRfr0i4pgD/
rmjFkFom2LNCgZMB5wS4kQ+NiV7MHs9hKpqMcrN16lM8XbBVK0qtOnEuoksdbFqAQY7qcTtrHUkU
3cQe6odSS54iLP57qNKWTIqvj51GPJd9rp9x5D9senHOsSgLblOxo4LAR/Tuo7KKVjP28m8RhGwQ
UviFUMl4Pm7b6Y+JbqRr4PKLw6dO15x10HxFKSTNBdSu/gjP9gmPe+A+oTfOavvdsPcM/EvMNaHE
KhiyivzYmWNXOgv/6PVXzkak62LDWBlZrREn9TVcacnZ21Nc94MEGGCdNYZKKLRV37sKHCaFMkmn
AiuaQp7VSgdjbBCyLJdnsfea9Q+G2a1XzNYXTfsoMmg5dMIP9AsTVND7ydenFaSk48KMuepoSWor
G84JPcEoHdyFUHj5UWx5e4Pypg57bfGZcpeJuDDBdl+ADYrp4+vROZS+IGFQjr2ltbUcc26jIfsj
FCwfb+X7ghO4vJBZlDrqZL+aQELozFLOgm9SmJBfLhVNQ32UG7L+Yi8ha8XOiGbVlARP1NLPZwbu
5yM5oZkYxgvm3Rj2+Jm3vtyFAL+5L5fakxujRnIQGpfN7CbDMgLTPiyHK3fGeQ+qQk7+UJGC3k3g
tA2IPCUWv1eCRA5KXf+zqJvDadEcB9lAW00yjBVAIxP6femQl54dN3eo6YwYB9G2p2shavbROgSc
Dl8MPvI16kVPS7LMV46HnVxw+Md6iyxH26w70JvPqS1KhRha5du2+P2Zl/vdZbo1bMDNoiZqmIxL
HCmFnSoVWuVHh6b6/Q76ojenTZ5+5k3WGySOA4lA2MtoObxC7fVqQ9aT2qStT5n51i0kHvcEPPcz
AQGhRGnh9hX8dqZu1i3HAPiv7dJi45p6OL+edeQtM2ILTBJpMITipB2cXcgPK0tnZyu2dhg6VSPl
D/XaCUssjHE5CX1fGRDLK67H0VqzdLaz81MaxcjQlgaNke/UkG+Uyz9yJSb6sNZmAeu55CAM62WC
aYz7MLCyzMqE2UAB+hCk1zOghQKsSI/swo7xy1J/s6cjdg4ZdQiVV8uMtaXeqGnhXWDEIgWKJgSx
LfHU4xsZluihZl2rzO9e5ZCMubo04MaPWhuIh5xWe/g1AOjFwfE2wldZGa8COf0EJqO4BkDxvjEw
60N1bXwWaVcqgzVpZSKFFm07Z1EHgoblstfDkRpEvB9yiNiQLqMTn7eglcT8Llcfy0Utam3HSrfy
DUNvx4SZ9cdH7doqVHGWaxsbDtr1m2FKRodzILz1CGahEm5ZtI6njODfKsxH+sex1J1Cw0jO4+J9
AigjdoXhXK4LhN0LU7RC+GMKxwTBLVO3USieVcErcCI0Sirq/gRG3+di34+NNwjP6wJ4khm9ARiH
K//Vxd3P/i5eh92+hwsbCDYr8Rne5MTjuQlrUQlj+hIV/nPa1R6hXexZjYI6XJrCYz3Z0CbPakhh
5qUq/Qus2caOcFL77fklFKmU3Iw51ZpRYgiNLraaYH+FAtkL/UDgNpV6/ZR0t3l5SmQgR8zBS+hl
RNQ+rHWA+jS1/zN9he6e403UOrEqSZA9kkBv2G/bxrUWyg6Zgdi67vi9/WiVmvDflpXr1F1NPFrI
j/HyGt1m1sOTv1ByL4RoRpApvo6tdH8mcu9iBnkBb1OZyFD/ucPSo9Caw9JXfDuwFSma32Nf6Nqx
ZOWX//ntIEEBAezSX7rMwav/oPpyJOzBEGV2bBKlt57fNU+1HBr2sjh6O1mV6k+BPnB+8+BtPqf4
XzMf5GgJfKh79xXm/lk6psR43A3JorUBdkS0gKpaDuu0vUIHJcxz47ej4LJROrx9/fXe3OkaMfmH
K+XJ5iAnKq5+EBMPGiH8OTd6E7x7vm+aNkq1314xXjvKGKuOfxkDUKU+Nikws4qhIJwfM20pT1cp
e8RiwjS1iiYlHnWsxrKlbA5l/ThBCOcYyF0Dt83eDfiO1F9HJwb0eBHmLyWVow18UhWPjW+4eY2G
JiP+qZG7qEFAkHLo6H8+Tw1s3/DQ/goKpoKVvp/K+5eB/bznaz7PsA4eHPwvKUwbAfpPoWvauE2n
DTFLXoognRh8DjUPwXF/Pb0VrZA5uBIEJuwwBGe5uXRNbHltURvqufo8E3LzUV+r1ubqRCczua2g
2KJ94Q4v1mH4LY5wcg8xlfLG1GekmdXCstgbRbjdpic2Q8qQxWmdg3P/UIweR5UWJX089Hq4iHtF
B4dDnk3F0Hjx3AIRsP0Zj9FpeK/Y0mOHhFISWnO5sxV9dSIHn9lF3zGYaUOHHPNlNxWmna9CqjHL
sUUd7Qjh7vifRsPDnJ9UTKd7lKvzkFsQsmQKt6vak8nghu7FehxE7vhLUL/Ec0ESZNZDuXJ0Xe6L
UmhdgUPpFJbemwLKiruexs3O5m7c8RUTsukjt99hKEaXDsLoTVqFW+J4sAJX7rqhuy9lxPRkaAev
eBifwdmy+V+fVBlfPTEKuxjWf7CEwy9xmIlzhfhQp7Uf0H7ScPFzEAswANpv+iqhSXz7QxQVZQgE
/fz4/b7LPNTFY270UtDzqu4FnqFA4uLZPjz+6KNk9E9AAWlnY8CuAuuYSasCCkXbwDkAH1TwPuZM
YukhgE3CwlyeeIanAIwRflAYsnEH5DU1iisV2AbcMtbbanHnOvJGGBnRUL2hnWM0aS889astgQx+
z27FKMcdU7Zt7unIL08RfSA+39n8dtei/B+aoJCLbHSVdbLxboI6Fj22PFEEW6LwGEn/YDBmOL1Y
8VVf+KgKO5g6J1o62m8TtRiCcYebS8qbl/NvHehvlNTtfi45Li9JFCYwRn7ObC33QZoBSTDqMdg+
/FsKC+docGwZr5H0K/TV3sTdThHszCxM92yNdwUXPJHZ4nOdSYNP27R8spxJKcUPj5TKstiP3Jes
3xkPli9wm7UQ8TkAZ5gU4cirZF8CDVWlesgomdRhtwjvVzPulkT36pRSEnqAJ8/RCEkM5h0JiO1y
Hef9IJyReoD/dhIWEdRL2VeWoibBTE0sHMNxIsCidycqrtqGHGm488ICND3nXD7aDotyukQzwbvm
h34b/ND5WdTTmtOi1luizSQIxBUQLgQQ+4V0Ab6UxFbXgoGfuMfNTX2bh0e6md9iO1oJ32YAg/yY
NxPbThUKekdh9t4lZ668puV2SHnvH3m1QTSkmMwSx1ZBMx0qFrKjAVtYBjp4B5ouf1o6U7wXk6of
oc+J+K+5XdQvqAB1FY9BhSHIw1gR5o7dsqxxZQ4AnsadRgc01hqe7KN/yIOYjCYtiy+YHJaSKNWo
wHCxprEMZysle3q9VF5LrNn4dpwQuHPxd3uNqLOx02Wpq2nzYbbhePIwzPWBWME+BruqP3ppkOkd
7pN2nDRAUqc/bO03ezvZyuDybfcq/uoe5k1lZt2mGFkyXqgJgQQRD1/h7PNHf3yUeubzirNI+QCk
rxo960MtbEhehQHRDamTgupv4n97JKPWzufejdkIoEImpAtQhbI9EefcmFIGU4UF3c5+ACNec48S
i/uOYLik965JJdq4bXEDh2YbXS1maXtG8SpB2n4cYGo7lFk4+YR7cCBgxWJ1u/AOHUcrLmcmXI49
XNSvOL3uLpuTXJnduwgvoFUev/OckcosKpIwC11yOnmY4JCBXCMHPBZ2mZdm3QFEfvLh4WoaoXf+
ah1yF4fJGyY+H4NA/EbUdYPkjhX7bNv2Zok8Gpeg07zMIccTR+Kosfs9RSy2ogZwSUcVycvIxPkU
MsAV+xH9f10V0ScV5XUMTY2LZpTNyaT5UDTpu50OMt/jAuyVbluc/lQJISQ/AvcaEx3weCy3o9Oy
Un0Kc1Rq2WOvSmrdMMrbSlro2tS2inUPsUyDZ0RX3dS5SsuV0x0LRzEac8n8kVEB4h6i4ejiwCN6
vd0Eo6bWZgyrWWVjUEeCbG9hAlWRSK58B/JKz0lbsRhxn3TPxfODsu2XUvVtjiZUYzH6UQwXibo0
LxyaGkfwKdg+HBcMAp5S2ajget7etXKlk6dbAAbuRkeQ/QMk+Oz9oUsK5PL1McwSeiwfwxr+s3I6
7NSgM6RuAUm9Yf7i0LYxCBLZ0emN2nQm5hu/tbq6eoZMjbgVg2MY6jJM70rnZvz9WLx4vJG+8uKc
r/1TlEZpL2bOnU00dTMN9SznqxkLvK2Z1gJNLWHjCZpXX2ho9OZR+JepuNrzDIkW+jGnHxkIuKKu
r7rxe4jFyYlKBEqTtMmb0l8ExmnUpOwcjHCObRZrLKiATeP+dHWsg0ZUHOlJc81pFcczyATXeRNk
k6e/FdmgSk6S5+l6ho2hlw9dSqjLTS+ki4AfFGFZZEzmAEWyI5N7UD7FHCg+DE4fmmmjcijhtePM
9xleqRsdY/kBXq9oG5lWNURFkgP/Lg1yPY4qUfMTmGYdFcVR4sXdowLTSbiwvq18zS2/b5/Ryu1n
86AAx67HkbDnRhkSN0OfJKUlal6iKb6d4RGXm2nkCd/hU1EDRwVAucevAcQsFPd6Sq6RYI6nH/K3
kh2xAiL+JPj1Yx+n9JYLCl7+uu2NtWBevrKT43nnHALx0L1QVYDCbSBCgZQ7cRP8X7WBbwAhlkq8
US0LSL/vLzAYATTl9cxfrkJuvicHXEytD0rMIYLkLjGT1fxe3vC8yRbuJ/JxHrItDeKmclCpuK6N
NVbFblTY5DqdRN9KfkcwxCM3VQJiL8d1A1mJf/0ohj+9+BGvtAV0yOjFiEMqI1O7yW6JT38mz3It
Atzdfh4U/Orqggnbr/LvvP9w+zljWdsYOFQy2H89QKkGZdEyQzIC/Fvnzix3plj3pRapwgJc+oKh
iOqjo2rAjEBMjmNakE68vUidETzODa3l9KfSwKxmLTUDGVq5x5nP1kfG5qgHgvrYA/zN9YvGgrBE
+JEKV+Jmb3KSALojsVdldegZctpQe/mBZSWfEMIo6EXVtM2y/VWG8Kgu66IQWZ782rXb2FePmXP/
zkFtGSHE0fnEHMgLQR/Fh9vY6Ds1SleWzDJo6wjWKHgwMBm5WqvIafAO8lFnYEIOKSL4ay4nlyHq
g3CTYMVQgn0l1/OY/C2vZ4V48THtC0TrWYs2ib8Y4Lh2/R90bpofGFgKeu5JEHh9HAUW0lEEcxPC
7JojLyv4/3sioB3nzlBrUIPUK5GFW2pMnAjpRAmFtyr+0fAvsd0CdfGIlI9ZjhHmjpnH4YRWjAqJ
3BZGTLTrHtGO3LXjVaAXAs/l9YDNuAO/Fe3iKZkIHxTkzzZ8yRZ2vicmun2kWh40uTsQzc1Z7Afa
4kOhEZzWXCl2JLT0SsawIBrsemEen8N86Hbwb/1Xrcz9Vy3qn9FcsccWke7GcGUOEBHgv8SnfwBH
7lPtGGASMuae1SgHPOwh6JoiqOM0Pf81E8/+CsCABhM/w0kbg7mGbThcRjZEYW8DEWgcm6bj8Yd3
tyTPg+gF60vwcsFqmwG2s6aZKad/mYEWaEOC/7m+a01YOvEgPH9KPzQA+6VNp0FuRrPL9aXREHUR
aThSFKzx5NTk1gKPW3EtaLTKZC7kLsCrEfWL2fzhuNIpXKQsciEV0NInNxJcyk7/sL45ov923UPh
26uusGFi7iwuGitB4VPxMzelFTyeJDYdriX6drEjlZiVvV+xgMAJUQufY/vR1TMn/dLG42gLsJ9/
6qw+sVc4DynyqZ8ndNNGlgU91GQaEvITKpbi0SMthiQCxTyMLXNmi+okoZLu8GkAPH3+ue+NWqnh
DU/pRibHpwPnih8E18I+PU9h4LvQ6Xt87k8SxhK854SQzSCyYJy/2sA3dcDKd0ncDTV8JZ9s62Fw
iKIfNamwz4uKwC29b6Xu1TJ7HZo3MGG/vLp72sCcwinL1JQUI5nIooz11fcoAzlU2gPhjoRJ2SsF
aIxxpkaNvYLzbh1ZsNG8nV9H5yRE0CQLrMj177UUzWHjc3QjB64uUU1OujoVisyzhyj2E9XTmcdn
jeqJnfKJxCZKC2NNND4ukQv3OYp+uCdF67OGkvq58tBnMAr149XjrPNk4Ccti2A9DY/5mc8u5ExK
m+lMsazoW/ld23Y=
`protect end_protected
