-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
cD1WioCIFjEb3rzypC/FNw+SEcABv3TwyZlK3NMhzgIKw9mRFCowmhkQ5EDm1gv4
8GvKUIxqRW7GVeePYJzWp+qiTxprEMmReCTh5JbCW1smVORXHMI8eVgYIt6G0y10
0L4EwVFunhgfwDcDMW8fkpoK1qL7KKiKvXexIYmiCVo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 20072)

`protect DATA_BLOCK
B7NVCJylIYOaeblb0JLKpyoXTpjh89gLyTl0I279hXOuskOLtAFA7WFyJiDJoW21
R7+6bvM3CIVFjX3Iki2z7UdESNWEU3JIslVDMN8OgC2gytLg+zaRJiqb0shF4yVC
+rzPy08wnKpf7DjafYqSMLeI5R8K+CPMWYW1WuHjoiJTZ3N8GEWdtCKyK0o4xwDx
U7dmrCBS2WlQoumUJRRO0+ur74f2cmDpmkehQYz3jvD9bq6dDGandfGh8jLFiW+h
EoXa/wFUPZB+WuUS8nMR5XxY3l+ZzGFc2KDA7WugTAQThjRyaCUL+icIVs7Dylkg
XcpXvbVreczMHsxiUBlilAVcq1rzEZLJ6ybDvhOF92L4QqLNQOqRH7qgT2gybRes
Naxjz9N6Rx/9lsrDy50Y02apGojH1MDG/hze9jeTbNTf8Aybl1AjumYaVckxJeIt
nASPWNPV0KysWuk7GmXYF1upm0qMNOSUvRy0H2C6iHjHEX089e2UCBt0kalV3S+n
kIRHB+vOKx7WCei9dpEo9HHdiakcAYxSuGZlwIM8fCiDo3S4AEI6Gt+eKcdJVf11
+BmPq/MyWHtAuDo3VGi8TkvnQ3Yz36J71HnoPkewdu9NMq9XiZfjDMlF3Gwob4nc
2AckpMC2v8vfbBe23IXxtWX9av0efbgn+nga8cs38ngYpRO767/ZJTyOoCcTnCKF
4xR7Yzcj300RyykkEZDiBaXxEUTPrWkoLQBVlFGcfhcZxqLN6zF6JHoZ7SEyEAGA
VyV3PAwnFZ0z3NUNkaRUPEgCJWS03YwXS3urvdHgk/0tvJWh8MGLHEU0gv+tEYH4
+5kxewEfjNfBJbdcXX6cFYh3w7Mf3LI3VXlKciNIA+a/cTOG9Ofqfu3FCSkgrnRh
E7HZ0r6iueTqZTJg9ToMuj2WyvDE1YDwlhke4bVwaxYPlYG3WEySzUV6J1S0Mo/1
kE5vuoECY5bhpCvDm5NEC5ALChEf6Lx9jKxM21MQdDxPHh/fr4CpUJ0SjPowFXw0
2Ey4i5VfceqX1i1WqS2yOd+TA+snlWDsvmO2U/h3ivfJ347e+jz6100RW0fXHTx/
JWtPRI32FjtApIK7lGw1KlfnuybBgrMbxjdjuRb4iMzib9Yry17ON3MxHVlIKd9f
SPJdwq+BLXxWE3ag1kH589jjS2x6cB8nmVJokHSoPAO2UxjDjVmSJ8e1oHY/Ukhu
M1ylyYP4BTNg76JLGAuxW/tz1XTN5baRzAOJj6uroJU3QUFAE5EKk32yPlbfDFAW
PsYCj3Kk9OE2T98zhkF+APLwOsuoJAsrmo8GAValGxtbrbc67SBKe0MtTwk9J2gq
IPJJ6trTpFBJR8extu9PvtCrX6YAegyv9Er9llhGExueyyKpjW6BsNO7aphzGzAN
7LkjL+YpQwja6z61IV5zNjDIC71/zjHWqqZVYatbHvYd3d4YnwVGi+gmzd+AW2FQ
icfgoWWwknClRDCZe7E0ECec1KNuf4boslPp49UwvGrbLyjUY9kajIpH2sTJ5ofI
JOLMuBgER93KjbTAltCQ0Hn/oPQbqeuFQXEnzU+1VkRJEoZ063sAY04CogmxRStU
k+irrkZwcWktZyXBoW1wlH7GXJgWFUYGgAzKWG24zhKrKnXHYkkJLxFqwVij1B3p
yrYTEvcFsLW6Nqmf9HPhlPGYSe2HIsYR8W2vh+XoZsFp2aJWxgy2iEYeKWcHSygp
JMdyUOFjd6We8ZZ4u/shMZjZMTdL1iuIjZjngUo7phJGExYK5enV+moLATLJ7PaH
gg18M3uwzE12NIWW4g4ASSd4K3uKDotYTVpRIjBpbfJkhQltQXZ9cMvFcn5YNiPy
CMj6VI322ZHLa33pE0JfrGrDbm4IVQK7pV/oRgR8tJVFG7bHQGmBUXEXfMMlYt7B
SiDHP22cU0qRZviATyy4bBAWWH+yzVj4J3tKEaKKfllNDmZBjX66WMIHBNrB0Vji
ad2E+iYoM3AcHGiD54kPvxFZl4+EtMMRhgDj42W8W22VnoHQ25jlicXiQRdqqJUu
+JPHDkpDk/Wa95E+ijVLz/qZE4qru81MQ1qXVulpMw+G2BbjJ+kZ7UOuqQRR2LaK
Fnca2d1oXMitU6m0BAg6VUZrl102uHZk+YRRxKFyykQbXF3KwvunyZn5QtM01c4h
Qs+dBaMG6W0PtoSFqbVmCJ+agCeKuXw8Lrfr4S1g8z6XY4XSUiSwJm5Oachbd02Y
YHEF/IFzmgCPfDmrTg4ZXPzb2cfMWWmi49sUmkIUdWsKME/7qyAcnxveMESEHs+l
T3fHJb82XQCaoBYQerwX90iJ/rNtTIquGLIID94+pbHhtcvueK+/LwlovGmfC4UF
qN6mswjWO12KtPmwqu9egP/DKemLAq5Ua9zdpDhKOuKIJDZexH7/7iFAH251+dP0
5XIiH5XpPNQAg6ZfbKrh9ApixkdSls1PNvDJJLweZQrKn+7NjV7H+FlnU7KeqZLw
eI2ZTJsgIPVaqkiuJRFXqyS92308Wb/08HXX5a5JzFr9+VLr7vfy9Y8fQL5ozsxf
0XLy4lET3VLcqSuw/jb3FHWmLuT48yAkYF3Gf1I8utpnn/JXnNxq0cgaXijBPalQ
hT6Ujq9VsRIjNU1g3V/yCIrHnIc8SdHlyESCWc3KEqN3MiyfzXBr4LJtOFmUhgKk
2ejPi+9Z8/uBnZHZcfrBAPCeWzctrjLCMWltC8QtkBQOprvP3d2QDGhDE4/Pf2ak
wHSxODmAi2CIgt5YQnVA2JhoxL9KGYqiIuKFjfX/gaQcHkNTgOFJJ0Bffq7JSPd5
/m8z9/VSR88AJIHtb4g+SuGJigerSKk9Xk3x95u6VurpPQaDDRjBPVX9DEFRLfj7
GWoxbCZ92bhpTyJUkH8pKcyGqLuylS24pCzBBZVMDy09UA2FYzWq+mDG4qJaCdoP
mIX02mdHFpyM54FDbQCShSPtgzoVyuDhOi36+MYUqyrUHFjpewZoJAutrL7pPmnD
t3ajoTkkCsocOBx4lMuFaOBN5ayuf6qOauvy/PE5I6zRDNTzLoi8i7FoTEfuDmJ8
dxcn0zkGpjyG8PLEQJeJqchajHYGDXPdZV64L67wFzTfT45xlNKbpZFT3kvog/Bu
zqcryOeitufnyF50LfajFixm7pp7yOAV8SoDVX2ZPQVCaHtlb1etuqUWrejYNEJN
RD+dR2JU+Yv9Zc1saiGxaabKILDjPgCEDafhzYAvwx1R0gH97/yriRhfK15N+ifh
yp0RPGfigqAf1C7uPGByajXMuc201Q0bXwfJ85TpInk3IP8b9MoZQIVfXGIJ7+PO
ra9rtemHbdWpfumeHEN8RPJh/czz15D8669r52kD7xRdURXJB9zAjXi+PIHqlIyt
AovuJ1e25KGQfNUtb5B2KACN2p2uoXIJwwlVmeOw6Gfr0rcRwuPTZ/Y3+hzBfNcz
UK2jB08rgwp1XNl4iscAuU2JCE6XM0ZqYVsufhelAKkt2BRBfRvPNpJwQZ5ONwo7
IiSDaOXPvp/UZvyPOk6vPfVudq9mFs1i9OJzUcoJJr/d8qk0XjRsFZlHLdYUXJYN
AgIQ60Iisfl4JkK7BOt6ACJxdccy8zn6GgVLB69ORRP3VHU1DKbVswmBNU4jF0FG
RuMy+M5hp4gAomI9chMMUs6+KrcEIgiVi+lco9PtdJWebiKxoWUOYpbiTTN29N0N
rpgkI6w1A1emnsIHALonStmAHn3o75hyZT6/AevFuOhltO+fC9c1oHVSUtXNylnC
CWUNjM/YJZwNnu5OmcNHNNJMH+89M6LNBqSyHdHU4ZKkjId6dCYtEs5nQn0UuTnr
z/8GLPHlL2xsjFopNqdqyj5zieEUb9ztPt5n/DReNFs4U/RX3c8uhSL8vv2BVdEH
7yeJQcoTmOO6ROKYl7/PfdFQzWIaiNGPHDLuPgpXugMFNneK6go0KF13jvSVQ9CN
cXzzobgsL+HvRwbdqTPTBkYpc34CjKtEnvs61Df84KS6Wjwjb0CscRQ4sC9VF3b0
yasGAXH/Z+WORWFoIb4/Vzr3kRGmYwnIBEDbe3Msjy9gVY683tmATm6HVpGxjbQr
YqGeZ6WYoWcrdtt676tXiaBFEKZIsE21xVCK75X2syyw1SEswLsxYy3k6UtOvLwH
OmtangmWHSHOIKgRaRGeimqxiVJVI5sH+MoDNMupF5tFXqF9ftlkSO7Ilrv6t2e8
4RsXbArV1yl0AGYTZ3OjGPowYBPhlmQlI+fZWJT3JvXaT+xNU26SFo7CDfz7AIH9
Rtl62lQ/4kPoPEqUYXJiRghcCVno7Pw2TA4OpUT2QyNrXNGGKZ10dIRnSLlr4Kk0
eV7GLsOy8J9J53oNXHThZwJ0nHCGkA6qthugL4j77iuLLGv7zxt4zA/C2tI61Yy2
xFUVxwEDR6gNMOVgxYtrZfs/UV4OrWAIOfNqpZFTNXPdSnCc0PeiB7aLFjlYXIQd
mAJKJcRTO0bnPWHcqHz/n3DiLnkMq1Skh2QbWcr9vxEYv0fmglzVM3qWX4dfldNb
LWy+vJXChq8J0dZ7NeAhRIp1LFXIBi0Sl0JqdFFZbGWcdHdYagkLAItIJ5RRmPPP
s+diPeOzY7eLpukqq9yMNCxW46xQXTgDUoA0qD58vYBB+XjoV2gbWQ9YXrD8cJeI
4nyN7vvRsNPe4ns3PEQFPHErupcOPwGSlXE018/Ej9cGdO8sTELHpwidPiecMHF5
7kL5bruzcO22l4V9hc1Da7suWJgAP0V/jM5Fr0FaIHA1Ya4WZwrx6IJux2qeix/6
QxDnm3MuzSZ2wpDFRQQJAZnFoWbUMu0NbZvmS2AYB82LB3PbztD2HtIdpZ7BtHZB
QtLwlFp6Y6oL0L7sUlP2wn8sxFfu7CxlnudedbeR7xrabbB9VcwbZ/hSmV5H9mLo
k785fQ+bITqIIAu1h3b68hZYDiJsVUSr8Qf3SKHD57+xluopbCilLpvdL4gTYhDf
Rjf4SbrIWY2mvgh2l5Fnzn48yAG1bQ5vYxUjqeilkJq6NgVKpA+8f5ejL87y/ntq
sWqh6GOPOx8YxycmD8FZrwv0SMfNLEVep038EGpR+xpngHuZMlpI5ZNqcU1HUopB
UaVBndgcOgB19m01Gq/VV6FbRf9p5tW/S0GEiHaozfDaMK+EfSFvnWxeVCBY+BtG
nM6norznwqoCvnjbK4mZ3B2fmGxP5rMWLupnPoEs/pvQmBpsjfk4R1HX7xNN95GM
tUE4GLnehxbIkBWHp8paJC7tuZlc2XFvB1QoaawZCUjig9e8PMi/C0+hcWjxUN4k
d/3wZQ8h2nd+kxumQhub636MMYbV/awHiiT6MEhqFdOAzWxBgP951SeDPDZHOABB
fAOYiKi4WpIHSpv8Qaap8bLhCHiI6PWMrwTHuNv/QyH4V1vG2LBwpO7lZoMPuntw
3eI1zdCNWJ7+86cJ7bY+JJ7AJ641qGQ4EUOFLpDMstElDJe70cV8ZXK/ohsrTvv2
ksKpmWg7RtrL51LouxedecTKGEoHP6+se/gGmLsTyNdq1ChrKlRXpDfUxh8bnVGs
JYoqKRaE+0Z2eLUvCw/2Yb4MXQUVThGtey1uRQEAFCqo4FWmjEl6Lq528ngLDT4J
XsBpyzJNN3MIWP8Kgb4g2+0kYkl6iroLk3paU6JGJVjXJlWrRCcJv8/dJSVu5lYG
m6IJo03itUc8DKz/+7Kn3/HfIBoPg8FqBBfoV21cY+1bQZq9XVLw9oZFtLgL5Q9N
chQldw97vLB4uk6uurdiGX1MAtffSTZfkmJ8NknLzm4kAk1gBRU4mmR5HMx8dZaH
blxcZFRU/TLui7eiDY5ZWyTnlXCtIS/Xi0GZUgG1mxDCNlcqIlvfjzNG0U9G+mCT
/0SlTDDldRWgPtS7RsofVIDLlOIDw6waTEY1OugOqqcSX3UNG0quc4ot4tSpy8q7
XwPmWR3n/EtlwL7QTRLMNKuw0jb8R7JBq1ZWr4EjWZNYuGOBGT0hVRRiC3gkwfoL
mL7acc3JyDpINgpk54ljWoD95w3uMCHq3R+9Zyb3MbBgE8CYZPsfXPI33bEF1oea
a0DBklwHONvDiENvC4aFSo4yaP1EfHrtVfAlYYAOhqaabdgYWoZC7RJlgzoTRuAI
G+NvrtdI39Lp/L+banRiVbVvDFnp39TSBmp6H1BXYUGVhujXptsV+TUhB8R/nm29
DsonUGiZBZzKQ2aP5PrvNrcTqpGTl4/+Jkv4JncrWc2CN4SQwpXC74xKo/kqxy8V
C0and2X3Y9dM6I2xDwkqaPPC2rWA6kJ2s6PIjMC1fchtUDOtTPCDdVtkYR8m+cka
9y5o5uqYGupHjNE3cW/3VMnycxo27b2Xv6b6GBZ2d/HIAUA92NEDibXC7jhfWmF+
lnII7609qLawapBYZWzUOwAviPz6QPnk4RBMDtxvgf9eeQ8hH1bmyo2HlI1tBZmm
FzaHIAzxUhul3gRljSShzpbyrv0M7Wwmdin9AQqKB2XUnSU1Xm5TXxQ3x06k4JwN
c1InJJonvoPB88mRtkSYBJf6mNYsheYYRsda85DFxSVVzS5oANng37J3XO0iGSag
qMB9Sd0a0vrvUL9dt1RAEXCheeDuRTC56ci7v7O0mahaTu76L/7LFBpsWc2rtUsW
Jn+D3NpAkr9D/sIoxB3ef7ZEYXTQGvnD3OOqrKQNjO7kFjr/cDp3NMpAO1eEQ16O
N9W/xWeGovOOUfrbLMjMw7NQcyueYZ6tQcYUJ2Cjmcm1uM8mAcaZHsnHiZ0tmOQi
LW7ETNC+ykl8Gt8W9a9X/2xJKU1KN/3WeY1ujGWhi4bD1sTXp7vjmV1Lo6Jl+3Oj
KvKeHgJBSQAd4YXJyVl8k6wLg6PPhgY43jHWDIRksitPwXfkCei8kUbgbqlR+Xkv
Q+4rypv3fann5vu62m+EFq25v0IFYToasmD5Fe+UUN6iTb/VbA2IYzRqpSDUfmOP
NLEqIgViyHgoVVSklWXXb18dfrXofReKS19qAqZ3D5/mxw9WasyYJSfd4BFKC/00
RJeuTFPnWjgSrptolmZRDqCnBxbXbnANgQ54eA4fSI3qORh+iqnBllSuQYcBL//K
ZK6eShj17hCYjvNnJ3ivi4/b/pVPBt83nwmJzWG5cFz/YBKyd4Z2ps8AlhyOiji9
/Uys9YAslEJup+bEU9A6Rn/xpBTaHA29gCJzQui1Z3GAveHjS5HCGEQHUJhgIcm2
6nsbLHsMWY5eRM0fT6Jn0yJ9qW3bNknQmYWUxnf2kFHetJWiGzsivFaEGFP/dG8d
tc0f2F1GHRC3TM5YeNL3xwuf0jsEV+CL+V99pOMKlwyg717zGQsxra3PPlV/8tsY
jovoTpqdPaT6RYw0tLN+54Nq1ByojiE69DkHu/o8XrtwhRO06lc0MevxGtc6IbM6
mRO71la7GNqcop8IRUkJCG8xBOxyFbQeFhrWUUFmvPp6XYWJNTq9TxKedSh/qGPr
8wUiia3Ht2oYtAeLOwE6hgE8E05kX+ByjqjtKHWejm8RkHPfgVTDV6U6m6drvKe7
Ka4eK+6DQkdyoqwXXWuOjbEz8IfAHbzZHem5H6ssNRaNOpNLHW3N/Mu8lKtAr3v0
KEaeyJIiXGlnwANyTWWPJiehFVA8HlOailM0fS708zKGIl6YwieK7UE4+VYbcRMB
CDQTJ407ndTcATkZztG1l+DyT2nKulqYLsnD3CG0MvqfTc7J7rvF7jeo0LQ0pk4a
H2y+h1BeJcvAs9g8OZD2rlmKntzAlwpyA1hZjqnbkJaXqPNVz9ETv3A2nwG3s/Fx
Rnkvco3dWeGOKfySOGUJY24eF8KhUOJfMDulp8kzJURJoulEv24cEdZESN84rr8q
FX99A57GaeFsizmfMue8+otDGX+5cS9rzi8OToiGNGXf3jJZW5nWz5pD8O4dbLO7
gjEg+3V/ffjRrlq2z/LoUw2Qn7wan7mCIGAm1yxzMIYClAYw6FYDAyuZpWKM0D76
TX/2xAV0jBD/DsQY1xn7eU9bSeLziMADAu5zZSDhKSKebuV3wOqQUo8zScp1+HuM
fmTyFBXaGssp9dnuDQsL9Kcc5jgEk5DtsTWusvkZPiow7ZzBnpFQglkR+jT246S9
6Vdrx+QMY9hezCt1BxgxNkmCnfg/i/hgAoE9+av4VfqysL6vw1tCYciRo7pYswVD
AVSJYuWqKJ/57O56Jdnhkshcq0UmIVr4UGAhBv2d5A/P/qUk937ZGCjIr/NrcgQp
in6N33qAof+Njf9ydFcg8QMU42Bbkos0I4XMUILmSli9c1oJgc01XHliyfPiv8wL
MnAChxAsFWsIndQkCWTRQaMBWErDYvMZR3ffELtubipx5nwN6lYfo7nHFmMq5xO5
erQ+zEheQGJP+ejx3QnwRWk8OSMhCVhZMkFyWbYyt1JcVDfwbxmBHpndV0jbAIQD
tsTOhbN4PhllZ34eSyFUHwmh3Ow1vCtlEYH3LvN9ul05d3TDt4xREyZ6xl2UiTIz
Z6L5ZG1swutlaacC5CtAfYvxEAc/a7TI6gLeSPQWiDFz5U4nsIclmG3IBPFU/87j
F5QE/dlGJWUDE3PLopUrX00ynuwrj/yetdFp1vr9S6z1X2MNpMDwVxuJ+2VBi2nP
rlGu9nDEUlfo38uy6CAB+EAzPC4RI9rfRV3nuxP5W2ZoJKfGIL/meONmRALWtJBh
aAsk5ZGiLLrNbJiEAsvPGAMLaajkh/6mrQsuLoXrpgQRQx4QazS4hCJGMmSnanb+
zrmzjeE31ndnXi9rxprg0Go4mRqnLBZglmADtn9K+C6E2JJFSI8RGmGpTSVLI1M0
FBzLS1GcYcutKHPhVftW+XGLmTmNyXK+iSdELn8mhLgX1IDU/0I+OdLD56O7wkhv
T96lernq3P0EoGZvkhFepdzDmUPGMW6zRp6rcfcVgwmx6aOC25dA3ycC1D1AXJlq
rPSmn1LMmi90QDWGci1lYa9a+S37miwFAEcqSl2M9HIXj1yy6fHOrreWgRE4v+yH
xVBNkd+w0wpUFQ0qHmKj2hjF6ZuRkmGZ8G+VmdUncR2qNlBcZbBB+dD9R3PRfDAe
fDL/5nAaFUVabVTYtGlDWW0Ta5E9OP2As4BJyfAzj39m2GQxRdlCb9oiX7BmrsfY
6GcYMnH5rWSnXa3Jt0Fbo65Y8MaAOWYu+8JF5KH0kUYrv5eo4viuvzYe5xS44ssM
MFJgPSqrmoaitHtgIBQhKdm3uhmz7gPG1v7RsZqj3fXTb8b8yOFlvjqKhOggkdov
zRdYdCPukingeBlFRqiUOBqqJ5GFyhWV3rWTW+d1vFvlctEeBKFZF+nuM07s33HL
NavDFFwx8Z3k35E9OzZlDwWUsXQqA8sC5WK48lNXovxTFMdaXMdGTe/txoVA/TGP
hFAz5o3x3KfkWqvgKliRJbPnd5UllGHuyHSXsrkQTjIRwOViO1x7JCo+PB+ggk6N
zb5fw3uY5c15LkeT+HyXZoV7Y65aZAHxYYHktELUopCzdX6Q62bkpb53OOqHbBBO
o5UgNVs/SuKIx/eAmJZsMVoUyxgZbXkSAmos85wiHobydevLZikKsiNaCLLEwoav
AKgOCIcyG+n0+kPay0ev+lalYs01PHW6b+7XnnXrnNfTHRRDvZjRKNKVsFlam+hy
ApLMEF8r2uEtAODXnvDs+HQFkUbaki7rHi7sCbgWWaQD1ssENbjV12WZot4OTItc
AfZJs0Q5iFDCSuZ0PC2AnZ0jK0yhLdx3EaVRdTiE6+pthlJHrinDsMEO3UIv2p5D
CNr9BKtYaz7H+24W7IKL2PucTKMyjh3Q1kT1GWtItsDWAY5AGvUnmJvkDNBo5l8m
05txykZ1A5N5tLf3KBV5nwfjwH3iMAFw4NVyp7cMS6nra3GSvREisujJV74b+9hp
nA5uIWvjRnpb/fNk+y/AAoj5yztTvR3h6DMJ988rRdU951ioerh1q0ofFJgfmBYQ
Ozgu8oB6u70BoiBbjjc56QnkLK57vADrTW4hZCv7eaKRU2Szjk9i0lkGRaYwGypH
oNmCFiytAaoyM5OWi8S1WrYOZcbx3Xw9X974Q6//vN2WNxoBI9pmWMUdWOCgoCB1
SckBX/D/tjOFcrXq3hqQiBFJyDw5M7yhJxdpwNG4gqcvkUmrv9aAxOjymNNuDpLI
ImVvv1wjf20tnU32DUxIKlE6GCDS91owcBznYDKZrjLyt4JsndprtasYSD+ndbSf
MVILtHVrPoLZqH0J4126HC6ZRBPa+rUYuyUZsUnaHMgv8FIShUMHMzwBSOyFMS2d
9vzGx7ynMkV1rmdkdjKcZbozQx4ioErT1GRAavYgEPmxgbRK/Oc/R1Hgpj4LQ/jb
zQpMN1JhIj02zuBXiyvVTMccFfqp4EpwABKgzlyS/c7uv1vY5GtMVU+hV7SUonev
Zg7wGZ6ppf37IPomTTsUdSBi1Dw4QL8t2NHLfgCTCCH11+EwF7v5FvBtVR3DnD6C
kTHGZyeQLVz68MNRcaDqfkpb31sJSRw0rvH4FeDPJi6S3hFsNylt+A+KBH6LNAWx
qdZrlonFKAinIrfDV89hRamcjVe1ivI4o221XeuC/mbIDOAGMEqav5ADL2eSpy5p
2acq9RCSsdBTOY7Ay3DQI6wxUB2q2t3xdIgcQKy2tinJh7hWeRH9cqcBWRb5vde/
Z/+dymbCJMHo7t9ZcPvOyd4mJ8dhTQ8lU9uL1UBB8j7oQUg4CqFT1vI7/LxMlAme
JmpPwPmroQORFuFDAViVesC9n8OxA/UbkUeUTT6qv6NW06QacBKj3sX99q7kffw+
NTWJI3HNa39CDPR3I7VfgygJtSm31Jkks6MZQbaU2Tex+RxBp0odX7FOTYBkXyQe
JSZ8OqNquDQIFdpdS/oxS8NUJ+JlVVGxu9AN49FUqclD1nedQGqkz4/CF0eRc/v1
/grtBouA3PnnwlEhR6kHV6oyUQJXHEE9oqYcPyxdsCIZZJVUr/PdVc26C0ysiVWr
DSZ0a12UTYBE+o45xp9hptcH3Dxhr438+O2+fqsvnQQMqYItO6YFbXCDu0BwspFh
kzebMM8sfMzgJDRKrrb8yhN3k9Sl4tRaoCHeIhElHke3D81HorAkCXpKXd25+Sla
7j4HBFpbr9ycRcq3PXBdbtOpqrtvUyfkIKlngMH/jAm/IVfPaOolBq6uQMCF/Gni
sZBarpEzs37iVPge4gXzhpgeEBo2/NX49RhSOi5GpZXYSJ+eCAtNX75Si7H+5KR5
vcaBwz4khGX287alAHNM80T9dO2tLLV/P4Iwi3U6NetpyqIZe6YOx3oHlYQn+AMw
RFcQzmHdaH7fDUkA9MyPv5I9X0sPOtK4Q9Qa5j6dvDi/CZ5e8OHHscu5784+GBX+
mcvdUBH2nB+xnxFYcI1CbMXIcnGaKlGOxrCIYoPrRk1fRTnnvVlIaLb9esEMDpc8
rrd9qV30fhetnu+MZgofGEWGDLbzneI0nkXWKyS0rvLyh8m7mJxmHD6QErrZq7I0
okLoSPawVyqcmL0/GtSBRRXAlPfIybIcEzbOwfdk+tjXV1z/UREE+17BipVhnBCL
S1fHIDoGd0DtBM0wG91PUyG9CIgQtgwFOMJA2Gz3nH6+jyBgvvdb5Au2ltRHekpU
z+G4ZjZUblMn2W3t6gHr1vtgscZku42JRoeL250VT71yqmuFE1EinqSQsovT7V4/
r3WnjnEu1wtIdIdEdC1XaWn0LxK62RK9MhFNTZ7IzjrmON851l4pYD8/iDjW1a3E
G9IMH1f21SYplIJp36ChdcNIFsCSZWbJE/KfQB0G5MsnvyQVYcJvmJz0wuMIyfmw
wL3bW7DEBAksOLZ5dxbbUhnTTeDLtEwAZjB+kQUkbbQdqS50SZ/iXNzRWbGy15Cb
qCxECN3sLBgbKfgczUzo+0pFTAsy9YzFp3QCFoC16hdg7eNodHXfHI3Ra7tSHnUu
vLpvbOx57Kz+WfBJk1hVW3tQA82D3noavhRNjdt3YHKc0+rkEa142chCicNjTSw/
bvPYk5vt5IDhxyuWA/Y7NAi3aCPRkhOZe6wHMFxjEHBb9ZpFgHOBlR5uuH4itU5S
S4jUyqzAA1SrlFkgXKxbmDKt038gf9sZWi3gyfqPPG5GS/1vcizcXXLFVAg6e10n
meuG0VJrzmytKFW3hCDIutRwfxHrDGt4gC7D4YxYbSfflWRbhzjTryo3NA4f6DZN
QDLPwXBe9thQAkq2+ZnlwiwtuNy4kXfUbKbPfb2A1Q6mg+b4/BplvN6z1dyBuTai
bf2/3hNTgblhdjbGN4wedwmW25wLJnInhOsSqN/j1VteuI3extRBwIQY5plkeA4d
3432u6pFX7G8nzuTRLGNA40phPQWbVmmgk6Bwas1jOqokjlhy6Tw8amLCrs9oDVC
5U4wsLgA+zqS7OzfPQQFqvWvUXUn9r7y9xpyf7pdsWISGqa3V/8YPvn3VsmzFxVU
LeYAkLs3oKNlUQL2Iy8iXmIDCV2tVSTKDCK/RDYUl1zPAcvHL0aVYIZMPAAQxbK6
BHzQxFtM100BuAAgM9UNZS5XygZScBi6D8X6YH2X6uYl1CWOU4NA1HF783IWmMHJ
sJfYVwucSNCxUH677a/dqZ6FPhTC8zAGZwaC0WWvHby+lcJUy6UfjLKZ33GBcADU
/7XWowEL3i3hsvIT/UsRq5wMgNe9No3W0hDJzdqTi418rIA4SO0riZxvGjx2vGMJ
X/7ll8Pl7wJAlPDIug1spPK9nUdP0FemutNAr9ivJpJp0EtgD5iq9l0WOg4QHTqJ
JlbBdrbnR2wFLbTumbGh8U0XIIJ3XqFWG3vEKk7ewDdNzdEeQtgRsj/k1+NcJyxR
EPx6x6eugMNg6qQIKqUBf0dAKiz7Cg3iQGCmaDCr8y3PV8f1yj3jRjLba8iZbhVI
SMBfQ0Zv+z0cI/gTPHptFyTvnrrW3ltjEKnWLq0hcGk56VSgngnq8t173rAnIDcW
JhxAVzKn67pfN2JcAf1X4AeoDTcqKm98qszjQR0i7G8t5jTglBU0Z0laTSfQDUDr
MVe9hZyXfNpK6dUavxFnzHzRyZr06BXBRWSmWZBzD0WGCuLC5B222tv3LUm9whz/
rP8Z2pbFJZWC15rCxsDKsdTsRo0ihydY+ZOnUGF00yU0MwBIOZrbZjTdt6gGLJVn
4sm78evSZfkeji5vKAKQNiyFEW2o9ZF6T9+VhpGL9h7sM7UFMZQ4J13LfSfah8sZ
yBGwoW6M/ba3k+f1k9kzqISVSvROpqL4UGnlxS/2KD7McDlmRAeBsxPexNjoZdNY
JLjyjQ/KmZI2TU9rhlxHUhD5SykEA5MmCuNraG/M5UlcJXUrNRwCmMylLaFg5bYd
RoDrdK5QQeRTcLQjewEgMFscoJ1uW6ZE66szZ9qEYDoCRHxg4DRausqCvL0vS8mU
algSjctzMryS5T79/CP8BOfYcowalXAZDv/w1qeYlhuCbVMGJZ4EExpSZzbWNuWC
PIr+2dcWEUVo6Jwo6C0K82vhNejA59ofzS071zpSU5CiAavGQ+a3Mhda2zUB241Z
wW63mrRIoYrXCeolAVZapoz8bTJT1E4xT95m8g/2lWA7EMmXmfBwnJHDGJnLoTly
0PK0u7BH1H6qawxGmKRsvBtOHYYwxvB4xpFI3MF+btHcQZPMZ9l6KapnhF30VGKS
KLkunRnmcgNRFyMcq3zt8J3O7Mhy6PycRVU+mLBGMX/QnuLUL5KLy3R25YoaZkb4
MIkcaW+ZKqHSGFTo8TRI+JYDe1nMExa+D9rlj+cevIJQW/bdEEryk9WoTctPsQXA
OggTkypslM/8JTJzgbq85uHFDwQcEvrLjweJvWYsmPneD+2EP4Ja+nNXVv0p2CVQ
qUUawdJTCBe/aMBbachsTeasspsjXDRfxjH9OQeqMkSvHVwUlp1iAdgAC00XWQ2d
GYjmlglkPsIJMX1KQcbcIEHOOFBgGFJwpxDyHn0y03+R9V6YB6bVZdAzHlU8sR8l
RLdq140M5C4Qao+5bdYTSf5VELeUbPquqAo7vW0NzfjASfbui5LXJcR2CdZVPFdb
yK0PjI6o6Q6oR7dII9MtuVEQndGybfcCB4iuu+UkCCRginDi8hKt5VBolIIMIaO+
SDnFdGSroUCQpbeFj+1rggfgbB44AlnAMhqFNsMQUduOhWPB9dTWn2T9FotK7onK
FiEj1B2WwEkglY6lU7IbWD/m8GjC1FNkI9yOlXor31hoVADk3rtCipxtglN0rS2z
V/ApKoHFuXpbdS3Ba+uiuadvAj7AC1eGwp2bcNGPSqCqqClcIDUsOMGbj6+MBwYR
ZS4Zp0bj8wpzKfeJ9PKGeG0taZ2d/LZGBLT+UTu3FGLsrLebUHEW1xkcyREqYkOt
Uz9IJoYi/INNKufVNzzUA7OEmPEvOCSsK4S4AixI7EQt3RRlK48BkcKXoGVn6IcQ
5im/VQbDI0c6X0I0h40sGsd4NnCMsqs7Wis7sJfVefAtAzG0UYqWVEuZXYRbodI0
iXmD3O4ELeavhcnc9oOfAMECvIZH4PK7zST3RiTGpgxcTepCZNmywr5InuJJMY9N
E4JYpBbqwcwpmpg3ijiBOuSzYuf52pQiy5zXi2JcsTM+Y75GqSTdbQ7IcW2yEon7
gaHKhl4biM2l8po/PlsWAfE6z984fWiVHipMBZ6DgPFHdZ2MSBuFCGF9OiQRR3m0
+Aefg0P1DFef0QKNi5EWXghGvI1IT4Xq0OjGFqkPN/YyxO/77FLmSPDJJw9ZyDMq
gA21sbqwM2alp2ScmDFkjXQDdNmdxPF0bl4rpQO+yNXU1ugiGQh50TGzQOehknk7
gCNgoWP8309BoIra/v9FW0TguWWylLBYo94XpbXw2BJhnSfyryANRGN9Ybc52Fub
ik3Wgr/H83uUc6CQgxfFv7YtCclKcpOCCwoZXkEUfmA9J0ou0O/cUzX8zrfZ4Z5Q
KyNjvouMeK5VIkYg8U1d4Lo+h8KxP/FBBsAEoA5XgjRa00nlWOYVHvh20MUgOKJa
dlxAtUdNLRp2ffh3vOiHNgFWdS3KDYr5Njz61tUwSurYAOTkUcY93SUWf/8aFGVJ
Qtdt0cSCn+mJPLqYpDkes3kditPWKhxQ7l/W83LHxh4Y7KrKPUUNsMkZ1F17fguh
qU1WoJMifC+04F69u1Q6A0tL1HNenMiMIgnlDFeQITEX/sya/skaHywSD80kWzmr
0nPel+LWdUfQHOJLqfRSUExAdHYKeDLFrTthQ1zJbQAyWDivQj6s2vw7noW+V4Di
V2A2yDhwPes/N0pY2ADXX1ZGHYMpC5pWd2aBnAIdDis357luhxDMpIrRf5yiROR5
jXWbpITgoOrb74QX4bF9BmXxOJiNQula9vxY7Cqs0uO/9+9QF4FXPJH8W0tRVOpT
qZbmLHjMTwOGifACQQEXLZ5YT1crwpFgNUrxxXDSNOPamdCXQxbDcp++9x6uuDd4
Qh9lsFYUwoNUIViVhSlgdwAHk8sL2GYuUsXQPssE6lzFqSsx2tdg0BelwLClRgzM
xfPAeb3uMqgWB/HCXGaRcb+0GQZheppCf1ltBVfWeHsGfSD5942wVrivoPJP7qFz
9n0ZpEdarCujNBIbJ6mseuATDvtRQ2Nu8YqEbCKdXpa2nwoTKSXGSag+LBecn3IM
YTwYlJU3LFhEmNZZ0caQSL101PShehKsOudD6Wxv+9jXE15m+r/CYbaoyWl64C2T
mXf8uCpqi6T1Dc59rexw0HnSfXVBvqoBPyutyZ98fQAV0tYA5DRQr3N0kTpoBHu8
kZtJgB/i7mw+9H4ZTHk78hyTCbebkWSLYdhHEeIu1XRLhKM+2nYBPxRXayDvahJ5
jU45JkuyhqDhSAelf+AfbKD5yR2HceWR5kCjB9V7B8r/YNv+WX7iEP36JkdZoUgd
3c4MM9CXEZSIa0Hr2iNz/gUlRsYyL7nNiEoDVidopJQ8mp70eMZVkQNpeVb/qdZL
wMIHkxOuN5ntHZZxXxWm9mwiL1jfpQpEfdXp/PPQx3Q2ROEU5oQQexjZZgeXkIn/
rDVi+C4833YZaDf3xTVOW8Q6Ewb5EusCp5hXaCJcrGjTRCQOUD4uLIzN/cB3SUD1
s9uG12lEQ+pb/Ip8/f/f4BzdkzG1/sWCxtR5MrhDfmfRwwvQN0J9XKlpSt+KzadJ
SfhTJ6dxmCb5fy+Ddv59Q3UbSPRc/Seqp/Bf5fLX+TT7yqTAWzHEsyLm/sDkJtj/
UoBcMB22PDzrrIpWt+FzlofVhDVdclTDVdvaWND+ZFiMpxwLdN3eNq2tIx5sKq17
gJoKSnZMaxkZXrbPWBFl1NotcHAFPoTnNTvVHcjlTuAJHrHhVpJIdka+OkfXP0J3
zgiIiXYiZlOJDix+h7ucdm2KhUa6/IkF8VfFZUWkAB3bFtJjtGIpWfGTGfaxpZNd
6g4AC1gQM2JgzdyyGnWr8eH5GojrIPMroR/PKPWT61Qm7B4Vrpxq0EQopTa3+c66
74ij/UC7Sp2VKQhDWIrYhHyhlSNe4rrAAaOENJbXE2hkv9Ly/Td0qAYseYdT//E9
GcOx9UyYzjCsPgxz6caajXc7CjhvCVayBER+GZJLRGf53eozYj9ay10qu9fezZ3A
um5O6vJUsaqZp6BeS5iSb6swecFrdtRfGDYW51batCRcNLuNvJTLOB4bqLNcuxXJ
WSLYllgRGrCehfZhoaWUqRb6O5jRqvv5p5s+ra1+lpV1RZJKr84gSchIUeOBDyMz
ZXvsSlPA5UjEFySDtiNZttkeLqO94hZZwi4sg8aKzC+Nq90TLJH8b/29rQUJHBru
+nqjIQibxNJSW9waF5YzD0BxaHl713QtrvUdEVlqcwcAVLSqcKmlqJ7II2uo0ryc
AonIlinA5158A41H1Fju6AXHxCVazXYlyNOArlXp8ENXdhyj7Qeg62Zh8DLRTcUh
ibea4r+XtiuthMi8iBl5EDuPPJtO0IsCgXmDnjTMjLvlNgphEa/haFpGoRviQZIr
aMRhDMwhkFqxxeeBavhObSl41V1+Sefaw2ymrUGcqg/tUod/pUg1G6VnpVbcNG0C
IFTyIgUkm85u61FKTiIs4iUy8FEmpbj/Z0R8jkEvThmkhu8vdGHODi/5+rCdE70U
eSu87l7MeY6LDGUmDZgQQo17+vQgK8Ux99LucY09T7Rcy1GA0t7CKuRFpayC+gyo
+3yiJuaUoM9crB0S9oWLUwvttTConUWtBzFQrhSd1S3C7KuO95Bo1pTR+zjV32rt
BKG9df8jhrpz5pAkNyn/WnxiLv78QVi2yKeZyWtmK/bZzZNjGlw9/45BiJKlR7Vt
UiL8QsW/3nhRTibxuAT8X41t3JlqC+SJvHNX0aee56a16Ry7iOt6iv5/x0iBNdtw
TYCD71+YVzefHXq6KowOQLDl21+Y9t0X39/O2NuwSs8GPJskB5LxaOgd3nRSxJrD
zeKYB5X8eU70u9LJc/Ny3STUHUoOlx/mtdzrHyvwgiRZyXp4o+W9hH8gTVei85+i
wje1CqljLDB0ZkVleaSprTica4GZTe6NwmTU/aqppuMLcnDeeWDOL3i8eQMU9ae4
NtCm66oZSM93GCcy0vc18OLZ0CbtS2pmsfh0YdMJMq0SwU31FuwAdoMLOywGW0Pu
44g3tCJemtyqn1beU5pPZOMCuALvvAYezqphSwe+cqXyLlDLXEEkzi4p41r3LY/N
E95YcgcOJXc0nRde/ra8KdwzzXTvefqj89A2Ck4nbI00YRahtx0XCstFbxax/Bs5
OlszuJqbGVo94nEWjKaj3oZKAZB3J8VcGFYCjvNDSA3TfNrMhCOTWS6T5gF8VVLt
mnDprgcv2GODzFSIxPJAk1McwTcfnC3D56miYw1aH/6rdVq65uLh4H6aHdEvHuka
OX+jkPb1VRZ0VPj9iESWYEtXm1SaIYxE6sz5H+2IiJmnDlW/f1C54qEahIEcaaM9
lYy5fjxAwoTBl2RAu8ZkiNGB/Pp+ySYq1ZFhZMrAAtIb1RsdHzzqyrMQ5YYWqAXu
kfpZF1TlW20oqaGQCEj+V9zNEcNF64j+tMKparV7NlFm9DCe8tdtsvLzRL7uFYFq
P5JFugulGl55OfziIwjYBdjCp+jxfI2UfxEtiNki0S4XPwJoSsbY2Afs0JArRg/C
PzX8XunLHrx1/sAlfN9S7RGd6MjPpocMklmPTgTaZBQ29m9ZMonbu937jW66gAzJ
al936JblQuwZ2NP0qGHQsRnKWdvLQQOS8uj965PN3l3mSSEFTCI727fBTgsuPRWL
HKeW4b5X//vJkhzlwrDkhCpaM6vbx/QMJtSLsI4PMc5X1ulh6fZzKQ/qZfkPgeIx
aLmJ2LKvamQu4JT8RckpWSgPegB5QksOwxx3WVzL2RLFkzUODuToFmbI6XP7WPiO
TJcApHWZgLVpOFdfsOndGY0PQLe8S1TMEAmfoCYOGX3PwwasH+EmkEjHyu55V9wW
AQQONOG/O+RC2oj7E/GIns6E0iU5vNHhYMUSR5lrHL0o1gTjAAryBmnVsboVI0BT
NF1GWooZK2a+w5ulqsZpCiycPakJx6IvA/ECcTjMRMxyUuMj5J2irAt42Z061b/F
wZXySHqEUtsSn2jZRMoGF+6yYvjsUa0LK29/ZIn1Ogw5eukUrYUFM71RCp+KnDBl
sKdYysAB//TuteBMsMoQVbemXVO9QhQEswLN0hzip4Th89J7z2afwtAxEAHm5NDk
WXmSTk5CQdxUf5qC6Pznv0i8h6hYHvtWIpXfQ2UFKWQMVA8EaJpAYrvVEMI1U0k6
X7CC7dmGeCZLPwbcvzWI2VCNevs5ekAx6u+ZhNIsV7cRDa7je3aJvWtP4wRznmb7
yqni86ATX/Ky7g+wOA2ioMGv53yMhKAt88S2ocr7ZXLABW4CSj2ZUEzQDGjAd7rP
OCGiDg86u2FLBjcv5FhHJglYRGO2kqmvH0KVFr6m4iKZgy4l0/VuxXMRGrZxdWY0
VSmwhKbk5T0DSTOyCxicMXBGCD5pxmKI0G2cc+0xlW2OevymuAlkjMjO1RWkpeop
6XXeH58TYMlWmthc+vr/CVrA7bUG5qf/8H+pHoYQ7Hl6MMWdK05JTN2KYhAPAqYj
bHqI83/V/CCsqU17XJdufmfegx/zH8P22WEeWCNl66jxmlQ5cGHXTGGKXv9pMcgQ
E66y73IGYh4OliAPGoYxyPKxB7UDHVf3UW/BFO3T1Gg8RkS8jOwBOv6WSRyQiGqT
Vg7yP49FYVP+aZypGt5YAXiYSja6+/Zt2p2A7Njr6wEisv0Ir3hUUcDnaU49hIZp
XIb2rMdM9hO8B9KsXJAHr+vEZJqjKDDOlnne/50KouHXbNNWR+qtkRuwKHkI8tCb
wl4/RKIXaRU0AhiTpWdMjgiqpRafsb5hwlk4j/4bXufiI3J4x3B7U7NKpR1AAma0
Pv1s5A0VoQo/jKbzc3HcGtDGZjoEWrhhgOhh4SQg1LDsG8989+JcTBqbODl/IGvB
dist5n1S4hzGqZfLWr8zLGVSVxR1YLgXkeDJbLcUvZGHiLNpV/ZlcDndRN0Np1vH
4pu2rYMwW0sZh2P/2KYhKqUmgg2q1sYpX2pIV85JeLJU31Qx+ffatLBV1rT5QGf6
ugkDzyYxBFP2LFxILhzL2xrkIgcglsrd81TeZrFIWGPGWy14k+33zdIrfLHeoA42
kuH6ltJP1vRUChsqvhcNfjkyA9looh5cOEfiw778P47Wo2h1bCHCgdUbdd71OrkE
271v2RlpIwCzsU5hp3li84pUtK2fKviRDB+G+qGZKOTumclNjWeCfr8oECSYqaj2
Owm7l/qDTdBjfASGxLitOFb5nmCJnLYmjoWQVCXEw+b1IOCi97bef7+vEaaJP/gL
61EnYCzOkooB2tYQfHHqWH+Cn1lgiWpc0WO/3DCoyz/cY+2mFCsj7O3dNgIyZXnn
dTNDhY2SSdRLtGd6dfXGtDbBGmUEBop3WNHzq2jZOksb87lFabYpBtA0aAszhNHa
Tf8aHye0CFjXKEm81wj3lFH9RtIKn/X6if7gLXrdrjMhDu98/S68FkiCXzilQnbV
tvNmMxOf2qDoV/YOAieJD2zbsWjiH5ZU8VZ3trel6/LSAlBtscWpwjD9RvvS5uF8
GsXzCHAgGHWMBN2WI6jL/DBKiygZqfkZjt2Gb2VwmWuc3jo9WixQRC7Yy9FCSc8T
j7fI+6X39W7bwOHQPGUn8Y+zxmme7tPWG5QLZe69bFCYCYgbAC1jMM5VXtEfjQIh
kWuPxfrV8JeHdYeM75aL793t4eGXzjY6xG5xZIS0Dfelw0Pp7t40vmO4mYNK5t6/
Bnr7HM3u14neQPoA+tsFAnBwkh8OfwqSak4lof4Olz39H6sVFcEz5Uvs++h/gb6I
XOa1Klj5hk7Ds1CoVwY6Xlb37xqjVxZK1xx4ZIeW3Zs+oWM9Y443TpiXm/Df22GD
ts+YDrK2j3d+BH9+b3EfaQQd0Ln3ftlczQ+YGt+/XUzYCP5ccTxx0QUKyKi5bqgf
V/1DDcB1t4ve/9OR7tdgVmuB2hYjwPMaYelKnrkSEq/cLolqMHhWUS3AUyvlSa9R
jCIPNlotyfesRIjXQZ60u1lBqHWmF9jsyegS+XqVVxmTwwSxnp9WT4Ta/q2cpnck
XRXcUUAkVozyry5sJColf93Ttt6Xu3PHsx3kSMhIl9zmhqNllgZ02yphF8E6sZYE
7zWzKsb71wt1zljA0Pzknxw5pJ6A7T4a9yCyE3cNHry5eU+okNFE75aF8JbNZJvF
WzNQcNQI7GQp//vrKfpa0GFpl2I5pZR8KAVe7ebf0cBwmcFu34SSAJ+K0SgoH/Rd
jEI+OFnmTRQSrJADgZe/Y2F8uLdBeE4hsIpXrGscB6i/aoI9+r5Duw3KpSybWWeF
41ocnHejB2loGT4G6OyxDVtpE9HwnsO2ZGifTuyL99Rpt9UUkIcGnPAugBFB8s17
ASD9+huSlPEZVBO/LhhVcZ1DD7tfNcdSirhtl1+ubdMG1BIbNd1lH0qOo3WITmYR
OqNq3VredGIV7sbKdn1hMWbfvVImbUl12q1g4Ku9kpBj3YbRb3s11zpDIv4Cwet5
IxCt3ftGt0Jsfsqa7FGhteHXMWaWL708IEx/0EQ9hrocymeu+P8nMGk1jNuJbR+H
97XgG4pHB1FOHL1X/jm0NkwFW8o+0fsxNReeFF1xRVTl+Pq/WEpz/GenI73DmDlZ
zfG9JoQ3mwLsHZxVCMqvy57QwgG37t0mp/1pbgWNYbk2BEdCBKf61EGJ3n1cCFyG
sGIWabm8o2T/Y/GgITSgBZLmQZtQHkGFQ0G4CG9r0WELG00NQtNiigsKijRdJ0UT
jCWWj95IYOj19Y0z7o/qvFBYJkWMiL7BrHsy5merRl5PY2EW9SxGk8OOt1YvW7b/
xAoobyQKidCd8kKaaqRdnj1yTlVc06+R2lnquggoBZRAUxLlbE/M8lB33nnPepkA
YbWTUv0wJlAZYdSkiCy8z+zSP9W7ddEnB7kzHiheSYMwIaVw8a4P67KCx/qw0Q0q
4CnUubRsJr+ek9YZ0av8F2bJYs26FkDHnGRQRbtsYL7h/cW/m/omqwSecFpfiPS/
tJGTty/2vu+mp6305JolTiw5+vzJ4Vi3maWs6oWcYqcBIMsR/WJ/p0S55Higt3wE
8MDY6WAPg6YaIVDz951vwsKG29XDWvWC0cgqmdXdizxezj7+68/A898plHre6GF/
LvTKyT4EM74oIiN/sp09obdr2VvkfztAbPb1JXH5FEtDEGCTmpYTJNAHQaoOEqU+
6sVWJs4XHiuKOeg2RMtIJpxLtgviJ20HNlBDXJ45hfgGOUVPQXV1KOrc8z0KpB7n
qB68gQbONAnkaXROwbJ7EGlwpP14SXtTe2dbV8u+nngxbse83Hn398mm667kS7qN
dxDZPQCcIiFCNozTfKZ8hRPDuHT+peJ67DkTzgOb0A6nsLnN7E6JnebD8CRcCrCk
pycglLPbDUBLjcaOZGwhUMO9oNrxI+4QV3NHaxdbFUOKWVE/ENceEJff4W/RrTGt
C4tz07z5rYQIc+NMcIYZ6mLyFfU98XVmFNl5SuGOKgansQVjz0/JCbciwB9mh+vs
8LV1GcjDeeY3d40TaEwUwtVIyLSSVq9/v33MKa/DRkEJaFVPHQywXMi9Bx0InGwI
VKA6w+tgWEks6EgL/UWcGavtCl18JeaPkXP9tGu9hMKVAL3TRvj5jsClSvoe4duy
0jbQ32bNjlUd4CHoHT7DD4TVtMQ0Af4FEMOdDQdbxK2tzqg8c3XQZ2my3GBuCrDv
MZcdbNhhBJ9UiZKDFRNcaqbSxAFSk+W/0Js5b/jEvEhArSq6Xx3LjvcTt6iyccX/
ERcuLtqoN5UUtuq++oa4fkNxpc4WGCeYnLSXrb09z9QT2QXX8nU8jmlj1B7RA52x
uQikEb6m86VotDjZOjwP4Nz4rIKq38fB2DP+sk24L5FTbvPvTdKRLrPFdZ6OJtfo
zgm3tke/+29UQyXQk3rnvgi+QPX4Jn8nJ3K/7S9rrGYSyQiKkLk2OZZpjSFY9F33
a0GQjf/Mm3yxeFYxqDuXE/o+Rc/4l8EzZDu69xVytF24b31E9ShLF7FH5n082kUT
qdOWiAkyDyicDKmZHwMl0Q+xsxzuewB5XPpikbXhLqd6CEOEyMTAhf/Foc0XJ5TN
cF5WslzPQpeKJrialxylhOHmJiyt8YPbOoQrLKWr2gW9enTc3oT/Sl7GvILN20Kz
1almAqqjGENXgQhNq6F/ppwUwb09jebQj65ap8kEAMwTueUsy0agHdhbbcX/OA+l
f9MXHSVxPBFBMalKGktLkBrHnn4g5EoqJFOpap0uHtUMGwZ/XSBoGFoFXRDZmao2
QzDNDBRSm3/I6nfpFQwFMs4lMoetMkHPVtHqRpMAbrZZZTxfN7luBwY+I/8fDwoe
9A2rxjrR9uZlF0urzPsDUbcehh4WIt64H7zKbcYhk2GlBqwQ/TTXkWd3u1ld3RLM
lrYZY3gp7EnYTaYt3CsFxuuUdQU/6o03dqH33Oy4jFRR9dnczkOtUIK8VsKmiDa0
LogKRjyM1sp4cSHP6m6QT/7KXPmp0LONlXTZ5rjGFU87euusW8fLpcjvWBCqZdMM
qQ8Ms7dzJCQP3nvr6MDUCnCCSNAW0puOFRKQazzWfy/50nkDhUvDCHeoDMTwsb+P
HkkYv4lYT/PHchG1ubhszj7VoSDo/wP9lSThwB5Iv/u/V4Opg4tOEcTNO4ie8b02
yADSHRlz6BYsUahP2WxQzw6PE+S6Z2PuaSeKLya2dCDrlnVs86HH95L7vQdM1Q4F
39IDYGnU+XePvHaAaoKCuJfTZlQZpWhEPbmIV6R/ntKMW8GRZnb9GNQ2YvQ+Ng9m
Dhed9B6NjS4nSRigVUlXsBB+DEvnYAkGRhyyiXs8MMjjOc/PVNflnfu+ymKzOn55
TijO9DOPYNFndHP2GgxvTA0GxGIZdG0SW0wk1aEhS9FckHBDEmRpchFEt6xRGnYe
jusYG2jAwsEbd4dlnpeJnu8NUWuM0nuvdxb2TxW+k2aT/lYBus3vw4BSNp5ydvwb
xIDnF0MjXUMBCgLnv7U8R3IWkt0Fq5XnhgSdZEHdpOlzc57uoDb4rO3g3UKhyito
nj/0+c0WOE2bIwiTkdUAlm4rkrY0Cg0CNhdkZwp61NTSfUDcLhb8VeT1ljgUdAQA
g7EpLYbTbCSNeK3XnbJQyHPGNbX8IXq3LMeJ2LUPsY0y+82NRjw7p+VPrsgkwOLc
9CjzrBdBNqPUMKny+jL0umVKGpXGdFS3NuBCo8I32RmhEoxd6FXyueMSAkz/Gd9q
Ys1ymyLRilDE9SInkxdAXnC6jVA4Ss21jm157up1FzvTQg3oh1uCFajji69I7mUW
H2So0tCM8Jd8/ZwcBBMD5Ap+ndCTRFWoyZkq7TvKr1/67nCC73omgOtw8/Ij1Guc
Rh3f52anxBe1niYgFTQPBOLwVkps5CG7AjyyKjwETgUixEmt69Pv/Gt3twwyNA/W
D7k5aciACnq45AN/undMn0LZbjdzE0xQw1z5xRL+4L1JGtURO8WplwaiuakCAytd
QoUUsJBE47Mpt/R/zuXc19LwXB4TvICMqdbWlvQ9HBu2XnOxC8YYV6v5ftxZDgRY
LkmM9wHP55xgJ66hPAUFmiZogelSiH/5rGIB10r4SdzEEVhGKuryCMD5pokiXWyq
YzDz7F2fbbgDPI62XBGYyjqon0OpbpTfvwhichwls+ONGsKK2W7eoxwDfR0WjOV+
8iMrZFNvvS2fkrgP8nvE9PpC2KGJaEiruuzhsMSDXJfNiOtnOdFJPjhNFXCWw+VS
9jp+7hLuignngZXV1CSIS+UQCK8UowObKa7A3kdBQ1QKaCL3/TR4T+BxBSNtz4Xq
eQKqitq9SqUB7ITXZyDJ0UTiVpxX5o1IlgwAUYoCUgKT6PUqMCp76K/tZ/ZsKqUa
42QIsyJ4ZppWxvsO54NFyZFhPQ+CrAMOPMDQqAaEcztYEVj6zVTGdiod/9u5W4U9
/6pflcyFHZAyXsDkRY1NVQAjpnUw5C+hCvhQe0ihE3rSL7q0jdbPXOz4tP3hcY5p
/jUBxWXFGK0oXq08qCyaebz3dw5bjKcXcIdF63LybHY8o/zUmP5T/qCYU3v30f3Z
6mrCGzVta8Tl6XNVdvZMcl5dqaegedSnPw/sPZ1zxhwbuwTjx4hVb8bZQZTNG3OW
pERaeadmA0SX8jgVLtoFB0eMs5bExvDtan96Nvw42EfZzyu0bJN2psdJjJdlCguV
QkY/pAy1GJDgHhBJH746PrWBN725R8YCJZ+CPkBZswuHm59/NvItP9CWailqOYo9
e8nhZRNQM1eym0T0srb0zeipaR9ol26+Iwq0ipSmVdQNLpHBxu60QSxY7eXZll4f
BkA7BEOPXomm77oGVZdunLTQF0NTuYt1lLaC7VO1hING1mFkzH4v8UjBixiyb/3n
NqLwevTSgeqnAIF/BlSW6TOnIH9ZWsmYYCmSU25Hhf+RpGjQX84nqQg3s1Wh/dgQ
v1YQKVfQhBR7GI8+c1DvMCcjx2eka6HoBkczZlSw4jbtSmK9uyTcluq/9WqPomuM
RJag/69k+YM8Unv35itW0pOzjTCXLz8boRqe7ZLbNUdLNGlkkTDPhyp95ugx9Is0
R//atbhAx6R1gd4UT73fdGxu3GwSH4d1Nw4twZilHT1K9CqWn6TYVj8HSKWrX2BH
VA4DACshglPWbamZLBY3hQu3fluHRlTjShsAMGgq2n2l+POFJKFCxZSV+i1HBeXr
7IWHiunugG+0Le1U9iOVUH4tcDoPFFLu7pncN4jCzigpw9rgP/a8xNjY4B6ArIfA
wdm6QGRE9GkPS736lzEXMRbHybdV8i9DpubSc+ouS5EX2qYeI10iG7a1bMcVCfKm
UxmmFYtriHxiIcVf6KN2pnJTy+tOxJUJzVig8p4iyc50gub4oQ4iekw12ASNm6eg
b6bfF2Ah4JQIU7w6U89sMqBlDdWcSmejDgA2LioOg+zQ+1fZPq+6LhTWV0u+1wFE
TCpR34w8SKPhNYphWnWGwjS4bU+NZZR1xwvZ4+9Mo0OFo3GGneEPZJR4VBxQQZKe
NEcbQPPq+LqKjO2d3TywdzkPLDadLdBDXPjKkSpDyO1G5wSUjt2JMRVkFJdcpO7A
mbje1/zqgHxfIwSKIWjhzl12krcGJDgdjG3GLJZOxl0yUMnihZ39cxG5GdvKpaQc
twnFl6VtdOJTJV7eNqskntletQFKjGPrHIFnx9vyVLKB+Czr1WiUxcJbhk+7e9sf
FemAvRmLpG67/5YuYc7OtHWe0vAoTLe/Do7Dco75aakarVqyRU1D07bkVsjIEWvc
doX8vFp7C6FgTL/GYYiF2hRTsIQjx+Du4foTjKr5RkYH6A39fFkyEpvcJhC9rT1U
tSTm2xU09HqvGk4G4jzxN4l+Z1zn8qFhaYBtwu8eWY7fmFro/deO/kjkamx6wnn+
82+r3Hq+k5cgiDZTAAEfBkHWpPD+0FpJI5KHdJQf/FfElvs9HugzzGl8XUOrR99D
SnPT6diOerN8DSI6I79MEaC1d2lUTqvep8fz24oEPxmCpqoYWzEekmF6eKnTnyui
Adb1WBHGFrfFEVQxRwlSUYSbYhL6SDh72WAxfU0EDV8UnfQ9UcVuGDXvADdUmQ7S
bP1miyTSyYDdyWPvzvl5FDTyN+XTPWWyyeiqFxPVH43yhHpki3vEaRfuFwnRsJaJ
2J/jM7LDVV/Z8+b4aLHYgSv2UuSn2Uozw9rYLW7BJUKXaejuiHYqcBRKTAqqQyJA
iLiyxOBFxeafg2336ENsOD73FVq7ovV7N3jp3UrAyvmtE4xx8DRdPg3CoidpsJ1d
YMyFnfNyR97+2EjSzQt2u37vXe1R4iUOnoe8vfQMUh4j1mh4r9sC/tTX5jFMn0BM
ywaKvwEyPdL0Ayh68bSLL1xFogLaXpxYr06ssXJnuuCyDIpKJcmZFOYoA/EXqIoO
BpgzcZpnsFSadEf/ApjSv8A//E82lbk1IdZ2d+x9P1CoXxY0vuf1y0fNaoW8ccJ/
aQwEJznR7zYyqZdY+B+9GLYzXSW4NoIcPgem7nBaF/XeAwLmVggQY661GL6uhb85
nLSt9f+cbVGNNQaOzLu5AKPtt9jY/EBXTZAurqcBrYAx2iuD9obF+q+uNSqvlk0j
93OUsMqjiAWPjhpvzCANvbPsD8moIZPYCsVXrvkNxpA=
`protect END_PROTECTED