-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
KU2fQ3ODgksteiUU42NdzgSJ6FoWmhs6RTeK9MgvIrd38p8GoecTKhCyk6KVyR0O
Cc9iCTFAJxEP68B7KIzFBb8xHhnKaY1RVoBzU9PyzDe1TVv0PdDde4nBP0W1VTL2
BVwftlHaKKIsQd6yeIUmJgX4s8lU2EmS8j6ZMhOE28PNbA3/E7PWEg==
--pragma protect end_key_block
--pragma protect digest_block
nhfoOnyR/1OEIWFSaptfJuLwn4s=
--pragma protect end_digest_block
--pragma protect data_block
xV5bbFc4PA59GLKK59ckOZldREOkyTJoV8xdhIVmc4+wuNkYH5eTQ88MhN6zPFjI
1qZKmnLvtZTUyTKwh1vzfHQ1SEhQaNgOJfrsjmZCZ+kPspngdN6y5sIgYRg6jCYp
BJJ0UXgGqVps9cMrtkgBMsPtlLgstyJ8wVzR3at0rMIJTlp1JBLgbJAuhpZ2neSZ
IZJzX4XJsX3Hgv+eYMRhNkH7GGJWePHIEobYnOC0vgwIuvOrluRHRN7u2zcgufYC
vGZtldyS/d9gJWPhy81/Yh1m+yJgooYMvrK0kWQgh1JakVqTRr9BSIcB47+FGQ/q
/o1vPCsy5EwZWr+Nus9npnQYriKIKCpvQY1DjL0X/i8sPzvn45vzWLC4VQC2GLPt
FSrNybInUbcBdnr1+uFv5csMUJEjLAHUyOGO9932Uivix0mb7A7L4IQ4qJVeyYmT
+t0H3npVliZtP7Jlq0rMW/s3oSZkYxRuRVr2xmUVqbyqJMkAuOlVmSoIM8Lh1UUC
YFncKe+2azzc4MG8Yr+3OmJu5ozohvEMboFCsDDWgvj6BUwwy9M04EsxpAmYOiKG
f9pfS0kBt6pfewHafkSkZGgehTXxUDzFj+tRzFfZsMvwPwAeJelNwSSTh5eSs1J7
AGw/xxzwmMLFydCvAu1NTtDxTVDznAV3YK5NFml7PaU2gOfpclIZUHwMxE6FIp9C
QharHwFPXFOiFlDqqLhyoidNxVqtG4bEuUlNRsF1GWBsHfhCRdfa800jvz7Ejqog
U+5Kgt+BZACACTUL/fAksna+9rJj1PluYAUrUvtpP2tNhFMJithKIiwx91KLUCas
SBS+v6tsxyAQPnWfEl1LijTo3rE/gpLaXNHJSC7eZVsmUY3XSSx8BFGCj4UdYfnT
mCjNkDvj8lMinlpZgYbu7Dkpaa7pvs/IPJuFfNeD849gzD+NnR3OyuKFCkq8iYg0
mvZd1/GPayWC9+xj5NkPm86GzUAimHBYwh3fWvcHm/0LmZBPnfaR85K082JN/SwK
5YxXsTK6fmFH7G4B3wz4kUzwdo3mb2fizb7/aKXYS4uiPyHxxBVlcUMa+rUBfv6W
/kd4sgrKQr30mPbTfzbtToBMIqlopBBMn+wMW32WejPROp/iw6p5ZBb1CY1IbSO5
ByoY2dbe3ECNstRW8SwgtIQfnrA8qOaTYaKF/4aoqqQPG2Qw6sXxtUnWIPLIodoU
CmekeOJ1SKygYzPrFHjUMIQiV9qrvW9jt4bQ4vNqYYGHm6XdsTCW8i0z3PBx0DAy
vAxK1W+7jNFbLG7GrV3K1okiZBuK1td7Y6sXriaOOaeUV6Wd5XhGAN6aM26CSjug
MYSqYzi8yIlCaT02NDtFFbvHYM/vTJpFAFrG8/WK1FS0ZSR8njh58cyGCep3hSep
rCAjerw8zSISDoIQ8224S9gA8afEsDoeozavbEo/1uYuh7NWFuNv4vqDwV7/PXES
wqIHwo/zs/7TWB9+Ags3t83x4MV6EPAMf8ETAMm4MUkmbpU611jIZ88EcBSGJTRI
rP5ldJ85LA8PknbzoSYoO0/0wUbbYX/HbaS+2soc5Iin68eUSndLMHw/cspqAyVQ
rE2rdejEveYMUe1J0ccfNqPEKEzWS7nu3nRflo3dh+2xC8qFEOyZjr5R4dp8EwYH
nC8eGtI3tY+c7Tlg55crsH/lpPK8UyUsf/ukV0uzx3hLFWDMOn90AY+WYSrFplmX
n+fMCkGbOJOJJFLOVkBMxFPec3jqEmaoEukuPPgJ3JOrqXOQRjGGHF/niq2AG9yg
CsMqdop6OItayT0y2uzV58rj5LKlEhrrkgKo9qO81SlCcXvbZ8F+Jml9skK7U77F
I+WP3BcswoR8O/9F3FS+jikYPzumTe0ly32oW9bvuVKUqNWwZDgSfmrOcVsvjrWn
ZJ1U+Ut6F6/b8LnqN2Wp/1zPqCUHMkWI1U2/R4muFyPNUDZS38cOZEJWJKMJlwU6
acezvGG4ObXMdkKZTRiD8kUnSmUn+Zu5NwLkkZ4tw2X55+u3pRultPbQJMMf3yvH
S/jdVWjvxnIZqnSY2GVSDA/L09G+bPcS15rz144ZHadr6Lc7jw3KskW2GIoekq7F
RTkXrp4cg1kY54qBlGGWMoFjEE97LEJwpLanBfhZacJH1aT2TrnRICYN1XuSy0eb
M5kML3K3N96P07pfiQj2pm0Tua9WSRZ+4NSYD58pIHpbex4RO/QPqdOA2wfn6FR3
pKDSEdvy4AhumUyusj3wMtrnxt2RrYxUkPp7+7gxaacOD/c5wfsEi+R8p188SK8N
aGr2C2p/sfnQgCFLee8S+XEKFEPjjCBmBucMez4Ft8Uk1Z1D1OUotFzP9Sd+pIYl
OdVeKIQOWoIe00GvC0k7QLAeIhM7RK1i+hr2X13hqjr8xTwtA4Kn5Fcb4w9E01gF
OvgwWcbs5mNhq32+yiYz9I11J4n9fUw3Pm60sgoZLi/XSsQ+sQGOoOZy6lmjg4MK
HMB2g8GtMH3B5lsg87TM8rvs6XXp3tq53QZYbCHJhictRtkbbl+zNEUK+yxkwez9
xV2OQYaC/fEF7Hv7bOFDlt+GnzI1kgS2fjnn7wLXetTcKAISGyliJb4/pOYgtlMf
t9Fc5+tMUyKzBfz7zmngfa4S6rEucdaCfyl5d9s078iJ9VMfusaveVbk23anlntI
cTSJW6PGbZYw/8w3tkpQy1JaP2pOiCWtkkZK0r5Sy0y0YMRrvTajC0uyl5Mqos8t
Q+lllu0xV1riSl99sd4IbB2YyFnE2KclA+3r3JiIDZSRQCmDet6ZtaDMoojZyFX1
j+c0x1HH1jsqA4CLPbxX4HlYC1qCsiNLZL4EmkyY9MXmFPNj+aXp2P9NGYuDRPme
k7fwgYnpRCrXYRamuPTqo02g9BZKtizdcXivFR7o0wbR8//F1satr9ybwuCUcC0R
TRotSYNeVmNjObgVY+PibmcyMhGI6O3m/8D0SI0Etv4fLnkRZNQJi/pZRqgYMv0H
8wx/6t1dbaUqCsKc9miannYMYl6KCxDsATUgXjqRuQWW9iy+shpa3/eeeBX7Gx+9
UueYj/yhRCYAYitkxslb7DEgErp36g0vH5MkT/IXDRqVBvnT9ESyuZpcUQje4ItK
xh8xPWS4UuyT9TxUHJ5prYWezVHG/WCrSlZOlNfdr8Cdnu0NLIRF43ORhk0sqFlh
Z6gWC/Vpd1bcmhuyNNavZnQazidUYTLZnbme1MTropFk/nsNk7YQ8+ntwGgVOC7h
6HW55VEiKmRQY2IUATCjVMsIh152xaA7vHoYg5tJC8aGyMnkhP36F9nbO6A+pMpB
QGzgne6v2G9JB6xI2FNAfm5yQUXPc62aHDuW4JM7uRwPmDUbt+uRl9bSEfvXri48
W35Cg3fN2omEg+SX5P20PwK6LGXaIsp6rFSBe6MoWN+11oPyoTleC6GOqj0HQC55
GFJFn5cV4sQr2Brlt6PPeJrtWf2GW9qfECi7HSMOuCsQ2gOQiqE/ArPVTRBwRDSf
mn4N2xWg/qIRfLAj02e+DZqrCC/LcFEKcjkZfAWyfK9WgPhTrhO1jBxQ4Eq1NJq8
6V2jpyjDtVPEj8ZnN20bMNBUdfdVHVQhDqcYfPeK3kYKtpVP9TO0b7U0mWxEPh5h
PylYp1bvtqmL6GNEagajsb1uZ8G99l8C9YRzP6qZmz9avggVr6JHOUO29THr2Ksr
owxVyliWPTL7Vj6g1KpoMenIwtfQ81RW+TprtwEmwPpNN+pToRUQEnqeOq88Z8ms
jyUAlIvpdl9sLUX1++DFsz4ugkGBDOLG7LAiJ3bu5BTPBioDSewFX+hSiVSpAGqx
J8a4vhKFMEmum28c/W5hj4TzHcPtFi7ddEAXoj77WPzPyO+ruGNe5OsMIc6ZyW3s
pPhY7c332dYZSH7MhzZU3ndGLVBr4sb7sz9Nd5G78OVMbr3fZkbMhMsW0E8oMIkg
wt/sAuSWxXkZgEUS7HbK40mDXseKDUTFhVZF6vEPMDBEIdogePxnA91h30asG+9I
OGQXnfwG7OarF1/eaSkDfaSxK3OO/lmZkGI/M+K6picGVoOUxK8VNBjxegEr0dyB
1pbqVrdEuHlp3c/9C6PCi/AdU3QzXHnjdY0P1SmoQdt/9iEEb4+H6rfOArYuFwtD
NPuKUbjlFmTbHhHl8HDMxaD39VkwRHXrOlKlsfPwsEadlxfRcfznmFl1J9j/DdkE
pdLezlbjDQrKEEyjzBEmH5gBHfbjz5kJ0wg2Wed3HiT2uuGUaSLeQmUA4TrFrowC
sr6taicOxI+yFCsJ0CnL9bF0zvrL9GEDY/sjE164z5ETYb3l6qoz1Fbif0nCTN+e
XwlAlvi0MhXn4Gy8EnR/QFH63J7L3mD/SCXBmzVfx9Iy/CUd8QrCJCQhPrczwVra
+5t/itGAdPOeMkWyfts6xCzqfiPBVVGIW4Us+vvJs5pgdb+M/7w/F+j0e0w/dTnT
KVmJpfqWh22bsHJpCPD+YHrE83nOoq2l9N4pqLv8cU3oLiEMRDM++qb9BCTaOcAN
wm9rGPyrCZsl/+BQhTYscrXNCNv3R9d1qxwAqY2tNrDdC0HBrjBnTKopfcvpVJQn
raZfrO5XVo8kFsibRj2QuEvYnBA2JdanON5tmohzy+uzt6RfOE/A3/aNsiwvuO+d
9PcNhJRRY4sAIJSnkHoYZssF2mZX8st3ClIVEh+gIGXSOrQx8WyuEsK+Rl/zm+fy
0jvL/IiSXgXNpLOzLpuDO5j2W7gcTtt7yqr0WcG1E6k1sgyEhbvrjfJJH1Ntj7p9
UXi44laGjdS6tfkBM8rcC71Ao7VobgCVNHQFJAQbhktiLnEiBxHHNgBNkQwiOqEn
yPzRVTD0G9eq3IgFq9pNnQXv0hd4FddKyInAu07jnGk57jtozFNyrdt9RiJBt9is
pI2eVPx6Y4RJ+UsUa1snCL8HqWXpzGqKTpHgmSxsokVed2zy+z9E09bdRrSY9uqh
Fx5wmXfT8zYGJVZLLx/uObK09UsjZMuqeMRIigTwhV2+bqNHHVD8BUPw/ZHmcWoD
fzxjl2MaTwNndzyGCTeXukfTCtrzJ3xNGEDMMMY2v7z87H3jGm05SMC+UTLtis60
zhHjYFdlhXhMWfgAW13BrMMPye11hCYczgHyOncNtCeIMib+c+nKIRuMP5rz2lUA
tzYesbx09UgihffqWKb6LMBHCGYqYmKlxIHoIEMpbYIRf80/uz7guDIzIhZPHXND
CZ/kXB1Sd9qgAdzzw/0t/h0Tnry09+fvNAWoaLvl/7XCWZrbil2aH6ysKrSkxSJs
rp+URiJoyKMo9be/n+3/lGoGrgPwrTQG4/wggYn3fiI1MQc26R0GIeNcwk6moEI9
WyPskMsTBrYKH7wG1/185HjoHQzOmmo9ydX18irj9EXZFZYuDpu5nxoTVjmNDWLv
QqeKhuJwupMdcOt782g7kgM4lSc9ySHkh1ZrBdfe2fyRlGgtOT+9xWbhBJ5jPAKP
4Z2xZB+NDJ4ZJrb4hQgE6tzMQTs1uCfwxPARUp/9llHvGDNJk3fEhQ8ojF84hS8U
277YGvwtwbfT1YrFnH4qAx8v+3ryWNMfsUMeJW4KNizO9qqhcD72Ob7cp9LkP443
k49TjdhaDhRVAZizZ1bKDcJ8xNZ26lgVdzBOZydoKrwuu6q/S04WnNnGjhB94KlW
8kJtunhIUOb6b7NjpPTrSEp0AQUNXpLyuzqqAkU5yRrPgnNIoYusd74RCkdTM8PC
ggxOxPfC5Konpb7BFdcquefapglM44nqPnS+PP74t7sdyqeS48hFNAuBjbTXGJBt
bI57611R9hw6BP/fkKN3PulDzLaUpbcD6RW/N1Qf/uWLilK1x830O4pdNZB7LalF
S8C9c3FeyN1aC2TypwWt5LWxMVKKmusi6r33gORBAUjm+yfx9P0EuFN5/59QwJom
kPLwnKtJDoTsIvAHBBjls204/sVZvkR8fNHXT/1aOyPLRqn9hJL8JpIim1wOK7Xq
wFIJVfayNtwPNObSXahYDoX7xe4RUhhb44YRixUgwSK6AGs0tgLtWJNiXUkY03oL
7bIVkoHHRdXyhvalQ45hTTBIybv//Oy6Q7LT0z7TW6MN2T6wis6Nr4R5MSaOHCkW
m74KMFckgxdXZHj85r1iah3lU5s+ZVX2ejv2sfsjaO8ep9k5h2un4M8z6oHbda32
han8QSXy05C+M71Umlv1aygIir5h+480zn+Fb/jnBrNH62lBCJn5K/K8uvda6lLU
FtT64Z+vPIQGGqSB6aKsm5fuNiMjBr+CeAZ61uBYmGpGc6KNVtTJraRZW0LsOpkn
cf36c7i3SHjK17ob0k/kZcl1t8YW73/PvrdElJcN4jPB7QYLGCjXLNas1GoPT5mO
uuqcFYfmibx321GGol2lbIZnwzqmG5tFpmoFEUW1pZAhqnql4L2D6D9nFIe7TlY8
oDFEfYET28zNe21ZixXGvYvywNSXy4IuUJ+e9RBkzUsjjvGl1/7GlCWcS7yiPDgH
F5xo1tSKx16iSnNh5B2ITvOLMY655oCaC4p8EFFjnXJsUvO0Gd6WO9eh4KtmYlUT
HIwABiWRlWFAjXmf1nZ7LKAgO05DLEmEowxQHKMAghjCASRjonKXndII0LICNU81
DQAZ5oh7TnJ9lJ6Q/RhD4ojwvmruEwkGvS7NLAK3cKzs5qplh3BByMM61LXegfl2
JqUY8tLiFxYeHa87vi/G6kRwf4BJHA1vC/5olHaXQeHQQrxukVcP44em4T386QJ9
byGTaqh1fyEJ4Cwardf83hmd4pjPKbbeNQQxbjG8wb57NwjotE1bL8SrbWOUWmCG
/8IwWi+lMwGLBhDmtRlAUWxAhHleqVeeN1rlqhZIcco2d+N6CPLjZcwwOVOPdvqC
42y5ulKLOAPQr40wh4R0973ofo2XJCHfAlqEIDBdixZHvp0Aj/YfeE12oQqlGIag
pYtuAP8FjFdggqyaiv8p1jT4JhnKCoNwCwjq8xDAnCLmrklsJzoxZrD+lAkxwpgJ
4YGdbeYaOJT4cDCeCwPo8okjxOgz5PZvnlmPed3LQPQ8ti+xDerNVUdavV5PKTRR
/kXtLLZ/8T/MqHyJFa5zXBstscQHwisAY0HeK5eHVIlzAeCcqfz20EkpUSuQEQdQ
fbAhbWTzwhDTZF7Uor8vwVd7kpqrPHNmt/pBrg2440EkRaTgXh1o8wUwB/Rt9KP7
lfVldwm2FGvlfMHZyptZaaszReRUSuVLhA89TNmZaaFl6ggIo19q2x0Ml4VianxT
alr2ihH3f7Aa80LFZazeJ7GZiPFqiZXFwWaqpYsiP49k7q2tDAjqH4JcHAn0AGGM
pVkxJze4xnTnGNvyWrm/KM5d8dc/SQkvlshJhksKIlzB5D8fd+2qPBDRq6LfGOlE
4hdISGPx/YH4kkicXagQwyW+7feVmJmtTWAsPdp/GmzjuU8fOZL6W0mZYE/795Vs
aYDRBF4pAGDgpY1aPYj/QuXlGyE0+ccrYbujBpPonncvGsnxk1NwZ9Y4FHtRnvT9
/nhuSyjJXLGRq5VXhI/juUvtfGpvCySj1mSbQcnq5bbxOHWbIGYUSVNAXtKF0ntS
9y0f6GlXaOJbE+z0qXaieh8VcWfWlCjUbW7nzrevbkRWCoZHh8vy4R4Eb/HpfP+Z
8jsfNM1bV0R30cvdXEvYL5CJDogDg8pfSnYHCE6pewM9ViJCKD2bbGyTGBdYBtmt
R36O6z7GVot+Vv5QL4RsibYkjzcJRK/qr595qV7sD+uXzCAPAS5U/k7e/6vvGkXP
kLyfpgwbYQtOZqR/8Fcvrszc+UO9mv4SPucYclDy0mj/dGD3OGedzpeMzZsZ5qEe
WKrdGxG2e7QwISiKmCO4xLKNlA49SE72I/hLv6Il864ASsKnTaEBGlE4f8lEvY+u
/iy4YFAC5D5UI0aU5+5u+GGY4lCJ71RAPJ9RPr01jmiJ09tQCHRRqAqPhZ1RZs42
Q8GCsd/JLEs01emJMxv2H0UNTSCjYPd0J2kkZ3aX+9zaCLEPM/qDd1CfcjEGbiPi
ELt4O/u60cMwRDiPaaSFvkoC/Fl9LeHiGENw9CSqntSqy3Q8ogYhosGeepLlNrJb
KtLq8F3PYkcKsdUllIdzOuIGSuRPR0Dqe6h2Gwmk+stY3nXGdj/U0BosJcV1I1pA
IfMjh08Itq9LjIgGQ/fdBlAyt4VAVcXeLePkZE9fwBRkZicWemTM92xkoxlNPWrP
yl0z4gmfOLuxOj2Ns8wRophX7UtiRcG0LAZ5nSnmDTSGXaoOVGp9vYH9/HJyc6+/
ZF9ke27/qhzJQBbOXBd0QBEp9THwT2rXi31ZMY1nRHDhXbjqbDPSFvtaNock8TmN
ba2eNOw2B5W5vd7UpTZhW9D2qJYEUj5kDzfAtF2UX4xuuNVCiPsEH8AH6QxlSKiG
T/WchGqfGDUXgZlKCo4U6VXKrOvUA3tvM2YX621L/Jk/T7xVws2cFvshoYBs+kas
GWCu/5c3siqychJgKzppuaaBy+2+HOfxwy3EmsDqdqIsIlUAJj4BhsQ2BhYxf+Lw
BmcM1rBJOO9qwdl2gW96caMo7N36B4+0dJX5TvmXfi2zcbYU4VZko/SuOVhRYmEp
hW5sfXq8WQhFgPkcfwPSZaEg1JSWDsbPHUFpi0BoXtKlI9EitqxWWdtAC3Sx+88s
Fs0I0Bq4LpnavfrX/WgM4Pi9SzQ22jD2y7Ob1x72NGKwmuqNMUNsfo/dKyaBdFAH
5RnZUcBhJRG6xHS7h62VTHSVwsdQ3P6iIZlUcg2w4Oj/0uy+FqjKVG5KC0jy1nVL
perISm0LUGRr0EnDvDa6A18+kJ4q6PYLZG+N6FYF/mJ2qT9p642t8KWXjyc5LwRI
uT8Pe62lhm4Teq0FlROpmeOUPD7SuzC2QvEX6P70FZ1B1Xtf7Fzk/epDTCZV/9DL
neBBF3c8iKvlSZG0PmG1cm+t9ffixe0sHbcrncbSMM9sqCE+nG1qS4CWMmC7Ajxw
2mUomiQP4pW1DV+2XtN7qM8R0hDx5NZf0UFRIhFQJ0I+qG/v3fWg9SbVQULgkO2j
4N4MSoC/dapjaBjwIY1nUHOzMxbW1pEPNy02x1oN30bbv82jFn68JYVCXmCAOfzi
02yoEJ4mUh8Vguu4NY993c1djVAp0gmYvi0KQOVNkIh+bPC1RKbl4P9NXwI5jX57
042ciFKbUQ+qlzaLP491KHN7QI8ceqAbguWO7QrS9CXk2TSAUdr7zJSlkoGieaRp
J8bwt3P6LFAZy7dYYxJQVJBhJ+2NPgNYbOV8GB4zPi7mK675x8IWF7BeGYvUWevX
gmJOhOf4vzPRVjgsnxAFs/GbOwr0C7Y0vw0+ZqWv4iuC5GYJrWpF/lI+KKoTYpUP
/20pU7j/NCKzagzyGgQs9w==
--pragma protect end_data_block
--pragma protect digest_block
9WxofsrPvSRq7WBy7SyWEiRwMEA=
--pragma protect end_digest_block
--pragma protect end_protected
