-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
j05HCfRn/sm3eDtt6FE3bVPAoO2e4YfMiuUXqomiVHN4h7ZE/4PqwrP9njVdDzT9
2b36kEkyZsvAwy1qCcLHLyU5Os6xotUvu2ECIyfBxRkFJceMiKqwOvIEkp5jRvhK
qNUccQmqCq87eV8+HFULnmfKDxGGrY13hPosQfGQIco=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5155)

`protect DATA_BLOCK
Gwv3tPpcsCbnZ68gQp6lNt0qQoAm4WNc2NQlkevRGTaroZbc0PzuvNPwYVloD2O3
lMTkFnCB1dNrnOQopY3V8YTD1ZYAH4nHQ4Mf5MqQWxhM4ofX9RcUDsZn+P3Vb9de
IApQQL6oMGwVvT2E/G29vSJI1F++MuxrvqI0pWwGRDcxIWuI8YqvdztbqZ0fU8Yi
kJXXXv6S8HGchnqYY+Epr00IjtWttZZJZcSeA1dEd1PPG9DCqvR9LxzzsjqmJZEF
fvcW/FqHCj7i+vWN/H7FaA2ozC578AAKMXTrHjJ/ZOaShhb1GG7hrPcl2phZVUV+
CaCqJeX/8ctSZBRiklziDmeLq39N0e1wG4gF5TceFG1kq2TL8BV9RkwOeJm2t2Rz
6zUAd8NQLui1YD0u+8v31nZY476uPsyXcYqcfw5gwgQqxR8eeridxVTXSj9/SPGS
CLmTT6OGkMZFZzI0hyjXvUdvwCP8gqrIYx9DRuiIRzP2PGn80hKtU4tnd3yRBfHb
GokD0RhW3Yijc9tTQyLUPfGGrr2uvnRvPltIHzezSXu/zIV8Nof9hsViiq+8Ym0O
lYmu1dk4UiCkq6dUjPZ2y7Q8s7t9oZMSCvn+430CD4a4TalEfg4Yj2XYWlx22YDT
RcZEwsG9YI0Ikl7nimiisJdV13BIkfobRU+oCnkUAf7/VI7fBN/5V79MZoFpYpty
bmcSBYAap/ZRFrryH9MYK+c1AIIAGf6u+a8mOkAWS6hz3laqXebk77eFFQ1tlZDl
Cn1lKqLL2bs6HNz3in6wGXM8/waTcYIPAfakZCE4LTIP/nHhhDuG3tmntyi3nR3y
TPLyDk/Q9mgiA/jY1xL/dzodrBb5vaBQawuCRchxNPT+k6x7MZ8XafxfZ73Jn1i3
o0WvG3ppnVYQ58pUeT24R2XBWgdWijM5PHSL5sKXnNwHf6CTWOS2kkyKvUpooWNL
HV1jcSimjaSeB0cALPh8E7vgmTO8e+H50GvFuLL/ibDrKSXv64m97mxzBtBBnTJy
EcEBvtNSHEYTAg5yJRy+uK9yGxvdzCKAm9wBuINxdB2FiuWiFTdouA/4eygPgWGs
x0qMLl8O8vMxvubjqCpiSgCGGA4lVsZni8Aj1kDXGZC7JbiWMeVSNoIJlTDPAtmX
tsBoIYUPAtvyc/Vi4aAo+oXbCDGqSAuh+eYxIwyl+q4TxLtZJ0VgmLZXK7ZXJZuN
QqH8FM4B4GtJmImwVvOFruQXaxNeUNQfRG8PGSeHIxJFO0nRNjoPtubTwpLW32X5
SlrD7N9yDB527xlLQMfs80BCyWwRtn0h+xXHk53eK0u0o98EMeVmrolmuGlGlS6B
YumPGOy+u/J9rt+XfiLQyefqfJHWacYvifdydgcXtOqQDFMrezKT4tkyCynwd6Pn
Qed2by/DNpA30mkxmcWt3/vs0htTKKKnemYglyO+sSf8fAlOtVCeT3xl32qFd5S6
x91jWnHOOHTp/aTOvZ7oDZviev2jk1F0tdmrkXsTR6DvQwi3tFFX0bJAFnS6yPqp
/pb4+PFAN6mFcHk2YN65ff7O9kPteqiYeoERpuutM5vY4VCQbPsXhME8CFyNNwwk
Jxw4XKAJ95FT71uQbGdX16V1oB1jQ5BZ8Qk2CUuYwHDKdvm9WpdlTlkHafEu15ZY
ZXSSGaO8/nqnIRqYdtAaDyni7u3URDlrfVqGePA7KWGhQMgNn++u7iL0dFvG8IeE
pc2AhhzpBs5yCHINQDisvfGh0YSY9V43YIXdQjj/Bs0LQuN25s604LWKw692H6ef
ItLNxHFy/Nan0r+yEE20bD8JiZejPOAu+gzfYDaMmzcckpgfkLquAY0YhNqcZsP3
GpNStIWDDxSO6gcrqsgWZRASon1n2ue9NCmlJhA3LdgLpObvv5hxoc8fUD5T3Ktg
cLcL6RDLXdxX+nFJgjJmIOSYKZnjnZtA0CN4i4ZVdqKphH0BHkXuE6fBPgIR3XjA
5MS4e8fUyP7XqTqFgXkQz6eEMTKrxl8M6ssCuyqr76DkGpUQ9WWWnIG+Xz60j7oi
+b/mQjYVScFzL4ukO8PodSrxyxRkTxCnZTI5ADQ2N/ByMMhrKxWeP/hfL/3Njojp
flYQrkZKiq5sxuDlIUsehICUkDLmRcDG7v7jFgcC/jzzPjYX1u02zJrz65d6nA6C
ShDF4K3VndCvq8EstOcNEBzYgUwfgeHb5QhhJU6OdiuC4RMaMGqs0Ev/+c6fiyfA
1vW5PnvT2YXSy/VS9CtXHameE/yRzEKodoE5gmUbqIPo9dDIdYGyipVVQetJ4jid
N6vgucBhnxHa144InsFv4lPe10+dvmRzcK04QXETd9Jly3ei9RnkPtX+Vi0iN5Eq
+6hLpr5pyHM8AaausKtdPizUEVoWUT0lVnTqk4rjeY+n4Lpmta3j4hgQporYpppe
VtK9FwwZEfCahkOrKJuYF2n4eCdL4lvCWSPoDqxMSYp0oaNvxq78IW7AbBeEVDco
lnp8K3NXCCru82Xtn3JQYMx6KkkLxJWULb5C8eKdxVxStbpRT6TpIIYI1G/T/rXj
w57BvLqgPYgaXZwZ8rRGGnefA4z2tQ6XGD44WqjTiYzbNfVXlZhWH8gKerxM45ZB
r6iHbx/R8LZTy5YacB4g2FeNwgJRvG5VUUNQ089rHheXqNjNe6LpKWb5eoYOywoe
UEN++OAEwaIkAd2N4UlKGvLH80KKOGxbbZRxPhNTMyu0KCaeo/Si+XYSBjvLM0Qm
wqr0cuwUwrIqjN/mSkxX8DWtBryQbWWEic9lI0wSda9KgbKDH5PttA8Y5Tz4TQOi
RdDyRjl+4OflTXsIk2dekeqGFgdkiEBFmU3lzLm2EVAYjrzkHDRYs0aexpXlHXZ3
Wk7oqDQ44UsLq38gq9dwdyrwv0Tf2U0S3XCqmyjhGmqalr1sIiCR8gwFsCQh9qw3
gxxPIJpmnvxIfPkUFjA2mHfg7IXrJJ3yXLJqpIRdFR+cw3E+f/MQ0sIRxMl/ogXt
turQ1K8t8ea6510pK6wyVXaGaXrUZ7xNZGG+JRu/SrY3NIYB6+yzE1wSv7QVxG4P
jtjGLcVr4ofn7sDrGAtbev+vchujXu/izbXVfFC80GYg5UCI4xMGhkxigPBCT60a
YIxYrayqB2t5p35IvU9+r1XYeAdNdRgzM7rLiwprhDCnzIj83xmyW41qSKDHuw/C
mZFIB0uqdrQ1FvCZdkbfJJqqBFwmzo/5oCTY7kU9xdPv7T9y7hVJd4yAr+HmEncK
0dICaJXoYodrAP89XrhRe6YhDD+mQHGEcicbq6RQdZoKuE5ibLdNBniTzEqXxu5f
Z+KtxGSV5TycJ02h+dH7LSY4g+P9+BtW8Ou7+bMEgEm5YgkX4NtiEVpkYM8kYHt6
xH9ivHMqfbP/3COqdCHpmSwKhOMwCn19lVGhQ1fSrKut/8aFsDcfJfl5Y3P8z35T
E9AsNlO8lNcNt49nQAGgVZK2Kas54JZ6c0zUt/oN6UXxuPanuUTv45D0HfxLfRKR
4Mg5ISLR22IiUDtfl3gP9CbtHBWt6KvmoeQLp/wUFwltV+i8DwyginBwJaxq9Cw9
O4yRDYmhe37+OiZeHbhFBZ5OOmvw+jAN8R6y1Dn5Gdt7ZFb0o2ZTDQnxx7ffoIUY
0RHuke+R5DZqC7ou3nt457/s31MRJv1hQsZYXqjBHgkBPtSybwf3Ymvi6V6+blBc
nty29jbhef00D1GqhaHagnHNfh6ou+t/8zbS86DHxDIE53Y0BP8ptyL6PKHA7COf
jKDLM1tXoezhIU6+bH4QUc6Kxz/DdX7guXvTBjYT8Fm3l18Z9iJcXYFzr+HNUHw7
O7BJLtRaAqXK+GLeO7YlO/kLfYKam77sMcJBpeqqjgynktIN6VaZXD7yfLjdh7Xl
50eICHygkAFnn04NyHzMALhssFSRw7ivGf/DRQ870cgHunKD6F5IdeuxI1Kmpzvp
sCwY9+czatG8pWW3PByLJx/r/BbX8O8pYaId9H+GQAJMox1Licp1x40Bgdwys8c8
Ua9TQpTtwcdlh+We9+h2ZOqiwn/r0LoibUpwrh+h/pMoabk2uAPsSsE4XEsUG5Bm
r4KabD3mNcjU5AbzYfEg7HTXFaXs+h4WnSok3MZHxoPqmnzjQ3wX0lG6w0snMx0E
SKmHrUZuW4LSvkMNG40CCRtZmPFGLQniVu3IGwyChmauMGMoOovd5oyI/mlrzq3Q
8Gx05bNcjqKo5ik7J1dzrpsr14m5xNejeG2R6v//AFFtkChEN33qM7BzjGrw/7tH
r+Zwifx82VMxUZakuDP7YpRUKODQGwsESlVuJWfyEwzljTu5mjf7xlivi1seQnOI
51fUo1IB0/M/zotgotf8F8MPdUnAhOC7lNgXubIJ0n0tYi/7XZ7B79rTEDvHF57N
jGQp2+c3swyd90zpQS9EiAnd9TXrHaHXZ7PfKudopX4Dny7cVN2bDdEAzYwoaEYm
K785z8wmsPoFCIiDcZOXBHJYyHUeVGYt/O8nXqab/sJiRVud33NOWYFBUA2H+iHi
9OqufBUCIyk7CQEI4nanvYXgi+M8IBjgmmTOe1MnOealgcahQUIUo2EaFWaIGkG1
sgSKJUpjGwEwjwYMHuLNvOdC9ZyvKy4mEcLVKjleDy2tgfwcVhWhNtZ5O5JjafLF
vziPz3+GZsXXmwmSXqph4nfzipwRcT5iJDVGM/ZW7u00C6Vk/Ii50HzUz1H+BRLU
fhu4ELmKKO6nB9Ub5pTY5rpu00t7weYgTpS5LoEFkAfVM7YPY9UWdGREP6zztQWq
T8MkQm9jJjmVXR255/VUeBqsf2TUGAWls/ZuJLMjto8S5J1hBKSTGE3i62iq4Yom
DU6ccaE1yAz68zDwU+6r83imO2G7hH3ZHL8Nw4bVp+Yx9VbK8PxyGCND/QEdK+O1
HttTx6KaRrEtCEaYsRauSB4CEtPQHg8TYaTsSLcbIyxgAbw1FWnRhyMrfWee35PQ
T4Oflr2+/TE5lJJy1Iv5KIJ6vuuTRkALubjKAr76i1qr9n3So8LUZSKZO5Zpy8Tf
SkVaOSKdxoZk5OhNpm7r+bRD/HlElfEVzm8+TSwALlcjQ9mBqOc9f8crfL7/bDjt
uYjwP+GUWWFCLANxoA6Tz7aEJyitA3Qrozfz5GWegvwzKmZsyhnRIYJaCuK0cklI
puAdMWbL8e2TOtJG1uVn51hCZkB4KnzKr+/LK0xK6MJGC0sxtVbIIlpn/d4p54cb
9/SWD+iAD1BoYZc5DW4pNRdbsBeUhRozBLMWXWISegLWdSHI7MUvKuuxVRFRLb3m
jNxHzbIl49BgEmf2WVEWEQu+XRoo2qG8svvVEWfQdCWrKOyqUEvOLE2vUbTfrNZF
gEFXQ1cDUodv5ZF4YuOeqC/YMraCOTABbecxtXRaH6SEOLCuN9GVT0rUfxBWiJh3
dzhh7auSQr4SUUpBmUGKVugtc7y1kyvs7hj3cvT56U04MY5rZpXK14N8xXFaBPwt
tNoN76x8w3TExivAwYU4yuS0kbJZmnXPFHDl9K38QUqorncn6QPUuGqwf9/ia2f9
CKgzYXm88I8vbs4iJMvKMAHidTAkZa773wabbAe1tplwk+POelB2YXbLBt+vOdVV
atMoQ/TGe7DdWYyE7XWPnhl0XBLImQM7VBHDfknevyKgHEA97Bce7QKNHXsJhRfJ
CjZmjcBOObfOT6CYtFJLGTMoqS4K6S4dJrCmrDjtKeKjg7VHyKgQII+j5YbTa8c0
zVqCh3FUTCMtfjx2VbTK7N1zU20vko7Pced8B/3EDczkuaiprVB+3w5H7MowDipQ
n20/jCu0L74wd0gJc69HxkIBbG9bB4GrPxDECXo50at3ZsLd1nONgLlc5ypS3gv6
K8TRi1479cT1yrvxyIlAOHvMpG+Jch4ZpUp9UQlNZObQWoIIxLlZT0viHgdbhCbv
7CZbwAoxJVFJvdWXEdir4p7LO5cxS3mC/HWfaQALUNKzYLO1V1+YFAvnpj818Dpi
rWwNIPVuNBGU9FbqDrCC2PsTTVx36YQbX3BIV0M49cI1dZVSurgRmy6iV5FWFD+Z
D0pICDJLtV9hc49vHDZfK5PPIWhZnhe3rvLSV1UGs7PfzVnJ4qaTIf8jJlsSHCnP
WL6z20DIK8jVqVZm4P6wBD+nYbTSMpGEgRvJdmBa+H2ijoD9CNZlWczf8WBnoWTf
gVGXa/z9E+SVpbLzsiel4sUSDzvzDi2Qj53+xKlxV0HHsdF6cdQrbKZaY/EARfcm
ghu4sIokGWtiIwevBUqIQLUoSekH2FWA+OVysndcv6r/Dw+A/r0C/0aykjdaRQcf
zyk680GXyhocAtzRpCSp7ThmmMFCTOnYU4K5hUdFXXuZiJXbeuP1elp0bFGEYBbW
7LUP1VrLe8plm5gufALbse/zJM125ME54S2lFu0ctooTMn+rndc2zl6cS7vO5tXJ
Bl/F/zUXP3hHJkDpWJjw3+zAUVLf8oGuIGjgrUf6OjsyApxPghq0IsYdqqs9Au+e
bo5WP+r2Xs4eMO5SjjfbhQs96wF2z6D69vMsxi0EOLUEvTpmH9roAy+6DSVOTUpp
R8t42HWdM+CST4FYh3f19aNw9nx7FyoUhRBQzWtp2ajsALKn+7xi4gSplydkT31q
bS+i6GMwkVDdZfB8yJtrgPGrn24/zkp99CflzsitCOtkpHP6oZpuj4d7Kh3yRmbx
aDwn0Mh8TjlYHl+K7WbvEtV1Ql21ft1a4AyuSSqTj4Es2cAMBdHtQ3Y66nQkNGEL
Kk29BI5kPg5atAJiuNG1PcLcVt/gEyB5q5dHUDm+KxUpkT/MjdbNpL7ukHvA0zAv
ipFG/t0N61AbH8rWNuntZnMBwTleORvxC7gtp+v8al6rFMDl889wd8L8kPs+k0iW
`protect END_PROTECTED