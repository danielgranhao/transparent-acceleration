-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
hVeOiun/83Nsp8wogzKud4NKXolrpV9oEqBhA+Avn3Gddu90+5TD9Y3bPtsVXO0h3Wd0wx3CXRm4
JkZjuU2rfUxIXik3O29GyWfO5LhYfw0Cz5HjuPR6rRju+BwNWKGYDjpXFgIKQjn8sEJc8+U5FV1r
v/HoaAQ3aHASS5NX8fpiiv+NlPZTRuCG9DMTIkOuPk4qowT1i3b52PyWHdJmiWmzqPD7gZYj3sKs
2IKUN5L/j3G5g2zVi7O1UMYM1C44Otm3c/dAkXKHuW/9LxbcMOH2rE26upYZlHgACNp/55OcozB/
ZpycJVhraSZhumvCvF58Qprg8QiZKM/c+8p+IA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11552)
`protect data_block
7yL7z7VlJ8T5xtOBGBiGMYGRLzH9mh2who2hSK4w9T4/7SVW3/b/U6ZmPHxgQNxBAxsQvvYVllKA
q2CFkPv7nsNePqrvMhZMHIUwUaAsQogcV2+T+xf2mSjNDXtldWUIWtXOPCUlW64nOH23eYsPxKTW
TPYHx1dVg0rjTCsCKQC4cMmWH/qUz3+3/tsljOTXUWgbDDTworlT5gcg4QxU+RoHo0jdEqoU1bg+
QU1ghfZ/8Rcb4Zj/O2Ku0yGmISL10/t2evhfXEVkXVXfVdO8oUsYC+OHf7M53BPwutlImUlxQEAS
ltHb2EHCydbizioHifvWTZz/W6mruMdPd7fZlpY4npSgBUvCv8Ojbp+FeYsRSkM5mwjAcyu8b5DU
a7u95XPglG8b06R65Cq01dBM5rDdcLrVvNyUydQNfqUuJVkzPl0FXqEZVlV5UH7tKWogGzKCcRiL
a0DR6LsSif0ObjNhe0rt3QKQeGX49amIe+rwW7tVfX2sorCN4OTva8GSW+vM+soMm+MoWnPa+KTn
evuCs6O6fxGZZLcJeUE6nzKx37LmsTLLgAwSH1PlnvKrkTDNZqqh9Z6+JW329d8o9J72zUcGyBja
GQBMW1CShjWHA7ZzN0oQxRXYzHmFO2m2aAEFKVnBzi6T5uD9K2cm+dCnfDTePbxyVTkSjzig2nHm
3MpOGRltadwWNzLCnwOQCLbXDnwAEb1O+ypYo7J1XccohHD/pXVYSpnWP/JNTUCVM/COQXge+7/X
Rj85IlhH3gKVU+72edRnB5yOQOMnMpftMrYGQO5FPQM9oXrmcFk6ldgLm7mFeyTPvWT3uOP8TQin
FdSTR7QPn7zJi7KUa9ZAEENfPomhLChBzy/2RFsacBlQOWnxVsRvMMK3mHPonaLoTu+Oq/4J8Oml
0rhXChH3TPrs6BxSNKiF6umrRAlKaluJ6oTAIK5o3/qtk3b7MQD4alYb4eaZ0zynceAS8MlWz/Ir
1EORJM0oshZWE+EC49g070mxoWJSdYrp2v7O3Wp3pw8uwKo8mfoMiKMkeshAyzkcMzEi3vjQhBfB
Kn0NuU3pIpDehrUJWOQGczLeoL2ykpw6QTyGvJctCta1bp2l1w9YoLoFcwt5f+RGNArwscFb6Yfd
/SIXEYDOhW453h3vO9gBx/DCCUL2KHPMu8LY4kaJHdzzsuOZCB9x1d7cgAzMG7jeVuQFYb0w+Fpd
N0+oU3LEeW1CXPep5pTlwuX+qz/xK62g+Iiu2jKRcngFiPAJTG2/p0lqgMi2RIonxI4nUT56TQkZ
1H5jGvb8p4xKIW5yE3oSnT4IgmHnkValb+qYXD79H36Jav9D2k4WterRSNQxqChczv1SPvTVlKtG
gZr/vUOSU91U41ZP+uJB12U0/RsiX1/OEOZ9Ne8lhNkNO1/fi80KO1mo8vDSguRn4yMngeE2LeDb
iiZpPSTgcUj/u/ZN/X0Kx43ud5gOmH/NH//DT6yqvN2JOHKOUN7cWjEJzg+P7HyPG40n+k/kzXM8
cYvP2nYwyhMFJhW3y8PHrLKbcTduvq2JXJhz+nZLvJRF7w0Cd4IEFU1TheUpZW60AWGk2A6pKuPc
/2w0NwjNvuGQzgsXIH6ATI4rMeJPj2GdaCdxsblS0kZ8IxWxl6FWzoDmkxbalc4Mjp1qHdCkZXTC
di5e0oOyZ4SVDJlri7feYwR3LkdwipxtsIVclUZYSZUbPxhvukZh0cTRxubwjy7+stsCvevZ+qWO
8FRYRi/LblNH6+h4yEXRTlsekII2hcua6y0cNIyFOOh6I9fa1RXwsEFj/LNX46WFCDi6SBRG2VrR
AnENfqdNnVF+VJ1bvslHL8LMZ8GojLzvb8QnXRzIUPLfDZISLiXvuCysTXyCVIjpBIv9l4el8Wve
UjEQOMHJ/Ke6jr1TqaJYnUYB7Gxi50erCY4knGwnT6JbufSnlrqG3mO9Tjo0JMSAnmQrjLTJMKEZ
D9M5fNr0/oAc7VET7WwmE7uRH0TUF9asnZt9AOSj9yqUE4Whl3jlqHGHdEVIGbWucxf133Dq1DsN
iiKXkExEotezc+/bLZmMhXewqFrGIsW8/wQvMc/9q8TXor2SJ2SyiE56ighXjQE43alIENzkbaMk
rx9E0S7IpXQE8axxMrzC/zrcrYqN3uvxKgFxCDrS8JvJYZRNSVDbs/vklZ4NVJ6Tm3mxfkuok30I
zJBHVVgYad7M6Qv1McuWbgRCOs8Ygars+hVwe5zZULlIL7BijCQJfkAxKyGYC1eW42pHA3OpTxJw
CSvJNWSJ0MIkubBLYvfii+35vfy75qfFgkIoNhI+pyPn/uClsRegYARGOOBtj3QWrtydoNdey5sf
CqOw7T3eBNQYYxlQDXWIVh25KZ9Ecg1KJ0b62EuXJNjtxRa+jK+WI70J9ROjrkbOBQyQdDA81Q6A
IXraEBsHMNM31sDx8Q9bDxxfKXBIYnslMngh6MqHESAVM82j/rO8XoHJ/mJODl3KbW2DzF/xbSOE
HoIEj4fU7owhEKGMDVpZf7rol7/xfmyXBLxn+KNAAxHnAdc9sfLmflkPYOoilQRyLFEzOwYU6BFk
nr6P4LxJZC3L5pybG4wKrNvIgspDZGVDD9ZFkZMAe/DSnNJey4rT1kXozLky/Kg10W7Qq7dXV6FC
0/Jv/x6r/g92q1wAGVpbbJgHNllnBfn/Q93YBMAPIW+pec7UnB/DFORIxcVKhDAWPrc1emsazgqM
1zmJaOWP9/rJF6WVqqFpwoww730JlL8WEU/7o9Lw99LvtsZf+Cob3cZf9v/UO+weM+ajHwT+0zVR
rEGS+4AquH8HUWDKNDp4bzNldkEvREW1TxiiECF1cJulM8TKck3XkFwasQQdUoMs9iewWcZQ/5vU
HXKEITbhd0kj95cp4dxqY7v3StTObMiPAEEiHlLoagS/fD82CwiPxxHi3RpsRonLKhilaq1B6XmT
fhlQVmrdR4+v3UUbWLygYQRvlbH9mvF2CR5qlcvt9XyP0kNY1qggymD6W2h5vqCai++Vn5YR5jk1
4ASooVOxhg6ziMM06YR6SAruEkOBL6dEUlve2Xm9DRyovWhEReAUJxrx7f5mKOPrYmgGvQWQKhNH
yknZcl/SnARB5+InzYkb43BrpGLFWDF9MNZR65ziRZX8C5qzIpb0520iPFsolOFgWGU9484S5eIu
jD6fUXGreP1hE9kL42n1rdjeYbR9CReYoc0WcQpEYmYC2gwWYvucEBnIKpCi3+y9HAo8h6kHLZzS
kkNZLOIt1MbSx/AcrSf/XxAUN9kbvTdlNVIEyRgVJxwmY1oT6dMoVsuridee/6CW5Y+eOJovLgYE
XwdgCsEjXe0gmi9wVIaJdtCOEgxskaHa/+S3cBd5ohiRSEMNeR1Hi8f9KmdCWmTxsszEE72Paxm0
V+C797qCI3nmgEAAoO10uzVvRgGFutaiaBrNGvqOfPdpKQh8cPkMlWYC+Al8oLueDHlPf+27fpkn
qHqGrCSj1Ktx75OONvuYIJej9O0kP8NTzdY/jrqEtmSsuY15BATRkGuIvqSsjHebtQgz09YwVmEe
ptbTJdnMWbcP6OBHUgJvoCi7wwkMshvaoKwsvasSQmdP0bBC56mX40OcARlhJWfA2vWeiUXQqJVK
Fph1nxgS4hIYn4Z/dLInG+hOgEX9nDf8iiU/2WMpAql9tbhmfLoZOH0VkBM8p7z0tcnMZLVY8cff
vtE2OCGZIo3lvI/Rpty9F5EJI5cBxzeaNOyq2SvXmWwgPUN0dxqMNNM25SzXPDaS3l/u19QhSvhx
f12fvtAXWyxEwlhIqUJU2jWQxh0S691lSOXHEuy346gkmteArKAFXV6VWFlnARcK1uSbVa6uaYZ0
c8Egj1mnRPeJG+VvGeX6kwK+lZRJKYFxPfjznKvk6fECtpsEQkfBZTUXHBT2RklEfOR6CHBjLbBT
nIfzHlAT7mc8TMwvNzJ4UnZHVsd91UR0OfpDfkwtnNVXvd+aCp6kewrmlf13ZQWBhEjkXwmqU88u
IwPNSjsUYVyaDY+DsIDYnW6tZwFUZpDjFLH55ipCa4iZyhlO+kFRXFPuFRjYPttdXjw8+D9iRuFp
LprIMmUqZsFZhVHA7GN4E1NNagPP+jdGk8LEhzEJtORtfAAWahAxakBYtFLyyoLfNqCcanr/vjYz
qDdb1QjbG0s8e7CJoA1MMhugzv7SY6MMc53yGEkauvWq71N+ewycgBHaalVg5/ZMiFncUJzdjxJG
R9crd8Ix6q/Dk70npKvPIBn2yNjHGz+yeuiJzNLGMJDlOrGBDPIm53CDm/RQy/qJX0d3HZZqGVkI
eiffuVgoHK8xuBmYZEG10/aI9PmggO7C8WQla79MExGGm1LddY0GsElp9CQK7bhjybd7TqmmsAhy
A6/WmVvnC3InbzBJ/dpZzniQ7PaJmH8vXz1RQIyTxOZeWS+MSfhhrNIjuhj2Va63IVB3XrzzY9r7
tWRFxXDjltFxz5WRET+c/l66ySypyv/UU0HlvANa9hz0qgwzPZ58sRMz4SIpdYZTjkdvLjBYBUzp
iLSAtjj/rdH8RbWztKfqjfK85XWV6hgueDUS6Ye56DN0Q5D9kGrmHRXmHc/vId2xpxUsFFdipuV2
auFmv5t4vR0U4w/suS2qTQ9GmNDm/azUpwQhWoRjHB5rfFmCB7AsBphjfq9z58Jn8AKOUA94k1bj
FXaKRTzTcdPG818j0V+1tIYBMrWvxBuLUiEBZV8uKyWZXNdemxsXqev6YCxkeHcDqOHs2Sl7pcYa
wHF2EkzKLv0CO8LJgYCKVnUU0Cfnv4kwEcMKNVSmGuC25A13EHgdBVI479izzGRPMWqHfSejYd9I
xv+KhaI32mjzKCvN4kF1f8/8dgsDXvdag2355xnfmKliZik5gAABm8tWXEV1dFfI+Sek4dUqNHP3
P/8YVKT58Qcqevb79fGUNrIACiMafxzkNtK2xLS8IqaoJwagHOTStCYbAfF088wLtK2pqnMrtAwC
hJqJUuzJPH691IzKe/VLcBrqroCtssCwWJ4B93Drd5baWsZQdRkhJtZiRyEiAh0aWj3OmniBqeC8
mGqsIS+SxVsKJqcjt6nSsdaLlKlVHIBZJZRgUpMjAnUgiLgv9gSWwQBdaAC9VQaU4nnD6tOjmrnN
DvevjjmsfP8Hjl+2g1u982iJQglAsvnyLqj4twI/5dODjdMqgTgo9OHDc0c5A1Vf8TnkCEFDMQmU
i1MsrpSmz6am26LiYpe+YVTTX0e9tvNXpxfSCDer5yoFl9yKQONUWb/U7orCcS0yEhrKDG9QnuO5
JGgPRKj8CcrmNa2AaUNgjQv6bsTx5igL4BfCzY73dNAjI+aT6oUf0nJjPMA3XdzOEItPTNfFaGEu
rqZASqzD6u44vDjPHPDsnj3yrCwdyuhIeThTfwDLdXTyLaAmjMQ3MXWkT7R9fDqdAXUOY66NiEzZ
zS78At7q+N+Oq6Q3Mo4n/Xje29ok4v8eFOJytsNUV+CS0WKffZ5BngZRvQwBF+bFkmuevGOgCrL6
9laDMGtjg0a/4idyFjUCgd2hfZJethSG7N20m6so/0vbskj8MgI99SlZOdTnvrbMA/shGvnYJ9s8
2qjbbu8WNjhC8rNZ26JuVe1dIWqv8xKpH6cA/nQUSYhxIAfLcpisbEDOjHJynZLRCpE7muLd1okK
rs09b7IDufAahCnu7N/LP1vOJRM56chjHc6ImQsrWm5MfzWcbWLM5vPm7/J8MlCZbf1UFBsVvW/H
ebpY1rDMtmaDxyIOlvdVThDl5Xta7oNuS5yDerrtkHa0UmsyV7OwBo7ydw0conVglesTlL1yVjQi
SKzRavrfKxJvh9/dEA3LNTUAPM4ukETDENz2pE5vJdlI1qKWTV2OpM9OFXEFZqjLCOuZ8rZTBphc
CUdA1VWb1FgGQ2QiVfSWs2sFOlvMwiolYiBZKUXbHbSh0r9z6pyuxrzh6Twy4kEFi1/cAEFcdj/F
i8jKxedc3bAHe4ruiIybCHBlSpiVqfQr38uo/O+WmAqEUyfMpdgGQK4V9jmy6C0QhzZqqsBghIZV
FchzYqcr3dfeDS32Y+ajdf5QwcGyYgJLfbTpKaQqXdLf3VYRr0Ed/Wtm6m7ylhjz2JmGnJ1MvKuZ
lgBwnt3VyigyJTrYLyt5Fvq+BByM+8iRUqKA09SnfImUY852hCP22JUVYv8UWBtpNbVXn/b/yksL
hJPRXxj1959MZTXGS1oivhjEIEEPV28mRHr7eK0wzolOuakuVKWxxKPuhQx+bHFRbz8kERnZIlM3
h+kz7nA59Acld/JuqdaTVOZazp+0WWUwh8wrE2BP/erejhHf90fbuQ/n+a1eiRJpjD0WaCj9DwI6
i0R12tREj/EswI5heDMFNzA6q0bOSD+qr56/LqxuyloznnpvmXv6YfV7MhGBMTYhEMGmvpkNs092
BmrFb2HQAoQKAtZcrDA2TufwaLtMmvlOdoS89jV0s8iAV2oGciAwQVWElcowyChARM2xzVKvBfx0
zrqFx8luisDfDxeiiW4omq2ZhJ7PQW8PnQtG8+2hihun4JFWq15Gl9Z45QLoTn+14/6K9AvBAl4y
9gKWiLHh2195noRuEXHxPH5h7k1KNF4KObeGrURKVZ5G/q3pwwIJv9YRm+DCoNGk87yYbsPQ3DLL
KNVY0vnjPkf+1QZUrZkbF74QNvI3C/RWtwTdpqAa3sxX/DiDFImZeTu2XamTc8V/uRtDst/YP/2C
UYof04Rr4307+LDR6NlMDZumObmo7sS/QJgnBCY6pRlVvPKGZQ+B5WEnsr57qKJZcdM305yFLjSu
f45PuAKAsIEpqa2e9D2AB8DSkso8HxrJxwzmDr5G0tO7YyE5TGryqNVK0ssKrJZmJ4Ch+OMY1nHx
h6Oq1I8sSGvp2D75PS4eGprikLFwv35whrvuMnc2xCEYXtzp/TMAPoxqfCOefGHPGlOcV3m4bnTh
IhmrE+VRi4suoCDBn4DmeDbBwISwNQxekEEGzHKatAkq9Iprxh2Ow0sxPRvjakutfUKA/lHFsl96
xBK/hhTPvF0x3THGuPpibRhyQrhN9KDma+P7chrvxtfO0J75knSJVOOnb3bN069yAK70+Xzvb/B8
q8rsg4GtDozf4S+J13GpYbYJD7cLI+PGhyq3VxmlaE64uC36Cmvjylpepiu7WaV3bjB8gwEnuAJ2
14B/ShpuLav4T574LgNfT6LiAcZMqrFwWg7HQouYwqo2SigmQ4F9ngZ27phTFC3ZhpBtANltZSir
b273TFzbVHTvFt+Olsizedi1e00TPVMn3XpSpwLbXlStpBS7GVQqCHN/Qdt4QRsIREkDBT0GKxcX
S5qL0X1Z5CzD7k/9gGLCP3mP/8DMmE2a9QyAdbESqwYIyAX/e88LOtaJ4wBO30/s/yyNVRBFYGda
8v9KtoUhQBCdxx5DKegn44zkN5bkNhahFelxlPG2c9j5qIYYo1VfLcjWQgN/XDNka9X2YfQ9lrwD
I/J+8T2n9uhk81lCfPyepbiEbw4NdZ6IsTnb4jlfWa5bGom37n1jHkZVTIT6KdoS+d5wS1qxVQ6E
SvCv4AGv+5BshFmAbz8m/A/IVYFUZTmKB3XjsPHN1nYxDhooJL80HA6UyC+tjL7qHhuIGYxYz7bk
A9EfHu9Zuj5tD6Anq0AGpN8RSv7t2LKpXTBVvt3cOZqp6JwKGucvW6bpcRIpBfY4ujxb33a4+hlA
vCVwJpsO66u6RX+gxb2Di/gzkjc524/7G2BBR+f/r0D3WYiOanqFh5T0+znoXRiMRGVLF5x5cR3F
Q5kjWT4ajHH30ZaXfvvptK8LA78+YUqPDUKk/2/7aLNZCw2suf5gvNBddImrLZONJ2xgx3+gRe4z
5kMnAZv9QGulkLVaky+amA/Z1zydkOrI6nry9bAyt/OzuN2t6vdfOjaNy4VuX3FVkEbSA8jHhAX8
MzZn+T62Y98+FskyqacVPgn0VR5kA720D3EUrcrXjVpXxFqq+2ZRqy+VUqgxHsqVxsWys38abigM
oFNDV0WFUdlX9wh0TK6N6OIFcig0M3lM8QgMQ9F6Q3E8EXaokgk2BxQqNQsyhW4GKJZojwcJ9Pn2
ZeUZ5K3pWe0DXvK7ygZDJnLQvHSCShUc2NDUQWivuXr6/fH0JfZzQrHox4k6uHjJnPn453lzjQrp
RkxAy4jmGUTzMwox7huxlNoneIyEVWJYPXnNYjrZpi1zlOh+TIxqiiki1C2npOMjTx53cJHTFc1G
gCGY7qI+kHAtFSFFrctrnL89v5zO9pnyS/GB3Jhiu9cZMUfLPhKnwE6DW01TRPI7baa8Dxkb4umz
zB+rVjdOX9+UVyeDxu4p54S+h4uGeEwRnVWx25ZucDX9DathQYoHLBCh9SUb1gqhncDDCZOTSlXq
DCwotMOF/Z9HaIoUiM2Y033RoBXu38MSGl18BKKePrz72A/qUBcsbwt78RMzrjxgwjE54gTaMIxo
W6089n12QsRhS5h/hTjWD6hBp5g/rDVFzrytb2lTLxfNvz72jfQujS0ASiGSG59avSQatFvfmCZI
lgaN4I6DPp7JZVszc9OZsOpFB7I7OYNdRI8Hvd8FQY/8eglMdMJ28QmDGKNKW4bUzClvvZDUfbo8
dpcH+n0NEB3fWpZZrUYeOn0n0/bBTjB1TbejU7hueiuNYJv7y8dLhn3OTVlxB9ZTeM3EzZ1BaSzk
83G0ecYJZugo7mmXkM2O8lXvJmblwUe/svXXE7UAlWBfTusvLTUaVCn+tQFzeNiOmjPuz2yghnRg
RjYN4S8/mPyzOyIpnc/czH3kqQRJ7kMxb3mnCbTy2x2qN+a2/zWj82JV/VP/y8GK+5PDnm5wx+tN
AX9y2V+GBckgpJbVVDC6hzftB7qAygQ6z06AMTyX2bQ2cBzpGuRH29oGJeqsH+vdUs7/yrzIHmq0
b0a3B0MwHwJBCNEXNoPkqCDHj4nY1Mj7VTYurMJn+fbVkfV45mmDxAVSfrpEyn2HIL3jniHNqC0l
GmqG4bBUt0Jr9ozXv8j4MFvoWyUmvc9u03ugZU59+J0FZ8iBf4pK7hCK1yIAqL0XnOjAb6gcjU5Y
yb/vE6ZDmqdHAUmLNr0bozf3pRfqWw0PrCkdPKG64DAyn1gqHiObNQJe/s3UTIOf55h9OGVb7A7X
k6saHaXzfKypR2hed2WPhLXdj++ZY9d2NLmruhwK/mcuxYIiQzu5TTZqH6Z6ONYdS9lLfnoFT/Nz
RkeUddubZKWE/rL+hWE0j67FN6Na2FrBk8v1dGxIMilBlZRNFsMplfYvYak5KVj4wBNsjE7khWZN
FV3NgvH8GKY8s33HL3TxK5YK0jgNAE40jyKKr8BKUxKG4d0FLgMhXclgRxV+BDX8dYuvSgLoWxo0
RRJjDSkqafEeIyaPI9ntcef0K16NbQJHTUVgALPGCoKtTxdz9z4y6uGCKS/ZNEkVKT2shAlAciyO
9caHj9RAyiXgcnyEZ/eqUa0ZS5i9ZmiCUV5XWLctIp9UyGNV+PuHYY8MlRY6h8QvY8I4uUz2sUJ5
HP+CFkVNL4+JXJUFQLK1IHX+CPMiTWk6Aa8IXk4PekBReIEB2gjyLYfy1cvYpPN9h7Rj4bptrUv4
y7xoQy+aG7mJeKJZmA9SPe46aYsHwChZwDyMvxgVPpkfXf9Rzj/coBjVNRvntZNfcWDyfIHFbRpj
dAx+bbz/8dtr1Q17sV4yPv141j8nvz7iKT9v/cjrDGNQpJw6g7M5IwwGI/+91SIQ9BCn5UsBqvmI
K5tPabeMmtwNnu0n+ZRSXijuEAmVlswsKD3dwaJzjIl9E36CUyDYbLPwWQEPed6glDJWSa2c3p+D
7Epx36zpJ9J3rGA3a7SM4JF8iaCyJtQ3ROwD3XGqooRCG5pHLkNmFHx+9OP6pJS2PotX7reCyTB7
QyBGRyEPooHB4D2sjIf8MIQ59B+1bBNTTXRhUmSxj98tioVfToZLoxIZSrlIkjN07zBxRt4du+wx
uoXLgFsEZK76+oWpL0QkfXGGn54cTOoZvxZJrTSp/cwFp/fOws7Q7o5RKxupZvPlmeJAN0Rp1zZe
ZeuuTX7GaAwig3Y9XG+hIC+CzRa62mH77CpWjF00Jx/CKEOYuCL3cDHFxayJTUUvRzVXuPDWLM87
rTgMhGedEuQFtWBUxqEVX/12H78lqZBu2B0aJmj8yZpwC2gDx3GNwPznRYq6E4/+0DeUCCg2Vpb5
s9+HxFklweZkt4dR1ZwwpqGc8rb4dnDB5ctQmc5VdXTHU5PJNsCr0hjO+ObAoUPj7+kRUIB7ujIw
WwEpjZFsFfDKqgIdnZ5YpyA/bH6KsHYXR/w0I18+m1KxPHG47UlilO4tIZV9e7GyiOnB3AvHCskP
3QkZvFSuU6xnE8gFEL/DsKZove2lqcfGmNTGHNzC3WDqLLNi8Xiht1khh6e6jHC9cUlz2ciePaIf
qeeLXnU53kPDPflSSWAbMbj7A73LTM8BVNyvUx5ezt8Y3fjqD8UCQfXUaWruijl7/7YzeiP0Y0tV
QErRPV2q+M4YYysvZr/H2GlB9NTWDAVH+2QhlHsaAMXRjwXz4W4R+/kwLYLME5rZueG+cyfiMUyR
LkoUb/J2irn+i7r2BakxGpeS8mdh1NwxOqD2EzY8bM27evW1Jl5UZP4bPb3GNqJ9E0UXhADzE0Yu
JOdJ4+SuKumyBdYCtr/qqPg4z+odXDopBHhcY+FaQ+mhGoCe4sASSfPBhlrsPewZ/0y0MVcvmkB0
0nfKI1BXiZPNQduxPdWR+QdiQZUUa0Qj+BRgDORL7YVtvf0Arj1oFMThR83SflCg2ygKp6AHTI0k
sQHdbOmYMtTb8u6YJ+6+j/c3L81h86VzqBnSnitoxv0ZSSCv4AqVJP5wFVGpRbsqGKhxxF6gbvp0
V6L1PniRt6SZ1fvc9kvQ0J4DVzH7Wdn281av+nwAawR5PvIjlYmM8b4cvpBtNmuq+JaxSDh7uG5F
yHH8D6A8/6HaXl+Km443xhX5GMzu6+Xcal8xjqVcY1yGuSr/UIvpg6HQA/id6cav+aiOopnnMwZV
xiQbXGUy6VpbdVnbZGAzSudLP1UQf55P2SZudKutjAAh3oomIJl4iudtzJlzzc2CLGpe1NcQ5M+X
vVSp0I+CqamJ61uHmp6Pst9G3hSFg31TwGbZU0saxORTdGjvvIsMnBHC/gIml8Yr9b1R8tiITWNI
iq+9nAogWhfOZnyMEW2yZp+mGfh2Zwg4boqO6kZhKLHK+uFzjHFr789gUg//y2Bm92NIvrcj65cJ
XuGhiBT3V+pbLy1dC6DyNMHfv5Df2xi53kSX6OBTM6Bpm76+okLdI0s0Fnor8rFVK3Rotm9arTV4
7OibAXpOaiyM1QRYsZp8vNonjaeKOgRriYqa90W8FB722HY1qYG+s488bm+k4MiA/fwSINuUQrc/
zDfVyct6dJb6F+2Zo0+0POo61Da3x7++SRwIA3Gh32f3v6i7Gs0Y3iG25NYCqLHjnN6xyyZplp7A
jlCqN/jb6PuDK3eQBcz6IqVqSAg8avUOeCENNlOEZHDUUCmb9GC3cLMVqHEya8g9gUECI2jnI+5p
nh6sBEWmS8P4j2iW5BBCWneJhzOJM4F8fXHoaffNUT6i1/4JZZ6P3zwY0wmLlNODan8Zw12AsIEL
34VKU0+hbzzCqEN9J37p3BSS7BTbONIyxxyCt7fKlT4chGmGTYIgtsQxDXz0kco4aztWj55zABRc
jyws+OLGSdvg4L00mVylZUjSZ/8Of3BYrPVxWgUY8P1FHwkgWXta0QTNUXrnwXxtaWK5/O3Ovedg
8Q15SG8ydQRQsFSZRieIMw1/2OQu5/phUOpza5yQyXwXMmVmUPjtBnmn9p7v+ARXQcF9hIwYtUzs
8/aXFTZSuZVgZHUHzGDqQ/e2pW0a7GwhDxGKySuXf3DN6+wHY7ZaCj/VlQJFsKShTicCmEE3r38d
Rpdz1Y195NhIO0NKInRybxGFbzoUVmU5Hoi8VwGyLhDuTWFMRTyeq7lGAKiPwm0t4E6lrM1W3XeP
wkuhi3sV9VdPxf4nhfET9Rp5GCwkbSqrzTtl8bRHKJkiNvi91RfVk04wbSW+J+5BKWHZzbWhWEu3
+a8u70dPbkUIE+EZ+0LbcRxb0e37WYqO9tZU6859tCJd/tXkWX08Ddvsu65uUGRNk4w+ub6FLPwe
tfuzGBr0ysqbSmBhubh8AggQdcEpfPv+BbzfoDUGZpgj+5y4N+f0eckV8j37NKuGVDfeQEZlF4le
cjQi8XPyH/GLeXQEzXazfZCFaldmR6r+d80/lqDBeEZRhqflwZLoUMKuP9Xn0C/kS7wlQecPLsTd
sVPP5bI5kKdO8dcZ3NnwuCpv4EAL5tM7lq+2B6mo2nX3UM5V+9BI/S8gRoCqKIfr2JJDa5tE1niD
BEE/ZEWQjSX/olRGmaJ+JmTzP8kz+awgjQHaASaZ3mgUmFcnkBwre9LlHKoucWKy0tberL6tzTbJ
VmOv8OKRbmjdnPsZY9uBs61Rtyub68FJN1GAkJCmINNw3nj/FrwrKcpV2gabO7WSBzfu5NRkejJS
i1hlFMa0BHkcCMKZfUqev55307yryFdFeLiVkBRoKwIHvSazfgLp7+ytujh4czqTYPWclbul58NI
p/ZFNHDpMH/2lKl7VVs1aJ4YN2qCYJchb86WfAYshenM9IKOBASCZS48k7Wy5e0bnxotZDnQ727O
DQ01kybknIvs4jakKHnXoJPfwosUMHAz1f2czQ+yUYG0kpJRs1Dmffp1Q+7aOyDOPZmYm4fG8hnA
PYRtAvgQkc2woIFvXKe/k2iFn6rFeevNq9/hwwMOm6OrXpXefbR4fFO2z/A8osJ5qvEYN/ewfQCL
ZiBV2LJCBNx7JF+Tw7vxMJG1oBZwSUWTIa0B9kht8R3XC7ebQ4nrC9M+cjuSeXgrCu1RiR3cN7Ir
FRgmf5P3tVWmeprvWSP5wX8Br/LWXLA9jDEzZ6rwC4mKuOUX/B7OMqNpDQoB9w4xNZfP54A6kLYT
gZ1MKl8dLoJTuIJSNamF0G/nWzioOclnMQkJR354hG0/C+pcdrSpidVcFw4cXPfiBOiQYcrgN1kB
B676fIYLF1sFqm+d3kiYGN2rfXv3X+uzoqmtMKn9RxhEl2uDsnYWRELuF3fQmeYduJT2bROSMV1a
dAvlM5m/geuOHNy3QPYpxpZaJMVdIXyVdpSLXmfI1k5WgVRfTnlz2f+bxtcAjDVdvJBSwTx8uhTp
kPvHa3n8E6srNMBdo+3aCA9NnWEmgGePbWbGs8uD7e49wQbi7QdW5beiJEp0CsCsOwUF/nfkIFD0
IuJxhY9XrbzadA1jXf6nbRlgIIy02qZN6dnUXOnsvq4CO0745Ko2XEswR4nM9C1gipX7NCP/Udlw
X0khZ3U131pSUePSDYa5qSWPiTpHupTdP3BiLx8kvBYlmCkMMk9WvBES4OG40nnY3plblaFzTa/1
SfCdJdrl8onVHhgejXmiw7Lx2l8TBcZ523B+FbC9T3pvupVOscvkkXQ3e1zJvKv+xWOTvINCQ5DD
ws7CFbmN3UwEy6NglYThSvay66wXXABo6u7vKol5/gwyzxWiZYmgQprTh/FaseN8+5doh+ywrVZF
13/QzUpJoT/x8g6FbT//BV70xyJtst+qt/dXEc4gn+s3M5rmzOR4y4WFpxl6t9jR2l5i3qv0AVn1
I7/Vz5llMKQ1DTLoFSA55+eUViSCII+PwbKLs60Qo4WhFUQhZgq5CN+Flv8tcCEwg1IcNeG+gCIA
MPI0uRKVX9ypVOmjYP7VPtEgdKsomYToZNXIaWOoGUCo8CVM+qRGUjg40Cqp128/UHogQVsQ7MWW
lj6Ou7Wcgdcmw5UJBY0Uj5b0W/2EAl2PO31sBt0P1AQ/6h54RBJ8JXuR7uuYJXZ6x41LF+V8/Kj5
ICEAJ0xJa+mT2nxTysI/y49dmTMLH+pwG/9L4a80JaxSG/+MpZEHvIgMd2l8oh1pjp76KUk062HT
UJoeu23jN3NAr5N4uFBlcVx41t3FSMYBxGlDLRWDIdVXyB335yptozEWOYMNCfButsRncB6xNoRG
dJvingTrHPrqjAf1Z+31sIiJfM3EkTkZpJ7/58XFgzDBEpht2GtEvMKFWRJ979lOcVZSpckcWLS4
7JBVGm+gcuADKfttgVwNnKVu91AyujwKihdlLZr46+9ytYHEag0S5WE+2UMUuGy/2c3W/Wjsx+sK
BEuiqRy9iTMw3LhA3Bh96IDoejznJSWU37RqIk7y/BaDJ3hjxv30cIe7ORLsU6VPCHcJxo6q8JWN
hzwT9FBA0p4XCEDfQg5eP7Y7dFzrCK0KQiHRjfzP0uxuJX/YDZclh+kouXWRO3SPVW1IjYBOvr13
SAjsvP+1qrbrc9cdqwRs+2iWBKxpbfg6LpLLkxuDe1sGBdfZsQYYyI8VioouhbGcr/zYvWtVaXpu
to7f9rmde76EShahBsuBiRuLGafxNP3i72/1QkzvhnQ9OxcUp8dYuQnMlbGtmfDUVQ8xqi6yPzfC
+rIwIAQrOtzPOSFpND5lwmKc7KmGuMrsn+TIwdWeD81VX7sUDotpJLu5yVtocF1OtBmzkAhULPzC
gMZ6qoBVWiwMxpaVi6VUdrhFCA9q0Hxh8minIN15ogTeiilHa6DbO1zA3/0/sHpXVEwGJ70CRlub
Mv9DUib+V4X3p9NsXNotHssOFHCPpVb0gosUR0ZwD99Iarw5SzxPJcsu9mjQjnBXtPO3nj9DXV0l
HnKQ9sAIZ84vmAALHg4ilmlIETBBEGV2kRK3rqiiOAKAmQpeIjWOMey4amaFUdCGwCh+coKRdaIP
/Dpk2ckJxdzlLpALYUJ07tw1uv0XQuSQpA/UVBPu1C/lf9M8bKlx09Q+KqHEdwy3FWXqtNGx/O8G
HQVSD+/hziBcBFK14c7uk1zhZVdd8wOe819BQbHo80SnN+esfGuV9CPAOptG307mN+P1Za2mdpWP
bu9igdEXDoke6e2/q+LYmhX3fCmDkEiti3wnwNL3qcQ1NkKPRbs5KpbOTF1hGMuIqaz2xoI9xhu8
KoBOu4UDMT3soSuCnuPnMnJMepsDggNtUgasz1IpUbYy2UsfbaA1sak6aMMc7nQ4Kg0gaBL9OYIy
e/noFFlWpmmmOSuvH7xMnTxkK2uNBbeaW/Ehep4dciYUupSpMj0QVduwPz9CoG43+3rkExr2KRRI
E2Z4OprARmYdhPLbswewS1dvb7BQhml5x/njMv5EvpHdHH5suK54SObwug1TZEXmKUFZPsWItxrL
L5UXCsDfsHD3wbv1yBPD5GTbyMb4qduXVvhiSS2T2czcKRJDTaI=
`protect end_protected
