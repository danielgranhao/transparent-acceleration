-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ClBpJESc7ryry9qKsEfe15CwbN5CzKTgTFGMHaugBsbt+IPEmTXeoBn/x551TIuI
HZvzjzF7ul9YKIvz+yX57NQGxPyww1/W4nueVRLb3giZxZgX0y/5dllhnC25qMVw
tXMO642kAOzMv/5nTFd3BsR+K+aak5YsZ7aP7YeRK3YPUiKYRmiq/w==
--pragma protect end_key_block
--pragma protect digest_block
xJA02ZSd5dzsudZ8tjJ2gtRPoEk=
--pragma protect end_digest_block
--pragma protect data_block
BNE65W6pEUGfBZYIJTKZ38mCKMEq2pbh4CgGznauQtT93F6iX7X5vC0mX6MqwOAG
9/EbiNeukSeciqcfofwuhsruEGu3Sqr4BY0OoMmzW90mL4e4j2+KcDrZ5rJX8wDP
KgTz+kbZbdhnxcorrFLcOzHpRJBwY/ddUetK6A60jdfYBbgCoWH9fB7Kl+8kgcNu
nKMyI9XYP+KtujVHkdXOba7sfCbjmUHXhwddUQRR1+dHucbDXItfwtQ9cfyVlCd8
pk88gea5W/NkZ4KuyrOUZJgc3L3hnjk7u2C/uVGBkWYVmarxl8dSzvxQEnc230qk
1oZssbN0yNHzNJOT1rv+M8fjknlVR92DbyQm780R9M04hrS1LFULIfLsZZJSpdLJ
A+kcE9mRev9nyYSLwahYBYAsKtz1r8JYv+ZbWXzo54o81HeiXvyZSqPOMbMEH4p1
fujKRP/5AymT+4VcjxnfjcV0flcCnsUumm5imIJdrivD+AmYpY1Zo1+H+b3eH6EJ
zkjVcFMHU70zWhFvz8UmQryWNFNOvYql9+L/qzi1JZabbSGE6xJV941LGWPG5vDY
vx4h2J8l8Wyz0AT1x3xu/qfmPv1DlSeivwz7J9SbIKwpf/gpHLrSkQkTLgIB666u
nFL/q8vvg974Yj/b8XGCJGPbocqW0nSkUVrIAwg5sQimteyB1krQNBiwMqa7kxYN
OIYsCnHdfZkIEqXvJGwPU9fjSmzORYQFjH/FH3uCyoJdIa1fcSRH2RXFPJddNZcR
LreFPf+6NQUtd3IYSyilvFsZ51sgspJFQgt/yZNbgaI/ictQAuYJ4X7bj2IQySo+
VMPMoRkFGgIYDsY/Hbv0yJ4ojxZQueO8EcksKlS4yl9jHN4Pe5NI+AMN+waoMiST
C2E4fiSmLFAKvyBQq81bZsSxMeAV76fDfFoWfNtb93Jld8OhQrIoDNpfoPKUNrKj
xkyfdDcgtJzRWWgmcl6Cg8umjzd0T4eS4bE++xW1MGEqoKuPua5F/jBHGU1alTTA
tQVbGBVyddgZ/h8XbO82gYKjA2NHuIxzCuFfBgd3cWvOnt3rZ3tKA3QSXFy01c2B
zp97SeRPpm669cs8vgr6xsTFEwWxKy6CwKaIhMEp9rWOaFKNMCqEcsOhdvfAmBEB
D9KaUo+fQrTWY35JA6AG6nYHWcVw5Ce366Qd8bBOanlhcYZKpn8efBtNu8sHTlbN
+w4oBLbMZdmmS2CSv7N4hxyruNmR59kwxgfaFcRgKjNxfuyvdwUzA5mPhS7yFcuO
9wL9GsI+fWj6PQnE3jGN+zOCAaL414YeLX7TcebH1kOKz+hUGm6/KD2OkBmbmgKp
4/REmXwtlUDsO1CBkz06ZyZvJylI3raHhvRsVXb+DwgYYk6iUZXANAfNG9QXvine
+z5NrSTkrsu3I/xPB5SPLE2T3SSb1sZ8SDp232Gkzez64pYg8Xu1+yRQLIopMiwg
I4l5MpQzUATXg2ueJqugyCAAOkU7eWybf045DgXq6EaVFFLYLqUmdzvZX5DAETIy
4qQtAZdFATD/8eoTggtKP51vRinF8t1SmU7S4reXHI649w7CYI/0yM4DxFUciP2s
09DQcyjroHEasCgD5KCfoeAG90DFOYPGO3S+uG+X3rSQU9TRhmppSBU99dWYTvAL
RzRpwvIP+5Apa35drkZtNNUtMxtajPLvPSncVEHzXsT8659VJKrusFjPqUxeVRyO
tov/2FOSrbVKGWMC+MjwSD3PvmKF4H7o5Z97Jz2IW8aJRs1WmKMH35TTvjDcRs5X
HTrxzsntFBXyqu2PsocwrqvcE8V1EwceuoaNW8QqJa5toi10ME7P8jCmAY78WcQl
aGXDp8CiqvxM2naFNv+g87+Ie/U3kqeVRo5AIyNbSOslhmnIA/h80NC5qZEvYdSS
TyYmhyA4tLSo3HBUWPYt8yE/LPn7MKocLJTOb4MkWOPuLFnabFOemMp/X9MFhMDN
wO3TDagZSOMHtBAGQRV/QfdzXqLtliB4MVyjATtEKhkbOY3mFY92k4gLXXvtv+Mm
l2AbYjOmMCKKJgtvJ5MsI9smQqRS4i12kEgUp3g2U50RKParsryZFvRaZCkOelNb
bGgI3zL1PEVZvUIocHCa0JrM5jn1I30Vl3qFIqz3khwcXHvJZcxROL4Ot9WtPEj3
friJZ2AG51zuKflkoF0zCz9zQ3ax3Hggcde19HI7/VVmNlnaTJ8iXtBQtQ8I+9kz
/QEiJnJJGiYw2/qtt2FYyAfDWCRmcrYYINalyKXHWZgVmSQ26B4q+0aHhKTN3kqi
1nZ+zKLgTBVh8RWnrlyxp0xoAaHPGbPq5sJt7qiUOosP+5k4YORCoe8rapI/2wJD
S0KaqZXEkFddMuF4xNDrUTJ+MgEt1+xD9xKvnmEA8eL3U9Rq4Sr5mgOHCYm3c8K7
ABtIJAGwuQE9XJIig3lNh0tLQ6Xi03/gA1HKjwpWoECszJVnWaXtF2+InlYV9gu/
NH4LFQ89gRWEewcBrJ6Ou72pPIn/F5g/DqXbgrsps/IxRRLb4aJgu14wXjcn8mYa
D6nhTrIu1IPrEyqsTuRzMI28mUEEZCNkUE1osBYQfk8WRga28wF2rpz9bfa4AOKz
f1YIe7Lg5O2ZY4pBkjHKUUC4yR7ayERgaUmcwQULv7MxXKJAfhMda+/tc+AtKR+4
ddZYdKBE6viIF9sJVBxFnExJe/1idl2SahJ7No14AvNMKX84UF0KHo89OKVGN5m8
064ZYeQjhTFqc2nG9cuchAfVq1X88CoJFzA5ryZ3csY3Eb+c1ACqJ8GPtUMShKa4
yEN4/XkfNs96Uw+9aCB6B8jOBltoI4h6lkVcirO1Evt/hVyGXHNz9IC/LBrFG25+
VUHzh7zI5qiocBrvTlFb6XA4fntiCgWDewNO26afQzrtqbtAeOWWPDK/vVheI8lX
WKv2kJuRIn4Y1VBSnGhzZaXlTzAuUbSyYezQ6ut8drbqDm56CSfMU9EsKAYXtxxJ
NqCepsXD/mWxscbhwHAHYTIB67QJnVPHUr0rT9vrh5vtRsFioqCoezR4E62KUzei
9ps4iqy6SykaBBQE0XSomiIM9tgVAegUEOGBO5/YeuxWzTvVogcOWnO8N3HKgAxg
9BE9BUFtkQBG9ItauWIe2Qlcn7kRVAAbW3h3eQEI9Cyb96JrUODGLJpn07PMokL7
6/MxBxhAUBJIWmYXym/q0YT5lvUzITezlQuL+i1cqK+z/ZzapJW3r8P89xVdAFnC
0qe7lSa59JDjfy/hAk8mi9okyNHkG1TGN/sJ2LAbh5rOLQ6mBmsVb90k8/c/UpJt
j0mR7vOphmsmMn7QQ6j8tpQfKFxqFR30iwfIwCO4QrWfdQ1JKBPmhjzlroyGX3/v
+fXzB7O4vZp0mTtDejQTY+xngTWdBlOWLQAUeC90D6lHUW7AjpEH/sQpSyInwcFL
mZqcDvCn1BBdjPvNdJ8ORdoOyLdKBZd7nTseBuJXa1TKGLZMBIzF71hKYGWc56Yu
heQ5Z3auMZLd4pgermmRlzUzW2SBi1QUDFD9TIRbr61FKqpukTGYxYuLSEJBxVWt
9zyWRPxKcHdEQvST+TH+7J1bFrhjQEOHicwMiYXIdIbBzSwFpeYvNIyU3cZ7xqYQ
fAiD7/TuhVjvM/FGuo0IPJRNYfCW8pk26xh+852aZgZG30VsHS9hcYeLuv9HkXxu
BRGM9zuIJ9XhNX34G2Pfu8lVkOORnECJFJDQcgeqOSggzE7SC0AydTTFaxwwavB4
Fd+FlGmIvG3C3HIkOxoMj/fykwyIUYpHASaPSXgMuQ2kyPZWiasR7W5ZGT8TjgrG
QiaWsYUiitderSc63MuD95T8fININOIHzUUL5yqEkeLHjCDBdB82CT2OU66EgNS1
lague36WKq+Ep5d0s/Ed/blQdY/Ful0mhDbFxjR04KRKJ1/FJ3LUMFjwegHmbGQy
/U5aIfKP/rzc3RCDo60X0x8voLpe4Nv+S+qAqKDA/U7R8+N4PST2BN8V+W5hsxjM
l2ruOH8ZNYXunRpwDTaUBfAhVgnH3bKUODK/IjlJx7hDanmRwWfyRJ4DVpAAd9sF
UkOQNFX7IxJsgzS4+b3GCeOkX3O/3RbVhC8s+Zj8/YcEGxo5mpQ2A9D3w0dtsZxw
tqfb7eYFljrflo2dBCqgjRA+TG00KJKGdpwGLA+Hj3u6uQ7pFbxP2NCatfl5j6/P
DFhoKJ5T2+kj3lDF1nCD2c2KVMbCEDx96VotEGt6uqHw6uacttx0t1igorQdPulx
zexELN5+77Jvxmu2kTub7DNLapzILj5qsqmBFksO0YGrozJzOXkjjfmEUVz33vKq
dOvWgd2IIpWca8mlp6bnMOXM54I1hefcEdAkJzrJskT50LfS72mZMh6HtFUqbSDf
PdYIIVKaSwqGprk2xwzpLKWskxYJKTY/Z9gYfjBX9pEDqLQ75EPJzVDeyZobg+0M
u5qu+gnJnbX/ug74kVJIrJxKVbEuvIu6jrLrCcqgR9RCWI2xYSmvOiv1jCD2LbVE
2ke8JpDNzk3ptGnja8Sla7JyzdmeuFaLb2azABUMWxu8yK+rV4PCKDrOyN/zILZG
goCpaocuAnh4uqjI4zUqPiykVNquTVCPB/4FDt4nu58bExbnOvkf21qV3Eq2Iatx
rU/anNLNS5268NxwJnXLPzDlJy+8xpHWYxLMRznqERSU1Eq+MNu3k6tq0+hMKaSA
loxWaONK8/gcEJ8CIWSKVz9P1iOXoN0ZH4F3RUy4WEizPQrQz4dlC9aQ7HjCM3TU
/5nkY7ezhMUzuVxqiJghWp6vY7dnqZRlzE8arl14afJ3yL7xGae0YGPcqrz9sbUh
zSKksVL6dX1i7bYpVPfRVsmSNRfCyRS733dK87mMUHgXBuzcZvTwWn3tcb8Cvq3c
DAY4yP4+5EWESCH092mhkvp7DHY5v0Ixr1WSr1Hgby7IFcYEKFh+2bfPh9/EA89u
Ql4vwoVbHjBLe3Jub1SK+hKcRiK7yaKv0VxTHpSnbD59WQwxkpvU0XOCCuRL7YoZ
+xUXjPYSRxNhMzS49xkhE9SWlH/MH4DnDtgOZ4quz4LUBUWnhYE4TQL1Xjs/CN90
erVXcpShSHMl5h6OIQFWBx2yigQb00yuKzVyqe+XY9nBazcrtfs6Oa8g1oR9ux3M
VkoStoJPZOt3eXZ4BTl7c8kfDrqkjEIMz7KXyHL4Zmb0vUW7O1gXpfSEvwtzPWKP
agR+pD88TzMkySDgrQkSE4w9QLhfJcldEM3KZasxHSsk2+EdNHnd/eM7XGJvACKc
EB6uqVxrmp4JGMeeC7bSuWV+XI7Tk1tCxnfHArTINLgZVzwEk5yfCTxprb4InL77
SU2Pdx+2oZlc36VypgG3sRRV0E07WgYxRuANnzJftfpWoa+GeTRAk9vGOGcJmFuW
huj7RY5y0ZzGTi/yFPfSCo7ZVrS5PMG1ZogozbHxcy8eATpn1m+VARITmEagGMbu
7Etw/PI0grW3cPOai/lwXBbz7Ofk3zPeVrFZ0aMix3rtwUn4ztwgsqzG+LF8Cyn0
HqlLnjkNMBGsEZPKtAJT2rmf2zjNAE9se+MADIYuxGgjfPvAa5+MDGD2r2FEVdma
b0hG7JYPOdLoT6yPYCqOI1/kpzVaGOBIVmLR9VH5Xzt75UynPu0wbFE0iVTOs9Eu
ut8b9g4Qjne4HaS2pdJGlXJNca9gmDtI/YTYUCiK0Ie/NBDs1msUa9w/A35OcYQl
ClNQpC1RMGy4eb4cimzgLg+wLGFezENy96oZfolsbKoIYK5eUAePPnJIznw/FkJQ
9wZzyR87s7nYzaYBAo6JqXXju4LV/6PdT+E7rxvsK2c11k68SnelF9nU3006prGw
6giKqM5X1mbTNn9BpOzquajVMJ8UvNwvyh2Msei0n/mt5gebnq1Kd5/W9LkgEWdo
9WTGZgFwefmJ5miKsJJoKu2HYrbdQkbP3mzXYxyKy3i/fvXqiuMk2qR3rH06iOX0
8S5hElyb5om57RHbzWgpLm1ICNSAvAX9IQUUsTJRW3Mz/u8LyPiawdv+Gm+RtZfY
wrc/3H8N7F01UEAt+WjubxBwCdx6u0yriGy8bbhT1EoA05dE4wSvUHUHzir3RJqK
hiPKrmJXn4U4L7t9ODSBN4EHRkIhmL4ad22Jq9KNR7GivxL2dfz+t5LF+kR4LiY9
/T5+7wXpClz8E9GfeQ1bl8Kd48Vumj3GIS/7lBXNV/4jjz3hDbWX7F+iN9vlR3kT
ny+eoGIwlWDgPeH5pmoVK1BwyUiNvfVylvy9DuCuWAkBs91Rx8bSEMNU0u2gjOwh
S5Vn+H8YfNUkuliSv3pCTYZHo12dLIyCFSRUkjfNbjTGKwuqM6E4+aqLPcnhft6Y
Bpwz89rnaQGpO9dECh5RVpK+qL58tTGadFoFh4pOi2fjfTmlc4t0QTcxNqzBvLwt
dhW4LUdzZPyZlGfvzu8ySC1t88YXpmckiLNoEgPmAtSRp+xL21vdKRSpY6E5/qXo
zziwQ4ZgQF0qgSz3YUZi/nXP3r1CdQcWM7yUQs8tKLuu+czWQiUMg5NB4JC2l/DM
IPs7dC/RDoTOVFkFlzswUQeLwMcNrhXSStyzGK2mKqoO7osHKPwtjiGu6xs5wSMZ
nL7TarHthoNb8ivmU0QLPYCKhWK7g2k4O4JqF7TXhri5eFobDl37aoU1WpmqNKb7
jcZm2tjfEBGIQdIPJkUU3yRyrhYUQCXomxb17MzjrGABFc7LGRzzI/FGUqjY2aOL
Lr99DGK4PQ4oKrhxdFcNH4OcIqQyp/ZBU8H8eQioORHxKnv1nUBD6Hf+QrFfVnP3
V949pf7G5grnon+8RH98UVQKCdVWu1bHoqT713T3Vt6JUOs+/VLMGHHRCoLM9sMK
ErBaqKpaIsSW7sACoyGBRJ9THnzopsoGmuKJkjM0rg4hD1/vdXIwcowlxRV6vzo7
k04pkSioi9iXa0CSIrW6kGiiHfR9DdnwePnJspUs331Wp1hvPturBMu8wglVrjYF
97JdL6jAGr2EyVqvZSiOpaBA7+tBl/RWdyszJ2LXpoH9hpiyM7hHONC7VtVR/NNf
3omysHUvv8EEHOQHVObjwoHOs6ZGzrnkSOo+/6qZwwrDCnz02v1FpP+kCQel7jdT
xop/WmiOHKJmA7Kn9LlYUIzbCsRtEZM6p0KIx8GyUam2ziFIZ4c09Zj6auGAMZQQ
BcLD6QkrUyUDr8ZI0qIt749Hbr6pXGJ/xTvMKSMBi+3VrJbHYT7Rdp/ruTntoqUh
a+16vRxUhWNfhzHQZ+jMFw7NHGJYn52W5Tmg6ZgO5Z8t2eCBbMmyMgSHZeIIdtuN
wz4DU07vlR0Y/YehqOxKQzvt+AxPRYSM/9KKN3Xi+Lp31I4ZpT8pOADDcRtjsAnI
1qSUY/vSwUWE6OdtISCkchR4NkhdMBca9IvLc07YQcL/ccVzQR9XbrVold90ykc4
ovHqgPQbszoOzSQaigKiId/xrjX1BE7exOakjNyEtWkAkDd5Nl7iu/NrNC0l+Lgu
7cQWGfH5e/iyUU+jCMb8R1lSDiNbwHFEuOg9fji9HwwdTnPDHFv0+Pbq+A5E22l6
NrDcFVBvPemCoc1Jv7HwXyZ2xAbVIlzHfzYKkuGPJuX/rbetX/1BnMjecmOvo9wQ
uhwG2HJShoHkagt40RTZ0Vkyb5mmQc7F3ed53e+frk9F+FgHAf0M0CsZD6YcQJC1
0xQpG++ne7cdNEYiW6d3KZrDqXGno2lXy1+pkygbMqsAtMkzie8et4BIN3Y+k0Gt
vJKOyTTvuR5NcKGhCstGhc8bryVR8sq8HeKsL66F9D2ArBOYUvGw5lRnhG5gA2je
sNGjwH9D0aei7xu+7FKjvGNmdp5t9rOLi0OahI/uwYhgFixphgkLOnfKxnmPOKaC
tt6cXp0ElZbRrOXdPFjSmnvH3bFTn54k2kCylIgh+Ehkvpk+EVOCCoTVNyxeVs/I
i2j8SyhGNUwGoAshRv7YKIGdJuHQ/BCsvGU/Qsp2s9M7deCMHwbYtEoUUixd7aBD
lEmk2METV7zRq6jFcNX2TDITMEz+pqidFU40chrhfkljPXoc2+JZvHHQaJaLMq15
8H22p2H/MI6mu0BCEMozzI+F2mYkCzr6V97IR6zENUtBFR6SoZ5GO5AfarHAKoxo
tjpqzhzIlx4eXaHdAatu2RPVNVM8mIggWBwx/AKe13/NCoOGemoZ9B4EDEk5f2WP
cKoEchjEFNCkNosbbDsHuOQMq0ue+JmZuLaDM7QetuT92peVVa2DoDT1G11jjDwM
fWH1YBK+xDtfc7Jh6Dxd3nXb9WrOZrnbL4hkEmXZdIiyBMCsrelL9TTrEHMpa/El
koeIZuR4qJDiv49VT0WQNbBCYE7HTt3wUZfDy8jJiba+gbYCS1/kV5sLbH8BbJav
IaR05hY+7aqa3JM6qzm5Ejjg9miqDBIyDBKX/1oOWVVBA5ifAoKw7sC05DNiLoi6
mFTkY7YQtsNaMyEr5IcDf6f+EWnYBFA4IJ3+bx0TkaNMsrJ9qTUmImvTVddwm19v
jXr6fNWqOEiDHt/sQh688ouYVhipWcAKlMKKczrilESFve5qNeDAilt7NIO2sr8f
kb7sRjFiR+ua2DprK1xGlIxKCRJitv7oRsuZmCZxlNjC69lDgv8+OYIC4MWZuoYz
1Qn9620BFCP2qmq6U+a2BRbdk74CvMcMFhYpgXEZD/mVyvD0uxr/aLDTdLO23C2o
zB4elnL/v90Udipeo3D2D8WjESn7VWd3Qsl3pfFHR49lWEfcjgPY79ET1gkweXTA
0X/sDfInPHvdwHhUeh4WCPQ+hBaR5DxyFh1uKBWisYT0AymyvP/Q3v/o0icOY0I6
ok1WsTJ6Zo1zWSt+VtM0hqdtDojmJo4yZjJv5+BW04207sCIfAgYVkzoISHsYs4X
I5OCJHFku1CskB1uiswlbyZwCXFpEhbgfyT7nXY/nMl2BWOvULUKgkCjQML5RwUh
ZWAMV4IWX1UndcVoAqizYcRxSqeIk7Ik8pjtSaD4vnLjLpiUnuaF2XE6zGg2iPer
SkLycmmgJ8nZSMYQxZhoYxtS4wa9AHaOmgnqsTfgsjxx03SZ+rIsimz3323/uxvm
/fkTIcrFYYAHjyMohdRfty3+yTdvqczX+EsTSWXtPqcF7uUpeSeyntgyQk5XcdTK
cVzbjB/z9l1j81Qh7DI+CGlrcxX/SRR+gc8nmZ4aqiiW0LtikoFWzd8Tz2exDIWB
fntDtF1fmZF0+UEmAxqGjRcq3/1yc2exr/IcyjtcBXtC1pMuD3zjRXDYbuVEC1f6
X+YeQYVvm3e+3eqhnjyEY8+XHICd8XNLzFhEuYRN8qYT+cF+FAfvp/8DfM4e3TSh
VZi3S+PhQS8a4TbZ3hBUk4f6H/U/NxV9pUHCR4iueEReMq9dfYsk1fQzAHjnXGwV
x8puNR+o7/og/5PcthyCDjtVQR0n/XIr+J2AGnA+BpjApbV0Fko8ZcPzFDy5ztgo
o/NQEcLV7t6C3FAQ6Q7ljwYo7yBEr+DU2H7ur3A4PatsYLsHeLLS5QPWA3BNqCEH
wShkTKjwhY92Imgz0/z1gQbO1SiORDQHka9rBiLnMKx+p2Yxf9lbG/FxaMuDx3pN
w6XIzGON2YOM4y1fOgtPRXI2YLaDWTJNSwMyxlUDczgVJrq3e6QEwTIbX/+7OdF2
+Uyi/i/eU3w1ZOF8H4Yw+h7pxA6X60E2O4kwGxJ7Hf5f5OWpsrVCEMwDLLFvZNhe
uk8lg/y1LcmbS+RU6auSD5pCE/1yxlmEHJjT9hL2Q7h33n4/PyhZdsy8yeEa1tzM
yF6N+qZKdUABvxt8UYe8dPkbGV+wjlomLbuT3GiFXL7HuMY0wtZCxQut34Xk8t+w
jQdPLY462mPENHial/rTiG6EkmDoGdifUoxiWzmtFRJbovLOCF/4Q1lK+Inn95sn
iTj9SRNlLoJRZwpxML5XNnDqPzpNzmDHkZb2hhfYXdr2hwvMWYSqwvogOBmb1Udi
nIRjrfptLbEFXwtxMfFQUUEG9P/050S17rEwA32O5/jV4aTdS7LeZReApQiCygJH
S2fj47e9BpT6+i/HS2vgD4MfRf08JdAR6hd2GceMt7OrzIgFjkAaSs7PZkOTrc+Q
g0LdYd7GrX4njgccpeOMWsYZ8/Iio/l6QqOLmuNFFQttkRwkj//5bGNrb6B8AMOg
8NKF879oyDEECldDUzrtyKkMjaPV11Fe39UWaQnTkkEflHowoZULKqa/aaKWODzK
t7QK1N2VXfnsPijAnnjtnhdXHWdbDBofaEbyTmGakb1DQULv9Q8rHWEEoEqvuLYr
IygbJQVHVdoKiAw3K40PjxsIxQRTgzBCxL5+a8lpponQS31dqxB8tK16fcSB6928
9IMBF2nrreN9BWri9gFVRHVFK1MUMabUbdSqiNTkUm9dMGjiPU6+mRbsgWcIQax/
bODb/uQUI6+nVW7H+4Wwij6dstZKMflP2Lc7hBn1V5PHws61YFMxeprtJy+ZZlwJ
iEUcPtrTTHDQLBWtGmPQvBaewiumkN7+NQwAdDVIwrWTSj7nHmUriMVwCKL3VOJs
NHQCY/3LUfKgzOrSgsvC6HWsBYoux01FPtnA90HzjIkc4JBFaqtwUmdAmddsgXx2
nXfvmD4rIHh0JYFgqCizWklRkagBWYLz9LZaYsgJ5Mt5+Wu99CvKTc1d9rg7mDKe
x6xCrLuaE5FJueOxyu9KQkYxdZspQ7Ha8r1Jiy1/KKGJcPxdWAO8dR6bxlb4yWlM
SE0nvFTa+IUkzf22thYwX9UwV2KxV9HT9jxw88sKhfwOAqbCaqVQ5MPR0usjJV/h
ZizSUwYBgbdfkx6iX4dV+USAtBzB1Vc8zpADhSSh8pj/9QAMlg03cOpex2FdAx72
BL3AISnXS4Ichpr8mLosFSWB2489Z+yI90uJd7Lizns3H8j1KqydPryPrJXfwjRV
FwbEpv/Th/Qg9LPJDLtYGVlD7tIs1TfCL0JeN43DVLBAl90sqs2CucShVXwdbLfw
/5s7u9iqL5wdjhyLOzxIch/p2elOTEUDbzOLgO1xMFif7q1E55/J3qDUiaOjZyg0
EM/7DaVOHWpOrUophNUCd5bvQ8X8p6KdCTf3F9Dpe6xdFcq28ZuNxt3WufLTbQGa
0hM/tpBK78Rm+brV6cvUtvaX8HgV+OZWLBPrxviG41+4R4hFUjLYPhxktRgkn2c3
zMbr+x4/UVL0mnmV8Fx2/CnpQ0tyG2MLa4iwNFwhkHjqcqi1E5Dw5gW1L8b7XEYv
Sr3hb5h8uMoUt1pFIRFRQ1GrtP4vsqMm0uun0kG6P7hfKGW61Wh0uuiS382YMZjR
wByYUQ+ruLrOd9O0eEEWjXtOOkTM/Pax2bk9Dto7WIfaEAFriTYUCDvTuqUanjd4
+FlF8GJHsx0dmZwQHknSsFZwr+/UoYDcv00kXUOK+HY+ILeGzcaAY6oKptsE+NDk
RrORLTMcA57F+5ggIHd2jCxKQX+SnfpaBX4dGRUsr+TXDDd9qy6CwylalTmt5OnY
BrSGU2ovsT6IvHz0Hd1VpFi1/Tcv4dLH//ED/xAtJhLa+2bjfq7D8x6qsir3QGyZ
iBvaeD9Mb0szSgyqX9E9A+aKBqIGiaJF1vI2UhwwaRXbSzw2ktyIDsIWvqWb+DXC
1igr3QbjFd/bD//4spK4yaTesb5RQta0LvZm3eo3pt/dMMs3XpMH2aw/1Ll7NjHD
t1cGUYKOc08sF0JZTkwFMIPHdpfPzCZVge6x1PjfZfJOtCfCeaZF4esqhJMkm3Cq
yLiAJdRxVqobnoNyuhQsrMYzHoIbkY3S3JMjBZwE8cjBPGEbQv/f5vugKTqFWSgu
yf9YvqF+6WCr2OqwiQ8Dulz9ozDRfYvLkTlZVcFjttr6ZVWibdoumDd1f/h8mS4q
6s9dHBr+ZPJqno55149jyJ/uYvmXLUhGCBegnqXoUiYzsg36PbuUhmpoiOnN3iu8
YSkD31R1U6lp+tGXezScui3R+CD+QzNLMDPK0Nb7MzsBQ3T5LiR74gSFgCnyJhuW
0XRnotgbYpu23FBKGf9r2FmlnL/79PlrcCOWLkheDONxbqgijkcNpY10H4Z752Fm
UV43Ya5ixUaezVD/GLMMQx2vtNfUPaDrWwyj8rGSCnIhXHc3vGenWI1suFTy2hnR
u2YC+1nvy2wezpp5eRLIb+dZFXQwXhJbuok+DWe2VQlcFt1Fz3qv2DK7xcSShxmh
DWfkr3XrJMRUoKN/ZAV1Sem5uPtPDRrO/rnTjz9+6UERsogkLa2nS2es4uCwKmC4
SXMKmL1RhmhqyenMOofPiho2mDCzVIXbaj0k1YXtW0mPzVMIMaXp3/3RlcP4jw8j
O9idmBqiPdPjlIN+LHUPGk27UwtXogY6IiapPAgm+s2vHNvOdoBFwuQXSORu6SqT
NnX9oHeLTpzEBUBBzzCLDXw4muNhsaBWbMUoe+G6Mo0UwUfbTf7YDbXqDUB7sq3y
tU8/P+V51O/yaxiiOIVCBZacvRLVkT2nnFXIuJx8ulUNHqShIas6SKniN/9vXXud
UNLyYfl+pFQKa9Ocx9QH1nZrA5HcRaoeGI990UkfHleCp3YAtfrWHMLO0z5zI+m3
Ft6hYXBm1DIjKox1lBApvxdXtL6spnmssS4uG6F4UpXZI9zNcAssos6jep9OYs7Q
RQCyYOOm8ocbjObKG/dw17OG/uqHZrWhSw457d8QPf+hsJCfjYlpNb9KqMewL15c
nVaRAjEnvIOcmbMqUqvioZTO/lI7eA30HvOTs/CF/aRKFLNSOI3D9+TFfbU9ywMl
nOmjXTsomk95Gq9FBm5LnmTZow7cPOs6MdYO/hNVJb1z69U2VCdsWGKaB4xEF5rs
nTRWq1342/e2wc1NklhZeN7MhyShCNWnSo6FcM8ZkNTzch1i+tru9IGUFeevgnWY
+wGO6k763+cwBKCPW/QXdyRkKLyK+HN1imkM25towQJTbNWAxOoSgQe11uy7Qys2
TgTMkcaRejri9vo+hwlIugLkHN8K3JGxxmZ+i6pvZ1XqKz7F/47euu98ShvXQ0Kf
V/vvDhRNYXGQHsOx4dwjCachV0ucrrcvwaKptt1wR0NnTkGdW6sww0yPogFxOtSe
1LcWcImf5oZcqLjLAW3P184c+Ml1cEHMXTUv4Tr/DqHMa4PPGV0NFzZ8jAC1irEb
hLrze43gRrjDxgYG8M//1LZ65FsJ/Oyf+/NFtyQrvWVwTYbKydhY7iqZWCNyaluU
84SMbGIBUIdNqUx59miBGdy2PkJ1HNAoxIhUraK1Ds3VW4VRnuM9KMikK+bjexf0
Z/ihZikzGcyUlrQWk1U+JnUGYYyTJJWIQlXRYG0I8rClnUB+XiweD5lomA1guEUh
TaKuqRtXw6T7stMJbq/T7PGpFWagEwalQIqXE8I9KL+w205JZD4I6D3z5c9UN5zn
4AFgfKt6Uhr6IJjfvLqawq+ugCUvh1FZ8NmTNxWT8YcAGnbWOSg13nvnyVaWqkXV
BgE33Gs13Vy3EwiHibCrYv/q2ihwk5kPjf3SHpEURBB1bwRRf4SWzzf7haqghhCX
anXtmx5VxVUd5WB4ZhG0WE6bBRW0+2i1rMRj/4ehvgUYX7DeLWUwfVwrTKwcctwf
wm+FFWV/TjBHPYFPLXBTC/eH1eDQlHPOZ0zqbuE6gOWzKYM2H75NfQUszcTmi/1b
w+YnQVoM8fqGIxWjYabGcRLD0O3Joyf+4eGjLrSKDhq0szeV+96u24o21oRTE0lP
MIdBPr+LM/ov3zC2hor8lbc6g0dzBxQspJC9CMbrBhbAv2nPRHBJjluNo3H7MV0V
7Fn48SfoPbP3NFQJV97MdiWxIT1R/r4iOh9w6WxmAytznE6qxg/C4ntCbVRsP92D
QUx4Cm4F/9YVfQugB0vks7QXCLTlzMTTL9owpxRc8AQ3FvVf1CHZ6IsQLsUErHFB
hNaQYUGjoLQPH+FOxPHdU1OCzB6ksfAxetugMq+UL0ORz1FPHHq8c+dWKPTTwVoQ
EgEPg1TGHQZMv2axSaswuhn1XoVDHK9KfmzYspaJCvT1cQvdi2ElTQLetHmZrvXd
0ZBhjHIRbZr4grvzbT44ms6v87KhcP5JL2E6XbeLbDxaBOZoIK33+w69L9eSKQoO
sXHGEq6S6MZBilSZobNjLpj63TQ6fuI7x2OEYFJYyFebPMnvG0DzW7upLXcTo/ZB
N08PnUlVWh4cehskEaSif4xWhCxHwmy5s9huwtTlZCBAsZ/E1iz1SG4lYuuhJjOF
Kv8K0PvGoTLoDCvJxQw0wb6W19kSGruAkjoW3lQkon8UL56oLyaJNelhTuvTmOpy
6s2tbtJL2ykhUG5WnANqsgoHWsajPAjujX6Y1Hmd8s2TkpdqewzVC2otCU8r+ASV
xDtBNZFoIwByK4nLe2OvFGRtqBQwoExOQXydGUOI03hbm3ddWNvqyV//4+NQPfqe
4thPkyjkhhP+rAUt1o5dq3APSKR8RyFhpQNcYMt46XwXau6ZIUMDuU0X7f9eABoe
6NHjUlR4RzGQQwbOiu4ppA+BJQtNMP3GKdIC+iCKgpol5XwO0EH8B9P32zEEx8md
jmTFqjyDcYnwaPC+SlPqmgF0+4JEqV85GvyWh4DIXm6avjvNgE7zy2vvExkFlxct
Kd6xGRqjIiUyN0JNwpV6RUBkeTdnvhBAEHC1XZ/LSKgv40xgiwFY8ejblUQpxfjO
lodv1UgiTvyTEKk8Dg4x3w02Zq6QKV42wN/gJQnGoJgdYLJ696wrmZKIpcqEC9NQ
SMpDZegb7hF0MCa5kWbonpb7/+6jyu1CMof+rTbcEvT6SznbSOuNMxn94aX6E+1T
o5n8RoZ/2iIBcCJTmv7Ry8fFGFCcM2Q3s/O0q9sh5CoWKrLABTfP8g9Vmf5c3GJG
3XtT0iujaUZ+t80uBWzWeKXo71qrPZEiUZiBHAR4E+rZfSqUs//e5A1eL+ONaDBn
mwcuQgzTA97H/MI9HdQfuxCoC+0FjLf9Gl3Lg9oR/1NaEP7jXQPoxjjBr/l82oA2
cbrk+DccC1ueYVf4Smm+ICJHQ79za+whyFcpdtTaAx8627Bd2rscm3mTZfixNUNo
FhhYarrWlnr2DKBQKW71RrDOmJh2umQoqqgyP5+PqVIGOPPLnzjTAo/jo1g110uc
z1tiuosdxDMI3+3EbbAOuBnbrG2Zf7ikb6kvPqqyTFN/rUOy75pQwrzJBnNYEdxC
X1l1Cq7WWsEWqWQ4kCFuc1SJpkmpBnN84dCU8/k5dxK/njMJR7OypMd5VDP7fiiK
D9Reg5s+isxrNblFKEnmywWy77cgxueryco1MHeHRR3qq/QgdokcTf7TXbsg25cF
nPQNG8ohCp9KBrjPxpH871DbEbksEZ3sk0kuURJSwYpTI0YEQT/XxybSW0FdkXl8
Q60gL1XLJABq1vVD8kn3LwUcOtcJzfxfEj46sl02IfJm9GpG/ASVzUuOW3qy9fdl
xLf8uNrO7QTr+o+5hLlXx8vkOr+rtrkG7nP34O4zFtEFDCrj42nX/qBUma9zJOyM
GbitkLhvZELEUbDTXEJBpXRmuEkLQmlyiSUy526vjnJLle3r6gAHLFe5RRTnh7/Q
EuDVVFAhbbKu9wjdDazp42ArbUK2JL3cC3skQccdM0HGpBbmrrM4kl8olR8iil2g
MbemxZ2tCWXGx8vr/Yc8VQOk4Arqu6w1GQ+HVcNrGQLEaY5DUKQXYlk3BGhmj3kR
frGjespnGQovFYGbwSg2NsiGlWHKUfuiczuB0XouSjg7Lmr+jb2tk3osX8vrr5ZR
wAIHGcmsCw0qCPwrsCdAiQ2Qaayw8te1TQ7W/8IVKcrBHNthFNF5DWMQf3ioMn3E
cYUHYI9cq8bwoGh8cYc+VFO5CV8f6c3p71i/bdiBUFOB8+yJVXdAkiKPkxDNZ16/
dbBFAzT1tkJ/atMECEjdCpomYs2lfQkOw+xru29pUTS+kNUIBuuIPexu5+AdHzdf
9z3YftYNBwNRXvhbRlBhxxslvypI2ekPCw9+WWfDVOJCfcfPR4rR6Zs8KgbSwHSi
JG763oOKVZCoZJgAGTGiSvP1zIUCsV33kyMX0i8B46DOYHXy9VJ9d7psxt7dqeMv
ZojMgAZYi5K0PRhpJ2OK0/UfV6gCBmDkC0QxV8TvcebGEOxcfNIC0jm4E6CtVOzP
zVu1TCNmSPeUYjBNFhRian5L/qJX+IqQyyysiYNITEkV40K7K34ziODWh4j8380i
r0d/zOeEVkv4Ver2zwPBKeBwavsqdfzQuAb7LC8KYeEW6QWkgVFEzusOInDxZ5GU
HQdy9DL4bTfX2Fohs79cDIOKDNhZA9bwA1D9mQLJYeWMGsyARFxtkol7jz3Vn49g
qllKEbMYZyE62Mg1H8o2NFAY1Otg6MsUN2YjhSYgFlIJa83l6QkLAB2CnOrCasXd
Hh5Vi6iQn3h8z116fclJIO9xe1/P1aDRj3VNQa9y+/8gMsUFW+67ygGoCJlEGR5N
uvdLwSPP+QQKErH8Ta3cuXOEoFDP1oPZ6sS8FbUKubZcZYsgwBfWUnGmrf9RbpkG
IDL6Wb7fxlX15fln9+4PTKgipUAJOlHhgbuIRdgOU+eJn3K3XoffL7K0asN1FU6/
8GE+mo88CHOQtElIdi3BgaR2Lfmx0OOS7+wVFFhfJUYLiLruhaq8kSBDpmXB9vcl
zszh5U/ODLFVW/O2I5l33+ohH3Q9+zgVftfeL7aPU2HcLlKBjxPXgEb77nEtCXwC
Mtflk5gcebRBqQn6EecG6OPScEH//AxDJMgQzIf7ruPxgjNkqbLSIHNXelqB4Klk
WhnP23bskhGqyA51YkQJ/89rwIK+b1M1nmeXMlaOrehA+lQ2kafLGHoCu57WWZqU
yG0mT4pGDVKOVcsVFtZVcdi21RfJCMbXFW0Y6Xh/5ldhLu6X2QIYaS+UubjcWLXL
cpYXNAYVal66nPmLdPpCLW08uCe7bMke0HUG4z94OBpSMzh2wu+Xyv4+gCXd3O7U
1OWo0CzBC2Ixsr+DLEOJSC5BPw71I+23mW+jaIW3+dEXIq6lga/KnYOJYGrHDJzu
StaTgs02ttYhQ3xq98wrVIdy3wNascvIbPau4tW37F+rMZZ0rm+U48C0xcpwqC86
mmcTA67efMYEDbS1xAKdqvjOxJDvsfgMppGexhOL5Ouy6b6jVgprqb+zLV++jd64
z/nqUI9D54T62nY1BTmZh7y7gYCJXKHzkJvWXDBlYWs1ZS1Y6I01R8vyoO7SHQZ7
PIZFEGCX4az/Mqmb6qDIdOi81vOlc/uS63awFHure/n/q/kzzgQRFxh0zei6Bm8H
i7In+NHbrQjYyszL7cNb061ObgiXRsVtj2Q48qc5PJOOcMca2qflZo+dyvEjnoz0
n9mo3aIFfCnL6A07QD1jpcnnD3lgmL2CmJ/bAN2UMINItfMACamF+jHQsWCA5zkQ
jbO4wJSkLBV63biELGDJdBKoGzF1QZjuEHbtlZW1JXeMlUSsrXOFIagmvcBjt2hg
4PLDrotANUn8OwO3MV7uRFnTkbpxaWS8TJsHATB5VFJl86T7SoRxqxK886jPN5Ut
DHbgkc2yYFgsbToBBckSJGJ+/8WtUjlRHt9i4Fp0GryO4Fn1XedAsy92eWZtxgVx
xlF0oWMVdY1bI+9Z7gf41SRlWh7PW3QX66g09t/5rz+Y8ODKDEwqi2sABaFCuYBJ
V+YT1ra/1gvJoxi6pxEU766Oors1nGhHRdWSaqgw5WMoc6F3bpmgtJ16ONMOFRGU
VlfDDa8Dr/QD37yIp9xjeUO9SdRjtL75GJ5nsRuhmYdeJtwVlO9+pg4JAPozFfUZ
HcPCzEDdz1wHzAEOVRWXnxILK/Jz1nM2CFI7ad9hVsPLYsbnGFohSuNtDdN6aKuR
s7xiterXVfxhBE0KRca5yX4cJkex2yB1g6K3JukNOcqcbd9SKnuE1Hfu7DcP42f1
jDraNkH/H1/1jpTDYsK4PtLgfzozp9Ctd3E0nZSaES+IxGR/wNeT6+BWt5iKfzki
KFkIFJwn8h6mrnyAxGfuzgyg7RJBIbkJm0uletBqUUfV1ys+Ma2Rb1W2AK42Kd/j
ljT/QEQxFEP6oJ8SzDgRevOchcMg+Uc6AKDsZ4q4XyxH/ELkIvcxJv/0U5lySgmb
4q5rOtSWvjbWDNANnY6SsM+6ZYUCuLjX+li5cAn2GdSne+bCuOogFTZjexRH27Nn
VPw++BBYacmP8qAE0zoHQeqAxG7ityhWV5+PE8rLNhCmzTvNrHJvPCei79bY0Wcp
NVKtsWfHqQDaPyIv5Te+lSHEXatREzOouDmswxGDVE4Q14T7r1+p7qu3tqhbX7//
c04Un17cqowmkhX7bgXBPjwxaVDUkdrIaVxp5/2F3a4BB5cvsvNPHnmatYJA5UpX
FP52kFIxvveKU6lzBHUw79YZmh7+pWFEpmTiIYYmydqYlfsRrKlpP5AXrXRS71KG
+FkFQ6pN8ebQkf8tHfl/AQG8WuAWcJINnux8JJSb7A2WXm8Wat290idMpUnwn3GJ
NerqV8MobWHg9UIxGSaa+r4RS3eYZvJjJBPvyeYdXEA8qR313Pc8T/sbmAozSutp
yUrKGN20d1VADNuOhNXJnkzGG09w6V1F04xJXm9DgFdt2FQ7Oxn8XPoKiYFT3oOd
Au85dzvARo0MRX7cA4iFhFMld3tQ+ue5rWLQOBKyy27U9ckhPoMKsOm0i1dbKdg0
sbQqaPGV7TBs5yTIgPiIs99nQmUSO11K6di8Ab5tqytpMnS+lwHqfu+OqRmKib1H
STCOYoWyl58FTcT+sAqbZQaTVuE7gUJHS/Idi6NtJBuAUQ1l6lM0dlHQG6iwfbMg
hg/XeJB65783xnk4gfj6lXx97j8L8WlO/T87hkcQBzYOxp+dA9E55/qBMyJpv/b6
47jwrjfeOfFqJGPwCgieQPpwF5pMprUkIxlhTMCcNBcB86Jqz/DxoDcIIwBFlw/P
G+bRHK3MkrmeeiVzPJIYnWW5idV7DUhZwQZuc3YYWpRn4c6bSCanxPV7yik5qWtx
9z7MU7ysRqgUH/r1tOdTcAxurlXF/FJe70EtL60d1LgdNyDimclUie2ZU+yPr2wJ
n0MLF4FZkpZoWg4OlwmbgVyLayA55N1c3s9V61ePdDGjDV3w8zBSXm5v9ll51i9r
IVgvk94tufBRzNkAFxzLhfRGYml+SHlnm6vCfW3ZzppM6eJFBJON2i19/JVTw4wc
68Pyvo8wlRip7bwgq4s0M7qIUzIEZl7w0CHnlSNIVMGqIZ2B277L02j2exetu1wJ
ZAzksY0axa8oa4SdchG8lvKk8SlOGyfKaiy0yqeB3cPldcdpwihKz23/Tah6s9ov
znX9H+ilaVmqywpt/ApjuEqHb6lMC/AUCSSQpBLNTI0Y0gfqc9143dA8ZGvidl9t
V5kPRvFPuaS6GCPtr+KsKo3rEEsET73rrjnHcYC/g5DKCkIVcI5K8EfSG87pWXH6
7/FcH/VwgcgDk4ndXRdZQdi9SBQB5DLttt/Ds91yDAjLMhuDJkhM80nTI6K9sBRN
83jx2Rdtp9hvQGoJ4ci730+yJux+iwYrX2fN2Xa03AHcphLuoh1yLaWgu0c3VwLA
Afb6dGIsRiv5LaMa9U/tsQ/Ec2lfFzE1wnzAlOhNhdk6Qz1RcUEPxYCwbYu/5pp/
rigV9qvk5Wm552nGcVDW5xwz5c5dTmZZFfwN3JxkzmPaY8tv8mRdKTAm7hwps/Mz
plka2wSPCMC6UkWOi1anLrZ3fL0sCUMgU+Vu2k/2DVKmaBNDT9ZYEhGP++M/O2yN
rTkZykIG9IaQqM9WY6/x1LyJcWP2gH3e8BX/8pZbtLgnMjIxfT5vR6iZyF/88rxe
UtsHyax95PawOuo/qYrI4xIQesKDkSQeCQJi5if1o1sYz3Sgvs7gjEKMgHAcnf9d
jCPwc7BKJiT9o+RpxwgSgRZI0E/jpEc6RQrQ0MA/olDNzrAH2Qos42idu17PRs+h
TJHj4Qtdqol8MQcpQSFBM+QBhA/ijIY9WPAP6AO4O6FGNu5Ky66FU8F0RSRSfOpG
nK0k9a7R3K8uZfOCTa0sTSbWb+sYYS6pAg/fhQDYAQiXO747v04CWK5kKlUb7YOI
4/uHb7gnAsfCXwKVl/10Udp/BRy1SiYvOi8eeoGocqQa9Li0h7RGAuED5ZwF+VRb
iRmlcyq1TegYsvydophudGWjEdTHxg7U4++ovQi0L9+opYpU7uLgnrkHm6zhZ2AM
jtZPlaVbfyj4kLv8PL65LZhJ2U6pUlpMA7guMhehiNvUJc9yJZNQPunRybXGBIBX
ObzEEyKMSeyB+cnc/7Jz2ScSiq3m+YJ8rUdJ13GUQKCQciV6InbkVxdR5EMpESID
q57osCLEoOU1MZvbItDUvkDwepmWlsIhQm+Hyi4DUtG0dRG6vZUFH7nuYciEkXeN
w1RqgXWOTEQnOP+rOuClK5JE7fuw6OnDBAydWRgAbSjhq1kjFP2C7AYB8OQ/4PMw
fHDrTuIMrYtZX1dkD50pjSFezwjVzfenxWz31Pkr0apwcbX8FlnjE/obwPaDzOQp
7fwWuu1+07oVFAunDjmzuZrYNVg8ynrWAuDv31bxk3aMZx5rJPh5ARUaNyRQYJuZ
5tdTbKXbXdZ3QTyx/7lVKWmr4ujQYIPDeAbfQQMaR2pLlIe6bjJEj3Yiu9ls1ayX
4uCPFzdcIwy8090G7ca2Uaj4FP3nSxbbTB7ZRiywMepTTac6k866UkwJ4td/5l3T
NeNH7in87PJeQ5d/zp8V746ItH04hVdvygonlmwqH5Mg5xwpVRNqzrvks4vtwbL5
TP3A2WhVcFzfTYhufgBhyVLz/kZ+nNNVbu4r65Aa7GxvpB1aXeqA1MguUJUfR8bM
gHYIdIqqer78+K5gwK2+b2cRV0MndzARWekL3xzw9/PAx7Ahk28zAZRPZBXatzgD
51TCG8NLDrOr9Qa49/LIOp7Le9X3uInk+PuDvMYCi7gAYY8CXTijSbD+NeMPNMcn
bvCNHWjlfwQPYXDhu5PjGV6zdPfp2Wrw/tCLBno52xJDINC0bhWcHehfG/ud6JOA
4eMZ5usLlLY549rxtiQypNUGtvL+p4iUDVmlvWzVntSASBg54a5p2jNoBIFlu8bY
Lq9vwCFXIH0Wz3fI27nOMs1o3V4QgXE6T5NhXX43/zvtXKK0mIYjqTJWdguAsYdN
imDPTRO58YTU+PODqib01oBl1Xz+1jFp18lnIbYVp/iSX4Gog4Kwzc5xOR+0hpvt
xg/zX3XI7Y8PUKwJ+vKrC882qPhgn/yQJ7YjW4xR9j7CGNyALaIALyXr5yxjk62u
sBsKoBDfKqaDekPVgNOqHLUfJzCSxQeu7B2CXBU3Z1/uBwv/DGJ5MoX5R6RlYN06
3LbtnoHQWgvnjxU856lFRbihmmYFmKCkLhURytpRGIoFXCecvC3pi6m/8AbBD2wz
pqDHc6ichLmyBrsFnzKr24oq82G6m50Bt9FJXnqp2PcVAZUDNEGarmoqT/pC6R+e
yhtnBMxBogXl2+bSLHlZqkCY0rC5xuah3hU0WkjEsfpj6SCgpLwnE0apcZ5V8/ED
7HkkHTHjjN8vezuFwifA0u2sNpNNvU1hJEkE8JPO1p4aq91Cuxt09uNIc1eMp+va
FwH3H7oyNWg9Us8vkGFjRIF/PEyAf0vvIHU3pmhI16R/RfS2+GSzsvGugywn1+6m
vx9Wr12sF9TuZCuvvo2aQT77+rVHH9VCLwBGryIdd2i7zD4POGaeZUx+/tQ3FPyi
WS8ZurlWbGP+voYKEIM+TL3kT5cjoRKg6Es5cpOvFr8UVZpCqVGXx8nvXhCejLQG
NVBp/+6g8i9IPCZIbK/bD5eLk584p5FSOtceoIqd/ArYtsP9Kfbr3wsMhqxUrHBt
U47hSlCWuqL7CoAaYk2P+lSndb9SHm4+8bnKJlyFT+3tpwa/7GzDcV7PgOzFTs1z
rYey/sa+6jUhz+k/DXjywhNyweB+UUhU97kkAhhJH/lpnmkO37tP1gz2Q3Gp/3Is
S+Ugry7v+VjKlNvCaMKjzuk8wTu7mMJTG6B8Ho89z06iZ3b1tRMs2sV/sHw7Aa+y
sYtInRamSCYGCajtbmCMV2MuHrhDEvD8rY+yjut/t7qjBJlDr8HrqclzF8Xq8n6q
Z00tjZ8mcHjzTXSyjHCDe9xudP+y0xo0AOOa3EBVyAY66QUaMpNbbKziErhz9AHz
gjD781gCcd1wooscjhAdT4oARiaRjp2Y9OLMLgfxPhSogkhDWYSVQTz7b05R8V/O
4AKx+pPIvttsV6b1r0IGsrIZpTOojb8FsyVAZCyzGb+CjbGm3OWjkD43ZhAA7VPh
IoxSlqq+p5finh7J0I7QvBXCQsHfQtPjqi8AJUlclJglqzwNjToy4Tb0wXixrC/3
fPXqIJwZ1X2VZ2auDVR+Ogyzu4mKfZvIVU/ne3zKaCQ5iUxqVlM+JkkD8IqBNUGh
C0SpOi8Yk7A+3R5Qnrmnwv6CuJrUncyZ3mEiFnaEDWtfX2SX+zwEJkPfOTgFcNLk
tuxjA65ltqVqsm5kQQTKtn4SR84PeEpAwAbL3sVn+BsEAtqPN3T9XYchfnvm2Nh2
veLkYwFb2Jg4wNbhPSUviLgglGTLVhc4zbPDSEJc9cFh/71l67qYS0NlrbXGryKb
sqj5sPT6OvSFt2+4SXC3FFudVGavYC9riHrTXBJEVE3T84Xktt8nH1uJwcwiJa8I
hcIyyatQnaT4xoSUeZxLXgnep4Ky+sSW2BCDQJBmPAxPSwA4h93HF4dudOmGOYj8
YpqHFxNTgkyQGZIRAH6OK/qsC2k+lelZ54WWIdjn0pxpCBPhpqU+d8+/O9tRD7EU
iZGxxBRuQCmaVy8VAnYZsa1KwCN9gVB9JYZAgNCHstCdHetNWjIj6PWnsPMQEX0C
EyKnVwzPPHCHb3Onk5NKstcaZpccQ1ZbwATmakTdxsnoQLL2JPLOYzvzdkkVhyq1
nVz5r+1BajzMqSS8JGyIJl3DAIkd675QZnkhw6S0mmHRbEk5+gyFkfYWxCwyxyK/
LUYuPC71jxYsLeo+W24ICHxkClV3v26c6wyL9OPwdqT9EMxLOZbyuzLP8AlnZGd/
oiovdQmPvCYvEviRg6CG+o/GYtc+sr/7rQlwRmxtzzDEHEsLJ7f4Nhh/EmVeFM5y
QATzKPgz+Td00iuLYkcylCNfvnEOiD5zX4RgBXEIn5ZiVFmdvzNuYu0BvDE7NzN8
BWfftPK9g71dV5EM72Q/JMnqqOi3f2oXBNy49V/W5rFXHqlfg3LnSlkHiKI0Z8TP
ifLIeKtbPTDcz8GAXQO4utWfcySC4f6VrUnGfR3zjjOTpepoyvIVI5SB5hrNyA8p
/+AQgmudlziovYDssbkYDGJjvtT6IVt5f3lDIdXDtpBFil0bnfecWVRC7NS8pUnr
afHI3WSqC11IWFBzV/2epBMbLpJXfL/eDf1TNdlag9Ru0z2/RZOOszINmx40fSPD
/9+Ej5w/7sWAnqsCFl6GiHodQq6dTqWvHF/3C4783dn3YIHPjs6WXxc4A3XLOhpH
I0UtQqnV6tNf6n2g13lcCEcG3WcQfBG79rwwpfqUuJv/Dx1CQuso3X2TaixaTRJN
41Mj+L7csJQkvWVVl4TnnWTSDQgPCvFuEvQcEDLXE+mH+qLFc89DNLAi/Ko4yI2d
MIHaHBWtTPHjrq04408s9/I1/QkC9tYq4lnJHAJ8eZ0oE2FKTaEToOLOn7oJUr3n
Yu1y+egnyN+/UbY2kYXI1zWayirzrRzPtHhkqRJPldwqYcl0EDBp1pK+LLcWqVld
izE/hmYsXsr2I+5lGcbNw45Pce0/NsXufn35hxBBcabnRF4nfvfZg0PROgrwzXbs
qSIawggQDh5SCtRAzZRHiBENM/GWyck49gqkLj3vrNUjJRiSZBxlLylYZUN7nO+v
4avnkDP1WOzfvDOmMsYEGF6jWaSGQy9oYaPrYdbaquy6Zk+y8YN5Y9sTVL/096h2
WVDXtBB2wJNmXOq1o+vLcX9ZyUHi7b7xNg/VrCU6rTQZs28vDrq6iOQmUaeOQoyu
QjZIybfuHLb8Xfv7JocPB7hKJsHikT2VrAgs7jceHCYopZlk0TOxKNzRAntCwfYQ
jLsiFu+xwCqgb9GM/FkHZQl7J4mcoko5/bgtDWv8lz5wZ429cMLcJxJAlP76RZu0
AsfLHobd7Aoq2MEKCl2yb/kyS4u5u4F+f6k60gQCfBNVXf5OqX4C7V2KsUqCivKu
vNFUGAUUTTpTficzzloToy5T9or7C/GZziTk/+TZhA89ho9yEDIlI5Ph0q5VqolK
ga80Ke/DALldkDCgNsQB2WNvcQEBP0V/JxTBATKaUYdKlR4jLt9GVRLZmnCH/itP
VOH8KKtQBW7nCJqNoko7V8GCMTuT3Rf5aBDsUU6j/6ifbn1bZH4dJcgyOx9rTcu9
qZBxy0DSuYmZlL9PF5/n2jmaRt0ZzHdZ9L4lsRfMaZWsFMJtKSxWZUbs0CAFHRno
SalAOezuE5lkqOC1k58VGs5bk/C3yDhB5PaiPKCZ1Pjo8wo6lOy24dJbLlxH17DS
0q0tBcff7rXMmB41Qn+IvxFAQcXbBwcZbaGm05WTKN7XnGh59vuwPDN7T6hd4gPY
nfldaL+9Gzik/8D+GrE1W/Rmb0JvC+ku4SQ0LYApcPM+5O6N9kIFuaIOS08ka5vB
W3sSdByh5wiM3NfYOkHqUxZD7Vus0wchOQ+TDW9Hek038a/X+H+urLhVY8T2NvVt
2d+EPYqUw/z43VlXHZ2u4TqZKxSAQB1e/M8pEE1/9YRC5Q7ZnuV+irhwNLBr3Oln
EKcEB4VvfiNQGtkW+S2KI1+VjBO6JyLv8HPlKI5qOPIZsphFtU2w/jb08RDWOub/
38mUB0MCiMUKE3d7NJ/vt9mcQh2A79G1/Obbc4UoZ0Cc6Qd3dL1b40/q2OcKyeUk
VCygMJdultUkMW4rUo4vYjTyynrUypD452wapPOppr50pzvvEYRDp2JQCMKqfWZn
pJ5AOben+fq2l+WMhkF7EAnaQSVfHITArrDa3S9ArLIL5Wv1ooBLrpEb7T5LHdDj
V1d3aqaI1qfBuX49iX7s1OodeSEBQEm+20HOPFIzUowvU2ANweMYivgWZyh081lG
AH/ZJyvxzC5Bv5djmLIgNQvk3Bk6Yza91GA4Jd6mjVhDs+W/GMXvLkdjiCN7RLf/
Knqfy3nHmvUqI6+2JbvxLqB+X3cB3G0MMEVIzZdLREbEf/0pDLeEE08QCJzdplWx
TOr50uic86Rm3Qz1fyX+EHiD2bOyUFAeldo0wV6zBTg9lQGxLlNXcB1xxnrzRrh7
fKTJzxdE28Lxncy/4hjjpfbyJGqD2+anQVVOJzhWdgz2zUF+fRCdN6MozZfkRJQJ
BvAeOoyprHPxzTG/1GZoddmzXJLNJvnP6+pQTta+TTwnnTIkD6M2q2jhrMSMfSaQ
KTVDM6hkbL6blKyOhGW64oOTX2GnUWZwAhsaNf5dT6ehm6ZhF5A5BCDJQ36I8z5i
aFKC2LmhHJ7TI2eGJAtaYmen+1LRg/Exg8md9DGkEUcwA7beY+S8vPOXwPHpNy2+
gfD0Dd6/0xmq6yVzcw97ITn4Woi6NgcBbDM3e8Sqe95NRRuDNr8kWDDLMwvY2sy/
zy0eJzocDZWqEK+Ki3eMEZYjGJnM9LlZA1W6jU3wTdK2HCeUjbyu0KPNm8Wbmkbo
4EbxQ9weEnKco7Zks6GMVlkJtw0A2n0FROjTBP1syoSJCb4qosADuAbM3845iosE
2V7B0fdbLYt1Mun/MuxGF4AP0qVlTyU5P2LdRrbBi9eZDKOTwoxqtqgsn7ZefDve
a9Vkb7ED+ho5fdwCgUZ6Kf5e1bJpomieQZbUsa3VFy2oAvVcl/WQli+JlUFV8t/g
W5STCSPcOyGzcXQycCvM+ZgM0YEuQnzzLlR98is8BpwIVGDU1HAaXCr6B8b9b7cR
U1Wwoj5QkDeBKY/ipIlL9q1BdRfR7hMof9hkQ3DMPD4klzE7n2ffaF3WRodOJ/ZP
t8j2R03djm0XkIasr3Nb5BEW9Roo/QX5O+2AmmLO7wnaGQyvAjSHzr+BhrgznY2X
a0XVaxAXSI6lcJmrzQNhMVj3aUynsFDSCXnWdSbGhDqS04LfO6W6KXaN5DHUBjB+
xrz73QfFc51g843wXn7Rrd2EBYzugYci2Rqjnj/thl3stVHIfZCgoLfkKdDH4oeO
h40sQGmu+wMh99o5gr1jZeNCvvyAcpWzzOvEFYgq/N1efz35tfLCUhdYKIJJYWTU
q5md7bfe1OehCayveUF9ctDxCnZQh0AIwZyhb7UBwGzX1NzPpae1NPBjmw0uGIYS
Ca0MaK7wpZvpQ362+1mZzZk8eO3aHofikacr10t+SqqNAqeEAJ7wG1nvTEpQ/ohx
j5IWYmj5FxU4hYm7p/XTLMy2xvDWuUdSHNQuHZRRJ1DkeVcu6TKPOxtu40GfhLVi
wFfVEQH3irRaQkBNUoF1dPBHt51cM4Frg00KEkb6cQljF+JTsOPcBh/5I0vBmExS
M8XElGKxkdqJkj/DYZ52xa/OqAiUjoh4eTXWvz0coG4mNzxSW3VYqZ8B2PhJVAtj
n7qDVhOkYsNbcq2AF8crrbTKxLPcNWSM8/PK3st0doUSl+XO0/ysxLcLVn/nuAWr
Q50bu8/Dxanxvl0shMzFBK8JYAnN37+XVXYlZgLmRKiXFk084BHeTolV6uQ3jHqW
wAPppzuYyKZEv5G0oOpBxoh402522LGzpkjcTieahvgX5Ebp6UW8V7tXxhVnph+z
h8o0ocwA/yOGIEyEqyJxuX+F7nqYMFOJ11R6RSjASpAeyIp2BT8xztEHctPvJDNG
fkPJaPT7wRCipYcXqLTPRfwl+dYBLholAQ2GLznxl8YMiKZ/AlfaxYTzNwTXNZqy
//Kr5AgBxkEc/kO/dGgW+v+OlsO++N7ppMvXYJLjHYG7qRLFzIU4d4RJKkihLyWB
UXEkNsT3aqSteLsPW7d2V/kV+dvDGn2AkhBpTf+V6aWNFFVc4lGpGD470IFICpFa
8zPujxeqkSYgbnJtmmsQw2TrKx4I3GOfsDNr5dLsn3qmEc/PYQSflm9k7CqZdRiL
wuEM0Yi6M2j8lu/ubFUHR93QdSe3rYE6YSqg7k7CAEau76SHb/p+TMBVVrxhDFb6
jF86j/GHxfYidMiQ1lD6eD/alpotZmM0LcSOQzxjCz7+Dr4JF+hszjJAv44pbVov
un7be+j5cxC34YY6jRhawLQPdqd1IJ662eN/W2cp2vpuVgDEkyCliwOfFVlqbAeP
SaQZ7LqpQvtj82BAWKU8EKrYyyDB2QX991LUk68qiYjC/wIoMRMVjMdEQnoSgn7i
Vw0uMpo9A7IXjIrRfJpRMoSE5REc0OBUobA1ubtnieQhu0ZpC4zToFQb0RE81xmR
WFRl2fxG6j03/oPp0ymnfz/0fPR8LwKqWxzHjmeTT9qMawAbix8bMcpldVGoXkth
T/bwmy8SRX/KX6choet2msmBvYDYySAfeEAf6gmYwi+ceNNwvlt0IaprRLDj1pPu
DI/nUI1QB0rrWcx7Fv8TWLTKqdVtiZiRJyyk1zs1Z9me4i7uYIHMx7KU84S1ph/V
SkuB38Lvz5tRYXcY0LOOP6oUUZePP5ZMLALc3xfS0/oq/G6Q/xEVpuLx806P/+4c
BI2/9+tPG95VnpRnkLPgy+VimlEuH+5VNe/z5RJbDQayjVF4BUMy5so0ayDuMumB
Unabi/VQeRpx4yYZMOhQdsq1aa1I1KADJwCa6GdVTOAtmrmI0SH95BsTNCwu1Hjl
ciwSg+EWwl9fWTkZFSmUg1UvT6KjksyQ0r8Zyuj1q1koYcA7y7wBvpwwMo3v+igR
9bHsIJOSaCmpiHDpEVcnh+VjPVOjmDIeDdjJvZZu80Rn5NkVq6nkxasyhc/ABe21
Nd8fODx0i2rPJxwQzW9mo/wsN6/CpyNimbA6vh5uqRH7V/XC+IEMN+rkI0X0aWD8
GkT3nJDLA0FN8fOY5iy+m3ahZl4uBek1C7oGexq5V9+dllXYBHyr/fy9hXV69iBl
LBg1vRfJ53WasIXGsNu66EW75mBSgsRah0u9PlK3LMuOdYe9gDfeKsL06egnFQgB
w2Dm+S1OrTXKGTXqCAQ/GDzS9izpzbCOu6KMm5h37BC5GfIV7qTIrywkIZhW4M/Q
76v224p3ev0YIeiDxAOg+/k86Ywt+PdxhWefzw+KgrdtE/xPZJWNT8gc+pwpkXiJ
Gq+dzcRYLInoea6Wi237hxCs2f07y30eb4DSaKXglgiaizQBv3gDhAH2lUxAeS0S
AMzn1+zLX0i9mXJB2C50gK/MQH+Z2zv8YpRPdq07fSrv8yE51Db1dA37buTEslIS
171po4CGjUhA5Ns0HZyNM8f9t5sRVloNIRAheU8cBfJ+ONp8twuDABpJYpm2l57h
+13wZNXWyQY8iy+dR2vnmTcY7i4uvf+Mh2t9aLYuExUdDDTJWRqX++Yl/8YGs4R+
TSUYaZRZjDQhQmTQCdTzJw+wFUPhWVevQh5auattlTfpmbeFAmXjTa/L1DHDETvv
VysQ38AcNjNfyILRbQsbjRD35rltaTt3aAlu+3SsY3go5zrXm94N0hk9u7mA1B2j
Y9tlrbe7W/twBfKSOO7xpzRienBoY1TzTZM03l96DkD8NgXtGrg67sEcbWAudoTZ
bYbUgvhP9Xu6OWBfcC88tVBd1qdJA6DUK3KIShnbEB/mIGR8tM1GiN9ZK7mhbIrg
Of7vXBwlV/ynU9TZQM+OtSZzA0vrwXzBh6EXf+ZXCQ/dJxxwlDIpLHIsH8eWCSqq
URgZ054y2butoYsc0eSWMBsx43PA6QOJV+b9xHxAk2j6VJ9w0snXsILMY13vAHSr
SM442XAJJ1LcdizZR2q3OxNJ4eQ4qi1VNGufTGYhGG+uWiAobvzqlBwyvuIQriKh
JvnGtV9c5FV/3c5BFm/0+WzIZLwjlVQrueQpKHAYHLEPY4FjlY0v1OF1hXG7O6Wo
UoWycHyIWA8WHVkRF3lEuGzA68J7YULSQOSZmNxRyFepmvFY0DkjYLiJ/7FIsoZX
hTxtN7K+ZCBCRnRwHyNcFqSLB4yOIbvN0rvaBjo32a+omkM/TsGSn8HTyNgzAzwy
MkSN8ekVr7Gde0vHzmr0hUgX1XBP0S6GdKxaPQ2fsyWGiKumqHqyZ8LtkOTcW98C
W46JtKDw1yDCMUaiRio7NdVOTzS3ZlXZpO8cUGj/Sx7vbxUknSf0YbtmPM8pDZlx
nGsF7KtPsdgJhaocB9ZBY2JLV8Kaa4aJH4l7fmQ0+dL0jPVFMYG4IRNqAEVmT4BA
YytcLwn10Rewfck+ycj7VSndich1LAfHtIOMl16qqA2ouYlGo99vPEog8RaY79Bc
00yLFX0d4bDG0rf++xDL3UMFvCEL9NBdSSS5gDjjAFwNuvYNJ/RuScJ904gPYof3
aZXCLKq8GZU2BQv9HOsWoCxZB6aiwx4941SzzV83BA+nEAVYr5zId/QX9z5NF5/I
AlfhMke9RHLFn+XMMDdXRLiUEdodnz3o4S25DYo+I8T0SGoleVPG7DtaHrjUXlVg
1CC+JSoBnFFSXUDlG3k+m+2JlY9ISL4xNfHKX3Thh8A+jZD4OggTHELGhcbhAkzM
gOIv67xVDccBYrxtFX+AUAlpJkOp2nj1HXfoyZJ22lbZD6MRqzEimJrm39bqwQ8Z
8b2ryMHC3+GjXMsBKz+Vxe2rGKcL+Cbkpu9X9vkeoJQY2/EBIdw9OIemIycbqZQP
Bv3AdLQAK4pZ35hcSVEwTVC8efN+1AhhzMlBowBbULn9LaXGYqDhh70PCtJATOVu
W+LOFTSxxKkvzxXrM2WDF2xXGouQ/ftBZFYbaiFXMfQmM3bDY9YlcOyJAhkY3zcR
8AG8/hhG+VZjXzasw/5xxQD2oJQhGW+zIM/bCuR7Rqj+o85VNd3lars90OyBk0CU
9QKYt0qhhiy5+qyHDk9SmBV67G6aAiRffdoPEHZGor5wvuZHhNotevKaDbLijA3O
9lTe65GyQ8QeAweCt0OCIzgXFcGONRP11wQPbO0TkKUDOk2VYVJyWj0VShcAjKCD
axtb51sFnoNNBmd8lqTWOKYvOuGTWw41UDlB0Q+LL7X5sRnM6WU5WmNGdjdUps1c
Xr3iwq5cIlYRX/biZJc9IYI1icRVdUJc0rB+BdQmVuBsQ1JARWbqWsorBDHGIaIW
ngOab8xR6cpNQmQs7HyDT4b7fWMNMjO72fD0x9ohw7jF4EOsiutq6c0erdGs+wMj
hXuVqCCSkncwkQQYFJ1oaj/s+QoLEK5swH4YWsDM8Vm/UDuid7sZF1aCqsws9ofm
1QHV4Pj/Lk+GA2DwVa+pGr+n1carhqDP3UDSs1M19QiXL81oPpM6NVDRxDvOUZKl
EmXinKIxtwZJ2u6yn4jXxtv5//3eOe8nLU/gVBzVmrTpy0UbxrR+G4fp8wtHlMop
S5s06o23e8nvvFHo3+QrgPK8xo7YaWQMUUUNJxhSO+egdAl4gFhxx8J4u/gEmuR2
dx31VgPbEz44CcUdGlARPjdtSN0SUaFlBDKCIfnOYBMD4wNSgO9Ca1xHqkTf6DSY
t3KC8f9/dMlVp88FppQJcOFs9z99wMEvbD0NrcnbRvqPDNU4yD7d3DlegMCvStft
Ut3U8i2LAJrMpT7fZNJF6U/wxW6gLuLKoEJxs9sUKIxxS5Iy2vYQgnwmrBS/mjqM
zxGNe24HCTxpcPAVLkafu0PYnBS01gZGD7+XHeQ5A+MVBs0IOc3ODJXhTHlk5LqE
ZUN7HRA/U2/+hT/k8BqAy2tG8no4VI8JeAR3yGyeB8LXUwHJVrRoQxWQjBMhU/x8
EV4oXo34TpWExaUm1xdmVItiTi2rjCBx74g/9wjwUSYQd9RRrhOPamWQu041s+ua
Cyv1k9HpVQF3XwCp848gIi/nwD2mFc7Lb5nqmyd5FX9pfqqjW1Ye84oG0MzwwURD
Lht1DcEkoRgvvgGrlgNj8SADTO2mYTJQcbhLdNfeqv1XXFC1sw7dA9wS7erZOasf
xYJfSN1r0YnaKyjkOJcZ+TEnKeX3YgMHf6XxQX9TQ2PWYtl8Sb+A7Ce8FQL9COge
eYiTf0QhtgTTUv2X0yZ7D1wzkFpgtVDqzM3IxdcH/k7GLPniQEFJXG6s/K+WkAdD
bam7YpfLJg2gWj6r/Vg/yLyFeAp8mteFgHl3nUfZaBrBESZr43GQO4RqB4AeWZzN
SqHq3JuyC2kyFjuM8IHezAvEppE0/Y+JSTQe/qd4BWrozLQ1Af+ZhHK9vNlGF/2N
ERVGlv6APDti6Kn/ReEWONadhqVJ8vzcFSd+nrQJCsjjiX3DTfdHMSpO1e2Ru1Dd
bkXYrlngM3L8YuN7fdkZdNqrNaVeDdrGB/KOScuLBU5beZu1+ETf00cNcbE61/xn
epC9Nn44SUpzQqmXriRLw8aKMJg23S7jgjWXhmy/viiLMho+Tir2CTRTwt0Gjozo
r5rDDiDqiCeys+YFR0jEfrFiUG/PPW+MUwrttrCZZPjc5rW2nKBviOpD1adQP8CO
JbORHWKk1QKhN2MC+lV4S8X5/bAwJ2RhzTg6pbZ+uApLrXsDB8Zf0COriusEOD8l
C/Gb3HPjpJeqBd7FEsie+D0wEPeh6jk58KKit0c4IcloBaBXfo3OAAinWRt+UxWM
6EN8oef3f9AduY+lyc+qGc3eXeK7+hZyonezlZjzVrmp+w1n150/iRj0UsOO1CHE
WUtHhCRZCaqtl3yYTWzlSdc18GOS9TchfXCc9PL9cmWDYAFbtcoOeqDNm0U588xw
gMb9ysL6W4F9470abmtxWvO1hAls4DXh4BIOVFBFwI0aKK/9pEmz10A7tHE2mCpu
7dPkVLqznGEiHeBOwDH4J8JrmO76e+tiFrTrj5zAOo/2oBGR/o32fuBOEt8KDlnw
vBMzxMxZGyOvGGcca3cal2ZmPy++e619B24OtYJfhWW+D2Co8hHyCbcg0H0qDO7M
M0ywz7Z7p3kiYmwfY7rU4O6ix+WbdpQ47X8g318B1Sv/HUJADORd/PurmwmWJUW3
4gFb2H/7vVZiSocf4IpDg49ThGf+aFXZuRLJREXFIbflYjzWSnyrxwUche/xT4Wu
GeWQYcILrfL74ZWWAfwgeu1XIGt6NVxEsptP7h5wf2MddLNB7pFzpn9uHfZgg0lK
iqpDniQ1Ezu8X5LgTpUHDAmpKSr1m0KqwPrF4FX2OcJgNwDw/Tkr+Cb1JTlyBWXg
KnqwgTZeA/C2MFmsJX+a/15B5/goHPkzzFKO/B0J84DHp14VsZ0NDk1p/Tmhe+Uy
Y+ze9TVS2UoyvYJTz3qX4lt0XmANt2FA6DDAZQkT7jQ7jjpsizZV/n9AqKiyc0+g
RjC30w5NohVqQdW0B+GdKV2JHR9kTJfVD62l01Pof6DdGyBdcw/rhV0l5+JdW1VJ
/3aJgo7vuVHRU1Ww70ULhlLYxkvZAQG32G+PmocJaQaQH0jjxPI9O7QFNxa1Zpou
O97xWpfXZq4/zQj6bihPKYgQar/McFq25pmYCtmN1C8HQi/5nkg0misvkvDyl5cx
5pgcrK/9oPA6qm2dreQoZMtGR3apjArT+XwkgZNhFi5lSGkNgmTT6Ts24NkrgfGu
mbYo6qdmVb453C5z7oVkNXZTq/vOrLGTFx6qknNKBejliHbMNlW43h63dxWvA/oD
jXM7BYSXwQx9KTN+4gz2bFdnKZV49e20SczwzNLJReGDW4O+1LXbEE0v4wWw/Rpw
FY/lAPj4saJAKgaRRc9BcHFEqPnUJb2FF3GikI5qmUe7nw+o9urlTjUIsl3w9MoG
Ub24b+5un56Nk9p/llpWT7KfZ3ySkZ4m+h6eLpe7aEUhVEJXA1i42fqNYDd6YCu+
hsOFgK2lKAqevH3qcbFH3Gd+pF9PttGnA5N8nf3fAoPtv+Dr6yK7QwWXQcVOcIGE
Ih4KRajpCMeUAOu6KFGGNOOdooTArPY/3a+CPJ2Cdizcpf+wHe9PrYCC2e4VjsWX
GmyCMlkVqPHtgkLOhmWvc03buwXt1Kw05YFq41+fjCP/2ijCXHbEH7Qy2yq8CtGW
s3sMEj1XaWeEKfyTWaJO5rjsvNYl+lCGuBtJ0twTwSwa2HLbwj50fOHph6RtWQxi
29d11vfxKuQ5pNN8UQtJtL60mZG9KabRyi3svZiQPuDPF2DNPco0nEq7/tpN3/fH
HUrOE4+BR3v2uzUAEf11lqrnZgKQgTsKgqjSuNtUi5pLz7ULf5UsnlWJpzZVp/CW
sgihp141w0arKjvPzVN85rkOVG4mbvI1KXCabjVnbZMMF3Cm3AevgfDOZcmYAWEI
d3XmgskShRbvxQae7qiRNk2Tm5LnKU2zkBpzZRCvm/jQFRGX0mHYsnS2i7zYI17T
o8v0rWrJnSWvpnly69G6YPO+yAo7HMEzrjJZUcdm9kTq8Sn4HoAXIUvUb0JppP4z
dlxI4vXKwaWDE5ionrm8Whe+uYn+T50z+3usri14qzh+2nCoi69vykAWupNhvpCT
TyzSqnSMZf5jk+Vf112vWkNIrJl9h/VkqAeD3IssilvumivDd13DUvDZtsbnKLrf
HNA282/dkQj86allemcuO4DtIGxQxQeHXmC5P7emhj7LB4S9rDFeCNoITAl/6cCU
U7qnm4c4/LOpYY1lDACZlpL+TfwzKTBSSOGiur7UTQxmEOeKHtOP/cz9b2LL4QK5
bSQSJj0gnmJCTMJ56KMiqJlQaO+Nt4XqTmW4tz5+32Fw9KK33oYofX5y11kftcyj
pCoeZILEi2cevTOWaTDzeiJXSpcBb/1klAy24eqrTt+tZQ7Yg3K/0QtmlfGysyKo
DtxGWdKRj2DReYGdnjrgv5jbTI68aXMKnQ4z6Ki8LxiA/nrQ/KFZR4tB8IcENZtc
s9jG36ctH9ezXOyzx52iK/2P5IT6g8E5Kmk1pRxacJyCLELYUE7qaIe7bYJm1ICE
MCrVMK1iDD995oh7QDwJzNle/9mfwKFyroQEtuQbmPam6pl8VRE5JF2pmgvrCDu8
8ducRkHa1nEqRPGXsyKTFdR/P17rA0ErO4cuvmPr4gBoH/8KJpZuaS876youusHB
Ghs7QJOt8Mr7kdr+uCCq++davGC4ZxDRKwRJvQZ+yh2m8wsrm6BcHORyoQYEvcsA
15ULXBBGmQZlgkuDRupmf7FwOJb4LqEF1imUFGPJ26oMHBFefieVXzvt/ep0RRdY
Pjp67c3iCcTd47xqPsIHFLdZizIuZ1KEVVnRgaZVAT689CnjUdFl/TRyg/u8iCFR
PQG8chKa8cPAvIFx0sHXYB0Eto7z8DDpsVWW2aluKItKlVJcSZdEWMXv2RLA4FN2
MQf4VXMgeTuHxB/nwIFQ3nzHL48g27hMPweVb944lKz5Ad74l69sr9J+0RYkSeLx
1jjFOjGmVlURP8fHUDUlRsPDwtiCqpZO80DUyEaWPilbieWcDDi5ggivAmJYvo02
V7d5IX+hYswBhqndVn3TnW2kFjlwFOaPMCqbu2Vk7vFr10nH6dTfDwy6/JY67zlc
3HetHYFq1jFuAOFS6JVkO0a3LL65an7ibSCvBMdFinUvIar+Fajw50l50RvlnSQa
OYFvYWoakQzL5N84Ae177Mi/oyb4r335xYFp8qMHhE7GBrS3csdks+UPY33nk7jw
95Wl1VjWSYNJZujXvvp4yOKWHj72j2P6PlisD8/8J3N29c7LtBPU0OeAVLfLs8a6
5QXY871ci1AQUSxdh4FIib0b5NjJAl4+8TJkjQ1avq5sKJW5XaTAPXFh87ZUJOqt
5yQ+wCzycvAMipwMUYeyuLnlRdUeon29zLauMShei2HNrYx2jXZz0sJON6leEvXJ
3Fe24XJwmk2YzPKNP6QRVjy4f3Qo7jnUDB5VkDpImCVUIafLS70KUbE1sAoEDQHH
AG/DBkbpGOQAsp2WjiUM856NqZXEtgjWICxcxLTjEn16IW09MU8TLraf89vEAeRX
HfuvlJ+Vu9t0upD8jAzO95G/TetKNP+dCOwB/imDVKWnsIv49z8+W91f73bDm67g
IbffQ4X+Sm135tlxJ21rns/+NCSLGVR2Bfa5NTWspF2i3SEtmz5MU8PG2+BOTaUK
TRuUyQlRvfmHF2xc2btuaD9ZV5ZFlgPO1nVLIsjXiFLlPUHhjyuCm/k0nkShEzjy
vQS3Q+Rpz0gzfGIEwA9qg7Tgvh/hahAexGpJfPMFm+kre1KrwgBiDO6LQNnsukZL
7sYye3uNK6NhgUEfZ3KoeCUsmCfwV3XpnRyQjYlE8s7GObg9ox/j+kZb9mUnvSYm
MBBTTG3mar2i+48IIds5HVLabgGHlCu/30UwDtQonk20e0lBpsUjCdwm1dD7kRSM
/rcd8eX3wkRR3w62fcdcy1y8Nys41K5g7NcChdezYGYiB9tSwt5PK7ZVajIjPnwN
Vi7VR9g/I9vFvZwroHMEwTJuusN1nTeS36o9gric5CKvBhbJ9/Qt/tRVSi8mmcBy
+1ireV7hJT+6UVTHF9PIMoQYTZ+jjuGnkgVbilomSNGuyE3kmvpI4y+ZHWm4Kh2s
8dNZVHStlBNgv9hD1dIwu+Sqp8Qm7RFflVANIaOIRtcBkycIuDbnsRlB/UEn+QM3
JsHOCzJh6lr/DO6s8uHA+r9uG3D68iPZUHXVk7tUoL2s14PwhbrqfBfld4lTdqaq
ABQmTPR+cCEFRHmi85VdmhLdnMKmcGH6q8UHW/sy8s80po80mCkYMkjSwedYlXCz
/o3s/ZVScFUrFef+fZOs4BiQ7Scd6Mzu/s7b3e0x3RpQ9KJWqUuLBBdGHDlYcsVw
gezKDDOWhAriVUkTWzec844MstDbLuC6J1B8Q1+4ItzrtW6q/3ZSWzXQfmTJtfq1
PmCNZNGyPylA8ozgORRfH+5zm7zLyZaIzhZ1///9WuzsKCSTPfskSrTLM+P7nhSR
2psZWFuvWB9qZx2Nnd+0zgQ4jhEr5JVUZ3NigyFPVY6XmiQ5SjemsPuwwOogbS8G
9jXscALKgjMSYauFSsgbiUZXISmAK1AL4CmNzplwL804z8itYsCCUPExD8cWJ1x6
NKc9iJpryOynUMxlMMiYkkBv/B+0xiAANh+l7BfPYsC7p/jHO2dTFpANZZOKg0l5
YfSDFhxD7lUa9Jtg/vcjKEONhimt3NcD3YMsKjWxbaeiSjD5fNkavXZvjU6Wm8sD
Ezhfi9EYoR3A20eVcYisJz2JeW7DX9MfLLqJGM8XYk8AihFGbOk6oMOh0Owx14ot
8Zt6YyZEDLozSSH+1qNyrC0i9gULsmL0yk7+paWUKzJF7hRDi4nRr8p4uvAvDSY3
tJoBvQIQDfkpwiBtFi42gMQKjBaE0Cy93M3Dm8COHpT5Crn9HAtBUUNmHfjeRlQH
dd8JyhdznuKc1mhpDIfu5J7gIL1Nyt0tBBiE0wb/V7g/ta5CQAgkJbcEHlBZbeQ7
PM0m32ZnodIWBLJM9AGf3JJJBDWN8CGdjgd0HuiRkb9RjljFvw9PH+h6taoa1rrt
9o8EkPP/BtW96hjbp3l4hbaPUTusRXOMO0W0h3R6MtITVapQ1awHvz/apzc2Yet1
JEBXrkVCyV4gA5AjTN7mCmLQQvWrome/JUwlDK6RGNE9kJ3If92GvdawzxTdUZ+i
XqB1WgkQm3WdWyojMVZvRfXjse1cJGQu4R5esOsL5Jb05JSoVxrmf39zUo9075UT
L5+Nn6TrIxfSrxgmvKqlLmAvAVEFwr1AWLpTpzaLBBeA7pkGTwb7AbegfyxNv1Y9
0pSBsmzG+aEv1V99Rs5HgXFthHikwD2nrosNnFf0u3Hw9oRjt1YKRbwlUej4E9UT
ChNh7FbeqIL3nwZwdzlAN18e0WGwI1SzK0DS51uFYoSisf0WMQx3FlD71iJpBcC2
me60WLb7BPY50O9p7p16YxyhIgRVC0df/sTu7XaoDJac0VisgmJclfiKj8eSKx9P
6w3r/jqCRQI/kCRV58ae3qQBEbvuD+mbXg0Sb5V7D02D6EkpTqdzsQe3dvjBfTrE
obEFTM7h7Y9pz/ITt25SEF6mICfy4v/Y4V42tbXMCXon7E6fArm4rygzBBtkE5ps
VaaqKhs5k4WqgOe/v3RgPg8f0uLWd02dgAfrmHfZoNS+XlRo4SQfEaCdc4N8Nuak
H2RzIHGXEExxSfAxfX86qyVVjhFfpX3ZLzWm6iCPTa0Zam2LxhZPgN8h47mQZeGn
bpbBg0u6ueiFHKXDHFN1CnGeeq4qOhPhUswkagSP513ryCPDqFWvJxQ6TysmUB8e
irIzyArEM9FE4pnMIK428VCwnopXMRCwk94uah314k3cW87SHJmXAKn9fohmE44x
K5Ip/WuuBnJZ6mqlLfZoqHnhUt3AJOZNeXIqOHf2anNV+sMC/ckcQQ+JJsyGbRoQ
NbE1scT0fv0ACneuP7oMczrSLmafih73pcawNZVBhyjZUPZ0HIczn/X0ufPXp0Yu
RmvvirzlYn1kOtREbXI8saU0IF4TVuxcAPsbW39q9DUX1iLpo25L9iLVNdKPeVQx
Pq2v5EncOXlRWhxWXVe1D/hAkUq6yqx0LUfu4jXxsRP16Ssa7IuIqtY1Ju9o1Zoz
cWyglD84M+cmQlR+kDA2rokpFIcklnCS7e3I2SbVp76D0ZwVBfFY2OOOU1gKcWFR
nK5DbdG8XCfg3nZgEwfqjqjFZEfJlFLD+AL0lSmeGHVKL1+sfYrSh4SdcBo0vqXL
wZx1UbkZFpCV/qgU7m3IKULz7VjB0BlVb5ZVvRrmTcRS0Rm2z01H5QoA9A/8cWto
XK6/pVmwQcXyBT+MPGnPltwxTOwONlFbi++y1Z6iPf0gyQ5iaLFlfrVV0jBZL6U4
Vw4lDd0qF2cTnPsVcM2PVf/6JHc1IJSTbNjdtPWkV4wVK+EC5rG49Dl6ZRFcAq6V
XfwZRT6sNh89FJt4fir2ePjSFeyisHQEjxrVphCd8QElvkXOBFFNoaMjoQdKaiVk
iJllcwNkMQBmYDjmDOUf5yeTNePrP0Y29K/R55HHqdAOkEFxxaiPU/9BMCNX0chF
tHQ/t4HDz6PG9dDzyhqP4JsyOHNTT/q7AxgDetUToouGgPD2SlnidLNfMHtgt7x8
GNDSG9sf9PzD2KLNG0+afpNmdpIRzhX5a0erRlCly+QiTFMp0IgUGTJbRqb4YXRQ
v8WAemokach/UHjgDWc0C3Y92DQuRtTWNwEwx4Y3iBVY44vlo2NRjNr/H2AAscS8
tVtgmoAwjBfEwMvQ6l+CvvpS615waYUiS2GgrFYlQaFUjChOsCTJbUD5IsjYK1li
87cIPtnd2zs6Ov2sfZIhHRa0wnV4Rs82cj2e+4h924/QLkBT4oK0wOCiUzAboGZL
XbAVhPf6gguuyhB4bv0VmnnGxkdiX32byLBEFhZtjPov7McK30yu2iRKUsGGvzO+
oEGwoE5VFo4bfXmsPrA+MrG7gCkpxM0UiupjW0D2VldQHX/A30qbiS+PPX/ozOnc
i+oVM5s55B2asrBCsljQunQtlvkO8Xvo0KBakUnSQjtyWPJBem5EGysv0NvPEW5S
Z37pJH5jylXoDrpvq7X+IM5qaYABK6cWzOHCmy0HOU0RA5KAJIRlQ9BEFQabMeR3
aG6jVnX1jizwB1Pjc024JHPa52iQtwZCPtossjVFUIM5oV2NLlvUyD1S8MWdb9al
2MwO8pMj1EPr52C9CB8xLj4jQ6o1TkdYcZl3FglA1QHoWloBn8yUuT7TUbjAUYxl
MvFbxxFoHOcPZBTJbNgjNcYZzRRhU/A9tBmITfvv2l/ekpDKEqpD71uWcU+z2BYB
6hfZ2K+FuueSA9BY7WNN/DJvgWr2W/CYZLgyQ2zoHERlheY/GKB+QJ1BZlPOSxco
IqlJamw1HRijQZaot286DF9nNhR7S2kYiMUMVA8VfcnuVEKwv6stSkSb79nCR5D+
gVLZB4EsPbL7Pn0GmSYrAImHrnrtonDvKEQoeAhGYbJoGBeeJgR04/LDT+Wjw5zC
c3DC2u0X7IUbf3SmE1ywAN0QHLlOEirbEe6txkm4H4s3pjKN68jcSMf7GuJYGW6b
ST9PICSq4zyUXN0i+FGsPMR2Ct/PVojHxB/b+bWezPkjqktg9VTc3CXyfx9g3+Mo
SgaX5puFW/geU6LCIrbyeHVX6GKnQHNkuZkD78+t+Cg68zUYenqx+jaMrQnkROrM
DuwxGCqnNe5HTzCT5S7tlhbZwqieWxbQp8XivOb5XjWTSHWypQKMvyyknr1RQBQo
kB71GCClECrx4C0Dr2a+iJ8q8i5mrx3iLnKxyXk4o2S+eZDllwyuZEHLnYqe8mxl
1vmtKFjS25M1myQBK61oYQesmIDTPBKDN3vgr94qF023v+AArXJAyf5sQlW9erJa
pORUfJ3ycWAOvnZHhNULOHiwCoEDQC26OKhNgJiaAuHLxB6yz+QSahwOk+mbtc7O
0B/HcSanDkX8R89CoWYTz7eG270P/HGhQwN+BQZ83pFwR1vJG1qzaL8W707h90xE
wQDzJmsNp+pd6YAMtSM7J9H3diVGkyODDyPfeB5LYHdGdT+tzzBQ/hTULLMMzZTK
j4lt3WpN8hUldsyXf/KNo3g/TEORJqvhwISTtP5pwU4ls1+ekB13mMBXP85JefFw
ZMsoJvNrOK5JvPmtj6YYBccwFZtGnLpQBJg541YnDTX867aEyi2qHHeLri092dN/
hWVSXJdzvjg2zq+ZJXq2vIl454D/8EIiy2B4Iwg0HkhqSEFQywtMj4QXvWlaTfDU
/KFUQZv00m6Mo+Zx9DY0oiqQ0RPUtrUykNeXbeW4ClNBJbYvDeZCRkTjdiS0ZRD+
e4Tg+uXua7udf/iK41QTNJbdcrukWu/+/ri1K9Ap67MmTL8prRk1Uc/WNJYn5zqp
9IDUnMiGbuln1mCahOhb7FmQCeHEiXjUMRmakY64pUX26m0gElFxcFnRWp4V+vqY
+MMzi/3GkdQKypRug7VD8ngxXqVHhui6/T+x0aj2I5VwXfvQm7dbfpWmb3CO8DQT
sQVIReO4oAkJ9MZDV0VqgpAPfNCdz9IcDq4XLRKrEAYJlu3MMQxqYCw8eAiKlHc2
LIqC9MDTlv1Iw4OvS66L0VGXj9kBaY7YHXTqY2XnrAeRomVUUxsxGBwL74+6GVbA
f1wMSQT0KrT5+3wGp/BcYKcYN/7BoJTRX9pQno1HcWiCDdBpGyUjvRKUEmdZpffD
l3X02iFSGAI761cAVebzt57azqwPSPq1UAGR31MaUR4PyUwNFk4JgbdWbrOtbQAK
jJz9dAr4de9ocRC9MiOTyBoknj1exa33Mnr7ya+SkosE1zpAJpkTPdgVjm1mE1ah
UarzHlWAmRRzOIkR6U4xXP4DSy4MHoWu4kDtRx8xV4+rOJqYHjUyS7YOza1KpE0Y
IVUQh9TG2qlS3mRd4njzIUuvgLiQn5jYpPFXE1iTVo4gPHi9izgePhZaI6Cy7rDq
yvv10sAJdS6MYbHfMW8Pbvn9mEFhJPIi0KIcQxvzNDODBf2dVM62FOUyc1HBWs9u
Qpk+gtBnwVXOeVKnxBzxl05e+ko0Oa/5jcAg2b451LClZ2Ob5Y0jLEOgil2Wkxft
REzXoyxorogqQdJ+K+zdeBG6kPulb/EC54NRx9H9saIp44jymU8e6SxjM/Darp+M
Z63CtoQNpkByvV/V/677w4oi2koHphZtt43nEBfaMolnjSW+MfNOfiRRFMU66Gm9
eNVCSQDLEBNLlMSWx0aq0CqKiIpChny6ZuLaxAW+LMhJEhVhUck63DiAUxhkaR6j
7W80E5li4F5a87wCl/CJIDShcRmmaXPsx3vEj7/oMdHdg0NR99M/malQOU8z8AJl
cQ0538YUEI7X7ErqY+Il3jG/Q44U/U9M5c9xgPEbCJyZqJaMkjsFWjIpySm8eHJw
ZNMHaixrVsTXv8zEvkHPerDDnwhpYyVXiicBhi0mXl+sVAkJZWGWPJmOWS4/Tt5n
x5Jvkb503InmQl1JH861ilf4UXGNCfn9YqVvnmgccf0UCoUyGv4kkjpa4+W645kH
le5IwyefVnNBTiMAZGQ1z//2q7yZMQ28Ugt5mzhxxXejPphV/KwnNRPeQlJIJC4+
EsiqCegQm1KTDFQX2RrKg4WFwABlKNpRkTfyFNNtmqZPw3CUJ+ujLWWpQCA53o1b
VrfbJQ1GlvyQH/dy/FAytucC/63AY7UkoqOOFt9cBFvqjHHEuIusw/tGgsnNsu8G
VwVWBldlmqVRxveUAneiBuoFSxXA7aQjO5wOAvzTVZDPYBg5veRCpw19H1N97gIr
corSyISCJOyOKRMNTnIrpTrCHI7u0/yhIOgyiLHf5yYnwa1dvfOXhN+XvPO5kt+Y
3CD0tkwO1qzaA+9z3qIKhHnNKhwNYhwi7rtMmig7r1GVTNyvrFdD7WfJfEuR8hcw
/eJvgxhzY839gBoqR+p/Yw7/dfbsZd1QBvHSj17OJomqkYA66aPOLugmZpXHwJ9+
pmhxWbDt8LKPt/LMGJrfb44AQj5+1gqPuOP4HPUfymzwW2OrVBbNrJeZ0GDwZL1u
MBtPeoM4OFYM7NA4Vfaha0ds/2Btl79eqtqzpe+4E6H4gCk9ny+bnNB4oWooPmQA
qRkO+eq94M5aE6LiOpzpUNQe1YRPLS67i72jOTIfRnjx6tntVSl+Kqp004xeJKta
GXyv+KVl1C30RfNHZDIEfxQkn3IuiCCmEUrx1pHP1eeCDeqcqucAOzJo+Y4S4LQk
H+RNkuN48OKk1fwK4JOHceUuJF4MKY+EKhDHzyfKUmElXXYrY62xeAk7ml7rBw3+
JuFid3XUTLec7JEqouM4SY25J1kbLvBlGsRWHFrIdQqp4rMYJYlcOD4v1E+6AzfL
95Az3pGnuJQ18k7g/mZhB/elVzyCXnjdD0XiXnW1jTnJScZ35VGcGjAFjfiU/dYE
VsUXDmrw1bFoYTqdzdmOL5pOwaBd6+DkKhoLFUokhwS2OkREbe+q2ph4VcgAly/6
5Isq8aQIxP4ONgTuKQ8RuDCQEoS8Hp7h4BRlTzhzxFmAFPlxij3A5HEocAhWVVQg
gcOfwHbh+Rjv2qZhCwCzmLovoPkRADKfsFPAZaLN2BrFTGOzASoJAkrNuUPzk2Cf
doy847bPTY8KZ95FQm0l4oZcOUTNC9Acx4OMS2OUIZKxBAKdCGcJMKxT9nGQUWma
TjEpIzjPauZk+hPcd82bTB8IKcK4IREwPrDtAH6+GOI0QCbXLrTyaab72lDvuCH/
vH9vYgQYaYxFssyAryDt9yJMVfIofltI4ZDL9MhJzRvdaZSrNIMDa6xqtbb/375y
2sp5MeM24rLGuzdkD8Am0o1Jg05fQZbq+pON6H/FMRNrBEPAgZEqce0wjtKf1uYs
VKo5m2Toh54PRsuOM8Me/dsZyP3/o0xuKt0TmnW1+DPAwIW1LFUPEaoTsWq2019e
PsGMBiB9Juo2x7rYWMq4MSNPd61wZxiqYimhtD5f9Rj35Hx+n2Z7Rksbdpk0sftr
uVOMASnHdTmlyNIK21PT23NRk60uKcyNMSNEEgfsW1ju/7oN5haFkCaU8GsfP9PH
9ZCVkpQJp2NX2c6jBMEPNsGhxQAaoKixm6yJD4PlkCeJUjLpYAES2Ckso+9CGrsG
EBN4OJ52PlYDY4GXVd24rWT/sqz/mWRl75ZN7VRGrKIyk9xfzGPS+G4KR6G/Fcsc
o8LWv62HEHLv0vAVLxWgCcc7EOP/d9X5t3brQWgZ0NZVLqYu3L1+jXY6m6716Jm+
g2aO2PU7TVlMpfYJUQAitVF3NYDuWrIPnV38W5/VBAYwiAVeXVy0gUZ4obFD/12k
HVUP68jjkdg9PVUoeP0OQNwINqAlZW+JjA0T868luaPcUMh1hIoxanw5UawDP1rJ
gP0EixJEUq+4xzf+9ht/EFB4NzwNYwhljHfMvUMrqJhkojVe4+PgTa3CSdyKIELu
gJciFwDWm02C9fg0CAEB0bANUroM6IbRLjt9arTeQi3F3P8RLKVsnIlXpHVrEtFz
qR3usYoS0LPtDp/iLhuP7Uz4IxEs/QoPiVEDfQ0N3xNFce5SousOxHitB0s+tToQ
IslkrTe5tgR8KVhcl4iwdZnl3eACuyuLfbSSbbymB9qw1Bp1okjfSh4RWc6UWGRz
Z7wMCzja/6yhdrA1zM9V4vfFc0V3kHJ99uxdTtDS8ye7vb7cgZN7X/5AmYSPhPjZ
/m8SeCC3j3U3CJyu4q6MBdvqx6kXpEO5Ufa/1bg0g21D7QNMqhfYKGxU19FI6HoP
XStQ/fCuGIL5oO+o5j+4Iq5gN/JTyxib1eUnyogaajSFZBAMM8/DwmqHzsrPV1/1
AtTPuawiA1R6OsdA7/hd/IVb9vhAaCOrnp3Vov0Qox47JiH7b9/RUKd6uWgGeEM1
l28u5BLpXWHJ4VM/tExykNuHKGw8029aucwdCYJpvOZrLXcf4AfuiMAPHWZD9tS7
rj/kmfke7ikJ8wDtba71+RTZMuU8JO0XIrfxF0tNzTxVRHD7bN6nu49hXnJP3EMB
ayVVaskM1vmhUZY7C95qCUkoBDU0mkg3DccsIA55zM/FVHKABM/fZG34alhdh94V
FgACBTzVuU/upc0YCeTMAeJh/FgvGCEfRu+ZZn6uBqkRakTEcwaVX4BUpymtoJIt
PaC3F7g/SUx+2ecGPwCEgtMm9gT8cAaLme45l9PEWCoRzOTDeuYJCxWCvoHtA/3y
oa7n3JcXmkLqF4puaIwE8iyVm6pGgGWL4pDEr7par4ZSuMMg9MtwqrHIe8kklywy
Mm9jqzvOo3rTXn9kPYL1PWITO5pTYJp8mGFGiV/9gXO1ZponaY9vPurWnYlemK1J
RmzShBRKHZzsvhJdIJBMHocciIffa0ZKeQTPUzYsSK/xigh116QmTjasU1SeTk7G
SKvBD6wa2+37jA/++JRPkG3DEiUlLM6yNKHXdWaJ6eE2s9ifPnPPFZOMM5hx3Cis
3pXvzsPZiLJbOqG/wWLE0H/jAiXQuAl19XQCrEx1gSVqsRyqKW4tdLgez6FXC12r
RQxaMeOhbjHx8YLy2lkMNGv2/u6ipIOppmlPVBKmjE6tDvmmWqCap/Ud2CLoCtuU
x9ybWvC9N1KAnBUjL7h5sDw3Y1zSMvpsny5C6Y0uFzkgTfkdPuikDz2qciV+BoSz
53yX34bn6o+oNM/tbdK36TI/ih72N8qwurAIaY4LvIMS1xWYidS05t+lf09ccQbZ
jKAVNkTulJfzi0EkHjnvwprIjCEj/YnyIysaURQ2gMcyNhwJ19FRtd4/PfVn2Qpa
1mJasA3qY2kfRxIAdfVMe5mrx8hWhHoouXDooKXdI0eCWbm+BPnh8irwkJRaGBly
btAO66Vo88hI1S9gA8mt0ggfv4itc1ERv7Ab49vzFJZnkB050onGqQz+54aVoaeE
l/tDSXhNyZitE2ZVY86YlW8i4UnYxufm8xpneNAdObe7AYXHX3h3isnNJAF5Dn0o
Jv+FTiNL7wWRxeO6D4qn7AmqXbj2wGZWE1AH1OR+rr81GmgnBP5jE9d+wJFJoSSx
KVyTo5OuKoxDcTFjR/hrbSIKUeHvV302jjt2kpJLFw96KRHenlzVWtDs0+5W7dAv
DBJZ1+N3aW+57z5C7synBmETw5e0bbx+eL+w+ubyXaF+GXcdXCx7ez2r1xHMtj/J
aceuFn81jnQAbFxKWRYAoWP3L4k7hrRe+BhtMOqtieCLJCPCHJ5M/0dGFyvDKpY7
xOlo0H3hFj92NV4GgOylBIJGL/hi0GFmvjrV4sW8KHwPaOWkI02xd0EJDuzl0P53
wLfQSAAo4xw2ZlBwfRjphMuPH7eoNnhpqp0hxB3VOMDoP84DKM3tj1P+uZ6wglXJ
ELe+Lqi+wCt8kCrzI3fHn+BpJ+Tc+moJWKoJHOFtUncTWot6r5K3Dn3PtPQFY/pq
85h4jhX5W1jQXwYuCAU5VARkz+aisW1i6ffukDpBUfRX1L7UsgWNsE+fV8gAqkz7
kUPr002OPydoaT9pD1zfj1mYI/nw3rqTEqjKUpnhDJ7p4EJ2nLiei0Tajaj05UWS
6rKW8LEKDejYSBLHbb4buz+dWLXjS3uWAs40/ScSsm06s/G7EdpcL7lKuN84xbEc
mI6SVme42bMlXy5WRNkBJvd+mTnIHG10nbn/lTzuQ44xBEkyMj16eB6wzpluYC7J
WfHwk5BfDHo8txFy1EdDqgCLJ4qE9EPJlt4uGUqiAmGmwWYXmuu92oG+5yCAKs5G
oU9CWRWHk8ctMjCLEwicFSHgY2/fTiXSSj5a3kv8FqouoGfe67cjbwEE6RBQ5G8X
HJCZGo1hm2/H43IxJ+HCaLv7Te6xf9Gg7mlw46jlm8J4oSpF5puUjVWo6Ur9b+6h
RrKiVO9ky0xbYgbwO46A1S4BrXoJ0fza8MNMOdnyaMpr6rMNNBX2x77c9NEb9EZv
xRaXRAKnopLcBSsSxAKPDMURLXpJDCmtJImSlBRQ7WFNdKqLEV14l3yAjJp8z3B/
I0xRHT7M2UA/+yJsQn+3HLaPq4jb+DBt3nBvhvJkff0S/SPHxS+GTP6EdWcoSND8
sFIvo86Hqj77UKQ8cGH72LCu2KkXjKepa189djkxNyOVF+VH2DeMFmBOecPER8i1
0YUMItHtyBzyalFKQLk0Mkt7T1R4riU//3/dPEygv85glE3jlvxji5A/sFbbtsNr
d/g+pZCsOPsImA0V/NMf+5GK2xn16j+dwx4aI5/9aHkTOeEfkbvYKv2mciTac4mN
4iB+0pty1i67BXT4szv+0UfK8gfbOWthALn+MXMr0mkVrlqJrdrdsI/cvjmvmu3v
plvj1YCPg6YOOBlSCcqrLj9bDhYPlUQuY9za8tG4f2zZgPCczdXu9SOXhcHUXKat
pHJNHxlgwcdUgkuZHtRALbBGPsdwUPl7wJubrSJT+LObFY03Rp6hXjPgZRZEcR9x
NTIgTTByetTNZc879dgWBfSklwAB9a4h1p9KxAQSN2dUlJQNoUaRmZyMkvaf/JKx
aD7KWEqijrP2bJZ7b4uebx/rEQDRUA677pSdFE+lXbfWJlu4Hmcb52icLrIkXDHM
UrDbR1ALbQicpl/zi2IoeR2kNob1v5ltyABlSeujLnNd/IeQ3tNwgSeJV3k5ZwQZ
eWZ/1OWj4SiB7a67Q27ouU9jh3YY0iT0VsrJk0Xwx/Yn/4j9Bog5a0g69RdUEJNc
XwYAhwMp2VFV4Z982FoG1BEnLkJcJhAEpwDsA6TrWyk3uGiD6SORE5QiDQ0EGsMr
f+dDXHSUXmsYiPhiWeF2OCcFg/7wxnL7Sr4AJI5sFpOfTgdW77Lb3N3wDzor8kkM
wdv5OskPbUXXGQefQp8AZSc92lJ0wPyact9XQB9O70gVKdAp/fRhn/QKi53TfjEh
gUycgq63jABneLthsB85q24QDBn62k8a+i9Be9bSqp4GE6iVdb40pk8F2QdGIOVY
ovqaO6YTwGQCqDigrvDGgFeQm/OeWDWCdMPmmZ+rCtsUdj37+LTq96p/7gVc5W0m
ty1690c/xDDoA5AJjOh8ouMTZr/AiIgHb+6myEoFl+VekKe+nTlW7iTR9ui2opNz
EkoLxPKu8KMV/Vv4JwSCcB4EAahp6NpL0MpsFg2iFI1fesYNQh8qifN5dsArP9gQ
xkgNyBfGaTRIGvyeWQYVhNsobvcbvhRR9Ra09rPpfli4kVCbuYelzf6VOXWwPDe9
Vn/EkDDe0lih11eB7gRHuQT7nnrqX/EBE0IdYfk980Ca2mCNhJ49TbKz/GEGMyKY
LM5sXxVJ3ucd23v/wJK58sEeUv8w/5lbHlzxZ2h/3iknCFaCP5MT1h0CC9pmh5II
6OzjN+k4wuAM8yHH1udtmnn64oWD8B81zK7MJV/3M4wqJIysTqUfI0HtOsx7Lmx0
cxyP69n0KW3XnCPEjUyXUXqSEAs4Y52N9d8fzXh71ByXzFEcAzH6N2B7jysiQUGM
yjSrG/30H/a1lPXOLx47jUulNc1jQfnn3fWqUCFiyxO6iXKlRdbXPOD075EEJQuF
4yTaG995Kdua7T2QqWh91ImAF+2T/HBLn3S8TQp4ZqwhXMqyOitpLp4Hg6O5dFX5
pQ+W6IJPHEp5WgxP1DCNzcGORSbriLP2dnA27XR0UXTUA1U7EZRyOCNPr9HHvklK
ys9LuwIEohrgW+u/2kGUFkaRRQhlxqRxx4jk14XYdiRlZmBSPITrmajPXCHM55vI
IeCLIhT/8Tcifjf5Cw2zLmwmNAn0p8YfcsfMSDj061s0/PsesqXMTTLmj2CGaWhE
ZcWWgYt/ybZmWIKuH4GmpZqDMmkpnBiAR/riaoy6BzWGVMf0+rKiGGDZVJLrtgGB
fvETy4pcWYZIMdD1S0xGBHEfMseccI14qkC6hygMS0SiLUBEMdH3gAJ1l5ssSVEi
TiRa3AYpmoYwrG6MsUjtJoX/No6vtVX1b3wH2pPmm5qJIt8zHTMqqGAG3EoY/HkY
yRhUt4UEBgf1rKciR4rPLpU3IqFKyY0MTn+30iVX7eAH7zUlMXdDx9+JEV8DkRmW
R+7cv1m0Y2m8W67Oj0EYzee2Vp2GXCrLcUAODf8C/pVwlfSHrDleiIqwUDGwLnLO
m0uUbpGX1v/MlIb1eNWrirVkFwmkoiFzS0xSByYnQGEW5jwGXyqRz+anGbDVuA12
Q9R4V2xCYbsa1HyL09XTKFBBt8ci97BwLziR6A3Zw3a/zPx36TEsp5CDsEvuaJTS
8y+Ibs0f99gwVSqhGoOr2NQ0xH9CI9Jd0BRsi5DEkPkGT/aQKDkizs59HUHsk5wU
Evj002iBvUMn99GPDUGQOfhHw9GEfUT25z+I/W+AX4Tj4ItqTeLRNX0zg5g58lgr
t0Wo5CAd79GO+a84bDZd7lCp7TqHgwEJFTZoy801W6RCaykFXQ9WnIpYFrjJLKKi
w7sNrs3DgQjEvZLfLYS3SKwjrdZaE+NG/FhnwYYD6iH0F1jMLOTYIKAFx9DIAv1t
JKpq9BNQJd74A5jgfqHqMGKK0JiE2DWJh7+UGTZwqa6GICdjbvFUwnPFyTwYBR9y
MrwkIFB1fIGulf7Z8Eitvsj+yO/+c1eLdhETZS8E4GrV4XAcpzslhwl6M9XIPCal
qBDy2GphrSaRSGm447vtOG2YWwawuyGmhDhIf6lbJ/73+AvkHVaMRu33oKRURlly
IDqN48Khlq6oLNcC0fPkQFsFhA7cm0/wd8dwRGwatRPDJUK2wRaVDDConCIi2dBr
cnvLGM1tfYlH5gMZbHgmC9llmfXGT4Z7+4r43oqxy0pa/33tYstoFBZBHTicfHgz
D/IeK7Mfb8h2pmD1OgelOMyImqkaf5e8jp5RXK4IRHWdKkbSDU7xMvNmvWJhZ8aQ
OGqx7405fM9+Gqf5nr2BFSYoRXxhR73loSyf3HmpIkWJ0k2TSL/o2I/NRnN1xQDX
RgqUE/AMJrUWxBBh+4BKqkRvZabeBOeEdhwT08gHq7wGjKorFGLTO+8NWzdVLluE
p4tYOEu9ym/XEnaIiIwvnIjGLzcfa6M7PUkRy06eXzRyIQHB0Dd+6mUpkwVeUR1d
lsHtI0i3k4StXNX4e5stgfe7IpyTz7BO2tzil6ERzEXER5K6Ras1QVj2XDxrnU02
kmHMhpswA2FZ6MoptUqr+pCKxhkejOwjjUI/0PIPUS8HBgtQV4oYqbKYy6qaP6Sp
b+gcUlU604Sppq4rJG3V/kKybsc/snQPEzlbvayM6/gUMYSKc1a5T1IVCxlTegcq
Vq52wQRv3hWlJzlw9IfbEKn9JchXgQl/f1ILMwx5lxqVT+QmtQdTMg8YCkRY3K4G
u6brHMmLT4CYJhMFUrpcl00RAteTduQN+u6XFQMO60KCpEZJntJAOSnV+Ckq3Q34
c/tGuU9KjWsgzftmdf5jRb2xqfARTLcLtvwW4N1itDfR1+t9bRb793wUzoaJm+kL
aMqeSYHyBATddNGNAJ1zzk9Kyrq+BmNv7A3oSUNF9bqi+yJaa83AkYKvW487qv2w
hWAzbHHQvrj7wQnhb8diJNq1lHLhjyGv85JCrH0U0P1YLpOX4f1b51ubB+EBayha
o1AYYbUaXSSTNiG9UuABhGEB1lwhy31sozPRR777R+AONeOLfPnoWNU6Cy5820s3
KnsPm3R+umAeMK8iAzYg1y7THDu9PhNrrfHfJvu9ISiNQEDKwoDQgt4ZmgpoNiph
NcZ72/KSjtUuq+EUO3RVjxDZZ1Ljy5Ls1xF/bqg8sNoRbrlTvArmRWy+/H/eUhOx
lulHtiVpTB6c5PPqzcUTEZOnTnaOSBCu6Q+dK6Njc+VIxR1VX+gMSe2EbLL+vyWn
CGpkAVyJ9nquM7jYGQ+VK1MsfOMJHZ7qLGoLdteMRAIli4voE/iPFX1TGH9rR/bE
JkyAboKFCZy4Ch0/Jni15SCd/csKVHQFIadRQhONJY23A6pMCEuApw//WCl5g7yq
++ZA+mZqJ51plEEwNSu2kWJK2kqA0Pg8TeA6sjHIWenjQQfHCnTNXMfyc8jpbKmj
c1vuG/ywiWHb35fkm/0S1boJIXVDalChLgD5CSSOLRrFqIBKJnxwnf3EOD6yEaoz
5T9IILRzNADq7RFctAF8EOKkGTgK7hob121l3oWgId0x2AoJni3opU/fTfzk575e
znPepD/UHaloc11YqeH9p9TgffDuqzb5NbHJJF2Fu1a/z4jKX7izHfmdkcN6oD8w
0mpbh2gIP/pysH5lGE4fcAHLB0cd0tIHRHVN2HRbOzx3UPxwcqD1nDC61Rlu2r1/
hSzlaeaV1hgXF6rjH4BZw0e8GusubSmTBqUHNJ5kXkegzqxWNJVccWO+7EH1cK5o
Az+bvjkY7HkM2jrdWvQqtUutOZ3OhwwCzjFlubYtY7fY4r20iOJjvqalZ9M/60F3
LueEruSbTu236Ygpi1SPm8mmaPzKxMkqX0kisi2PndzHAUfIZiqW0RHd1VN+5JLs
Iv1qMr/QdH7GM6VQfOgKjXOqOM+UWrEciYTa0OPIQQpi7JjaBjAXaZu/eQuJnBBR
u8+neMcDABPuaLASiCenIZF7ghDo1MyXp5ypKM6OsdiZL05VRkaumSg7CvgF5N80
+2va6ujWpO17rMizdOVjCINVdF2HeE5474w6nLYmsl7HkoBSAMHIHAlSc4Ei4lGJ
tzHs6On7yP76STVMMpCxiQM2YVS+81IJP+Idmdibu3xGX6sK0aKs0tA9MI7qMg1n
9B/fq2DflDuGBbQkCVeNbKL/+KkjQMMV3DOqBiZfkiXOV5N/CDEQJfqcaS79iec1
zDuzFt7JA3XRp1Vap4V21vl6dR9b2WKQV5odaO2YvehVJzI3gnZXm1+9Q2HFiwFP
o95FPUlaDxepiNLdCRwqMhaCwQxvyG+/COATXP4rOpqqmgvZzTTPA/9dEbPysasK
aD7/kOYwCVt0ScDHwOeoJaLRNSdXDslP5VKtsHLF7ennga/B8QO2P/k7Ks/yzbO2
3otBDQef84iMAWAzFFufIJuGvLSI6PMRw47WpCedYUCI+dUx9JE8VJ/eh100c+vw
v+szyC1eUFK5SV61zQ7IQs9kQ774UZ4iutcS+3pGlyXLY7+08SY2zAEdj/eAz5Nn
lhLgimdLdCBJXz0WxzoFK96Tu+xB7A7mhgJbEv0F4DJPrRNeFBlUsjyGtv+dQeax
vb4WTdnWMM/stSJcQrMTqV680xWVafZXx8ez4sEMztoikw4Ql4TS59vHA+psBp27
AJvOXuEFNhrfK80ujIn3JO7TJnQFVqBMiUWk9Mlgrzmq85YIF3rpHInV7rbZzMyd
fOSmoxNDPQf8yBJ1i45BdCwQxqY0n5Xz85GUsuSwjthiQfhYo5g8iewo/bSL14/F
Td1cMZrgTgPsJ0vum1gdh8lIi49a597BNiNNOSjin87qdM5UMq6W4sQTiFKZMr25
RjNwaidc2kyFte1hn/frNpkZ6N0Yi1ipsrrIZgkLG/7jTVaGiczPQ/MAiQPAtOlG
7NS4HhubC6YjS3BlBekp222lmedtUO6C8h2d2F0u88/RYjK3gRrEzGSQvzhTSgsS
Y8XdZcFiq1kx3EyDY3Gy4l3uK/KfWLB3o8VUwvBsi1SCMxP3CgrkVYogpCbzudVN
vUA3hC65TMrgKnHGVpd9wGHjArhar8FFoolrP/BeLcmT7IOxFu8rNn2vo/H7xUfK
B++2e/r96TQrrEvVlCEJQOrlOIdl6+v6E3lPOelgs9RyfRmvmMCOannissEnvZn6
K4gQdpQDmrNGQ4eFG2Th/YtmRdBNvw42Uv6pKFrDOD+smytwZzGbbfsB5cR3DCBK
ciT6VZ+BEb2Kn6gZhMCY1HTZbWWUE1Mi+BPJHOEoKrq+cODExv8JdfaRZphTxquZ
MukEZ5vUi89IxpD1fiTZPpf6rKZZXRlRiIh483svmofO10Hujdq98QJcM0moaRzP
Mqm2kf+PPqHnzbcqUVk0tjD8MroUEJh6OQEi5FBBDDOMMjtEw56FcLRGEHH6ht7C
NwPL5JN2z0f5aOP5XWO/JpyeLEFCuQ+qIwL0GBiphpl7kKLnyZcgdMu8AoG01dGg
zepXACAmVAWbGpNmu/IFqazcxDUu2NHEcVcFP/DkT1L6k3dkNcKIq7JtBT7MFYXd
uhFn2nj96MDZrDm8IuOLdgWU4XW+6iadgVnVkLOy+2RDQFb2K0C0u5sISpi+i1nM
1CbZJUHeXvwwdlwB7eO/+VF03eXjx1X3V5bQtJKEpyjCFQXEaEcDLi59tYcx1HBS
nGMtdlf+pT+KKnpSobk2kNWPXMBYMGwFg3aMgMTQsF0ZwLm1dJ2wJevJXrXRJq1N
CKTLUo2qlKMEVVVWx95nRuP4kqGuvHGcT3hwIOjksejTPc9Zf33/20SXUftR9Vqi
0YUUtW/rn4hc/t7Y45RiWpqZeKougHgWrn5FBiwWeGRd5i/A8/SOuZqsA3/1i5mK
Ks5NFjk00j52H4C6cxf5tV/4VIpHy12kgBS5DZHtC4eWeF3PrLa2YGMEXO4Mkok3
iZNEZj98M/eH4s3dU3CuYZwMDbSHrNIdaXDYpwAkBXNnFLrYwC+oS3LLm2hDost/
EuYy/1Xc6EdySoUGaEyZpcabPOOXWwMOsWHWRtJhD316H9aj1kCZrfDP9ggrTvQe
ys39ScbR+WYK0Q9X59kN8JSy5llxqXKT6adG6b0XanF2tURF38Q64N5JU1fXM+n4
bJCOZ2Md+ypet8OLFBX73DBL9AkSgqYRX+QG0P9pDO+/M3Pm/kXoTkwjs1+5DIf3
5C7qmYoc7NKu7jxLRGry9FCzu17x3/XOuY7XNxZcizqmzfJvdKyzGSGSme7N+44z
dyYMxZ91178zQJoSd03Zb2Yg8pYYNcAIrPATiqLyzmQc0LcNqfF8WZM7Dwe7sSQb
BFcrarGIMN3M/tJLN505deMpK1JyUkHRofOe2UxFGHAH1oZDK+UMeSK41Ex5ozDB
nGtnGhy2xZVQisTlyrdudedBHy/ldb+db69glAp728pX6+jrw2YaixVRdvh5PpFu
AS9472a+kcSOM4bf0EctqLlgT1ufbtY4jYHbAsj7/4C5QcQunzXdnELQEzZGgX9M
tkeRyod/ZoWZanWVeitcyK/vZt2SR2HMV1I8yjMOXBQrOqbxWV3zn6e7XHI/fEQs
+zd4xAkX2z3QS8G2yc1JuJVzFmSm651+6kSxvFRHM1OHf5lqN/Lk0Js0I9ilo1vi
6FOgiQiwwcCVYw8jCN5BmUQXQYdZ7Ij+rC5yBevJNb5YRBgLFqgRLyDqOY5gcb9F
RJPUzKozHvO9Wf8kN7732a8tJyVuikIyTe858DrdA6vERVm74XaQKjXnNxCMZWSp
1O3lc/wMBLI9X5mLm7edvnpFUvQRTPvjxFSMeukh8TEYEAfMP2LqdPUO0kjuBW5v
5iDbzUBdxViFLrE0MzmFeGKzq8MXLHf8JjDP0D9djWQJbzYSgBzapHI4k8Ozq/jl
PgWcgQ9fau6K+Ky5DBk6puv6Ivth0j2E4MyOyYpoWpzCZKRXs93U/g6rHdDQbrGI
e6ozai1Ac/IyuVYDNpLPBUrI2Qy1TPGPk580GZDnZaQw/6wB3fUa1/nYQe+oXyxs
YWUn23/Un+KZo8lURKV/FgWxP/KxFpq09M8H2IpFO/VvQlmMpRvheJi5lggAzJgO
3El1k+o19IzCarRu6BQGyi1Nd3gLtQ0i16KHta+LFSDW7TQSNp8hQreLl80J0hHk
uL4UgaXpjuMRRQ2uQTyH6NNM2EeiB0gIW5swJ/9X/21XGr4njdIgX08HtTqAF/78
KHaVz2s85FkAtmsH4nJcKay5JcGmS0x+whhioDU/+uBNGWJKTqke2GKBiIZrXW0v
nXCeaN/23yihP9v797gO5ESfTUSxGrt9YxPeD54cWMNm5df9KFZJVEQOzcK6ZHpC
rtjQV8/39XXBX/lmMwd82LfNerc/ThoeD/VFzLNn1jh8OyesOU7TSHgmJT/lPBbn
kY4vACKK4Ys7pClV0rRWMn6awpff067RTwylqT8uN4vLIGz7+FeJJzEv64ibLt3k
SLqblnDZgdi6P2jQv6fOXJekoPojZ1G6Qpro+R+nnVSAJfMFXA6LZrogYwd/eUDf
bi7e6nGW2ssZRMIo9gMbZxdXZdpkhpZbzrzCbuadwg5P1IENURpSUjaWxz2Q8X81
mz2be46QFumQzwPx58upn422Fy2uOqPw06at1fwIONRS1f3wEhHzMVEM0Fe8CkPS
MW0ReKyZ8368BqWbGHbaU8M8/Mtd99sJREY2a+qiyBaclpZc6PvUrIltpTd7JQml
H/aPLadYIh2a4P6Dot47riwUOz/IiG3BFM2bYxjK0M2/yrv/JwRx1l9/qLkCpL7r
ryAqF/OcY759u5YXa1qIejGG2HQL7fsMu4tBHLK/nVJo8+P5elWK7YGKRoLM9Qzc
ldaD2e/b/5C6hfiF+EzcXeuyBh92+Hi/xfT2Iwuk0sG3SDOmaE5/+pU0/Jw9bL1f
TCiwuvXdJjtbA/GOrZkUZ7vdpcvzA+HrE/qnpvYimWvOnx0mbewQmZlEQFCG3khj
G1Y36Latn8qazj+mlR/pRh0Quc3qHZDsiIDZo5RsZT2lfHw7lijbg48LE3xXwgPa
oTMi+hUPo/k7whbjwhHv45co4EoAhb0aHn5pc2XDFqot7fP4FZEyIFP3/84Adndh
dcck9dDmd1AlQBt5PzydmPYpTJ/7YHyj12sBtj/sooOsRqTOFTx0OFfOU9FPwg//
J2lTbmMIG0v44Phu9M6o37O32h/AFea37gySvdBtwfkVKKl3qWdCuf3OdbSIjEbm
0JFM7fTBLZ7U3VCm1kYFZP912r2Ty3oen6f9HLhtN2TLU7arOBUYE9gUmCMEQKv2
TUwT5Q/GAiqTZ8ec8udmcZHNs0FY7wpTN5bdA8vNUP3vNTl6Tscj8voWAUrRYTha
z/TT3J42veAYfMLiVSUu6qnddq9igtulscJq4ORcTZ6/tD1CGKXIoYg8V0g3aeLr
7RKDc1vVLUs6+qIsbcNnjcTrqqlZjIV6OGNxW6Wcvqw0OPXCWtCcyUjSmk0D9HcP
7XJvJ0qlMcg4brNNSMhP9nCAtHiSy8DJvRXQ8SVBlbydEF+AJwJ9x3X1iMOS69I2
e4uzTjVAdMYcvwNS6hYMWXvTnFKftKBqGBg/YJN6M/qaEYlyP03P4vtcHsC/S8Qf
u0tinIgItDzh57jV3kqehU5lHdxE4tQkn14s/kEb0odhR3By9QiLF/v0/TQozVZk
iS4XzZxlDJTEHzKuA9R6hKta9xuc7WrMN1gVpfVPU4hIFFOySazBvKb5gAiqH/yk
0GtU8tcwOAtmTCkG6qm0yJijqXgK1AtwXodmHzjsEijpaZ8VGG79d+B1a+UhlDtt
5hFGHPGmH9Lrh2xazYl5Um8ucqnsduw88t5+mZe194jqAnToLw2OKVZFDbwOwNV2
SYVErZccFR3WaLH6m46QNHLy6b/LO6bhHc3c9QNMeeVPSN+enkFZoj0D6Hg88HRm
JlNIY/ukL7+mFf4jcV01zUpuFwT97y0/W/fCstdra6mOHBfijpifyPecP+udqfsC
6MymcJkjFp1Ckyo40W/fPZAlyhz084gGuiVEh+L9xS5Jl+XA364Wr4zDBVJGmVR/
BnI5UWL+BI8zU7yLpOO95poymdPO8SDbUkLgKU389p4t9kQx/UOSsc/24BZtqZzD
c8Cwt9sD2O8PioM5DitcC+bLKDmIuyTps/YhR5lH/Bw5reIMd6puXTbXDXQhojaN
n7mjk8avsAFIF5TbXBu8693F4zXj3yEhLC1hwge0Y36UrXxOydbjL67IfEZZznd8
D7jcqV12zLL9ixcYujTP2B9AUvqoCRAR4Bkic+v/QZJ7jRZRBG73kbJmtqXJZgrd
2FXwzzOtyvqVtd/Vxrz33NmnC4Rv4J+Y5O7ufuB30v5ySQDu+Gwuph/UTmJaUGOH
92NIi8HOXf6NV3MmOFDvulyPH2J0cSIcRPOJHLC9Sy5FGWEC4tqdYKJav0XzxeAJ
cTupi4+t+7cJvCMNLJw5ok5hFiKBxGGeCUFQ1BMnfAz2uFX6vsYMnFkzuWlazxR/
3HqC+oPbrpKBd8bFDuDh7+zk6heZ7oSWdwKTDLTEZUhd338TWD4xNy3purbGcN6y
T7iFrzE8ZDQ+0PGF44gYclTis2NinuacUoK0jHABIBWY5kznak0MnPNfXPIJcUoq
0GmD7+PyHlP/0tJXiRe2DiDOenyDAdbXmwJulnKNosBplYZUrxCUgVg0FONd0qks
2Q8KdKtmR5dyS+WKoOWdAi75yrtnc+33Mk+nHHkWC2sqFIx99DIVA0cemWeMlVAR
slfztqf4gkt24nvORgt0tOp0+IM577iOYTdwof44ReU1zAGClRHtfc6bjiFd5Gcr
r/uWDsChEENUhGI8Pjh7GYSBuuxCa1K97QV9p6npLCV6UN/yFrQpj2zcEAOnZiQg
lIelqlXeXji7apzoXZk69d0LPU0QJX7cOSfdRS3zhRM3fTJcCb8txVNeK/MiVc4t
h59OCXj4cokJXcVToL5DWMGsha1Tt1L0cj6fBEyuc9KCtLSAih8+hwOtL3EYHhHP
1qel67d/NWjG5Pld5u9MCLPsvWsTmDp5m4eSIk66IPkuJwfGMcecviD+gfS1pnH5
ttTK8oCbRAQWfyjMz0GUN00/1+A3zOs7QKwiT3+UhxuzOEaHVjs7iTgWzrpPF/sg
RzN4jhormI8dqE8vZ1z1gK0KlszHBFPm4IIU2t3p02NI4ZxZlfIK/+z1EvpXQ2Uh
fE+GYAtY+pgmf3tj6kdk0rm15adSqrsmaALpythiuVLFSP2awyMFVMl0f1AY0Hl5
nIEUStg8bKn6XJWTwBatXQwkvlrHCeYjDCdXSn5V5dQzamZfX69HJHJhKsv9756k
Ht5dBkdkxvsN3dfluFmlK/DkVAbTY/8/I2RljTgbA1kpVCbUuTIxqoMXTpoLOrtL
YpzcVeHf2NBHhkZmmE3yBEJlT0vkfKxiOkg/LL2/lMscGVB4HpaTKAaIiFqQGhLM
SVyeQDyxA2Ar828NU8VD+WOLD9AbBA1BbSrvkkk67HOUaJokV3llk5w4Ew/t0sxP
tdrw1hAMpz+Q/omOEf2fgUqSO/Lb/77CMMmj6hUvovdur7Xn8a1wmU1VPwIOnJ+D
rI1Mf3ZN4DxU0D9Nyh91WxNqNrLXzH18PcTmW/PPz+85lzTlfSouxjq5fNImIXSk
lTk4QPA7LtvXhDzA31VjH1BhoFTddX+OH6DEI6zT8LHF1bblqVtY8n4IB8Hp5G3d
P79yLYEfVRPs6t5N/ZFvU+7FJtaprPN5CWusx7GGm6Mo4aoNHF8il5HkXpCFNh4F
Ro5VaVotYysUd5/PqnYcZuU+6+yYnrMr8f45fwQoijXKtPVzTHqo7jenTd51Ed5d
EInFg+fPRxA2shzNDutmRUmFpHdBqXtnB/fwXsTCvCL7p2eIaLwlX9sDnRFg7ICE
y6rzP1MJw+jDmk/4rNVRyzA89TXiQ6WzKu5Kr2QCFP4B8xmIZ9E5bqBoB+gY5QZS
Dt3yTKuXEX4IGMX80jgNFpkrnsRrZm/8fjZy3O2OCX7P3PjyaRZInftbVMV52gyE
tZP6lei+3AWgSu0jRItapzr9qqzrEwNl6l+OmHcqzO0fJTUo8ds3hYql1wC7hzUD
hgL6GkYQfMzqrVDMGeQDSnxi7HhGwj5poq0+O0H//T8uloX6NAoqHWhDu1w9s6l3
Ihbdnqv3Jydz7xbUW1PceIL98rihMBiaiuDSlKkfCsU76qJvEaOxbqohvkkmbgfS
wBl3iVIVBKwl1RPAFC9FBm6W27RGr81aayJRmIthZgqCzUdxb15tV/bNrF6Vkucc
wvJsV4q1r7N+mmi5oL8GQSIUSOKGiTs4nIWSbDKoTcy6udp+zW06dMGZF7mZgMe7
QTqB7L/R01nptFyvihm5ASuv8qgIwD/UAt1QbGH/x5vu6eo+W2lVu2gJikorQC/o
i21qMKA85iTie+vSLldZLnuw0P9973dIzX0VMImyS9M9dOyxEIVhe1Can4Em7kbC
w9wKJZWYRY5FpwLTG6emQ6VLNUSyg+YFUACC5Y2EwZxLZJUoGudeQrB4BtWCWmMP
PRKvsAUf4B4/pdt+fOWXUkpjIWRfOBghV2VQH34O25F66qMPvsIXJNtHic7m9fZy
En6xwJuR1SrFZCa+QD46042QGf2WaL8wojTBfIGYHAuY1buc15xTPajcXAeV7BQO
YiXwBHQL5vqpV8+TC7b18odONECi79q4SXQbq0rMsnYDmwhLFZwlMA92u8JGx9vH
TNNYQI2M8L07APxS9lz5b6Y+WcAxTQFHHVNE7B9acrnKq6oPUPY9jUR2poOhPEpz
FfKMrNxOM/BtGZfdcGFHsK18Qp9YNLcgT35jboNYiAsUqGW7VnbCh4en1ZsCVV3p
N12N7mP9SVS9ijW48Nf6/XMuy9Fq75Vg8vreK6sW5OfB6wIkPd1xiU7NyhoPg8yK
ogUrPgi+alItlwJeU8FD2laKE9E4/kXedtn9MImP+gdp0oGZVfmszA+wAPftL5m5
lgUapA3eCyvu35iIH/v2SPj6SYdYR7uM3QcXTyKRB7r4So5MYw3i4atSHvOOqryy
tou5sUQ7nMG6DoxS63VENkIBAzL19trZ6YNyTLMyE3a3tVhg2XhQPe75L+Iwu+BG
uXKwzY6M1ygXY2dn5IyhZ2tZuV1q9GmStxb8isbvKBX95Smrk+b0sfrdyVpsBNtT
Sz+Keoe4Ab3cuhOmuGS3/Pgo8yWCYTxEOQDS6xY+sAGUGOm+DCZxwxFMXLl5vGT4
5Pi+iifOBGNHjygeR42ID+GnTT8TwccgYLmIRSuBFO/T/rBsrTieO6/nWOZvpba7
pvu8W9c0gmTkdTz2LqhqIDZQqwfVKWoVVewznEN9AHeeAsupH+l2aB3ME24SesWc
4PQAxwq+ZqpJDeXN/EKxiWrdYFS59WN7BpTxpD88jRQAExSRBMjU1WdrQcCmX7ly
TxTdF+ELHxji3gbcwjkcQ1E6HBJypzw8VB5Ue1GJtC0AZsntMFcJUp1I2YkPLWjv
9nlLW+aoCPscuJpPKjMxOMjw97Bb4XFBCIdQISHXPKGnap8KBaEMoQYdH2o5AcVv
mBPAXGJUCcHrQt9Yj596WWRmFsU5Fk1d66Ako112zwZyxiSLWrmWfPiJZlNbOi5F
r84BPvQRPlx6iqkvvdyhy5wRvQOX8ah1eHpH5+n6MJMEOEMO84g5EKUnEG/3zW1f
fAWYMydAp9EeM6U0zbMqDK5/pzy8dJU9Jju2IJ2mv2E2EKokWaQQFpLVOEflTi/p
E42Q/hs9p+O60Ql025grr3wBz7y0vrrXX6XZHjPVLVUisvBwS1v4kh9zc4q4N/jk
O+fSD0copkgvvb4IT33oZmmZgkSsIXwoQN+c0qKr8Ip+86kaJJe1rb/QGmJKTYpM
SLeOG3DSWJyLdasgATxKY3baH3keCTih7exJl7fD5y6x7PL1Fz6slGk7alDfUQuZ
/wiLLBKRFMftlkQOvpZVFQLtL+n7oLUTZzVZHLZPOeQiuoDb3NFeZt2XnHjRcFQ2
T8UgEV150hrT0+Zo6S4A96hVtCmowhDiF1gzKLVuBWPqAr2Br4LyLloV+/pfbbPE
doDl+bEwFCVvF0vkScsxQGvFDTSqLRZtJVL2COOYQgeno21vo0I+arowjBQiruJD
xx0gTdy5QxkZqWTkKvPpBq8cLzmqaD/rlaOi7hJdldSz9Uuh1yA5zOiplD0qKgku
ATUMsMEJm+IGR+g0/MEqp2UDrtnZ6yWStILYGp+Z540vvFeLeF2WkIGxKoDXOQLu
/PLz49bYTTr1fCFwfQwr04GASD7yITUZDtHRgnt+o8nSD7kn0y9dCiqMZiUJLRzi
JQruoMoxAVtqxF3HK2yO0pBu2+TF8KfEdENekiaXvgmCD9FmngVWGvdXj+2W42VL
k+nd1/87zdUnL/a0By38v9Flyp4M1nrysNJ7D7T4csPIucgpnwU+yUji4NK08eGw
AdGI3GGd4z8DGiwJf/L8zi9/AlWaVNMePgMkHdNfMQSgElk2Solzf/zpovQjwgCY
4rRxLSWdlfhI9ioaYqSUSzFD8F7ZI4qC4iCYVtcfK0QOXZhnTq8IBx8u2Y8b1F3Q
m7ybUV91CerbJMmqVmQqytw/K14geHwfnlcr7phplxfKgOOmbfLUTZpMeaPWTIvE
YidCJO3jdpw4vemMAK6vgDFcn97hT5fNr9gyjaAdAt4i0FP4QYF3BImgtgAH3InP
oFredcGojIzsKVSv4vZlq3epaCTX9nq4+ua8qQFsfx5I4m3QbeTzQOZrTXNNvmgl
1BBlrNZdRZUHWf5+vX5Vl6XVDlcXXgFOwdCzunm//b4MP2AGPD4oxJM+QFiScrX6
3uUWChb1ZvMz7tKmeg6j79z9zkTUBJ/OTEv4Rat0KbCMGR4AW6vg1dIYpXPpSKsv
+7Z1eVD5rKFV7bxp703gdKP/xqsibtdJoCF1hlkGYqG4CWWP77cUZrRi71mW+20N
lWRAtQs8GD80bRlF+JlQlMh9Dwl8Nm0I27eyti6W1jz4G5HgF/AiFK5oH+zwqjws
ogjoqxXu4MFgi7KfAv0mqZsSdf+Ipf74hQJB5ABi/f/XbkN8UTkst6lj2CKpJRJf
ao+vRanP9RS6oiUX1/Xx9td6MLJVdiNZixypxBkE7XrjroEHjrKPNfXE52ALy+e9
CqdemZTc5Fq9bO6sO5iI3vxJ77u+t5BOb/F6+ZKTTdzPVrKXEZN3hwsTsOGJ9d4C
fSh1mh08KrCp+SiZ/wmwDtJEw2ZBBe2Qa+NHAmtKbz0zPPoNu3Clddd77apjJYd0
gJsuExbYL68FNbim1TE0xlscsHrR0DLiE7Kq332LQwE3jLZa6ixHpvq5XSiKIdZQ
W+hg9LLhhYUr7WuFyTJewwj6VzFIVKf3SjEhna9nI6XaB4EOWVJCTRNTBKlnkQM/
QazROl1vseYrQkZKughsaGJwcM0PGfXYTj7U0Ou9Y6eR7lSifvTcSIqmjcRQ7PpJ
LJmi+6MUfjUhg5BY4lMN6PKysFENG/5wAGLRqMEoI0gj8iXnMALj4qGnZPj15rJt
vydCqx+xhmKidz/I1yqlmYhvx8Ba1kKaqJUVvceBRh3FDcac8fFkZQyslxxkvn7U
XOUXiyInabn+Zvoxc22mzBZa7tusPnf8FyQWvvkbmh82H0H2PSxcRZpHmxEBiu5P
vMlF0Q84KWfj2k3gMffAWy4S03oRgNXRXO9h3w5v1POansb3Wr3Rkqb8r5msqZWD
kAd1SNp6Yl+S0v91l7ihGKBv08b5q3FpxKHswby24vC9IPobfZnDEKnJT5IzZi7k
46tf6aZQ0Bg6SLTDEJJ5ZnvrG/871IoC5S2HPbxgyLqjV860eQmQA0LnMXiZa5qC
qwXWeDfqWR6O+NM95LM1tgHFf4jQbYouDmpLQU5N1EE9OFYm8JRP6ec+wXIJBaUG
ZgNxy7o6SQwB+HbN84DrjHKFSRlr4d5IweC+oKYfaTP7TCeSTfiSjzK/ZsdMT/E2
eeCiEDSPNeJUc0uTIBgXhrvQNpQRItXe8m5QTpRor68HCUMSpZNqcRcUR/sgiUXf
vGMRpTUDgUTNdNbENdzw4sZW+sqXnXnSDfKULpfgQ/B9uhbRWA0mH+ixJIOwY79k
bDDssgkUJTzitYOy5Jdw9mkVlaJD0UFgYUCB0V/2sTxANbrgMUPpBAqj4aj1NWyx
I2JXsPP1N/TLpK2Q3sHqD4aFNJXMHkfHAj88/E4DrZsPZTC3k0xwpSSDx9c/G7sR
htzPPlKce0BEuSGo/kMobPD8Dmr5jqsW7+z42a3s4u3zWm0WnqzG9KMoSzg7ikFb
2S5Jf165A1MePCIb0YUBTNPJha1H4wfnZ4jX0AUwKhA5KSnGNshDkr709+OI10sN
DSQRj2fFcUMJjGl3m0CaARTm5cpfXtiiwdfyyng9UWnzIn/jK4kFN7FsEU7OsRdh
yzE2bLB7VxWy8QQWU32poG7shTt3HU5u/cYnwn5DCuW8hlF5DrYvl6DtSjwXu+dP
JcrX1I5RkFm4lppig+msAW7t4OEba2980N0Kx9gQsoyi1zvkPQCou+YF5Wn8y0OO
FAN5M7LbJh6+0rBzRFKh4PPFXoLfpJKJnYYj/CLqL6oJ31QT7NmZcvGq19wsk/0w
/clyR7nBdq1g0XDDQOK9CmgOyk9SJmAG5RlgzFYhPJVQAKy8x9jfp68lAhAs1GIK
KbzIWMqxbdNke3AxU4cQ7NzeikCk3sKBAh0bTXnx2PZnfQNFTdLg+wrCFtIj8kOd
Me7/ju2RCfaacqlHUwdnpAilc2pHwR9Td8QU46l1LLKkyQy6sZouhWW/p85pEZDY
F6cwiql+BY1azFUgB0LS5iuD5+mE8T43uK9HQzIdJeE3Ql6jsfSJOHxXCaiMM9an
VIgCj1qUcvgHT9Q1sIFspHldu/40SXLL/h5kye4d7IKQJgBm0TKunmyEMAScCqDD
E1Jz0s1GHciRrqG+3lGGTuFgKDervscpgdafzQAMQjV4YulRtVbN1diTnEYPA034
OJm32ZX13k6vaVy1fNfkgCO/63tbZkPf7KSByL1Wq9RNYimJuCgl6+FQkzztwqS7
P7QwVvxyNr2JLBssOaaJ+hE7IEIi6G00CnmLPx63l3jBpTB2ISJmtjKEgMmymDSX
KcWWfByYiChphu8D57iabu2GDiqb0M1i87F7O38SLheE3zlyI+Cqf8tFkC4l8Kt9
kvUhWCbJFHkHpYzMKMdGV7VHDtSocxG1Vv456gFzxX+77KVVKrPMIhlkikt/jDeD
5oWvYtcNB3Qt+4OvdIEo8LX2iIWjPj/aSQQCIRWqkJmgAzKVpyumOuvogYXLS8Yk
V7NGzRxYICssULRAcFtjS9lNhlt99N9JuW2D/wog5rbWGF9uKmYO9Y8XCS70GQDg
iFJX32eq8PlrpDBJj3Qo7spClc7W+9VMkytTG+NBNe2aQSCx3QI5kf3wQK8t4hcu
HY///+DVmgAhmvc8ngLwhn6a167tzL47ecyCzNwkPqIjgyiPz+DUG6NDY8M2Ccub
DLWUjOI3NNuQXh0gMPHvBR8GwDP5Exzj0/Am68rttSuHWFN6YHwvXXe8/vEmQtwJ
oOsDXnq9pPARCwQGlpXWLZ1KZr5F/d63t6kRZWE2LwEbwWGyfOoQKlYkQ0UOr+Zn
WXsM/PxSU+HvpPv3MNeSS0J1n9pZHyk1/HTqtDMiZXLOHc+uOK/QDqg/GGuMPqF0
JXwglnCQIGl/x62kki9Ec0YMRpC+A/HQvMpPfiZtyowtgfKz8JRCVYo4DbFsBA1O
E6jWfRSc4rn1h/wQe+jg3IB2I7h7za7ATO4kNEwOcbS2+xKJWC91kIrOHJfjzCWs
vnnTFlqclpjmma0o25bSw8lT8z4/DF6mWZbNvFqG68tK1HUdirthW9lrGb8jhNdO
2N8pOSNuNi9Vg2mTfpWLCkB29dnIsOonvMmKu9fVcBEKmQ7AMGhPViL83mIEHt6L
/Spu54TJ7rGDUnSFkBKKl8A4I65mDC6aYs0Sz6RGeujvtranvd5aIrN+gHHBSdLE
odSrydbKPk5c8YyNL+wS0hC21io0+Nw6HOI7uhR37UxSnOdzbY3iZBYlM9lJbgB5
7kprYxJcZJnDsh5Y9OUaVGkOYl7Yoq/mMIM6QpknyjAB3wfGUZISzG61ecGIY4d4
fYgwXqt27GL/bCUlwhZDTTyi21Zkt360HfNlU4k7TiJVX2byvJw9P/j8tfgVklbu
e/iPi2D3pU3UYDPimRTjO1k+NWGxZQOZw+skWsIvfJvQpGcn8X3MlITfSqD3sW09
KpPsIB9l4EK6dVqwFaGVvKgGeDcbjnc/RSr9cm55nK8ud53YuDs+/9vXpEWfaGKa
9P+vM+s2SGl60EFP1UiIAcksoKvoWEuVZ71flZkc7AOM2p+uyhHFJOu6lHoLgUt/
fX+zWQJzsE7TsbXodksOZj7EyflG3qpB7/Ou6mar+X3D0H7pViDDjngxvgOCY+Tp
+ZpIRxXCGIkHBrpeoyy6MrMsheTAGCtnjMsdKF/GNXb82EUtQCRqr8l7pBb5Di5z
DWXmNSjsE/KG+sy1ytoJJY4IjEFPVAMTXq4/SJ5NWuvT7FbZBoJr9WNY/zRluO1e
Vxo3SpzA8pW07UGRnVOt0B+MAO56MTtGYfz0WSzmxoGxj5UQv/phvquagfjtDygW
4K1APZkr/tbWQnV5PqjvLqssPm4alnXbXVAdwhesHEqpPrP7nOq7uDRzTd124PUJ
6+fr7RFim813s0KHrdIn0D1ZhM7Zs9DuxlIP1Rc1D78sPyRDQO7TXDuOnh/0235b
w89Gd3zRKs8DU1Is+ZP+B5cAc/HzHU4D3YPgefY4Q3UAoyiHIQzI+ScI58HN7t32
xup9pg8mivvtSCMvqkxfTq8WqdYl9UKO/MVWiAMBMDU=
--pragma protect end_data_block
--pragma protect digest_block
1xa/lYbwkbD542YJ2WFyJcNqZq0=
--pragma protect end_digest_block
--pragma protect end_protected
