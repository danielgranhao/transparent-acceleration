-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
lPQJqXwxJgw6d/GqWjYY9sAf9UIJsIoFI+pQO7UBdylm+7J35OHutudtlK9mzO2JxUjpCFuuIr5u
81ualpx4fdc+Qpl2MfNfGx0zQoEnjOVdn73IiapreKvJ8nGOpaOymcskppYHgQEw2Wat8EuAMal4
pfTRihRKQK2m8QSz9BLycIJmV7rNnPVaoD4uqcNpTWqxb51k26CSyLE9wJ8t6QRjr1I+3ils3Xv1
Eo7pF76U+H9E7jFFu0h2VaLw2h3JNj0T4Q3H7PHu/rwEpAHNJGGt35iT7JNdzR+ZYpZFQjIhSgja
74lfCDTyF/isUdkkehaZ3Wwb2Hat5+QEmqVABg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4288)
`protect data_block
WW7QIOJ953C86GaKWe1IMzGWyrHuSw7iHV66zFgYJSzvm3a9DSI8HEvikA1Nkr2Bwpr6DmPqcMlS
bbvYKRn1/uhBkdf+NCk7WJbGdM5bdgofbdYoDadd3xk3mE1dPJgcQC3aTphY3St82DzLi9e2y5yl
pBjR3MLZ5Qz2VQfmPKP5xbOLEJ2YR05ARocVFTAjDxeACbysOaT+u/LUZ/4Mteb+4T3KgI5GPnVS
N1oJ8HtvG8x7//egZDf/SU/vcHh9/REl8pWgHbxqbW11NLqhpTSKYWK7f0XvmMdGFco1zJUPQD0S
AO8xNHpucrp1tIZF0Kx3BE6g3Tl0PPvgrQF283imio0nm5pYof/k0jbcnwi1iW6dCQPJpveppqJn
/DFUXguaN5I/Z7SQDUmjSvYKZ2IMZkJqmS+dHImHMRyA09x2FFsqieK5zTHc6e9UFXue1Voq49zz
qxtz7z+SRPzLtyfW5qG/TDD3R4M/lR0VdC4OpgnionHjy6zj/i44q1p9au8lAIjGAzj46NSiNckB
l3m4XHXgixQLAAi7o83cY3vuQ7L3bcWGu7tKNxWOSgtDjOElXOvx795sDbVslkvvcC+p2U9RLE4E
SQ4ObxTzORcgocK4da6pbtXwXfGo6N6n7LPCmUJR5IYFLaeXfrM4Yh9EYgSHkn3VPVryRraqg3cM
/hQiwm0PWC8KBSrhUGiT52weE47WQ7RiZk71s7HWjF4JBccqid/UHdhFMh7KneMASZk9wTZfiBCd
rNut+bWe/Yr3O05i9Kihg7D95Il0LKZw+xhvflk/XH2jYw83WS715K2Sbh6PESuFKEHqb8Y3+GU0
Wfv5EI8LXHMi9Vl2iYTK4ZKwqzVfOAt2GJ1UPNSNykiGfilbVxr6EKOJhBkafT7+BHFlavuNseHp
I6fArT+D4eBrRmNLIMYl/6Qpl9+ivlOtnp/aN+nhcYm+DAwDv52Auo9tUhZ0EbizlnF6ij6yR31Z
Kz1AcF1qxXvzy0QmwHHKspbLQqhxwlym3OyII+OkQD/JOexIiTwIznup7PB0w3Z05U0OP/0PT/5n
q3KV5/RGzDzDC6VERAM4AyHlV0zIoxxpNrzT0TDXXntOjtjZHpU/0ROmBXBjzsCJarUGsMsAiN4u
InvWzHS8LU/3tXBUKGQkl9uJb8IIQL7so+8txJZUScvjWv8m4kI2dweci7hbFak0uE7ZFTD9WnS0
eD2G2uYILJgvNgUfv9Y/9Ov5mO06G83nGM4SqgY2TuNk9PXyOJHLk3SvUm4z6oiZofGPzULf0eGB
c7gPj381D4/O0jZIQg6x3Pr7f1OZWqmgA1WI/4SL+B+lVC1UcpxsEhadRpUe9nnSnaunobULXYg7
IAPKREYMBfSoMijO9c1m1VNrd6CjnO3H/qS1AENrNTAShA/AFX4JiXv9k6ZdafebFf/RL/eERZw/
Vtl3KaChwVQFWfz0imiw6r7Nsh30pX2i2Di7bigiuZitKihhIyFMM+wmJtf46d0glKvGjjufDXsj
0fcDhYf6QKhgWsHJPICrdFaytpbpGvqvlsa3l0aRV3rkff0nR0+8732PZkyFFamaQaODF+VI1h/K
P+j8G+QEqmes57+kO5pL1V+otxTGId36SQxXGF172Pr/mmkfaYu2bcZKYNKLaNS2ya0SvlCkh293
IYSnePkBsrXoy8K1gb6SbpmT2Jc5Zo0S++xGniXtW0M1aIgy5cFCxTtOsULw8HEYJfo2M4wCymjk
8iHcRpeEfr8xjKgelm+5ZU7mwMxcTkv5TVYDzwOzKfU/2vzcHn1/1BEkwt1DQbRChVGxOZD+wbsL
h1UDWj0CkshohYKnIPEao5hVXGm2V+eJWIZrYAcmBVdHi74MAoZwQpdovJ/gZQGTe0RX3rDBSmHn
+G6x5svPhUZ9hQTkyfohKKYF4pW4Ix3phEDo59zB2UZnUe1ixhvT9xSfO7Tm9ZNQgdKwmpBz8sXz
QY42ZPq+nPaVadCovysw1XdnlJ9rXYiYawPYO9NcAHCYu4cQWhhDHdLOqBeuri/GkE6iJGFkZtj2
CSYJAtyDuWt9bWqzSzVPg35Q6b1luwsmriuo0Q/pvCsd1WphbyG2cFdLWcuyvhCHmDHV/eMJwruP
rskU/o/+zFcF/QpxylUgHBk6A/0QhKI65GAPCIMvmWkdVwjMTBDMxFYUY3xOQKM8wGtR5YM1ZlQO
/dhqAktL09YI6iqePsuJklJROrwyzcTvGhL3ny5ZVURYKr/Gf0IlC+AD1VomKOV9oKB3Nm2lO/mT
s8Foa/G6mEcIypGusHB9c6fc3pYslhwM8Q/h1Fkrpmm7mBjspW6vDMso+tjs8etnWvlJOL+tCOeX
t85fsE0J1lqLW3ToRj6Dkgw579MnpWwu9mHqjWJtFOmJeT8tB76sonvBcOOgcGxzG6DuuF2EtH5Q
SttmpTbgfqxJwKQGBRYsiTS8aKItPFZMaQoiMvDZ/e+Ztb5QgHrLFzdUm4Wj6HlHH0wC3dQe8TD/
utf/MpO4cQZLoY1p0eZZxDvqazhQwG+Vik+fidlS4BZmRCNiuM0A5LUYvXepqwnBQxZEDNfN5+HR
MVFLfpoj5XOwn8lnDkx+jZUuF8/EYPp8ptYpp0vgIb1lCKDu9AOTeGth3LRHm0ok6lWNCR4E2xqM
UGxFtEdQzley0XDdZmTn0Nokgg9dQKCtpyrMMPn+MqNHSMOVvz31ADoCSSv3Rr1XyOAWwHHI2U/q
gKjbQv7Q+gyowtEW8j0cYRazItYoRTq0UnJacHhlBx2RcOhM/OOAim8Dqq+y5/v5/soMvQCEMNu1
oRC43ax5mjl9xyHCOw6pYk5odsTzuSehVgZi+gW+EvBhNXrN2d8RxyZbM1ixS2hZYArYhw5BDLCQ
wQjU8opM5fEX4KPSi86EQ+CBcQ2v4PtK9wr/kuFkHj9i8bRYy3FoJ7zowj51M6WETSojujMzzuaf
y6b1jps1Wy9wqW5Jazx5U9TygGKoA0U0bfnGmJOIWGmT3dj0z0QmX0BdadsxuEHQq8FWiGprN3IH
7bfk+vRvspypPN0ikUs/a/4gCVOs9A3qGFZEyCBTK3xgcrJs0BJnLkj6jFjcybcH0Dk75Cq+t1gy
ZUOeS5P5Rvsb410v0UJyaj+zQUelKIQdB0yCPRiQIr07LfPFfh/gRwLPu1Fo4esyoJGc7dtgyLPd
chvzIWMz1kmc4k2i/rqAgt/yPHMHJSDOVpYu4xSLX9x0ujvh8emL6x4fhDDa/48kvRPUHxLbLelw
d5Bav1A++nlyFxthOZMiQ1R+eXxqtGXyHiGTXY51e5XR8+1sUkO4dMnYFsZJ8YGLSAbXhE3pJJ7g
rQ8kPhmc2yezofMRvfFx/4KgOZlIflkqBbGalxVYd/6YOOfenjjqDkg7zKvz8I98AUNZ0j+3rZiJ
XUygh3yfEJe5Yr/y179njGmHcuJeS9FXdcDQEqHxOZNynzs2iOXnvAg1crPkcKyT06TXaNfF7Zib
ILgf8DFaryjpj9dYw+n2KafbcB1vKQfpfxxXH1mE8Mthhw5Dos5WXaDxEkXx9LSAk7z+Wc7CBATc
xnqYuNOo7EV+EnDCZ/Izef69mOEDpoexqbeRCE3F3JCw7JrwbOwtyiverF6yog/OsxFHWHkCByQd
MIlPz4H/IlYBfA26vSSuCarZ9r+8t2/v5oUTDZSNxnjJ5yaf1NjLEHcghzotr7sev+YZFP8ygg8q
uzK+WnKqXLFoLgCwlzB4hPfvenPBKaIWPrFlC1c58D+ELKypdFIv1HzIHIBOGXq/9JbSxNA69vNI
RX3hVSCo18DgAONP5dP/rOgn5YMxQcoU2Laox9/1PFOz6nSomOZt5TaxZX+etSg5veoZS5THrG3C
zARHS79KRIcGITStg4qO8PGc8lsVe9op+vSrQbkORlczffdyZ17DUB6alRFtrom6UgiUsDBw7+Ak
RDfo47Hv26YK9ENDlcWWCHk2u6WOanVeoHoqPDBL5i8mzWCwqsa0YfnKb5cAurAyciFzRBFeDowl
gFaeBnezhEeZGnfthAA/l/93KdI4C5WlK4EHIgLbwi0fEpUGHBM/hwmXg5dzky2mhOyHlr7XP8yU
OQPeodVWOQsec1NHIqUAeeWnVEiM3o0ixZth7PNHwn8a36F0oCbp5VZnk6cyqzBhdAqjbIU9UmSk
TAaYJGhx7gsRApRdL/HgXn5a2Sj+t+5LzmJ3cZ3U0fe1HQi2oWd1LqimRJ7KwUqYJ/01R2MoQLLH
RypzTw56sr8pShL0miQZXGSpP2TACTiWsvHEvZBMFFHUVQXq/X5vKLM6kRr2P+pvxumPW4hTAEG4
rBYUE7A2KRgdRO/Gpax1oHkGuNLVxFpA+p6Focc1vuJm5l9LlQr4KpnZjXlEzrTL/rOyT/273avD
JuFzCJ8IKiWI71gZgxrpzZzsrqoYiJ9W+iBqhafOxA0GgWvVebWw8ClWKJK3hh+x0yNjwRSQuhMU
b6uqlmobp6FYzw4Dvax0GHBv42HznCJA+ZpVZcYaXwaHwa091kKxEP2u3XiQOxfI56QFvPcjfyxO
2lr2EGFSUfhUYDxKi7cXNl8Joap0vfrVHfWFbTzV1hNQG0o3oPpqnfWsHYltJi9HC7QbkWSTmoGa
In+3+DjI3a8GOfo1LBuDMFgQCpaLzxTvwWPeusUsENvtyRGOJDHPwuvPEHmtgfnAk62cYyod+Xlp
nq0d45PIXD4HszMZ4+trOz+AvU8za+6BVsjao4yEwdmtCOSnKB49Dk1ORJo4jXYwzAjutf28zDA2
vDZcT1n+YPyKamr55Hr/gAZj2CVxJwurVvcveel6w5+8pqKSGZhs9MGJlfPhpC/cVxD8PSI1PxXQ
3Ok0CTpjAPx7yEI1rxVZzUqfhETzmoFSmttoTSd5TOvbZVj+UeXRkrgfyPPjddJC8lxestrDyoq7
xD0Ro0J8xXNYhIfoJ9otHeufAGJ1puKD21vGOngTBb/VJcuam9wDwm6TrkaDNTL01PUq0I9o8bpn
0bae4BDkvozcRx4mBA3AQmVJgCp0LDf8AHQ7gW4B7ilyRlB5sLgJlM6O/Abxx+ACgbOXnWZKuCt7
MXB/OnTCkq/UkCWWf8Vv1hiXUMStmxpQtApt4spe272wGRBvYuEz9LuPIHQYVkWnrpYPNpkDEn71
PgY5YTiDJ6yz8v91LPtbcHh2Pqg8hxO+/Jr19ptbWspjt2oyRTnRLO8l8d0ZjHwi0JaDxzRJo1Qx
snsSKK8o+QeoJwuQIP540fRHGfRl0BvxwhPWcyUtlTOA1/iuTEfAYZP0TosnHm7intmvhOc10eE2
lwTKJKLeTcf5Z+u3T1FWzZkWyikRIUJWksSD7+exZlylnJjgnHZzCsPpcARoZp4bCwRpCEcfsWvB
9RArduB9nt0IIIi5q+Donvh39yry65JH9zm/00lh/H2j0w8DADOYP8Lh54O8SFWk6hC1/jtEardP
BhBxizSa2zQMgNfuy2i1okI3/0w9MgXrpCQpZUU598mb0bLtJTPM7+mJqyTwJC9/DpY1fZwz5PSx
w+xDgGfJDWoqvMJ4pvYV02Njq5gF6TK+GddX54zG7xK3ULmj/e4UFZAuqpPR2s81fwWJIQjeM25y
uzycgSfHCqZlgoyFFoB7nIurs4/hRkPJCALazQdb47vDVLwoCGWxR7Xn+K409uxbijCx0inq8UuT
w99JBvUe95RCMgdSxg==
`protect end_protected
