-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
U1rs4oApcp7tIJDvXkpcAfLFFdPkQxaCWkzIDaxXiNUpjHiiFCX2IA/IhMb7xwaY
XrEBXj+tq4LLrNJzpRMVur4zsShLFOZnssTD5hk1cSuNg85r0ETjjMod9RYRP2nJ
rHfD2ykLiVLJqAR2zmH453LWXipY+fxgYKg2FbF664I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13219)

`protect DATA_BLOCK
s8sqSRhwRQALi+0b2j6VHx6jiCSSRyy/hQfbTKhnKXF4yYbfydaLhr2pSy+up7k+
9JFp/Opz5SGKCd3REIwM9M4Bmi4lIS6/pwH2w3NYg4npFJthL9Dd4IkMv29y5Q4x
Jxnk3Vb2nWN307eN+PtrFb8OBooF2EoMSwgY6r8lUnC/BA8V3jVJQY8mJ5Z1BNWN
i8VJd/qq2P0d7GbFF0f9Q2tIZi8TUQqMg2cRX34bMLJScnOqYVAcwoigyDanTTlE
Zwbx5J4f1uIpKpWfZwXKHfiBy/hOX86EUJPg4mZv1X9pU074Vi8IAnw1ZSWEBGVp
LVY1mv1FNIRl9ypVv8HkvaQQcvzTqEU179Zu3nYN2mQ0kAWCphsGiXVGZ1iDJ0dp
yMg+YrbNeUjMHvODxmKBZeBEHjnJlbMP0madZeP773k1Ua4xyhLvDCz/CVz4uwVW
v/+ihKiPtylp5sUiUH/Zca1YeMatHPxxeqjrFmU8UUhuj2jL+XCYzU14HPSOlB7R
+7MUEAP9CiHrjcLOGww8P/LbT77VJ5kuSiph5opjbu0YnwUUB6ZiUqHhhCvwTeSa
0nv3ZgIsKcsMBNEM84oDvjEicM4egVuGnLoM/GIgRtQwc8oc3lyJXDIa9Yd9bVhI
Uz5M9vSAmWMIR+4JrW6A0qlghmp9fdgiFVUhEYyEjoX+M6Uuy6DfSMI7lTPyb7mb
/WBOEls2/xp70X35hewwCcGyekzA3rZVDg5dtPNcUctbeZ9TiUxdAm6wsmUHe/Q6
czYA5j8eHitMWE0ZDJAME7KqoFOMPwWCdaVEl0KT5YiIt5VDSQeyvPdMO/JuMkbo
qB0zSglO4pWqvXlcWz2SetrosNkLnwSvG2QBm3sgIwFHXI3JjNdiO0kAqvipyUYU
KcjmYQay0PhGwecc8+Z56pwFSblrYaT5hBP/fiZ0KiJUvveYMhT06ctzpgPRf3WA
FSgijCAKAqYydZECrho3PGLTxDwleHzI4mj8z8c24++Fq48InqzRzOrh6Uv/HKwY
n8df1UXBbTe8ossX4+C/m3QZkqNbdQ6Qz54XKryOrggJpmJB5Bj52KCXEtpVhV+w
3aWSmuxmT8qDVvL+fkhiNjv2cJt/QpYgb/dBNwj9ya5kJL01UCshVNJDdmkRn7qe
se2kRvg3LfI5j+0JC2uS3gb/J3O5pK4JezqXTR5sDk1NagjT/U5swj+5bS+jZsjW
/ttIAAdERFGbsOdZAP7fe8RP/bn3XcKtr1XPtDAtWuX/SwHnob7fjq2Oof4MzJLS
4O/Jrju3C8k118h7QkmcS+M90UNOXuqbB6zLShHM/MitRfLDg10ULBqghmeYkQrn
WAAY9YUyzVKwb6SqKBdaNDX0wUeE21G8hv2FqbOaMSirZisxhqSJdC+ahJSjvx+k
7Pt7mDfNbKJa1oZF77oRZ/Smi2De2vMMYt2MBsiJqhhoVJl5d7jB29CW2p0kPzmQ
2Z9IftuoASPzK8AcBU8MICfCn7STnZHXxo12gR+M/4Z2VPjbhEb0HQwIW3+oK8hO
xn/akkFz5ZMx1gAVnpVHHpRGodcn0B/S8pwhT6qumdY8ZHMISrJe2Bx7lesGsQod
dCNNaCcA7qH1VcMxm+VoCI54DX4vp99j61pzYiYg+Zj0F+sHUfIJ8sP6DPDx0vdp
7sq4mY/S09TWy4LOzY4pnYCC6aEV2WfL4eqgfnklDrNDhmYB8sH+mYqW+hBPWAdA
6ebJ2UFoWr3iYEKO2VpN9AYqIvG4CAcRSAnU4DInm3pN6PIqBkDOnDrc40otyiyq
UuuPaRMFam+bnh6syouTUNRz3oXMB+Gi4LqboCe8O8PAejgnkhsrLWyfc5Tk5LlW
FL+QsTLzQzzN8a3ULqDZZvu1cjQ0RN6R/W/weVMjKBpnY/jJSBR7H8cB/pZvZXm6
yIaW76XADlvuhCm7apxavFCuDxwkOAXN1T1yThdB1PE3IlRGNh09NMztF6ol+zDc
REsh1yY78kULBtXx2fBKtFeNhiQeUQ4wjnoijJSYwJqsu2QMImcAIP8AnFrwn+5P
oII3nMzQ81TEISxvQJWL9gTqWxsg2G7S58DUi8LERvohJugO7eh680dhHLRn9F9Q
bVM4MUhfpc8QKA2qI+nJWGq40svfuJulQ+lAYLSD1sRCqg3kzWI6dAauw2kRaENv
3rfMRC3sIUNjyVjyPVa7yCfxAuWuN4P1/B0dLYNvnbdeNnsZ0+VwgorajhhoUVi+
uTct9GqjQa/tjpHrPu3BTdmmZ1sgvnuZLddAHWnYh7iLlAne14J860e36H0cS74Q
JzhL9g/6tvEdn/5ULlIYbRMW7bY65geTw0I/kexlscgsa2r61VlcH0QoEtqNctOd
9zymJvxiw5V56gyGwIlhXOdCZFqqRymzMH0TmV4kAUJ62s4RoOVIIVPj53VpvHgw
loELaPVtZm3zJDCUr+BvWPT6hYXRscZMCltDJNvl3N55Oe+FhU1JHXJ/VzUFIFZa
lbvVUSXfihnLWYVpbIXc+u6bonM0Do9/65wwz2Xg/9mbowsnv7h9NKEh9+P/P834
h1+nIOECHF/WR4hHWLYT6/2s9ZTil4SfKeCq/8UyC7pR49gXiY6efolFrVOWDLJm
RELA28lBMHlIH7SrrNkxj5/qIf4R+UlnK8z3C1c4WvqrUnBiDzfr83FKkorZH8y2
VtSRZ6EOLw+BXml8PcwPKuIZF3wMVuCwRnyCGIvDK06Ybmq9LslTX8lPL3L82+xi
kHK6HF6qZFMiwHNBtG5zpQF/lj8RF43ot0nRnk8SD9Vj6Z8L5BIZHCIDRgp/GmlS
bpFmmyCANFm36B+u5Vlh6xefOLnGaYRlt8eoAbsCxtzGAXOk+d2drWnkoWK9EVzq
V9k/HxrZyAw29R7pRHWynjQuw5PYowfdzYm1avsTosR3DNkIFAcpZ4TXqA081ZlU
6fjm5T4cAmEbZLB+4kY3xLaJMDvdC/ysjvsZtp7qGTHkGo6dLWzmCDlfWwTEuqsw
3KKRItUaczwWJ/iwxFChWeazzaG2Z2m+NiCsRbO7v8JyFRNkCqlTe4O6p8WA3m9b
RZymGPzF9hZvJxCo3zp4iCcWxSmw19yoioiYSgNwBRYOTMR+em6MYFY9sO+T3khY
9oEGFtoxjKfytztTqGg+UL96EOHo2wksDe+t376deu37rdEcCd2cvpnEV955ISKm
0wJQBhKxgB4pzBjfBZXRUyxgBp5cM0OBhr4uBR1M58o7FCpahGiv+AMaLgzc3Osj
VZVSn92RggTqC6MpwdkPZgGJFjzptURvUeW2k18lrVgbqJm+rCy19mzy/dL6irTY
yML8+MqLoZiNKYjGjkmi/uLE9ptfoMpuxuDOtrOg/j1F2YuOF3VzZ5kpbifTsIaE
fyNSSdV4O344zX6kPDDNLwbRrAQB8BSzUgaSrMMf5uoukjl3V0QtJX95YgpXmXsH
RenY365NgEV3xkCDAE6kGa4gbRuzRuml7mIXyK7iNKHt1jkh2n+sH0FGwA1PAWjU
A9cV6VWPi7JyANh5PosQv4DzX89NHP/YE6my/aR2vvvegrjoue7CHiGaUKpeS2pS
pJDpk1kuK9qKjWqwwHAHoC2iRGOLGNJNA5pqjHpmTghwpn0ZU3sFgkHQwMPfKvTX
XGCjHztTOZE066m0D/asuzrWbtjGmGZ1xxC58lCwmM1Mt2otgKQL264fdBmJLM6e
6JK6oJ93t2uFnxlZOOgI9zqe7P0EU97vzMtqKVnaXQJAcCiuRVlm6Pfi9/5gcvh4
IBn0K1Ng/0lYXtC9N7GNkGW8cCj1aFQhL6iMsu1R4weAajtd8foLTI0Y2/brxrtX
gluJPehLHN2cGW2IO5N4qRbJn72HkFthSSKIpN6dz+W3fV2dtIdszoPXQNRDxgXw
US4y87+PDWDMrECrIeoyupnjqyY1TL8i+TRwaijbC877yQZnesa0SZkWFbKZqk8U
EsrJxxEN00oN5Fv2XeFPvrM6I7p07MJyWv3OlMXQe2LvTDVmjSwW5R0amu+Hc7m2
I8bCEK2Ih8MAmWYCQtyklrfckY8dfe1YgbnFHEidTPFi7HBvls8ALKMOGWvnezqR
jK2FJPSWqt8WNAIJ+LrYKDJUkDmp+kATIMW22QbS6/j9vxffrsUlBMLteHFloxk7
q/51h4sS5qU/PwK3ZM4xRD226sjwnqIDFqNBTJuNX0ZDW28YvJv2ox+UZ30DpTHd
y26fMRiFc0r6XGVcUaNllUofcu5enCZ+/JlyrpgcYTo9rt5IfoJGxmmSut2KQzJV
RZGFdG75sDNlF9w8+TW648DLraCldPg4ylkziY7SRPdNi13wMl+XOWq1M6mZm/8q
JtemPJ5mU+KRRGSlg4juh2W1HD0OWMNqNXr800+ULqxqDYY1Vu1o9YBHVKHd/rcZ
RVwSv/1EC+LrzRgdiHjJ9la0/wvukX1NjdMrlTF3vWWVsZQ3xMQdNQ0RouV+9PtX
XZFgNvoXXPUPOsup7yp4yFVugnGpwLZ361cCPageMEwNv4Eu3/9VydCcaaNSPSUd
eGuRBtG9cFcCK2NjuhVIR81eZzbscuEwxlM0extVOE0fhBKl+2gfzEtgIfkLAczX
XbIEwtGd4fOusePKbnxYUy5Zsjdi+Ox4ceugxdchFcML4/YlUCBeMcBOmc73PEQX
qLzGbOplDQ3jskNbNEPNPIJpfg1boVnVOlM59I2uGYVM6yQllk7Ev8X5je6DgN8N
r+0zdXhLWvKNuvPEa6NJ+FdNn1IqWcVn0FMDvdX64X1Z6ezj8qQMdruxdg8vitkz
GxiP/FktTxg0ctXgQPmlQnN8HOSeLevZb+hcSBwgH9H6uS9lVMfwr0UOhBqjfCcJ
h+aDs7vdcHrVlZCWED0BLCNwpK+xlEHgcVGqqrcmaz9wWgo4uzMiXNx1orGQ3fV5
49FS4/NbO1vNTLtvujGEcz01AtewbDLBU8osgjd+APmbQGRXUYMTYNNU7/VwDPUT
VtWftYLGpxb9LA8M830k7s+MId79uUxnzDbodv3eCzV5OIDuTNrL3+qkV7g7jIff
p+uXHFkYl7znciXEcRs1Vd1bRdlasGD2IxV41SxjiUAFI0rIq+6xj8OBID4q/wSF
tkUxYq0ze8qJkkJp9/DtKrFhvcEFHbLkgeocaHA+NHlVSqkNhe6KdyKVkG7jTHFU
PT0bwwb9ZUSVjm2Xf/WFCK157jM4i1yvx7KS/eSxuDyZ1VfuchPmn9TNP9/jrn9K
qUNoRLq3Asls6WmxTzdrBe3XGcnae+leXoKFDPpQfcSwHlgZOrKqG+v4zLOOvRTi
XnW4OzN/GqsRtRnsezOXqtnrQIBhET8SwYEJgqHmj6v/Fecjn4AeVw6RxqEj9n5w
VgCnhOLgv1aJExb3rRERioTXf0TC9JvLB6cm2ux/6y4yKW10UjiqsXkU0sYHs13H
+cIWxElwIWAM3R4hZN3RUJynziSMxq2NJLcV5vQ08jQH3w9kmv7lcjY5OVDywyGf
o93p5/KcgsUSVdfMI2RUzgh617zmR3kQiKjWlokPZz7ka5EjyLfD7pbMacDK3DhY
pQzV20aGMu5aG0BmH9KKvU2w5BeF2jYH1IuM4iOihasUi7i8gHy+CrDPcw5M5IVz
MNnL6OsNzOsk7K+NEgfTH8H+XkyosvUQ2qIpxTQg2RHlAXY47jO+a7/Jy+3lziIn
04B0+dwD12XfMPXB7OmjBWgM3Fx1eGhAeFXGkDSyHFAZZIv0h5pkpql9NN3LlgKE
D9gfsPGywf/EK65J+Ghr24/2T5UzyA+PKTyARTusKBmgnXkAwII9xMhL4mF1gnRo
FMzsN4kxgFWRZEDXNjepHoNok5I6lUa5c6eslzMkeq1cDTROFI4SR0fX/6juLL/M
NIgxJQ+x5/UCkIGLy9b2phaL7S1pVp8Czo9Dci7XTBdVxsEwLS5Mv4rNlTQVcOI+
s02JwvKbxtOrc5KxIIHABaNc8uGj/YhHsxX2UiKtqrJYSOKJr826KMH7lMYBNyUW
sPbxIYrTziEigQqsSeqy3r02eu4pYf5HBr25wRiNsWe3+uJg5Wstn0/lCcOYAkje
SImDDX1lNzgXNUhSDuxNv5Jo3ffZlskkqcAIb+UHmszpsZ+cMPKlw/wl+hZVpTjV
pmzlHGBHFjFlI3REldneKXwlUpTJLa3DUPyver5RX0XK3vzDAUOU3wkLLZufombt
8NCb6r9TD7GpcDNifRLccc+K3b7bZfLrDsgMKvCdta+Bw7HP49N+DC3RUcfXiJxt
+dWgoB7ErP+5hVp4adtw5tZnSZh2NDS4E1XHNd7tEAYIwXF7L9RXHabHHNoSeast
5mdtOuErxriCFUe5C2VP3xONpZkihJxYSIOhYya7xCZOEnWRaoS4dPNBDvd4GpX2
lieXeSYWUzZJg54cfAOwS9gOeAJoJe2+d0zHGwFxFIfa9sMuxPc35avikHgkMzxb
qlKTOV8YpOu/soy+fMdNEqJWdAzSIxKLb95aTTlPIOetA3vhunsk5uwjjZEp0I+s
bZCJcz4Fvx3EUW9VheQ8vTzvxkQYHCKCO8DmzNrnbFmSueziOYTAn6MLN3uneISG
twYwEE5gQS9mpSFqrGT9k6DSaA2+7b7dk7gBFWqj+n1KFoN3Vew71okPOEaSACiW
o8A2p6wgdDPIJk69/Z69uMZjRF3wP90pDBnIFPFkUyH9oRV7H9RwQk+zVKbUWFhW
4rTvmd8agsLhKXph4tlra14xNAav9F7YHAQzKe8Knn+lpHStfTBQ3YjRRi9uukdt
cNNcjH5MbC5X0kSAiuTx3/kErHzsiHF6dVAAkes/ByBWZx4VhMv6zCUfE6j532RQ
I+IEIx6ngPDLaF6psqnYAs3hUND7KgZei7aGOjisl5NA0HG27nW5h2WFg7RBQMGu
0FLGisP1ha+A7XvU5Rq0V/GGZD/dRalK3V7W9Cqck/men4RYUK6JQbleWEchpZTh
lboRd1gF2dUaHrYDKCE4afjTz6gSCjJypywho9q9mqAS74WBjf1Pz76NgQT9XecX
RMqoatFeBXii//pRr4bKyErZPmhjXThNFVnaXDBHnMjRE3PdB+yXnFCr8JQMWntn
sNB4pHn0Z7m+M7c2m06xjbBRHx1EVqVJeZkIM3iPOxcCpZXoIyw5NERgadyBBmXL
027isIylOJJweJ8LJlKNoBtz5bqygG0Uh+xsGLUIVE4IgzUWxvGI6rVfM30X+Qe6
SuW6qMgcsVxeUEpqT0aFrORcYW6cAzmrrYx8UgVgDQlNxy4yHyJxnjYVBZaYMbIn
RE4Y54olvtUhRNTbKB1jCSE6m/3ITF+JMzYcV283Os0Gj58kl6bSm7K0YSaMK2t5
T1xVOLSoePO7Aj9vseaB9YFPxMxBcoklUsaSm8f8sN2Qpwg+ylb1eji3lkvMCw8g
axm6EpKfclAKBGltFOido+PvWcRD0rnXvu/EMs940phNB5qTlW4o6FaEpkOpr92s
1SZ1EwXbZQomWle7yKk5H4MaGMCFpCRL+PaaU1NF394k/b3joOTRyyhJcmYsBhi4
akzMwqLVRUToTTaq/BEjBtlgCXJw59ZsoNrEZz+4RKfzwdpFh7pgdmKGYEqdoILa
G4gSv47floz8N1SV8oqGchtThH6XizMpVAA2ThMjqk/b3v/am1yN/kCOj66M5E1h
hACxMrhjfyF+mC+m5hCsJ408BF6OsLUBKKI/jzpZSaXw7A4kfYUchAWyHpUiYu+y
jqhPvQK7doAxKGNB+VwxZEQQ8muDlQIBSbsCZJ7P4LRXIWqreWjGa3/kQWlOdP3Y
jB1ZSc9cl+/5CekuFftK3WuBxd+VvtYsF7ZmV0aqpCwH7TM5ssuv0M+Vwb0YWHP4
gARcq+6vj63adyUGszYMl0KIKySel+EwhWxcTnzNOQtOvK3ii4a4C/REtuxN+fgV
Ryr1fgrWge+aD/xBHP7c7l/ArtIPkkty7fflPobimFgHA6Jt4ozT/MzabhtyLezC
ZvEuy3zpZ1ZxSkb/vupwKXckiJCu3ATewbDk2WLvEYr9PTyajZZ81v/hZjkb3E5k
FwOzLOpA906rFX5QYwpzwNaceS3L8KqkT+MvSQHmI0Qr9Ss4keGORAwLRW//rq8m
zCqj62IHtGfRc24kolMqDGKHEcA1n+g2iD3PkF8ErVYMdvpdxdxN4h3q/lF7M4Ev
55YnxejXg/MX8IW5Q3NlNnW0rdvqzyYMNKwFWd8rFpA6976GKgTbaeV6EibbLx+K
RSlyOskg7hsdW9owmecVkrzwtzQ3NKH6jrciuTixyC/wXVfcuwuKUjpCsSEXTH2b
bJRYEGZ8jnkN2RN4fK9l7pxUgw78u42j4TtFLmt8GsDDQlyQt4yQeIREf7rTAurh
0c78cHKqCL5uItVsrM0QCbmqYJni6pLKlFHZ9vIeFR/OaAJH+g6gz3uASgwHn8Qt
VCDRuv3pd3M0ngFs3iN7A2hobwOJfBAOUMbv8tvjXTOSTyoaAvoglF3rWrjZRPSC
dLX7q/4gTF/byhXYQx+xBgeYsmIaMYl5RW/eMTs1UKX95hUqQ/kigqElwPmZiZ/6
qVL04kF0sjspgk5nC26ZEeYr1gbpSaHQ119mkhQS2FZ9/ddgF6WAA74Q10VX9slL
gdGYVzqoxhwFF00qCuCPErBwSo+p5IO3g9ojHGBqD+8fyHxu/lbKHoLZdP1lmV9d
xTlDPQvh+EldQ9Ys3BJti7OhWQoaUujwmHvhghawiyn3TZ7dOxYNGW18N3CvsGXt
B8mfHMc8QRgIK4/us2fHgFTJ/AzACqUJPlaodoLANt4DeN+31oBauEqO0O4nih0Q
erVsvgGUx55LtipIEhNEABxJTeOzmkgV3QR/xZbMvaaeAKYq4co639IdNbs1Y8FZ
cAtDPxBaTboIpgObVi6/KEyKFrZtnddtSwzZKS3XW7CgtX1m+rRekYj7c4hc0NCo
k/DNjJSL2a26ZFlqEhHzQko4nLxRMxpcRahtjicHJ6MYWrJzyrgqL5eFhS2FnsDu
+uU7NiuPKTavTh8jt/KxWal9UWuzD7/qgiBhxQyJBCEYKoClsGAzvvSi7IjgBQnM
8M3LuX4S+rKmqtIuKAna3L2XZv39IANMRoyADpj9ZNSHHOCHQ2frXdUb+zZEzCVc
f+SibKSO+CLJMYqeRNCqir1Nvt0AXcyfshCM1mXkiywLMXc8M4l5NtYcROAFzKZj
RbJox+KuBlNGSlR8ghzuFpKkzycmOTVuTFEa9ryhM/KSJXHSx61u6+gYRc70BGbq
IHHRLZFYX2PuyH9d9a7a9tRFOX89EVkOiiT1dTage6d+kvOHaGizLguKDqXVeUui
uVGrjumZK9fXFiJsICwASlU05J0xE8qiva0JfPUjHfSvn6NygdIdBrf3nA8ocbFf
XXjigoDO+AYBxLzfTEjA2kVg985fA69+x+JJumU8enXpmc9h8++YK3xGS3z0eK/8
NfT8VpILlMw+MNOutS9YVAUlS+wp1cYJmLSY12eVFGIWJEoPwAYD5O4gqMYu/wtp
U+lHPv8uos8DoeEUaVFkWE4HJhut22RBW9UPe9qyW0h0bqmdhxABZnvcH5MAa1g0
HJDnjody/+aYYjFT4qSnioqUGEIoO/VHibmrwzHHURVXzEWb0aqi6K4U8vGz0jha
ekUkbGK8q42LPNLKm/xKfRBwUq98Sjx3+dqHf6AmnO+RZlNci/8tT0S9LQx39Fhq
jtk/LNmqZqz+5yl9YhsmD4tROO5HPZpBWMk+hJZ7Mk0GiKyQwrjG+qHIg6eZXPGr
sdGd+PSk3f/52xaUf/HmyTiKvJdW3cOUroGN+miKaEBj6wDkGMfbhkl2IYiWrYZ8
7rpdZxmZkjW5qVtBIaaki2cyG4eSEJ11eqhhL9x0bFBexjyUKyk1hvA749HyNbZR
tfhEX/jAo/8nYd+zVJaRjdgzzEjvGjY4rrXF7QaWqKOY1ndG6sIEc1NpIhTvaeZ6
S7AVFWYKji3MbfvfEsukuhNEEPtjIaG5SuUPQnrn2Cbng0xJ54d4p4W/50vpr28t
1nC/pINZv7iP3VC7sqK7vZdmd5bAUG8hPfsofyzojDStli6s26GB3bi/QrgbJINV
EZ1sxy/UhvxZSbRcpztYj0WdBUICLLUdJ+i45C4rHQJy3OiPuxe6Rvddq+dvl1Zu
P019xTDakx734DNEnkfHilcU4zZzdVzff779gIMgQLa1Q4o65/k/Z6P862fn7PKR
LipIfnXKpizDOxIzU11ySfjHhyJlT6j/P5525Kk0oAAGiPHFrnFPhH1KOlc06LGN
zWAtMu3rAaD8UplOox6VU61HNuHPOb/ckMiw3Jm6Cm6Y4dekeIzWpVt1rwhq4B8p
DaWYhx2y68UH0v8Vx0I29G43Pr+rmTufX3fnR7tOS3MpxV7c3LPFSlfthxGZXDUO
ke+P1hfUPQS7fQFAH6ZIKFf53lwAkSSB6OZ5CGcj17h4WyyiVjK4eemMZQvHEgID
0jo33GlxoQ71qowOOII2JB5G+NBH4YTXkF99RIEMa8DhNAnimv5csNFSf0OX1fcZ
yt8JhzdrDqBfyICpV97YYMl8LkBHXZED5N9jUaa9hn4WZF2bbdM+nEuv1YYBwM3b
Rvqav9RzWc0B6avL3R+DFbX5opPvk8wfQhdXCGLy6NJE+aIKpemnNlF9RozWGcpL
ksGTKXQCMFf/gc0jKE8Tf/4ah+kkY+2czle2CQ5ilYJRs6tkfUn9pPldiHP+d/Rd
HfQrldhC2rAI5i/PJqZbVRtqQCMrSlQfpXUvIgn1kCSfMbiy3vbua5i8M8rtziDp
DsPhd2K/TZK6vMHd8d+NQr4EVG+tA8M/7bbVkbz45VCACG2yb5H8bBCXWsLNXXBK
UgjzvvTY8fm9dfounqID7g7XEkz+64ZRyxQIHoCl3eS3fOtl/C4DxaTekLSWxhkv
F5Dk6vDW4T4tmYFxNN1ZGmjqr973vXK+cNSyJRyMRSvbN3E40vZH2WTf70jID9Q0
hjBfjIquvrpVWi3kO3Mn1bHVF7/heJJPH2RXc5v1hgDQDtQr/0XeJL8Xvx4Y9qgQ
PU5KS84bKm64JPaL+Dh3TW5Ol8HDdnbfmfJG0cx7dSN7AU81F0tVNVCpr82ZcJ49
3gSsT7TYbPC873tujadAng13lHSRswMwp5zzaaBKUgTzVE/Jura82m5aABwXOkJd
4SkEF9U5j8dWI1Rc5Zb12rguv9Y05Jf8VfoprXYfi5DO0xZnC7l9E9vYl3zAhre9
XB4s7ZkyX9lTzt/1YrArL63ZZJ94NnG8h8QH7bKl1VYHl4jJCGmRQwJ3STdchX/k
RMmXAXE3S/L7d36CEP/PIXLzQXzsTgEv1KRpVbu9ZSDHktINF/8Ri5cq5Oobeq8r
RTSG8A+gPG5161PwrrzBMv+77faRMvb1zNTcaMYURJXdbNNkgHglV1+doEE32+Uo
MqlH9cld5k4wWx29X4KUp0unJTjnneWm10kSOpHbQAim+lVtOcWr767OftmOx0xk
IcCidqHmQSaSUm6ZcwnINzhJNXz2FgSdV62sw9NmxBPgJm2m5XR8brFb0LQrvBL1
k28/LgHi/YnepRiayweEW0ea1Jo4RslAhReSI80aJ2ez0meGz2955wNjZs4+4yej
zlGcvo/sZ/wGdYwgrGUxMe/vw+lHX65Kc0IaROLKOIRgxdYQp4YogFwtSYxBrwj7
agRKZDBiEG+qcr1UgmEazt8aNF6vQ1CRZ6F26BoMjO6PAbvDFWF8h2AcgA/VpXA9
ONZRCxqMHGQzfdcz0S3X4P51xZsO3xDKODTtNOeyHrIb8qVwXX0lkJyEuvVbh3Hu
0ogWSskf09UoAWnwq+JZh4nMtWig7ldcsGrVz8fdgkUCDipmDQGKsr4Tyy1FyO7F
VoBp29YrFO5HoFeAQlx1V9JvVtoyXlcS+HsD7aTmeFc6sJ5rkVBzc5M6tsW7Y6Fk
54jNXYBYlJYgobd3DOBK/43+Q3zoOSMa2EnnlplbEwWVXA/HHKE5n0Kx2xRe4Xlc
qOUI6FlOjguNe7s5qrMIhlnmNP3ApRJnMZS4nzGAgxgYwyL4LnC+OtpFxc9my5UZ
HTzcIr78DiNkXVEX7HgiKynZqZtWnvsqYLg4nhgYbyZTQuVtes1ejGsAFuQS2KsJ
IDlxv3l7sXVaVtk8x2nQWV0z/0RtUzIMzgYwERe3o0hO8qt63AHUFM/GF59qKPVH
8bfVsjo4vQDUJDVFqzLQXoc5q29nnuKpjhtjTDKLBxlVuhFIl+gsbNEgy4eK3HlW
oVZ8WUu7WDOHmuhkly4QrmkWJBdXp+zQT1+52y/mfXB7fDI8VZv5pl3veK/9guz2
t1Fo+k9oCLHIOweot5A/WnEMUtrK1E379wVhb6C0q24mxhPK3gMH6WdkoRbt8Fut
gscq5UDdaEJjONMMyn5E3Zc44bIe4FAIIbYnmn/lGukDlqsV2FF3D47r0RP1O2lF
r9sc4AlKkZpdPK9k3hI4GZyzsuiClde8s0mfDzR3y0k9fV+GdHuDsvBQ5YNqqUBU
JhJSij1UTUg1+vU6Bbcg4VSpXfpx6MaFqAJPHZc4KPNtbEeJnWQknoIEYxInwBf9
OxRzkWkra4vXdc/OqbwqP5IxcaCW6z6pSyb7OrWwJvWgjGVIUPhGcE0xyX/utz0F
LFw6vh7LCTMytMkMeAnl8tc5mHvPZI211A8f9mJRP4tNTggW8xKRUYMd1mtMgEDl
URJg9xWgoxG9EsxsAt3gpaTTzEFyFKzkDCp14S8Pk8fg/H8dJzXLDbr9tv/4x6Lb
gQQfuGW2FpZd2wyMqR47vn4sIRa0E71Rq2sBGWi8GFlLypgrkpxwY9vB7Xcil0xH
so2AOy8TLZTf4jsEQvWofnmjNxcWhcYz3mSfsT/lPVS0V9SsqvCCtp4LDiO1lCAy
ijMB/mErgsPqN6y+4AUkcDTghonA2iNFfVep0VOe7NW4bADVs6uYnyb5pu9lFERG
xY1EKVJvZR+mtqwRcrJtbP9Ximtz2yUlTmyTVXGu+mr6cTWVn1f2owDLxAuSLzwk
wMzP1PKb11JlSNx/gDkDv+9/VuSDZ33CN2fUM6T5HvGF0+5cWDhJP5qoPRNc8Tdh
3ntmqvgHUedKJXw9Nyrx46Rc05NMss1EQqz3ECwHrgb6QggENpYcRTNBA9o0EK7m
0WlS9p0Ti/eP5a7yOM2m0WTiWbcQxuUQy1FkMXWlax/HoPb5YUHLBcp6aQHGdyoC
zQqvro7fu5mNETpuWygXG2auNPKIhO7wBU5HZVx3ESOa+zICP7QxLLNaz1KcMxVW
5BxkY3k3V735tcTWmkaURrHJuxSwWvCcHovE335UlhCUPBPNfF5M2XAmgmmwCQMd
oEM9s2nHd60FWYkazsUEj+9YowoRZQSZZmH+JcqT8IfVeGx0QBFAL6LKlaOK2QF6
+ehzMDJ/Zsv1pQYHwx10/btAMQjD3PeUsxEiFiaLc653U8vm0vhyfRIwYzTD6QKn
mFPvdXaopBwzmUPNf04CKjQm1Gtp1DnjQ7VLTPUpPH19PbZJbzu1GruuKXCRvfyM
HZ331rdYYxjSKxkEbXlbbOSQqKHgQSXiwbes1AEh+r8kcZhQ8SMoaiaCTnx1W5Ib
Zp5huqT5MyTJVQr1jwVaOqeSBbt25LhdSC28xEbCF0N7ZYNJv73NVrNmpBgikCo+
Mcr2lpujN98BAGBdILuZRfD/WB9GI+Cgh0tBcnDNubJfq8HCej8Wjc4Y+zlujz5y
jJPhIkCRoWG9eoZOql/ZUWrLpIPiE1J7rwwT1wrb81AnTBzpDz1wljjS6rsSrGh0
rQpRGOth5eRgBYcmB7iGx0QLlwz7TMawVFLvzdm5Jyn2PD4Il4zY57FPG970w7EX
Xavxn0G28iDPOc3FscRvklVLXgirOq8bijFDbGwbp7PMpYcGylFf7dG6fR1mMNBw
SItwLUso17h9ri3T5pb5zDMwUCIhv4n2smeVScJG48AKZezBay1LXHE6isN+mg1q
5HzBQiSJ2teyi3q/S1IKrzc0QUqwCdMK27cmUuHkMJ1CR30D1Y4akWEUs8kMhSnP
6EFDM2xpe+E0LhgxMhjRe2aX01CbRAytn3gUTe2uGndvoAPNgbaV4utcdC9ozWrB
ucWhKFyFFawf6my8n6GKQqZYBTVIo5YWi1gSe7dtjJZqnPez26VLOGLS8S+XJWWt
rjvEIv1g8XmIuW4hKxVKiaGr3vLNE/yI+6j3sBAhFMaiIu06aU0CN4h4mZi+aYML
htc+d21Kjb2waCcSJZxXqITzCVJGvPRF58WXu1XbeirWZ1Sw2sHkFtU/E5QjcoGG
5iAr4wD1q9x/0liqSHalnHchYwGOuOq2UfjP9CRqV0bC0e8+bVb0dQ7QAGltTZYu
vV6FVXu3r2jeXYLUAeGI5yN73roHsblgWHYz5GtG/jxngVf1Acknu6yfUSYvYmUk
Ks0SZEnBgYvSk+AU+y1D/EgePKsEfIkPvvVpo98x7tGy5vtuTxghsNhmiZifqQRn
EvqpkwizjGmxq0SN5aKvhad5HGMM2qXkhOWA91b4u0worlqls/MN771LMxy4hPAF
EXDZZLsq1k2va1eUkc9/HDcX2RqZNZUZLRf5kV7w+OI+L766JPrw+iXWddzZhmbr
tCbz6qp0zOFXqOJ8anYysiPq3skRZjhg/G4UjHdP7AK+0KMc5PaCVxA8USbHZl6j
VXd88tBk6v8sp8RL9Qyes8CaJQ1f4NhE4s/xAURVyX1K5rgrKqPymMarCv1l7ZtP
+tNxhh8xuaeI1wXCNoKGMPYX5A/lvUgEb+WGEVMGsOxQpXW827XWVzzZXAxlu+j9
Zq/6OLQ0aBflQB169sMW09fwaXkqk6OvXjfa4rwIIYVp7IwIflUd56fNd+JHtAhh
8+G1HyKDg50qLE0byYQghWGq5Bcg3/mVf8vPn1pROkRPG+16UXvMtK64bcT5nIaO
sb0FBIbZEAmnUSKq18BgOSp5YbY5fb90DKOBmXPr/dF9w6hIg8rDkXBAhoNmvTL7
eXJVYWoEow4MA8xZc1eSRjSdK5NCPK+43/7KH6BZFMiWeCcddkDU+Xz3F0GmSToT
4uQeEIIPhrmi08zKh1YCAmq5Tae6Hx1EN7H64iQYzrL5sj9IfNcJQhAsX6u4YpgR
hvVmBE35+fDAVE1Cpr228/IndyMV8pkh3B16MPUXrE3SCfNiY6MJ+RQ6FI7mXtl8
choLN7XDpSnpZJCa47FvhnirhXhhqd9o0A3ZSLt8hV6gXxkRnhk9knwhVTrnlX9f
GdKld528+ohcu9z6M2Mz6dSPzfb72aeA5qUCWr2p9uhoL7zjowJftOPogkWWNMYA
AetIjTNSBA9LHPbUXSzP+pJO1DRxBQxOMcncJChBvulw6noSLgrb4D3ujdertA0c
JTGTZPbmS24YVoe2oMTdu8BzylPOL07aaMURIjIMkS6C9Q97kMT8/eM+qVSulZEV
SLB1doJzcmIVcZYosl2LJYyeusFw4BILlIjdSUia/NuhyUsPkFsfKNfL/RodUXNL
yS/PUmdZ/WC49GedQiOthcLLsfWjM+/gEXdvKIkTlfy0CLYWCGJKPzq6kvKZu15U
il4XDli6remXNvnOA953SM/X6wBPhUtiL32rhRbobtFslDDDbUdxSjfEr7Iw3RbR
9LYqcoR1Zoahk7FHrh8PaYmTGvd8tY73Ghk4au1uOI5aehOr91xAgcdLTUVFq6x1
6PMnmaDk4xuEIhqfEZNao2Tg/rpbJATz2rEdokL878qBa9AdA3ay/fGpjZwZSKLt
rZQw1fU+X+MuaMca4inGkhqDXeb+b0R93/s+Ci+8MOA14RhDKX+0Y6GEh+gsQdYP
mgJcwv5FTZ8NWdt+PQLe5E9jcRRRAD5rkvIB42LOHvW2Rh4QYLFpIc81qip77cUr
bePyOhMWOXvv0EJbi0w1Veq9ouMWGZVWhqJAJ5xdB4js5eHtWsF172B9/rE9S6yZ
LNIXzdApiSBtfKxy0xT1T+ynJGg3H3EF+0BxRBvnRVAD371GlH0zuzno48J+sbqe
EnoLHHKUkZoIlQG9k0OrUEm1CV7Nc+sMhRQlboYbPcXYpI/JtSwM6RD9cNv4AM/7
E5zv4jOBu2zgCCLwJgqK4ulvr9uiQ86eUKw8aLrFTwqKz/GiJ0xE19c8EkMsR0FZ
DpJuKYkBAdvlPrBbsojz/yJhY4FsfKOBWUqaFjk9wG+BAP5oEzI1lbf9sX5LtCPk
D3HdeTJpw5OH9LoKOQI1Avbw7SRrDqQSfbU4G2Sk0OADbhSPWAQ36WSgVCOoxWXE
Fy2EFyzfiW5nMnVn0it5ienm79kIlEj4xvSVydIVPgwvQrYIt1Ru0KGRiXAHQwzN
cRpPTb5wUDgTADnNaVifiz/7Opma2345b9OvDFVD1+4eW/OCm/d3NXXfCvmrq1Qk
yT8ICZ8DM4GI+rV9EPk+WVvXrH6pSjcSmRB1HylZfuQrruekogzSj8yGILjG7kQG
i31sFKLTW/4MHNpYYhRZgGcZB7aLcKZydVKtKCTQbHKX6uvli1rwok1QdNhIwTTR
3dzHAa0XVyVHOJoub1x2NCCjV2XqSOtt1o+dqi0k2sDLSSs+9Dd9XZ7V+uHcKihh
g2FvGtk5DUKmELRuJVI+1X5UE4gnfy3ztTt3TuuCEypTvLmu8ek5XQV2eV0oWauA
MUFQxGOpvi4xB0yshq6r4gZHiVVnyL4xmVjt/O02JYSmNnqd4R5bFunO3sX2r7B2
6KwFgaSDWydbziKapMp7xXHOENY1ZDYu/Xbc20xAjwqkpp/PRY2QPeYtRwlnwv0R
BmdmkNPSG+hE9Ivr88evNoqJD7vYySqoJOd7pGKe2AfFbVEqXFK3RTxHHEIEa8Ph
XjsFbmNE+oiNwnJleEw4X7cC2l7O0GGO7B5Fcy24MtuTPmFKtTUDz0hbhgoxIy/+
ffCc46oatD98cpFdMZBbFvhzMwGiQD0BQPt/+hol+Hx2USTC9F1A0YR6DbVI/orl
LXk3R6QT49IbZRqRF9UIUR7y9xT3RRRGBUyplc2QVUV7XjD7iluwLgHqa0c1cl8e
4NYrjNaa47hUXYtvQSFgHE0hVlBhh2lnOqqyoii1eD3wdDL9X0mbIGA0ob2OcWC4
VSobYoV+XUumGDzRqtpkb7FXQqFmt97AcodoV53ars/jOJAlZLaHqp0kJaIEkyaG
pTE1wMB3og3i7+4rAVwB/yVVSYKzPzWMW2xPQHghW5lqn9X93rZLhzUk9xSQpC3K
6K8ckA4VNLMsjhwskVX0jpz9EjEuQlIiLIMa1QHbiJSOy8SMjC1P2I01aUJFU9wo
ZfGjtWwieRNNRNwfZuTui/J0aSfR6hLG32qbQgGrMuSGxflNOZ3+zMKk+JZkvrOe
QuRVGIoPCqELVWixm2FfBrn8vi+HB2x+V13qgAsRPzc5E+R3BqoCniy6TFb+8EAP
bIddifl3LYUCp90vtLh9L5q4FBer+T+LU0LQORABznRZ7cgGhlvCHvHqF7dgzB5A
EQerxJHlMR/KlN5cLaWGDOgiycJDAFrevO4aJSC3TBOkLnfT/RLRfEKPMyRPWjcL
dzAKogiAkKojbBw9Tv2fsKNdF+1/Vls4ov0XompKLQFresdl3atGQ6CLlZJ3aGJ0
`protect END_PROTECTED