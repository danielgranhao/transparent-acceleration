-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
EBNIqK45sd8Pg81sDsfaxklDLlk2qY1dC6BX4Va3cJSEwNLlax2MIa5c1mwGO2P/
aNBssfKFwEa8qvMUvIEQz0lmEx+ORiWxys4mmRmgVDy6vS00rvQ9OV/zyo2HK8fD
7Os1JV+tRDzHXBW3nFeNUXgncrAHDZdR7uLSQTXlfF8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 36320)
`protect data_block
hVWYyD6eqP7Cv136QRf3hdhFZTcVXsY+a1+uql5aaohQEQSv+h8f2xNgeidtjHxO
PN1wgkDLLMuh2TQ9dOnq5TU3eDiMuxGxWKbsjo6EDmGZFftHd+9G00oZpWNbiNh7
gxZgzssjx2kTiZFve3cdGIzSDYSXDpgLLpbxN7i+5uwLyA2uPDSetsXeUWBBUU5U
hbQ/DVtiCApo+twfk1fvMt2/ePlNplv+wT2vUwdBMl9X1l082z/4d36QcNiiTJYQ
ZVoCIoP4aIq/sBfQpKm3s4oVO5qL6ZQGqKuvptSkBo7SY09zKnKtFMALVtNOfxsZ
RqGjLKDrWZEu9soCeiJAmEWEPDFE3PQYkEFP5HJ0+fLOfBZPDO0j16zGSTzSv9WN
myuKy8S0r9qoSG3Xe0OT0DhljXir5eR0hSefYCBRWjOt/fX5XMiRI+8vpf5J7WLJ
iKo4mTwL93LdSGf/r4bECgyH3cZ8Gv7RzXV+ZPsmb899Ubr86DY62gudARP6Bivn
AMghMEZTzsDVLtWK7HRADmtBrvC+QXcRqhDvrQZjMPgucqUo/z0ojt3TESQhraCX
kM6z4dvuEyekVaSuafS68FbKYRHbSOyRiwA1NUTtDJetbPrjlTibVOgViwre26lR
QeP6kMDdYkjWzO4B6JKDjZaRjbjlpgo3ql3QOaKMsPmHIul8H5P+l9Kj9Ep5N8Hc
xjlbd/2akFjkVYcp/T8Oe6QWLfTqWFyFcgGEF8sji1yTo6iww10nuoHZ4zSmiCPM
a3MMjQ6VWdSvNBE3q/soYzF+ivBa93ffaovVrhJ2xf//hynXt9IoNiEnk08KheDe
5RstS1CidiODr8w6K0UMNyVfkWwL5gavC7ruPb6JlOdgIuMNkOSV9jL9OkvV6As1
8MBiS4qOApa/Rr4DcaEeixm1CZ0Q8B9lSLtIUMjFHqP6RfzyfaTA48nG8yIj6Qql
Xeo3UXxEfLb75rSPBZOzZ/BL4eta9ZYAkdNmSLVDDjQYK5VMVf5fwOxxFQ8WtMMs
inj3b8ChKO/UsjccIn0svV6MGUfewr9h/W0VI3Rxnz6UT/x5xi5XNth7a7V7I+hA
U6iDes7PnJIPyaOl7g/YuA6oK8S/pTBqUXlCkG/MoZ59VlaZ2r7NgNGc8gpastpH
EuY2F9w11w44K/zax4HfeA2+Ls55X21pzQW5RGuXYukz1nHggBBJS2QCjMXJM89Z
KYomOnokQ7jGyNYU6KK3mxri+EP3A9JFEJxj4qjQ/syS0K99YkHnQJZHuOOgZnmw
UHRTQU2xjNDRalcn+ZPOf4oI8rUMYOkj7D/Ve1HFUhqCGjuCGPuLY/fKYeHDVUpT
aandTYAZoEJFSPiTRwJsg1RfB6i0BEZTSO6Sm4yFc2mRze8ILnah0EeypsBtgV/g
v9OdMRKpE0pdEjYLA9DWHRZn5zqHfMT/h+9UQsbgsIQhho2IwardYRPKjb6cKlE2
RSh0wTpyStD4X+ayFlIV6p74I7clCXFV0Jd6keX/0L9EFdppjXnMNZPqrTCMX18i
GPoB8/IYPlw/NIOIUev+iamC+Qxt5RSjAnxd+7b9skuEPwk7OOtFe5LXtgrH48Ts
TzGbH9PxxLqkq/eZxRLq9RxzotYaIk8DQqNHHqEYZ3x1OvCA3APeBfLeaNXuz3Mf
yZh3QG79C/QUC9Prk2lOL7uMJSN2ziNV+hXkSkMcfWpw6E5NqVVQiu/l7K9KgxaV
uPKiGZbx9e0S8Yxw7qq7QlFWaBY7C3yBnN7NXQAAO0T8uVCUdGf3GC/gHvi6ZiyG
tOR19GEsgkycd/VvVfqXTOSU1Ppv+5KmrDvZmGG86tuoVAXTkci4joQBVlhzREX9
GaOC44MyRBRuBQccj2D9tMalKmlVA48FwY50HjYYPZ4zhXlERDZ+BzxNaxcZJbCa
dEGBUsQjzCYDyHyMRMRQmhPztIo7SmKh7b+Z1MT2QpC1XR0euyk4FlzJDdwCsrsF
YpKUBois2Vs61kil9eFEtJwGGCj7FzMh8nSCz5+r5xwyctBWNWcJ+q7Q3snxQrN8
M+GuOJ52/s1SalE6Pea7b3FYyQHC8v+T64JJ7je8QUD0yGEslj+AEWfn6Nw1LKKA
Q7oNm4UvEEwnw8A3+Gd1Aw39zHlRnJxVP4BlBmvb1N53024Pj5yrSc4nMlA8A4/G
b+d4Ihx3nNuC/i9ERnxlu3IeUE1wAlD0sgop7Jjt+5uck2lGmVqmrwBVIvfBsGRi
2xOmaupWZiuOtPTVXORDF/xno4lfmXoVnNblhhCyQ6ETmZNUYZGUgZYDKT++8+pc
RUeXbCaPQQTRo1YShtRLjQ9KeTirkaIGQM0ap63vRMzQ0/V99Q2EhgNwC6d3g9X2
Jjq+67ghX+aPZxJBGAZCaI6u20JkWSbkAbRY1B33V7oSNA1V4kSqFNou+5+7AILD
tjT1P0yXs7cif1VPbFnS5YRXj7lFTfdswoKef5dp8TkUQDl2xMJOntnr4WKGtqTq
iD/G/U8Aj/ZGzWvDUmWcAr8/lZJzTxoCbWCWl5IgbCRUE+ZROnDo3XZt0xhWs3M4
nxI+dAlAOQPpSqfH0SkchBHjVkompimZmPMz0GFiXued3YajVb4DvoKYIiUxrKQy
mulEpC64UxrmVYOR0g7OnEuQc2gedRPQfNK4StwVeJ2iKMQ06RVw/MH76VmsXsws
tm45UmGUUJsk+OC4vYx/n9Qo5W4tUpQfr2EjTUhS57FVlVhokKVItx4cw2ANPnaC
eS43X1Y9ZRE0PotLs0t/2EkJUsHjYTzyKsW1dGYdTypwAOWKHSrwEPipy20xfA5I
pz1cNsW7GM5l9Cz0xGWbcRnH4pY2rdKs1au19rWyrKD7vD5DY9D/jDw6Lp66yD50
ovJziFfGJa4zkFUcXH1RlZtoMtogkGmq4RL8VM+42SRtGr3tt6mN/3qB3Wo/XEbD
RF6/aSBFaQPDl0k31XcPmoj2vgJA4HPOGHcr6oMD31vYUZLTzFvLCGDIlQ9NltAn
AjS1rXQ5haRS2yty4FuUv+N53cOqvI/7XbBpvIe2NUsfu9+6bjgN5f96csBiIlJ7
XTb79cXn4pCiHXaBEUIgml1w2re6sBOD8y/Or67yhCmlccG86/NPUQkhys0Ri+wz
+OQy6Q37v6SKNFYGDzV917ysSKWcWt5Ry8AQCvINVsOrJ7OKbQSMStC+WcJdZqSk
r+4jIXLpBpCA0qESS8BXaF3nf2ouG74I86ZwLF5N2cDVUPip1f1DRnI6AqE/PJ3f
0yBQ8SD0LW7Fwly/zAgEAwSLPR8yN6twoRqtPwaZxt4mnDjkDSq0cUZKc2U+eld1
FKAx9M0sImDi6kHDif9dVePxADdt59sUGNTQqMSLmRMpfzwssumSe6IKWhTgG3rI
CvJQACeXS4l1nydHzZSAdTSiNKZqg027n/1yrxNBENnzpp9O38I1daWSVbP0KPyN
vW3WgW+08dqblmDCiqOLw/BDysMC9xgKXGM/y53kY//kN4mAmAxg7jvtmGFv9Dui
2BM9fiecomwuLY9vj+KIFDvJVgaiM1MvXsV8WY8sFi6c2mPtbUhbZzMAmTojSz24
zVBht30G4tElHurmrNw5I7He9zaCrazC2w4XzhMmGduZvdNAfRf+e9DMWIVN8sLd
VQnGA2tQT0pD/lqrdKe2ZIxnxNTDSL1vdkz5UG3lBWSRb5oJLyZsZpQIbrxLMaVI
H/LAuwfTgFUvto4tvS4PcsmqJUcXVjFdFieKieT8WiM5E3aBJNQbXkXOeVoDU9bz
kGz8k1LDYX/1TnNVHRIQXE8hmrREZn6aOYaUNvX1rHEUFq1vFUf/WR3AY8b9/vN4
n94JHSrpMqmRgj2uJLYxc1NLxJdBvAgYxKbfXygiB+uMBrCdwmWCcuAGHe/morp5
Tqd/WfX2hqZ/Jl2je7TBU22+r3hgnQxk0RPA/ZtGCaFlbtRn8Id9eEqmNJ8GNCCJ
Vfsn2vKNULKJnm2ZTRDacHSYDMidIH1dOXPYLWuJIndy6bE+TW1TNe2njOiuYXhj
7+fVQvNZfq3Sq0D57+B0ewMEnK5U92G+XtlKqZnxVvi9fPcYJdT9wwJqFXlr0kt6
G4g9HAKQ0vdZlstbBJQbCdWOPXG4eDqdmsiA/V4BZ/uFXoDgu85A8OCdthQ7A+Bp
M5+NQzJyQS14CUxGWp5r7gNpbLXfmajdene+E+PkSeDGH8Tc9GkpwvdubLgJFwgd
JR/HmFxN7wLjko1+MXGlqTkZ8PvYcVuq8Y1pMt/Og595vOIn7DPmRX0U1rpJ9QRw
7n/JJKVJNMYYYo693WLFYPl0RkHTLr12Syj4CmpE0WcJgo5hacq2sFndpIK/S8Y8
k3+DDkoEi3wTt3Kt+ZlSg7rl267yME3IUuV8A4dg3Nk1n3izb+KCAaC2e5TsU7eV
8GOAxwXmkNI2qBKucQq0Jw7EERynXZNjSwmzoUnug+Orix7Y65ky3JWRsPqG3UYx
RCfm/efo185qcnJ6vFpsT1w4eZD0VXo8oX5xoIX5XjLO5ggdR1mNCEGWvxqee2ub
YOEy2QMLulDmMTxjfOgsUuOjdx1WBcCc5g6Xcp2zMd22PIE5QdPPHvR2b6AwNssb
EOzZAI4/Ppbo3b2SEQZZuc0Ki+660FwZZzAzhIj47N1feaH6kmmf5TOz6Z8cvEoN
F3XX1baHnMpW8tMGFL0Fo51esYf/Q+tedmD1QfyF40omghnX+P4zAl2PmIj3uJ0J
wPICC+1wxBKuKcwyqPZPga/f0q45JPSVJCYQNOhcvL649JTWvrGVohWLTCzc9/EB
R31q7mMhyvFEDcjirDyYiy6pGOQ1Y6v7jAiI6Ywm0GhKqVHmOIfDiQasb6OrnRoH
W7DpKbhNjB67u4t0d0UAC+EckxoE6zBiLHaGEkwMiXPL+xpgQ/JM9+IyyjD4ZXxt
Ow+eOeKYjt80mIb80qov/gvdjz9VkWbNqRyWM0DqEXUPwLYcsmw0jD7p4xE0W9Ln
m+uqZVIUzt/lNUFafUkxZDO4VtmwrO1yrMglTzu3whxZm6R8bBNhCXxJqX3igOXQ
K5QU1w1UPtdubH7/50F8h31ry0cQoT1F6h0I9mzs5eRDvpZY49crTC/J49dypKmE
+zLoOIGQuxj/5fW7VlJ5mORLudzeHmm5rsA/IzSuwifzs9wI7HGs+AEX6AQs0KIT
ysMEaREeHjKst6S5z7Pi9o4px1nZ1F9fpFJushEyMptiUfqvKaqyRJ7dKjc6sBIF
eM+dzgki1+dK8efINRewQjoqkeMlHX5NAWML/VGhqjv6zfZiSfi2iuejKaJFdSxC
eXyKADQUFxSBXmJIyWnTwITf+h8p6mRY67zp5xe0Loro3NFADCWxJEvDGQhqFoMN
5nw35pvH0C5oO1IONWila7EaqSsV224xVsZ6ieX5ILv17HVHQyp0LDKOYjUJhLnP
6q44YNrkLqhwXx7T8qv2Vdr8Msmh8uVMKEP+qMPzruVdBZd/nuowSLNeRS+lSDiN
I8H+oAvCdejd0/Us3GX+qDan+ytDN8pBABR51ylHB3N9Z1o8RmJCKlmR6hbtHm+d
GWjRtvOKdaYRfUA9woBzB/VazrVhoHvBtw3wkK0vdsWfCEHsEIe7zu7xlsn7pnQ2
ae0CvOW/WQEuMNdRjtIcUwYF+Afrw3G/zQbgRwt9smj7TDAdz+uacVs4ZWmOLUvL
6lXqeb6oeqk8VDpTlT1RX9mTozE7bQt6WRhL3BXpYPzEGmtMKHq4l9ZVLfPg22lN
5P5aKhzthb/HVLZSObMUyJ6mlTyDSO+KR1oFl0kyxFzw9eHrujWy4FW+n+5D6DVx
gDO++hJlHsqqYQ5kbEEA9sg2429Wuu4e1QqgwT2f+6YAugvnyYXzJN1hABeMZIdd
TfeyvAgqNm+AB+w86jsSqcFEZDzHNlOk1YPW5FRmkiqAY0Z5I3Y//pMXFl3qX1YT
JMs4dUHXFhFpx5x9WrjWsYm9mgbKsEi44HfoBt/GH4FwgSz4tdTFmUetNGtuwvgx
1uOFXS5IqTQ21qxrOTdetDVCXXQvS6wloL0e4g1CdzyfInxlNFFrBAGC4H0BjlED
ihY9sxKrJTLaPGgqwkSQl0SCemqF3rjc4+O43YaMF18UgCiHUzVf8IPf71/WdCCL
AbXdFVJ1kf31fmyF6Dp/I9emVrVYEV5HipnZdAD8RuYVAPUh6418336MeADCBk1R
J3/1l7FVGXA/3SRlKcrIBN8Fi6GQn9Nr/Q+qc+il8YSevDoAGqjULOkRrBe2amy+
mMIvFR1DWC/07Yha0hagKsScJ7/VPsWDP01IpB0Q0iy6mb47vdW59De6WISnAldt
l2lCPwjKH6ouDu86E1R/FrJUBIHznwzefd1sEfw3WWWEl68Hm9OGLnW1843BSNF/
GNAA/2jQJH4qjcRwhOqOMIduXhM/xWzEPOPkc/qfTUrU2zN9wAgYkVNGUlugC6uW
esk5FgZpGi5m7S5iy8ahNEqbqV+AUPrJyhdsbDdq8MT093jKr7MZKi/lioNLzKhF
9a+u+Okt3FARN4dAvzNEr6aXCQp5dN53HAvcea1mryil9Jab6lGJl0bl0k1+kqCB
mfLXLhS9QUXnw/85IRLjDLdteUMVPLJ6GQuOxV1lyZz2lZOjIbjyazFN1u6yI+WV
1uAF76rBIS2NeIVGE1Vk/S3wPGr9HLYWnepjswkxk97C1OjWmdQfWslxhsE6Sjd3
Qm2XmJHLk3RtJD4NWza6Rli5N0DUuVpZ6r5ycsnc6hanMpTb3m8HmnBalDUH4VOl
o87zisb8BcPtjM76Erw+JABNtFHDRPbMVawrpt20QfkUOJlT3QNDVM4WGIuhdqb0
UZdFmPxH32qHX7XHZDbWyNA+IOyZKHFpzkbtWxZLSArGz1PKaHuC0TqE8HBKQwD0
gJU91EqQIFHgYXs47AW7V+TiHM1wsQrjAe3N9pRTWMooGpufSkzsPK23ZKWjgERe
39UM4fTpghwvmmC7UKStARLbPb/9muyPbSNRVYLS5HNYZGvtmxwCYzpSuIW7CCLH
Njs5qAuzpAaq7NmSBA0MYgXPZL8Vba2WAhZvGyTXG++gpj0ENtcHIoIrUKGaKu/y
fUCoCH9ZIhVK2Q4m3Zq7ZZxU2zj8yuSn4KgVenp0RUWA4b4L+qESsAY/SsIF5Nqi
2bt7ZMyRMbHDExvKbItO25EAGd4AUpo8VrDZqD5KKc+zPfrqATJj5XJNeMw9C5M3
Ax3796FW940cbuxjYa+f90dJ/OgegODxZN6MGT28FnLtt1dRvFZMsNbYkz3rQkE3
eZdzzDbjr8Agrb3G1rhzr0oEwdt/dlg5e9P1x6+rfeLqyoBrX61TMRXVQq4KBE3x
ZxAtvj4euNiuwDTEaCjsxfP5BlwmV3wYfcXoJIn7I6O+HBzImAH1ii1LBx3l3tws
rtWSS5bt068su0o6vGLhSaC9yUOBBPPlMMgWN1D9x4wDLR1PylXStu15sb7dtgO1
si8No4O8ypt5v+skFTBDCisPdjM/vgOBfnZUPml8kpt3ex6KhYsS/ni+CoWKiEuL
O9iHP8mXhNJUrsYulqaXKhcV2uLc3DPcP/8W3vBTAT74ZE5aPGSJX5vHQXNbJDfl
Yk9lShq74XANJiAp7NP6KRwan9C5HfQfeMPzdJNK9VWJeGe5UGRZMoPe/NCdxfY5
pbWf0FQtdimfMUixKLLrMAtTyDv+6RAlZrWEEZXu7AolSP0VWow044LAmGGd96xQ
ph8qfdkw6eI949maS4mXeN8znBSBe15R57GUKQC7SsPUaA4DJnjiIBgx6kg66EDZ
LbOtxleCg81OW1ZUaw72X19h/iSyfzv+ktOT01ejkxGgzvjJV93GJg9IGzvsKmvz
/vTQ8l4zvwj2b0hUTbePt5GfO8GEU/OT3XBhjeK4WNCagzyRe69DGPvWMWqGjeua
mJtSbFA4/KiSLsDxo1thyawCgIO14tJPwcA3iJQz00h0UQEOo5vhcl3qs5Ty8gQv
pwm/NkzYHTSgT6pg5YGogO3u0zUD+ZK4wUs8w5WjZSHnzv3/KH8jpEbPCR1NusQy
iF1ag0Y+BYPskik2xKEMvgfVytCLT8Ly72vzjsc5zwo9EfvD6mw1tOQFAWNH+W+Z
9+I8A1FM/icN6khGi1y7NH/zBxg4lm95luRyuegSS6Y4dr/uLA06avK72D7818vv
06UL1MyxfXVMGGZWOymW4QpEnwtBOseSTT6ZjdGoWGjWc3vSQgjg7zXxOaeT1cKl
ukRk670lsjqDAKrV+RMjQjTce5LNgehsmjDiJBEvYHmCMxrKyhYBQq84BTo2/WOq
8ztYszBE/+XmgeLeq/WBrtm9qTUlojunVH2a2aHF5gUgVE0FTX+el/IH0OyB0qMC
KGQLac3jcCB0t2Gq3jhNrjUQcGoUGbtTJ6zwpPZVi3PjH1wNYCHIR+rJT+Wgf87v
QEcb+ALHpsRAoochIlC8PhEGD8Glo7Q2f/7NyXnqWMs1l4NWwOLRfXlPGa/wsIwr
0io5RBYpVJnnq8A/gFDYue+5MGnSUDnYYjUtvfBKW9WpfoZWdVewBcJ7KJa7UFt7
iExw7rDb3Obv9nXYpISqFLH2veZP6uhGs8aXyphMrD9sN2Aw9/N9JtMqeCo2iA7Z
5s8vTo9+sbiR7cy0JcHU+jrkqWsxjV4xQWvumKCvOJrTqNC/Vqt61z9+yfZe/1Yw
VpBq7KIKl2dNHcsImdpx/DqUiDZ1XJj3cAMctin6fzYw+Qq4G15COELgqHfZ4+5K
ZSVHS3qmeE0IPazk7c/xNNEC87ARUjEREaclJu2Ubp9Tv50mHFNe3oOUlpP/dFsf
BRMYaNRV+GCjYxBczvRWTETCVW8zzAPr5PotOh1HvubOe57v1Juv95IXZr615Xdl
YUsQMOmgoCyX6T/otT2j6aA3PpcctXDCvD+Hh1xwRNJkBv+MRhCEfaWfI3gaUOrC
oE+G5h7dgd+4HAhB7WWGaXtLVw2MrLjHKBuqEkIevK/tPSp2HJTK5IYGtGFdJpZn
CBiBPACTL/ZTJH374FucSqAW8cIzFhslalqfurSwbji1qGqAxpOE3L7R5CauqaOl
9fyf/Y8vmdPgdPZjdS/zz7rscCgsmih2T1/GCKRFU3jqDWW88kB1Al/to0SEHJ+n
BUX/C3Un39ar+4VucUmQzmF+vDAxkEfdj4lU4ec5N730GsNZxcTkJ3BbkHW+z80l
eAidXjtsjNeCdCL5k8yZ+4qBrKtG/JpBrhh2AE49B8oNYlYxarlEF7lfFH1RC4Ex
KF81qEoqlEABVfxfoe3PoIDiO9HBC633Sns8/0eOD0eunnjgj8AuKlSJGg3qnk+J
HiHThr4k3Fc0zBPaSdYSXfzRcoV+uvlQhrb1Iqnf6Zs6GctAiKLPi6oTHF3HMG4s
7UPkBbTHlmDlW/ZvxvjV0PcLTPfNhLVfoi/I7G7IgWILhSFnBKqLAcLchPY8m/u0
ZbviuSHKRVg5ik98jAwWXefvUSqSJEgJmJkNcLlvK/542OEUj3WqP/9GA3whQQnD
Yz7ZZa7qcMGJF/zyjUdb3+rKJ+EGAGSrbw2sI0g5AfGgGTryy/0LuvmivN3Qxjge
DiDzcvO2Y1oJzYLfJoJZzyjbi9V5KJUIX62FhPLFQpyEkGVLMxAA2ziEfaVunYSf
/wxqX5jWJLrBNPJUZgEfmOVvVlEfy9ngJDjqKhfSiih2FfTWEeMChDNIC51eujNf
tBbL9ENYl7pFEuJewEkrnQL+95Y+5ySXCf/4Y+S1fQCnF0wh077bKwBKJGhNWmdG
xsgMKhLdLaOuLAz0MRWeMeeMqb1cqSeFI09CkquHgIxrOvIEQDZkFbJP6M4qqzuu
9LPDcrVoLqqky+7puuDsFECWuGQKkpYsE7A+EXfIFD92QSY6s4W8X/hkXaq32IRV
5HIOoiWUhp4NkMpvhN2xsXQIhM2rYFf8xPGWEyw8avdC+KQ0UoHKxKLL9WSOt0QB
3/6tZKXIus+BVpJrIIAitpWZgtg+VlxW0tJ6MzFRjMomhStVK8drmjPsch0N1K7J
F1q/rBQp+JAoY9iWhkM4wTLqEUkGZzgngqjNjZW0pkUZdYRsCRhQZCbrs6cLOhdh
z+h2ED2FKpmholtDyOU9xn6gHiJlLK+lJktw9O6mcoDDuS7P9Lw3dkqUAp7Qar8b
X+BrnXEN/h/i4yhe0IXzozjHfQafXOP9y55ch+0dKbIdeoplkPS+MORPr/bM7JqZ
e+xBHAAII/RdMqGd5+/29dg2cgON8gZTGog/ZyBNQNg/gNET2Lu9YQ55DufVK4e/
kE1mRcByfDZr4eQJs97mcU+BX8QO1FCcG+WnTDI/njM2OQC776YOuiVs0NocI7VQ
NwVVhf3ThiriIqSgUvOqc2eWN39SLMOqQYhiBK1bW1fapghd701tSSZ73wiHpYAw
SoJ/71eyRvkh36Xk6BCVD8rZTFrgN1mQXCLJnKWUiQzGCNq3Z/xbg49gtZKlaiIF
hrnZLdRzIybzn3dhj6YDUW2QvnicpIqIhABYDCG4OR1kxm9UJKaxflJJZZJVoYhL
s5lDR3rFw1myjSj7AxWye+Bo6L9Gb3CRtHqV4DYJw+/ITbvcoUKXOVjbctxFva2H
neAXhMpAThLVoGOzZ9xlGBdCLJhOJwkyW4xN83IiXeBDPySz/vpdIO4ESdeg1+ro
z0HY32fs7SO06+FM/682lVDoOcRDKZB2WmT6vzyJ4Q2eh1VhjqHU1dtz0eQ4hQ0U
dj1ulfLZa6aVHd+Pal/fUpBezLQIEYl1E1twGLgA+KoxT4zYX/dSbcz8A26rrCRU
z3Lqn1AC1mCYhhf2/BmDFEGlqfVpVhABrNvuXRp+UKcfezq+R7J8XKZECNy4Yj+g
Jzu2l5Nj8JZ0Iol2Fm8Uj70myJU61aG9LwP6LgC5lCPYofF8OkCfySpyjfxlzJOb
ci9HQ47aBCfxqied4n/3aNM//UV+c3Ep71vSwnZV786vbShwNtfLr3rKVmog+kog
je0dWAGrgDZhUaTp0+TBkDUaRZxmZX9RkWRk68E6t9Lt/QM9f3YgB7myDG01SRxI
JaGobgQvbyLtd+CZ4oN5uML84e1JbcpXS9HIj+9R+INdx+CliLo/NcPgYTnfzqZU
c32bL2AvbD1E8WcwVTJqP07xJJNRZUd61ht0J66qIzOtBABl0ihxRaeovAIeuF8Y
vHxkQ5jVBg/74UHYSD3ze20NlzbQkVC5LhRtfhiGSgFHpAtWfZ9zJ2vdbfNQQoLT
NhSxsOJuH+9QpjpD1mqGytfMnIjoxl59ekzv0BJ+7HH0BGVRuVSQgsyttGHmrp3E
Ueb4j8lpnBo32R9t3GPQpau37QDvbWz1lTNroK8YRsLATW9jHzNYAYFVoo8tjox/
Lm8ffpMieXf+qEsPGT4qJzglAQwLgcVH+KeR4VIynHeyZeGycz50PSqyrsFewv+l
D/lWD4P2lRV0dAHYVnqVtpSq8HWUTXioknNcOAFJQYpN1RBwuM4eY7g6KFP+hzfQ
KQ3WaySuDkxlgp6HvmtaC4B4TfEoaqKudZL7igHrxOsNngCROqOLnqhpQtMQRND4
oXvf4tUunw6r6he/J5vo/8usv9EXGvD52inVKyfuqfYS3KzA4lyq+LHsyfxxBEtD
PfctLoCQrIJ6z648AfjyKbcHooFano12159fvcHPs1FKjVMHZJOtBSJj3Bm1PtrP
b1iGMt3705coaIDPwMWpCGt4LJsOzzkzbaPgU9zzizVC6RX4PDeAXGSE6K3WozPQ
PIy1lnv3pWOnBPp25X4Jf7X4uTl+9TYY0Pqa8MK2pNSCe3Vv3VPPG5ZHjStTEnwd
54SZiNvaZnIyV4qs4sfx/WTCDWxnhuLtDXyGrF0yBVMJUO10EHyfnpxHiI9J8Jsz
NBZDMENEeZXdMexrfA+hF2ykzX+qa6FspIhGWss+gloMqg3cxCtzY0agP5ceSAZL
YqJdj+QUDrf7qS2V+S6pXPktCwF2S2GFYxVZcDGLsSau2O1iQsSSibRsx0RzD0Ta
t6L9PhHTmCGwbSu2E6E/X4NersxbYqAax36QXt+u30SGgB84vvzF3kofa8wSWMRb
bGLA5/jHe9HPBNbkqIZ+2TlRzeNtBL92mlkyycU4C9jFRczw3psgWhDqSLzqYFBs
UDfIafzjH3bbmUnAfrkd3NV3fIAfc/umLwiu8gF+78FtqPX4i7G3bqegQKl32ue3
D9obvL5thPuO3hx8GlEYDg3W6HzNRjYFuETjKBIU108q7JdlPpwYR0wa7tyO35QR
Ws9QJo4VdsMD/uPLht+Lfe0SCZH3wfGvbAxwwN7/SoeF1S74Sx1i+PuBACEw2Ng1
p3JRBN9wZ3wHjc2Dew4Yh1Z5OYaSkfTDurBs3LtoOpDULVKrE0Oc3KLyMAkD7dQY
5U0d22Ukcb6IVWgg/ryRCWvNKdQvvwuM9Ld86I+d5OpwwiFCYnfO8LDq1I5TrWPM
dbJ5CFegCjE9calixsznqX8IsxW2Dp+F2ZbnYkTY2ZRLgwqt/gTKq1yMi7kW59UE
7CR+AiHY3AVDM6zmAc5u7G2cEDesJiB70mri2T2uO6hk1LXXiXw3vDSw3GLaYQ1u
5RGuTukkaIrx9hZALOuJGTZcBzU7ObPOZO54/lkmRPBazbW4cS85WkwnD/vPCZMN
APsYC0p9w0mInWItHLcVG0KSUT8hGX+jANEn2Sq+g8zULtaJdYzc1GHjXlObBY2H
zs/3vhgYCaYjoJ5xAKYlXtmeqqnk6nX+QKtIvr5e8lkAwAUb75ksVJ2IBCFdMQoh
6dzhYOdq58F4xhbWpYqRIKrTg2V+XfcGsFX3oaiLde8WG55XUvdQulmBzA2dAzcr
iUDHc62FVK2zLSXJ0CTAEsgYV6QG/FdaBqgyaB5hIZLa3AQonYQp+3+S3BtAucJK
kvqHFrWe2i5m8ht8hLuGh5uuGN+VKnRxed2f3Q0wPviE95w5z9egFUHE8aDzYjnC
v8qfJwhMkW3taEyhQnQjZ33M8jQGoESdI49ZY7RNBQ60pskDboSbTyq8gdl7WpdZ
3gWHWDXZjRq0rJLIt2uLxME+Ncn/uxT5UmdLJFueyJ5WYec1q+/Z+qJL8TwRqr1T
/ZG9Tr+QjyBS2Ygpn527UWsFLJ6rt6WV0/uHbI75F9YxiSh1Whe/0ji2PgsB6kk5
fOwmmE/pqw6PAQy9hwKPo++1lho2GuefN+KWvcas0cDURyFY8GcdrgjXxTL+LFIg
va28x/eLCJbnD0w3b+SUWRmQRLoJUbzkkSkdTw74FqlCrFDc8f8ZUkUDc9JI65Gs
aeS62CPQH51SxIirhDMTZDhJxqsEFioYAAjoB+UDkUWdP8IHQSRTRCbre5wBPuhN
Mop9n8Nxt96J3gbu3unmH/xJiIeuS7DOFybkB1/gdOl/st0UBLP0cXrTaIMcI6MF
NAse6vLetkCrj1ZTBpQsp+VNvs5YUPUQ1vXA6AHuqOYDmI4OYsX0mhlmHisck5W2
u974JABcej/x3WqySU8SClK2jJYGGWqGzvpBjxQFRpWGbxax5eU43ZjjkWN/GDi7
cC0ezfzAf2xpjtqh5lypRAG6KUCAw/CXfh6xA8YWbabZMrBGydER7Zt8VwZboyT/
EQO77gjRMM9vCVTG5bECdDXUBXZsrV4NxNBMJ7U0SkERFON54OyBfXzgw2N0Ya3X
RtoL3+ctoy1/dZVj9QvmTLEtwoEsi0TeBo8U2Btdp98Zi0ScJjCSnazXVOBWfpoC
b2V6ktcAyGIrkR1RGQ14o0t1YH06H4O6Z9D6+AlK8mNIYKEHjO8a7ZXwd7ee2Q4W
8iV388R25s9XARFt++n4dmyQqoX45ea1Hkk4rOaOtwgwhx71qnLFfJmmotMDQKJq
o6bjVOh/9TthwZp7Ra8JKaDgRoRxi+/XrJav6OWBeonqe70/GnwcEIxhzHu6RP9y
nNcLFm+72kY7Q2fPzxw8eOP/kyZwsL217aCPwLUKPgqNJlNN4IsxCxdAw/qdlgHu
WaeRIFFZRLa+dHNMuO84Lur4XQ5tbGZDCE7vpF4swvM1wjs/zwHOjXxk4coZ2deJ
PNFI2+AKrBHLr3ozU19wsT0BOfqNSKoSy5jXB/phdpmhoUlA6GPyQz5BFtSkdSHj
uft72t16fuJ7FaGcYXLlmfv49Ge8FAgeUgb3tE8COTZrKy78H9aNlLwVkRNfcwIF
/+yy3dKyFn2s94/ToGvMZldTC6Kupdld2nSTmU08jIOZI5lbxJUHHK8rSSYlC6T4
SQw5xTP1O0b3FEkCoTU8MZ4+0jGLju0vQUwVZRnK2V1cAh/QEqesfrxR/0EHvlj0
UsHyVVZXVc6PKpnh2dYlqLEBQlQcZtmjFTetTTU6k3PHmNZuBEdGvKBjLE/Pfmig
9fslM3+JnZhA5HkUj0E2Am5oBe6SYVkb3JZPb+DmgPicLkfroNGrlxRdqYNw5No1
zqrfd9Kk7MajKFmF7s+Ovf8H7Zdnq/ycBm/p+jIfLF50ThnzrLpbV13jwMxugasz
zwXLDFo55aQ68ghRI8rF6CjLZ4egNnxO1yeCFgrC8AP7516ezv35GGogaKKRSDeG
bkST1rUtBuJ3JWD0jhsZ9XB9eLlNee+/MchzZ+VbwvLpRcyY7QNI13dEBobgixe+
RWx84oMXk0m/Nnl4+4g1+tOCTVJ3GONGwswJxhXMHlwsoFzDOnwHIWtSDRf/dJc+
WmmbCUFKJdI8pybZQBzBuayShCgFRLX9LYJkal2g3wMzQ6+uWVUJVyeVZ/r1B8h7
HnliuNDuZoinFI5osolXauQyfOe7AV4KrwIIwBr3SQv6gNFrlDi/VShEDg7RfMi9
r2TD0hxF8S0TPKbOsBYGft7EpUepJzcJQEZq73a/RZw7bNd/4Isc/kH63oJwmqup
N4go0H7S3kdZ+YeF6lD/bPkKcJ8F3B9Vf700AaqGs8UBeY/Ee4ULcsrZXZb43FQD
v+D6GYwgHnNEbOYvfUkp4R0RFdr3+fvgVlmL1YLOXYCCjd4JIuDZenBVdCS7CEl3
amvnKgFW9yOcexSkSIeoLAdvw6HBN3K+iUT6Hg02twyIJFqHBd8iMf86/29mWZMl
0MlIkm6dxmxg7kIXVhSN6IDQFk30FXofUoa2atsEJwpOOfuXTRmvnw6DZovyN8DG
M06dl44MC64rjRBGTdqww9Qpj77sppamQlSJmfX9V4G/53EEYn5ITXa29b6cEWnE
mwAPQqbQJfFsCXjqsjzmI8GTENMjgRsuGZ+zYKB9qqmrLm1AGONK7/XZ9HQto9m1
OmbMnFFqIxq0RudB1fP50hub+9rLJJd55m87AMOkDIOQ9gy3O1sG6xL5zGLhV4Hw
hhG6BYKZ5RM2lddbBmjUXkl/ItY085SdQZUDCCowPckNKkf2JWWdBevkx7M3xCxo
fFWCS4GJ/utzzbtfJtdo64w9H4MkHo/oOLQRDll9KSMB4Pr5Y2FIcO2oY/pdQalI
B2hcguOUZJuvGQMQ6Qx2fM109cUqyliyCxM7s9WMpAdlxJAqjUYloZ+zTZNheUPN
P5XPvN0LUmG1cVTaV6SfuRoNaGGKAxPEuC4BvZxI+UsnLA3QnjKVz2wcZTcL79sH
rghA/KxJhUiMIyzp5ghB/VzRNH4sUSQ7c8dFWb+g1Xf4YUmIjnkX2/2GTTFBFfnA
tyoJds5qqVn+FldmhIbr/AVwaZupP/5FB+GSLxaWoNBFOtflUWGSAt0Ujcj4zjwg
RjOw60PJjZWhRhvLjJ6kNPmmywBGgRXX+udA9QZzR1OwfA7SuLczK32tpDnVGsIY
1L/UVCctafIEYrfuB60hVjVL+ToDs4K1KmUV4vk6kLnat/vQyQCXxKL7Vbllw5sR
0o7oZp/pSL5MDpVB8aDRBip7M7mqTmQFc2TgKxkd2TLS2CCoDL1cYVl4kdJpM4Wv
Elocaqe4MCGgvonB3lDchopZQuKLDuqrQAlf4j05MhS+aGab3vrkfxRaQZTflFgq
6hDWiY4xRpc/dwTUXq7i9xWbAOB+zvcUFnzFCyCI0ljt5bVWckrthrNl1Be+2jgy
ZnbAqRUPjfv9WkNcf0GdJG0RRoCQTnImT4Aji2/0mqilKLM1U1DJkdOaC3QRiN2Z
StYim/mygr2rqvAOO/AzWLNwzIJle+HUNesuQ7WyFVQNJ9Fqz4utDR7YpkUQOhS/
mBYhTwQEy+Pm4Q3ldhdvfoGR6j7dLmOVOqGHNBkj9mx4cbRPslI7TSmYtwJzFhJS
kaUhZMVXq2DR45LJcrDh5XCYbfqI+oma4TpnWXDDATo8Fql/w/2eCIwoVVm4ljez
Oufjilp5BST3HYQFLog96BDoUvE+lNyKJ3h3EsbRoy3QlW9bjvlRaGtt61mLAoGw
+d7df2jgFLrzOqnoCLmS8GkOpvdsXmB3bOpNiZ8U8D5fkdGYVfW6J985mmm6j3+j
JS6GCWOu3ZYldcMvq8Zca7jjRnrtFJFvLXdXqJjb1eiI7v0VBEBnEGYwvgA8iu28
hOAvn/G8uZyGZBaNf7oChZqmHfEL39ws7Kr7+kUPI5tlJukAZv/jF6kF5BRI/R1K
PtKMy3ODXDkID3O/EgXsy7f8m7mJh6fZ63VFCPzjxBOu23BV/Ym/46rZ4CUOMlKz
b1zidX8vW955EcgYCVYfZinZEA2pwdKR0fgF6NfbQouz0d6iKJlQLFADpvqlfanO
8ys5lGDerJbnnX5yGlG6ub6reJciZczkpkSjzocVlKkdCrw3ZeHlBmbzGvsO3wRv
HycTqsL63UFVU8IzHo47uwDFB7EzyyG3e4nHAw+AsuOot0cCs49llFg2gyIlqYNi
UpjFiXOk1REiw8QW+Ah7ueDPntSoJg1dgAWGZkIvf1QnE4u8fAZaGNPT8rCZgppP
TazN5ESqEQLOmcnhGqbR4KTrFrCkuqoLap/fxYpzUblf5noQeBJz9aSZXNu/txJH
XJrXGEfP2qn5sTq38eQy8IN4PZJTdK5fU2PzG+AEdI3sTnlNCQzx4C6Dxk2GMtEV
b/xYA4y8kAZegrphhiaKdBf/+iZgugX1YEclzHceFYUk2YgBP4ShEdWLLKYR17ak
F8Sf1m8uuIj8SnkDbLPawULTCARG1HR3+Hn7WddbOwk9LUTxz5WuVkZt0jbD3K5Q
m1BXqkki3uPxJ4/9Mw0DIxlpOVGa5+fTcLpfwmAxtO6rsCy0onExBoc+Fw6Pgazy
3V6Nuu+k1ahtuwvzn4eigwa9wNGS73dykW07edzDrZ9kO2RvEDjgy0Wrl1lbdXak
Cdrq55Mm7bYHlfamzdYlZD+Iypu5+m8Yzup8Pbj08MJ2O52vBrIE7FELyslgRro8
JM9mTxjDJyrq2K5oMTjUvAfsfMqyR6+w01frGAyoPJ9JlOgQg/slUV0tKievudFf
/bf2nOc5sHYxkqtbucdvAhLuDgczpTVAfhe6N+PqXfryIJNLMqGFJ1Pthq+e33SO
CLD8yqBdlRftscfPtJt/AnIsMLlcGWUUzjPiK62oP4d+ueG5Krhz12MpcaD8XOdv
W7tPmqSjdtQszZ86tevgw+45Fo1eAm94lDdOgKuJXD4SBfEIPB50FhyTmtH11nGi
K7X27bZ+SNmfbH1moHHfWEASvHWKiecoETVVamwPbgXt4i0/1w1tj4NQ+lNviZTw
IXuFhqDYr0tGmFfr9bkLZ2k1je3xZjVH0mLMu40ZGUU3exiaEDM3/VYGyKYb+LzR
oozoyg6oKp0r1GkpkgQfMzMVOjLVtSLtA9BuaTcOcJGmQGI79V9m5v5mNETat285
BsLCIeqhZ8ppyMDEdfgkMKSd1ySAkwGPyHkqfY3Kp3lO8x+iDYQFQV026sBz0QyA
wnN3L6MEAFAbunzhpYcRBCygDNbCu1bSgaOLKYzHTL/ALythNcxi+/E5Qa/pN0C4
UFGtGGqDKN4eZhGoop2v1jkpBuRsdg3JAfhMxjy0TZH2/oP+M1FaIMM2B2BoN00T
2kpPd/4P4A92QjbXO0QCbXA8Afl0B7i40ltqh8fR2XCzOWHjDEXYJ16feqE5HRHA
csMA6M2l/oOaH7yFH3fIjguNdPOiI/ZUfpYMJJUambWKTBo0tDRUgZw3vjZe1pTF
asx3NmYwiIDLy9ILy1NOQfjShzlSbunnuDAw45iwIeOkLhWyfl2NS+Q+qA/NzqeU
yY1OztkWypT5Y4xCM1HPi6AXNThy4jhlJPXSUY/pukRMVzIyYjcD6S7rlsukx5PY
YCJfIixHYUawTn27gzSD4b9MKDoHryXla7Wnva76tDRevZca0BfwhcWpt5oEAjlA
lmO4I4xntGKSY1ylf6+qOXa0owLk5ZoFzzRe8BrUVLiMkw7I02JiB4a/CDP33LOj
wKCmLK+g9tnRv8xEZklPCYsiGQSmXNvHty8pjbtu8vmZJms/4w1VS6pxPFbEL+c+
qFYe4u+e5hBWUs6Ihziz4TEErQY7XCfeGfmulm0IWx+SjBuIGm0MtYgaeHrQLKI4
tqvqMTl/K1yFPdhS2N/yDmDlnpjAp27cT5inzaV/fjJe0RafGFUs37fm/aBDO4V+
z4nuYrmfRjPl+DRfGu/G/uUzrP/2N29B3OPGlop1hUzxBCNKYV+0ILthV4RFvVqL
oFAWjaIlBm04FpauNkPBhtzRNc0J7oZijcIdPPYXt3iwwTczOmBdMLaK/0TuO3b5
7zyjlnnhub6UOsWh5pKxJsMufJ+2j2+l3Yev93miWtnjaDSDp7KFhmk20WSAU7Z+
ECJX02KWwDUlHFyo6v7jqVSwd1wNqmb1g+Fvs70CcfsDoYWnkZTtd/GWSZpe6Dp1
L747MdRs+z79UGwyRNEF2Q7Zmlfv0Qxjy4oi+t4XcxkYSIuWYdlAiE0Qqld3+V1A
lvER/zL+/UFkPY/qgT8uEyv+JXWGQo9KUDaJVu5wcKH9Zg+lqoGB8E69N7LoH9W1
L2pAvKVMkLKAHn6ewQNXOk4fPzRzVUPs9Oixo+IZNQzTUwKWWTrCW4oaxrOdSbCL
w+6wNckV4yi+wgsWVmLlUfNY9Efgre8X8BCyYUrD5xSFNM69qPgAwnEoMR4onfdf
qyVMW4ZTDWW5Tg79qDIXH3UJALI0pWYo3emYYN/6ABhg/fnjD8MxrZX6J4AyFVGQ
oaQybFK+PyuNGOdfhWHTxz43djofPqq4vLFuerEJrdrBAOPe1q4vwQi25Qix40g+
ffpXicTWmHGt8ODiGNTsaez5ke+klCXvftDo8mlDNzqP1Plxebl9nfTEfwA/g/eu
wtkaaQ7dBq2Ell1WFp1HmBx1UTtJWyB0SSW/rDATAVo27u4S7uitudwEKSC1toI7
zVn95/Ulpq5dLmUiKegFfEqgbsoHhrHJa01yd6KmHE4fAe+73SQJl2pNkD3vNCOP
+hUoFJXL3/pf12D5H3ZRG8j8VAInAL76LuCUtwdxJKGhuRUyrUBvl+hen8HfLuFI
4ZbRpuo+oYmiv0yu4sDw8QDQoj9VS0enoqPZMGAQStBMo3r1eBQsEQ3SHb6+uei0
IHdATN7K87s2/PvKnu8wU2/s3AIHA9UwtQDZF91K/0a7QkSbH2StdikKFBpkkJhK
Zb/3s2tBH28PDZvrrCcwzYxPaDTSXlqJYpvWYrPUo3T2owHMlL53Ntf+SS0FOfhw
/TgPsjk6ne7mzU3NzwkgGY89W9PuzrJH5BOaUbXP9IB7adbjqbyj6U703qMlLmhy
HcpWxztCh9WlgSNIZL9otVO8qW+69CTneEKrbqRfMS47pZL+SZChBLgeBrN2fx4e
Uwhy5aYUxQNXBj3VNdoI3+lA6FhekJKpTDUCkFrEp+If3g86mOIG6YwwpU5XQBIc
Yc+xAhFjPQ5xEOEuvjuRvo1+CckTnvhpBvj8n1AzD3GYBnMwbXpSr/0Ehtv/nDeL
iGNngZJqVemW67wzgoqpllzT20DKJP0whDB/59kovuZVI4gcHsNmFtVD7shX97ga
RBddtTieq3Siiqctz59KuOzXOPs2jzmknvNd62s0QvSdZtJokVbe3IU0ml+Y9YFZ
D8FL8Qsw0Pq7eMJ38EU15g9RMyOG8hTD234isKmHQDBRQyuhE5aT2ym7843FwnLw
MFzoM8OzIVm+1JnhoNCnwZuY7Bc8PP5bnC3j+pGMbnVh2g4cd/s57nsqumkCXY0c
ytOsS9hx9scW0SpfMkt1ix+cOB7o3St2QRv+6mAZ+BvUwobJlu3HAbK3c8mVJgHY
CJr7WH3u1ODRITpYpYodovYnSE4KRSv1rs04BaRU18smEdU8oQ331ydFZxCK1Skg
fj7jQi+eKCFWU4+TXSZZl3bdOL/DcYf45mloYgIBRm+v0/ZVshSmvTPPsMxD5avJ
RfHxk8Tgp/cTV+C7nXZ6enA8MoluQf7H2+9y5U3oJKvzivAePxHz+A1z3eeuLO/y
dWOWqhLnUqmBJUJ9xAD+mYmRbcRoSrZ4D5PRXoK3rYyko4TvOLmlqOELL1r0vNhc
4bNrR4AMEdsYY7vkzdAge8BYKonRPNp4nBfOz6jUDjAgePIk1vT5h5NadNMRMIJ4
7V7DCsoLX552cDOszmH6vz6CckIGnvQQSnxynLh+IiQyN0ajGZOAGQqClWtdJFfR
qwQakVooyR77dMqkC4bBbF0IQkCjscrQBIO2ehxnqWm30/BUIjcXcmaFXWvIKxct
4UTHLwo7+qtnm253LRHQx5nO+I6TbxLqTbcX4NBPgx329tb2i8PMosUHUF5ZyWua
xH2XvJGbJWKMyvzt/AI5wUfZbpd6N+7+I3jG7/CpC+9cAMzPNvCBBdRoAvb7t+JR
05P/ibXdQNi8bplLAcZgpKaedkBavNS7jYWQ+TDa8aaVibr0eRyFPIiP6l+9uGFi
UECbsgsvEmbTVrVmb92lXpL5A2nqlaKofcKpIN91CVQ2Qerq8gd8IiKjydHI0oHz
fYXuSSKPiDOtyEj5+R9E6JJJMKHKT1EDd7EVFAa6A9GtyBzmvriQA3/gTBWvzevC
T27nx4/oejjhT6+pRgFu8NH2tneX15jlOtsG9ewfSddq+tIiTWVEVU9fBrl6ZZYP
/K/2iAI6zIDtWa72sYGZpnw4MVthVkVS+eUZcwomUz5s0JQAsvXZGOMmHH3RaOL6
41AmM/9j94f9dIMJgKO0+fPBZ7S9F1mp7KVz4IOb5yPHTnk4CqtsASgiBMY1SF5I
OQk5k0Qzvn6mueJs6TzYYSJ1JZxdRwfg/tL7XvSiIJjN5dAd2PBNErpmvs0kJWeN
1XCmK7s+WN8XOSasXAzoilDHWuC4n0Er3g23+Czaht0qr3ZKo8zG0ZpVsPsfsGcR
NWECNFOMK2hKNxmc3v4p/5fBSQF0Xql9sBcfKzZpujs183Sv2l9l3zreUzgf/X6s
9odlDLM7eNc10tsTSWwdSuE/PR7kLfzXgflCWv9eWuLTQpvzD2Yv/i0aB+W5FVlW
Nt0qc8dWof2p0EdbBZ/nvd3VICLN0ZHrP+1GqXiJ4fjro3ko9yW5UEy6ZyJmgGPD
Nrl7mlFlYuBwfdR3WmuZZJsZveew1OrUk/tZueA2b8E7bG4FzZpDaExbsdgV5woU
gnMogP5FjorrWYM36Y+lK29/KA3IuvDk/FnMoG76W7X84NiyJcTMuiZPCnYsHb9A
x8lVxuKOI9lrG8LVoY+1ckNoIJQcNqtrT3KY4Uq98PQcpoonKZQjTNGSKz2CDT2H
c5bspPx1MryOryywkA4nzS5iPKUBWEZcZfxZLDTr9Uh1cQJP8V4HxEt5rxm1nAAF
bWIXWeME6677D4svaToJJKyAKArAwIPsIcHFT/c7A4U7IwADlkcgQ/+oreMSmoOK
nN4d5rienr2tjG7K8tVm0vUlszwN7M93BFakarlcW+t1Fg0nP834rBHQalKqlRl4
rVM3PUGbemMKHR1iyQZUjzBey1l28cYRGGTNH3uSsIWJ8XHWRt5AoHk6i3BUFy1+
uX4UaXU2rb6pR0Zlfh+czNMCIsa3viHBDsI/4JeBla97tE4RgGXmi3+hbiftn4M6
9o8VYetiWW2hGkK/ML0IbJxCcZRrqcGJbtQKBRGFo98QOB8rrxQI7OkrrS+6Y0gm
uKjgE+SI5477mGWo1h7j90fvcqejp58CmXJzBPdJyjfo3XPd/5LDlEXrG8H0VpkR
utghXRoGID9bpkOOZsIHzKqo+KEAGB1Jw5KMuHnOqhqk7fQ/OZzsUD4zDLEc7j98
t1KBTQ+nOaAXcT2W1kys4zN1CoPOw+/ai+rqYpnbXzQnbLzcDygpwG+8x0pIrEsJ
MXlmkseAtLdbVVn2olnQJAF8aztvvbLYG0md1eVBzSSEWyvu0t4itwYMAAVuVIlT
cNgrrjSfNeurtM1fMcJgNkUz4DW+JL7Hoi1h9E5aSfwhcnww4fs20f4r+Htfgt/i
f0wJpCIwgdbdsbmwLLP5PK4jqCaUkHW3HU8nRkMrq8g4vhaewXov154deGOplnu5
pENtFPwrV1LIQcZtXhpdX3P/0BTfqUg2NJLOc9GZR06RE2xgCRzFmg1mp6YVFl9H
JQVrYIL9UwBZfw3dYfg6AyXk9fDrBPaTdOXe3OrLCLmeZzRlmKfTs+6pwNnXixB9
IHEywbHhZi/NQisRtjdgXBtQClmTdEZM2MT2WCDXBlmrXBD54ekpTlU9fOlGYZIB
Mq0kce2pceTWyXwjnZjIAQLC1q/YERGRNLfjjzKkzVQDNrx8TS2vr6M5Ub5QKnba
eWkk4QFw8GLISmpeU1ASJYBJ+u8nUT/quKrREbe6rF86mUVsr/185AT+Kw2L3RDe
N1ygGwbEC95dXeAgMPkGxmSLvq/gPfi1kGZ+d2SQn3aFSDVNaYGknbVm4gg+ZsCR
HbaWGSfhI82s6WlO6m+Kt6AnR6QZP+M0+/RCcHAfmClTmhtzJUXa3R4hYiuHpkcj
GmAMeGWupgnhoWHerab2EwKqWq0wMikV+Bk5PzNLVilhdGYx2jj+BYGOTTBN47+b
zOg+zTVwagUBzWnmHzH33/+sYrlYorezPsShgeh2S2jV5ENwpuxFLn6wbN/Jsj4O
YkPvyOmGK/o3fT0kgjNyO9/E2hhHzvV4+Ob6sk0lADrPcK4nF0474spkTuFcYlAs
Vn5MN+aD+JfaJYynXV15Go820hFVTiDhFXsbBeL5zH2baSQqdtrJ/RKy1GN6sktX
0ai0B99Syk5lcszg/8L2Fv2cFvtAC8eR3YG+zaynPgyIOBK08L4snJI6Ri3pTTl9
2527zdFurH0we/ROF1DvvR30EonuxyQrllM9LsQHXBTFWqApAlwj3vTZPE3FeunT
udZY2R7nswHzHCaIW2U9xR1cdpayvsKzz8ESZDyS62MMDrPlqSyiZyO52BR1GtaR
Hn3LaeWFeG28M7AbmIuUwhh+iazDZMIa4+Z6lko3f0bL7wJE5vi2mr8m1KtDAczT
s2V+Rh2nQgEY0NmtoxSa3EZYYItGNMm/Rojo1Cut6EpzDlJm+BbpkoZLSpPr7drQ
8kS+Yzsiigd9H3pkTwNJywlDGinIbHrn/pKdOK7kRKV1UkVdj9GtAktkt/mumt/y
A/EE/HEoUhXZNodKZSXL3xkwuBsWCZBU6kIgEZBiNyTGi/nPatsVLXp9uhFMQwk0
CJ6n747roEXqkEvS5ETiCil27fxCACHwXue0WnFmI0N3cOx4TNYjlz1UnGQP633c
YlmrqL4VQTkSBhoK14qfJGceAbvzQ8HwDV2rQSbCtBw4CleWmYZhIFkskRUVo8V6
O/n398e4gXlIFQwp29588WNvNXZ3OO1bUXiFkva1NMFvjxeMh40u7LHFpRXC4pE5
6J3O7s1OqzMP2wsWgESyK5kBxBotQxbN9FlOI5HCBuyIZx4eNbGpFL0DQqdOxEtJ
TVBgxBZiiKDiEZVryUU5xJQD+HZfM5Od8CzX3lBDeuc0FhPCMcU055gYqVsvCsQT
cVFeIL2OsGLgLZEMczbegfVA+XJG8pu6nRBr1QAZEFYdT9RI9TS8ThOF1hEZHSXK
KbXwA/pdaSAqm2bLIpViv+QLyTEhhk0AURjjMmU3gOLFmSrmMonDvCspPGSnSMFG
o9ZHl5dsfIbC7tH6HfrY60DojJzkc+BoOqNz/0pm2KYMmNR6MqXQj4UPPd8pbcTw
jOeTEtp6LiFdoXe/fGaSKZsgT4wQw05PmQ9PPxMFVrdVwOvxAxllKl+zg8eXlf5S
E7+LIr8mZyIzy+7JY7tqy3HWGTLi3zGps63YtuLhb9/EHSucsojnt//LiUiA11tf
9q61s+UCx1rvFzEfMQAD4dh33RA+1TdildWVGoPtgyYYW/EdOjuDhpDH+0Rzi4sa
SU3n3rux4p73O12Zl8ILv1AVbtyhyCWyc2gw46OUEcrtw1SCekMc1Y3Fm+bS2wsc
0W/kyTnftjd04sQMVMFseOaQb6N2XflffPEk/0OLg+oNxfKk+PHS2RGjuj+Uq/Jc
yNGDQt10/G3TSokC0Rmm/W6VJsw28fRE+hAZW6UxKfXCeex3xzSyEp1mNmSTUeqv
8j1jZrdaW8rcTO/SczhViLzwl+oNshH1Nfkmjb75JXzH01HAdT/mwAZaCdhJPlRH
8sZstcs2ju/FoFnJ03bc+3/SILvG/K0aQVmtWNhrqq3FiAIzfGuFA+ZFTrFydj+Q
zr5MbupT7X7y7W8HKIj/b/B9Pr2sXaRzU5fcVc0MOrP82YB2lEUXHFsJ65AfAbWi
DaLk3shNLsdWOzfJCDRPEi5ukiGiCAK21ribe6GNwxgsCRarwt3sjN/34HjNhQ69
Jr177KY91Wl6F2NJZZP8E+sSsQLvQWy79Ttf7tBVKfdbEY/peVJVaDj26BJ5eh+9
yxeis7DCm/7qZe0d8gkieAaEVKG/B+xs3wXZTOu5ItSKlvP1DOUiiSQ6iX0b0/JO
pqr+17YlsS5Llq3GwgtfGISVbKkNnkE9xXXX1bhcl3/MafwHSRX9f+kDvFK3uW4W
OYAzJpv2lon/217I+RYJY1+wOFtjCbF4vjN8dCkJH1K76tGvyeAfI8L8kfKLRNld
3XaaFTKw5JEbIuZl8HKzgsnAZ23jIT4iT2EA8AXRSrrVky1jAoTR9mGc7xpYLgLM
b/5wedWiNo5nHqudem+Wu1CPgjvwO61/KyeEg2GthNRztWcn0+PAP6Msu2458hFO
01C5eg/wWowf+H8g0GSKf6zphBMhvsKH6DUStPBkzHEI8AESA5053YAcxev5HdUA
r+lY1VsFtoy4JdN1vEykC7RO3R0S/XXIBkygSN5HbxIBwh0IRzGrpH9W3hw2FDmc
qYYdUrzdd60X9jmUADaxqtjDFgfmRzhRi34OObte854qln/pUxV/CXFOjt69OqqO
5Xi2efczmXSyiZlkOMINkBbZzI1tXnSwg+zZCZkzw3v5h0nafbfEzNhgBo9ExBpQ
cF5CpfLyE3WoJYxH9KcbMePfsTQwtRdVF1wNlggcX0MUCe22BwllS/CBe9YEXl9r
6YL2+gN0r4E718pOCoLSgMHwuTDOrkfnfJkKLIJo2laF4hNuVws5b5V+Jg1hooG9
H8lI58YnZ2YQXKz390qWF6EctFUNiLDIzcC4bis9U1SDZkQ0HUMPx6RIXybrIRUD
kUcHKZHAAA8gf4iLBn5oonWoQGgg+3HJc+Df6dRLe/Uw++h1K5LyfwVy+ago6c5+
iPBIoSfrrt6r+95f6EQNVXORaqobdd0FRJEB28M4aPN1llPmZcSbegxXz2cQ9NKz
rgdpMcgHX66BTI8L+11HPsLTnX/RUcsDDsuPl9lzwPRbVY/xTZ6OLlFVkS2eHRBN
MY5sSYDPc6D8qBD/eghRU/7mCXnw0i7yDQUjcVxk7LJEgtXx6EfETkAOYOQyCauQ
sCoNF4EVocpCno02VaoQb+0qWIgjRbcbhlhdUylEpsEo44c+Nv/clpzfqpJ2EY7t
2dzMBqLKcufcGTE+ih9foTYhOWuzENQRrsI0M0m2vIYj1nv25sdzx8FVyKkUFM0q
Ps5fn4iUGIao6DB3TxUBa6jbIx6ipQFqXWfcnQfTeT1uPuZz121xICj9IJDcicop
OjhAKmFTT2Vi9AVwJuJ4BkuJ6Bke13X20duyoQUlrO/dqr/aVO5Y4Gi13Klsph3a
/i8w6kIvSpaAvq2CDyJ3tVkT0ekso9I0vUk4uMQ1C+081l6tovyw3rEJVr4tfADZ
XGSPAWvMSjHQT0Mds+1fXfRURqhS+DUlSvniwn9+7nwKgC4WfVsng1wK201bnjN0
h6Pz2TQFKwvGZ3WmSnAmqQtylM2N+sIBifYlX7Tfh8PTOeP/c7Jsfg3ZbgutCB8C
A3LgN81ZUblHeN/3qmgDaW2jb9UBJvfnMKPBWTAf8Ofd5Y+tDjAjOjj4F9Atixrt
Wd5Y0CKIIdmi7TpUzbRJ1XhF1QzHtNqASMsJXuzRGe2fclMJd/JsEWhQnJqd/PLY
LEm4Si7ozlrylQsc8MhjL7mzw5K6BBeoStMEv/x42EGat1tBKPT6mkUZXh2O4fPZ
euvxAvvmVCC1+W2nQwz4+FgHrpW/Bo85pjF/xM39Gvcn5IgRWTWYpQdzmrtmcNiG
lyrX7Zmkg08TwbETBGEtsrYmf1PQZtDpoEVRDufze3URpewTxv2MTCKVkrIT2UFL
AdmSmJCa0gzUAiOZJXcldleB0KXAvcA2dIcFYN8AyJFeNM3TsJxN+XhLQSvYbFP6
vO+uwa1ENqH1qcdjg1vdgsni9pf/Qx1r91NJjRVdj6fg6UMZBbMkcaB6uMA44ahP
VIs/YD5jmkTmtDjy26b0gohHgNRItnbpXxD//rKuheb5jO1KA1aLpXrcfDHgz1mV
4lcjXgvOqaJpNWfOD959WFyLOvn49hsMBaw6/c+EhPzMSlZuLlSyxywQb1wsDuUq
YYGcFTtrswwUCzdwK0G78fTe792JrgUNhLAL8/q4bdF4tQ9M1SQaOWywxdw8cGaG
QF+j03DT8njWzdMFVBkaLNqv3v6sL8anH+pTD+qYtYZYD0gK5igEaTnnEV3xu6Uk
RPRlub6CDtXt5YH87LSvfiJAzim/hGxXv7mJc5K4mfmJY26fJLugOg/hLABAk/Zw
Sxwss4gOVvrJQS4QjeEEgCy9HRki+43QKL5rLQ7Pe2km0pdfiYDEez0CgIG/FmC4
s03UqN0bgSC/845Gg2jYGyanhyidsgjJOLMp4rrzeeKB8uqXmfl38Ocevi9Dff9D
5Yqx1bUWSBHW4T3CyL5VCq8OicOKMtIfwp7TDIPiOOaXePhtVivh804udY4+iLhn
hVSuLO/EvS20Gfe3V1wrAWZOZd8XkTrWbGHZ/zZAWEkMXaBCfFmujauebHmuXx0T
tXb6rXNCbJTC9mgICUFaMBqDcyyLbA7mLIg5j2z//hZKayNtslJm1iCv2RI2NsGc
vIvY+r0f5F1FmS+8b6n10Z19ozXwlqm1yF5esZxpNx9r8fpsOYb9BXRqUJYWfyuO
r/BtDC8g5z0s5fxTzUVggMKG7ZQFZwGUDtGUBImx/5qYPM7nb6b3XaVAngz3nOFm
2NYbQ/yWR0vBcKsAG6gqihVRYGY76PFvvYd92SQs7x3fFMTQ2vfCjevb/akh+Mmx
TOq0zRq8K48f5tIYECxKDaVmq+M9aOqXkN9eMJrgRbjx6omPYGsmjKzP06WkoFS3
zs6JvNPZ1fwF3PXtSZtkyRseqjNMAkD4RuSAqbupcvPlZecm94AygpNFBmhRGss0
zQVucMkYFQW4B7ScZa9VdYxIXu5ajcjAw9LLLn2qjmDx5J7cpUwcy6/VTWrlsMlj
l7vnwKdaefNXNEW1oN8M3OHr423ZL1edgZDlv4pCAD/lb5s178a/VVUgUtnyMzlN
CMbUL6fIZl082uYKwPRKwecexxezjP4uytvTyrouB1FD9oMrtOFRONUPdoWbq8p6
ZY3dFCzddRz+Vu5YruYDKtlHRVlJhTK2f0/ag2YsHmVgMJTzqlLNmGbUimVHIepO
hZ04xfkH7deTB0flWEIJ6esKXoPpEcbobDoOMfZJsQMHjb7NFmpamcRG06gZyOkR
yqHSXDCy/vsNzESw06p+R4DvethHEbYK4FMb5Ko0Xoa6lsvk4RBVWnwowbotjPKL
nAGnSTuSOXLpTY2L8kjIkQiCSzqRopmqU9wS5K6jc/suC+GkUJcYSPbZqTGmx1iD
oCE29hBTAQorqtTXXUAFLFmmbYSUpquDes1nI+idL9SKoV7zwKcV/NvcOoDpyyWB
wJCrMKt5IDxChrfap6oRWlsDEb6SYx0u7dGngaY5nIG+zDmve2Hnm8UP+ylHFS29
H2HrVXW2sMY/oD6LJnAxVvorrTMJHNlfpjbX84+HaJUuQyoxRnFo8/9vZGJjibD9
BIkHrnL74Zs9NxJ7WnFSgODgMX7VEOSFPaHFSdeWMeFh+1PdXuhe8ebBoc2aFEV0
9h1lQ9nMjEaBMY5zttiEwaK/BMpPIPC0H28MN1edoN5UwScVTU42NRONm+HFamDp
7VjjszibPeZUHWsPs9ubAipSmoNtjWBXUyTyA0u7Sm1UyeSLmT/go++MCGjmT51t
QP+CcW980PbdTm9zdz26o00Qgg1se6RiVtpC0J6YF671Jj6aXUf/2KNh1cPq2D9J
ZRtPP+3/3S+OVBTB8I8hYwzpynaLowDip5Sz2FQTYEc0b639dV3/s80Lg2mLWJLp
T1DfFgyfoblg0JXV6+jXH/MpuFIc78Mn3OWBK22Hb1lmASgibbNxPwbFDgZtSDx6
f07qKqoofQ5UPU41YnW2hIfoy+cNiEiOXaDseFLb9BToejr5OaQ/FhqJr9TWYiYR
ZsYTmTLF/BFkOfeUKN005uPjo9FKXfJRBA3Or6MotzZpD13q1wDTvObpiqiSMoYI
0XLwuqiO/Xd9B7hTIf+4pFZvnskaU0Xl9sautYJezQTi73EXEnOkholwjM5RdLvX
+g9B8X2qAtwnF93R3yyFm4iz8qMX6ioOiArDQ3R9DkU8pG6900XY1QGC1PnjBuSy
iN09Y7yDUHTXH0m2F4KyRA6Mz7E4p1pBcwRva4FBwzFhKPbmOefKxO5W/s36m1iN
6l6BPfnZtQg9IPM2b/wr82t710glBw5w4oBSTUJPHOLdYvyl+OHA/DIpJNvdjhf4
Cnfou+vLaRAkY54GksSuPvU9u7lg30/uti2Q8Kk3xuq6tZiPQEExvRJrek5oCaq0
OA/dkYNWIdEXkx79m7LnE8vtoXMfvg0e29PkF5Er8yZ9Dfqfo41lc2aLUMWgoRUf
VPFDjVv01vAdUVmxGSkyaB/prnEVnL4KKKi/Dp/eDOEBJIOK0hCeLCM+b41V+Xv0
kJci4Otq3sAXYxXTL8NZFW3KQdrHKcBOfsfmMA5pT9JCPTjVwxskYVnItBP/9QaV
AUgOLYUKolz9ihrBI+7uOIlxZDi1+TsGcKMDgeLtSeorkBPldFFTD3adO64z4qM2
07drTP7YlMnpj/xDNrqLRBIrHsaIzZ2NkJwMS4kTt0uHQ5rjqeGjDnV4ybbGtOQr
BDKQqnoEOWwbluwZsQ/8Wqln2KfNl0ASUdh45S34S/8tOcVNHjFoPlp/44402pBF
PbeIJdpP//Xy/OtdMbsrlkm3meverZfE0iIIfFuNXn67Uuz1Fu03CxxsRTwOrqA5
XE2OoKkk8FhhOhLHKFtFYk4K3/U0hcm70mkE6zUsYSyL1+6oEMNBxuYf67BbCR+5
pwl34S4ICOqLsGK2o+Pwh8s8dHNoRhkcBlMEknfXC4psTTcBFRJAXJJ/6QcStBfk
PS6FuEDMkL5EfP2zz4XyO5vv2lLUWZK/NlV9iWBvyHyPzUyy42Rj+sR7hNnL80k9
1clIuMZHw2QUXHG+IpcPgoNu0OCQ4PTmtg8yCUrGg8fYBKgzjEsAVEUaaWV4KHdZ
CncQYgbJbonPUS8y39ZVOPO1GqZk8B7tx07Jw07G4Wp/cW+qznAfyoZSmtd944RF
mxmHdr3bVpKkWmoqa4Mf3jrRbQc4AfVlIig/DbbEWKjLerwoVhVQtslx6m4XVKxc
JBQe4QmDgbCytudgfFnhjdAxxOR8d1h/Q8J6gmeShNTDn+wpBxlDP01P0RX3/+sg
tE5ypbOtYQYRncGAXFQlznhnT4lyCjdNbvKnstPYbkQWt/cboj3UtawGUCBlpNR5
MEa8KERX4wdPhBD5mAG+9lMce9/JTBGEzY2fNBNi9xoSHPl4bcmSgrQMzmUkmOwN
Mz1ke2JZ5k7KYqrZgsfpYyWOm6Xst0WZ617xa3oSo//zpN4pK2t7NMtMUJRQUrrc
HjMAsFDkgbU2I2Dlq3BwomiREcJzTzHnZtBZXzavslXYqqTO2yKoqFDaYOhlrjqz
WY26cWGhc8Dc1GS81GDH62pI2YATVhNpg/q9TxhrwOdrsHHuKwbWBlwuc2ZDcf9/
A8gE825Epx8wXOsfLFBrB+Nb2SNcKlGB+0W5bfMrvpBs6N+wFaPjBCdlB0ydD5hJ
6X5bASxN1Z2Io+//iO1BWLu3t1AmlFqwiQ5ZwuNSJKwZutd3l01sKr6padvlFnJc
ytqTc9TrQZx1g7ZIt5xyKjAdhtdqCvjT2DauhLDX5dtuv4HGHLxw/g4o5do7yNwB
X2m5Y6HPexkw2Ra+QXRiR4QxK3SZkgxVeAEYeVsbckiPlQg0tIx+fOqJsAGy4KvT
aXAcJ3K0fhAbbJhaSzFRUZT5jOD8JMnvR42OCWrzrhqNIbZnprbIygHFpY8I+LHZ
Cv/wT+SJ6UynO34JKMpr+afvD2NfCnjCEksX1DKU43PL1bKbk77PgGs3qoEQF0/b
FA1Of9yE0zrMIyPaFGb7fV/+QmM0pwIzrKoZWnenzciJc8HMQcIvEF4lztB8k4BM
cpBP3V6HaOMYuQf+5FZDyyOTbafBtbAuh8XwHcPfQcZa40GM6wK77Cph3m0+cVhO
nZa+xeDtw1ePhbaXHicC6EShnTwlyuhqWFsz4ck9KlFEm1mc0hrDA/kGyAKC2Yj1
UcWFTDA4aZitSuhkbX/bKbcfkdHhwo9XHIF4IsSGYmhs+YboSuNHyx9t9xfvJWFF
O0zc4oCY64jQheQerUOr7ytzxHSmkyoTfUIvkhveaxzsZqO4ChAs+HQWKPtEDhoC
wZXA/M01iCuv83EBZ1xvYxZJrzCYQLLSObVkSAPKOasaj+rasfAFXcwAgRkBX5PH
MsKVL+leaPTaYx5Fz5yBhvApnhfcsrGV5PY2KQJ/D8XUmQ7dSzeuItCAsU9qqIan
myws5Y/sAPdP54W1zpLGxWDMM9gd1HPhnLlWyHDcy7gny2ouho8zujToVM9lySqr
t/N3kVSMM8ivI4cIMETi2YbzuXKsuJTtNsTsjQ1zBV4+5TLYjxuDTHstPOmi+1M+
/s5kAQy3V6eW9g1JZkWPUTB9BHJy1ohXg5YSGb83CTfNcKaVofIg5vR6xuBh6FVK
Svy2qP9mg/MSZ3mj4lKiY7brwR5ugjOJZ9lU0S52v8XdGXKK38s+uWbLJFNisf09
3Vz4CsenNshzqDjk2np5A74q9AVy/6chR/Ddu7r03kyQLslnXBd+TbHqgHyqLF+t
7WwK/CwKYt53j9JVB3Pi58FATfOLEiHYUKcDNb2Wq/ZmEDc3woGRy7l/ETcM6rSO
DY+YxkItmXgkiS3VksY9wh4rYadeROuDb0k2Ui9h0RKlunL9Z2G2xuXJ2zxFnFtG
yBwJWx4/hEwcX5crNNRY3UKOcXE5FRlVtjElb1uJMCXtjZ5uMmz24mggGV066PM+
o6bripyZuU+xsSrFwekn1W7IfbMQcZLcBATL6sHm5vQD77CYpQBIy2KcEGuGdwBr
LiqXg9a9rES+OjeF1+miQyo/u5pLFyOU+fYAapPmLCktDko10w6gmZ4HKNFRFqsn
nVvSUF0uscCq3lgdVmE+bHkQ8TmDmTHiIUEZCoxjCGEg26CO7aYxSVB2vQJIpJgn
ut+q7qYI78PECpBwRzp+gHq5pApmeJIC8I4nOL1posZyhAmuSx66JNCrGWeP7J9X
jljd0wL+fXxt5CjwlZ5YfdoRa8/pGy3FQ+QYj+Ob5LroPh5782G6MyMfyS/pI/l/
uA2Le9JbrquGe1S3IRBcmU3Txg9dU7qiFE5GwvQyHePKFlbWApQLbux95erw4Lna
xkFp5sQRzaaZNLXTK8ijT80CikQqYdV8u35d8fIQ5z71DwysufU9aHJ2o7q06+kW
pPhQPuY6IKvVHRsKxoREH6SeuvPvy/LufTkgsAvzoR1ePzsY8czKKMEExRxMbttP
k7RdgtUR2dSkAA22zuwkcmQIg5bHuK+/GYRj0mfjYz4FuD3d2GQCop7Ta/4Is+FG
THS5ZC+w9bdJLsqxRtMp07RxbDAls4osmYS9uZvH+HYBfZ0XQl146XNoWZmy4KMl
LaMZvePMiG+SFgvwqIymikn9UFpy5ZUd4IG+S2rAsboMKFh1oLoR/wWBVLMZu55y
erMYl4xzer/X3JYTFjMTkDv7xh63MnyNv1PG6NFG9iJGlY/qgp6pd4OCea2YR1HG
RI4IT1+7oqO8c/1sRuC9Zw44v7AFTT1JYbyoIETQptIO0aW8LN4WfufPL87dG/8a
TuOxgMXB4cvKVJh+gQY1qyQ5gGLf23OfW2sMssqm3HrExLEEDDC0zrjdhUN+NFqZ
cWzAkzMLSKHSh56Y/HQreVKgBQBDCrZmOFECYynAjcb8FsEF2jmE8T2Wtd7Qb/xP
eb1xK3d6pc+M9q+e7dOfzTxJGU6rSN0ut2cK4Vxw6yk8yei1i9hI6MyseMSDWzMC
nRFodwKquFkApTAlqcsHzryKp38TNSYKpuwr3Lmv27/crEM86H86GBOLlxkP4d1m
YbQie6VZVgyvbj7BqLigjlv/uZSOmfic7Y+UrpXrj9NeJUo0o+L67CN64CS3nBIC
GhhLuLrtdwjBBcTTdjVZh2CHmBanNd9zAKYGHT2nnpBlyS5P5vL6yw8/SVZlG+HS
g1ybxH7IOguezVxL87IPPzMaKWB2te2iPdU/5JesT/HS4u3yAI86F3TGkrFSC1IU
1Rosj1gZHmniO9XXs08NpKLfCE3FwNPT2Zj8uTITY3E0zNh5HHpj6U/uBxbeoQ9L
pS04+jgA3iQdtyASqwSRIAC5wSySd8kPEW1SRfuXfAg0Jy3fdLM3vJe5HjV1mugJ
5t0AR5Edz4P3Zrsodb6eXByzeVTcYerLlsPa4VdJ4BmbHFXOcRxsctAa+GYW0o/9
WqdId1IADUsq2nMkSLcvXxGR0duI+Wy6YddqmwscAS38PvhmrFDtM1jjAzJ3va+C
kAApnmw/JTHnCxVN4qF3x8sUbuPFkJp4fUUP+58z2gcRyl+I2mlvkqDpiMHqZSyr
XlH1hkV8kaq57449TCUQ0rMCoHGEjoR/FW5AVaPcKTy6f9x7LfZGxKwU4asXSjcQ
PbPynMM8pzYqIIMxzdUHdbE6N+JKanHxWoMTqOjFqJzHGr2CBuH8fk/zFF3+BD3v
S6I1+lj8PybK3zNMmLosz1zdVH43TEgBAIB67V2yVM68ep+O3EIiqtOROTB5RCRi
su6NS8QztBetLm3toHLp98aKhq6BRNcpGMhmbiSzVkDlJo/zXfWTlisk0ZRdShsQ
c2EtfEgUy5YaeyWhObticBkU/EV1XE+tACp0H5yQ5aYD0vvk20N/Z9NgQZtdGUY0
ccqyWYaLcftEf28QgwpyaeHNsALh/x+8US6cPw35GMURt3AYMQbORE4/FQR5IpSl
Mr5RhRtqqzr9QiHW7IUADTiJ49sP8H1zldVwd3BlAgH7MitbenNYr5BUqC6KmL3x
RW8MZB0Bo/bBLHa8vJ0FHzgrtGZ1ITTM+ZTc6oeICYSf1irxyh9ffaxfhc1IKHiJ
7fa8Oe2lv3gycRGT22gE5eZU5bGSNER/oWBOn6ez+HoooAGGvYvktqHlXcNZHC4A
OKp9C97SaKyPnjyCZ+1CwplF+gF2f2CssqRsdif87CgQzQVLrRmxMTJ7ffbzLvDB
t6/JiQaQVxfLGYGkcVU81iONEM6H0sZSB/WcgIY/6MLdKuURkwMlBxuk7M7kmeaN
voLSpBsrwfZgMy/CkOWYd86NTRUeXlG2FIXoK5i3M2oKAM4JzDUQbf7+RRrCyu91
dH1fUlH4f+yz7Yzh/M3Zoyqv6y5tYt94UBS3/RL6IiVAL+468GHHt5sJ44WF08ln
VqYUjWqARX0qMo7fQcLnKbb8wPZNGbawPJzmwQhZLJyqWQPbl6yEnF6P00QrV3YT
jgyeeTgEHpJTUDyneUOK2sDkgzjQuzaywANmoP6JJqpZBrgvM50kj168NrRlqmQe
w7zC+wrSw14lY2runEMNPh5DQ5N++mpTZYg9C/vXlESudIItoQJUIan53UQJgiDD
g7klkDsso0pJLyqQZzYJO6oPxMFjzCFJCdyAE0gK9xzL+5vBMuH7I2VbQlXARIU6
4sUsUR9r+30tYG6EBZNaq+FGwCsnx75971VTCrthae68Q6Qx+tT3wyr52btK1bjt
CCvkww3D7Pyd98XryBN7HocDVUcKsu2tIZpYkNGCID5eyhKS3kIbvbFzpp2DZrd/
REhCAULgerHKxhWW1BECW4aFRC+uI4NJ8DYt4jH3LBuO8oBllaJH0i98Nl6eIAzy
K9yW0mx5dNNGj5HOT+wys7rdzIIGQNgH5GRESgHamuqB1iEn9swlVhKJSAdAsakX
re2eCuU0rSISNScaMatqmoxIn4FsKMwGel0587nTKMByVJo2w8QRNMPEYLvBdBQV
77IUfMn9sj+sPIDCp9kjrpE3PX4FgjghQS9WiH4BPRRaIDgXGTpZ0gS+9bGr0edH
YLKYohh1DkloAjPgIehnhVrxiLp7nWrtBT6zRu80rUA9StgG6eENJ5pub7c6bjiu
AoedEeDw22MRW8KTQfUWBnV23+roqAIOJ8HxS15NLQEmiCa+QCZIYCtm7gd0CTN7
SI7uJC5JGPedQi+NkLNdFLvnF8J5Ly91c8JqVhrIyog8akY9zPfGSozqZeugfXo7
gbJo6WDLcW1erdJ00LM0WiZYFJHF3HsYXqzUMR1wrN2CsFmqxjzoqG8rGqH1JDmn
kEIb6lBffOHpoHd55UIiyEYueldEDGfWp6ir10aS8iWPbwKjKGHmVuvU68jSuLQr
voQ7moTHaR6jBZqh7FOA3dZ5cpA36zrO7JlHoE2h0Iztq78hV4ijdGSkfMiYPBjm
4kMwHODvsIWLXoApHMaQOlPagEo2kZG25tmN8Sym4tqS8tLkmhnCXAerL6LgOgyO
nuTNMoz3A4LopHcxIgqKnRzrsLn6YkvSkqw1kLM0XI5QJKg2VW2jx8ZFQDUU7vDz
Xmnj64uExsM2gGq7O1JoRUOH/AoPfGsjN8wNNRg8LKtb9DcULb4P87hzBzI82+rs
dcNjVgtMYAN/zUBzZjcj/XvbXQWj7aXpCDKnE+hX5L6S/IBw5TOJZSWaGvdfqXxa
nYsP3bHi2g5DDWd7Zmkm2ASbopLCyXaDBvvSw1gkwmO4ywx6daZtrLm5nhWEH/bc
2B/6mtvDzS8t9lmG2t9WYlStTxgqulomiICcgyuHxU/qD8h5Hih44efXWapDji5S
lA9B7kuvVWlcmQadjTJIJFqkmLGhOfRyAs9x0qGb/+74gEcHSL6j+E2LdpNG6bW0
cnHKySmJRaQ/HSH6q8E/OBR8dkRSsQhm5HoBRo1+4l5PpxEMaDL5twAmsIn+eMyy
rDcO4cQf6cj8ZRsc2SKHaojyqYTfu3kC6vlTQ7BZF7Z9jQdguli1OnQvaroVDkQJ
+xa5VZKNkhp9zH8K09aPqeDE5VU6FTXOS3lzIwRQhnbW2KbvR3U/2RqmO++ga5Nw
s6LdYObqdI+o3T+MyrF685EhCCxVHmsuHrLhqvS3Es6eu3jsvYkQile9/MIxrq45
AGgFlnMGKV9ww/A1mvtpXExITKAUjE7dePs8O9ERuvmptU7FeSfI+Okz6BT1wYNY
XdSHmcpG2SB1tg+87uTO/eMpCb7ZveZGWk08+hvowGFBRGCtk1sE4bqJ1cvhh+WV
2rEu3EHUuwVKYKMMvqOy7Gfa6qOe+mw7u1uT5EyAnKtbpO93lEL2r4y+ivwErmvJ
K1WPK51ttiAizP+QXDaSuWS5J1jnYv649omNMG9pOIpLhIgsx4OFN32DlHOT/4/D
zxA/KzKBdeWISQDm/yGNP3aWOUquaKZaGZe6PKkHXZu1ga0zoki2BsSKTwMNI+u7
wvTIgU4n9x0xN2m0y4V4eX17aAPpIgVMQecGlz53nCDgGrHtrKdlzIhFZ2nlMNX3
Zdh17Mr/52QjhugkdLcY3TC3XcB9Q9HjnLc1iEyK1PDf2cwM2tbaphPVrgtOPkKl
Q64WoN6yI4dtBYkTmc68kKTFX3pFmoPVI0JmpeyBqFPcd7mp0Ybwz30eD+HeQKaO
VKKby4KV+g3EhZB5fRAhrstM3+DLABtvSP2RdlbSVSKWEex3W9bgW3G4VC94RBbB
H9bVlFi8hWVBepyJkIWkWawyDa/DZ0seOTejfwsSJB7470QlWV9L1y5hRHfbrd/3
o5U0W8FcIiFyZ7Ehb0+mWMQlSvvvG4gBt49LTziJxfFPN+PNHt4vTFAM2TfE3F81
xwwCSheIoSMco3qGD2lN/uVkXGRrmcuYaZIeQFmgnMv5LFkuHNjKq0HF21BZokEq
6sbCJoC9pJQ4PuLo9cUmMMfBrkGUWwEc73ChWdrl5boOnhQ4oCYh2RgDQfwQSm9g
ky0LyD8XNtLtTWSV4c1yBVDMIh7wqUVFWvPnragUIMYGjJoS3X/yfKctcFdTYqAA
QRVS7IaRv8eaMdUWazj+XyZddk9SvjlUxlT4YB5zYaQ2qfQSnoSinWgS0mHkrJGS
+/H7nbHH1at97YNgqpSRT8FtKKoJjWr/eJpLCk9jjLeVwhJ3CVFlVecgp5pgRj8e
+2h3CgwC/lLXxxNiVq2bW4TFe6DtGHgoKCmmgqiY7M39SUR5tZwjYMVNyQj4iodt
cqFLR72YmlRzF+qc1YJKrmjzW/AlafliHiYECgGEz4arfiDhhmfI5I88whsIEZm1
pF4mrjpF/21gkY4NMvX30yXbHA05DiJca90//fKYIwg56A8TzsToRzF1qgsYQ2z0
bRW45bCtudJ64GJc36NNZic+gIiyNhTSOvp+aAGB4/vzmsHhtnj8FTiMn7kW+g2z
8JRQGIp/L/H/bx3t8aOQuhhjT+vs9fSOIAcGNflm4Vh1zvuTZ8evAuYQ0TjNgRPY
72AlOaYb47I8D/tdkhwksTA7gf1feQNJEZV62OPdSZAumhsZPhwR+zhbrYdXMEzC
DTzS76Z4M3ZeRMvE0zdxXyFvTlnG5RPfZ7Hw4tu5olsV5Tri5yMcuNY9J8E4b7EH
3HGhjIgysKPc6P77DZWkczWjq4J6dKHVnTg9TLRGQK0/wiKclKQ/VNJFYlgw/IGA
cfuJiHr2C2jIwSOKjyoREz4CvZYwMdcnGHdGWdZtvHA151CtqXp/XqDoWFSUSnNU
OEcsCoQUCM9AN84amhQ9K2TiwlQsDdviRWtaCJ0CRt4ozNYXurEOUhwjS8UC6kFt
BixFJOsDpFaGzk/ESsxzr8yxYI1OU7+ztgLT3varFo/yC3VYTvjNknmu48oH/RW1
e+SL/fmWIo4iZ9x+TcCJqr39GF4RlTnfXcJEhfkpcP0IPV9EvhWv7mRwVOuKhfSC
964kKhI/lt1YoMpVU+acD/UxAP/oYc8EtmQjL/b4/dNiDL1cDbs6S2doHXQURubg
HdFUJI59ZlN+LCnDx3a02Al3yJkjEYtrdOgoCxebSYe/f78hCI3jVs7dopcM8mv9
Dn47ePpv+cqHjpuDDSE9IrtcewzFpQkwb6vnH//JUnOeUlQ8MIJlVmNXtY3w4QMc
e0ep/y8N5947Uup4+G+tarxizg7wxj5MSoYyRk+ChgsLvH7QWJyA9ER+KnoIsTPe
ZW8i0qtNyE1CjmQMOV0r7+0oCGG4BKU3gnFR+Jgt//xIa8WLfQCtwMdmH3TydYFQ
RxEz9Mu9LLvWSuVb6W183ywg/yC3YlnuZ9Tk4xqRYgS2wFWcDWAZa20M4xhP0LIH
P2For1YpmlfNHHwgu+utOVmHSaIHZIcR3vuX3WAepNVrKrtgC7M22jd6gMRWhM7M
SSbwd0z0Jmoku4yun2MR4J4fuLF9TdUuzqD8+H04ksgInRa18Hin7aFJjdZjs86K
ua97O5Tx8rgYRCphULE1IA85N+fqqgfYV6xM1cC9Yfys1X2k+LrmqQ6bMJ1OlGem
aOgvDdVGNyDnk97L3Bcq4eBjTWy1t36rK2wbe+C1g3V2r+lo6hu7CbiQgZnTixF8
8gjhuL5AzpnDpY4S5jMiH1BCQ7vDHTWR+arD7TXPwWiIpMi/1FBMov57f5PpQxbG
fVerS0t7b4Pwbz5rP01iC7HQgw0M31rd7uldCo/uYfpnbzm6pGwnveC+Kz2ncAZx
GYKZpYi4l+nTMAKv2AF/MTCohefdS2F+b1CD7ZrA/YRO/S8nLA9B1JCnm4GpV0aH
mqtkgN36nXSsHNQuY/DaFgC2jBDGgCGDulqsFP0J4QsiJFwQDc1qFHHJ2ZJrKO+F
PkH9juVPNWgAK3bvaPSvzWqvPbNHX1W31qZfRa5Kk+BQQYTndEGn0MHdz3iqNrbX
/Gi6BvIyz39FnVcVNsm2p3D8ZATFBo0gQDi4bNKh0hMyFkABzc7ULCx18zYjWGQV
drNX1RZdeaBreuxc3vWgwP7GtsHNhLwK8oRhSXURNOztUyOX3LE/sCbHGmvdZQ6w
djxFNNrRkP0wTNYTHK46qYrJpFL1qNsAXXL4ye2rWcTaB9z+sKft/jsRGXk5WMWX
80Q9bLx7hVyPvMaNtNX6eSgGQ02UG+ocq/AID2mYfwH5HeVTvT65a5HsIK8i1ItS
eFvunj+2UKlCdx0sRUcp9JsdYXzN1zgLxKCwET++9FAxzmJJVRrlxszy29uu0gYg
wm4Bk4+bL/8gj4VAj1i//DDLB11HTuTU+u0em+/iq63Dyl2M9X6ZEnDPQMECrdbt
DdmxM6VKlDvdzDwS3ya7xInJuCDKyivdnmhjE+c2POFZA6H73SmcJFxshnHmm6JR
6BQc/TKP5MpjuTJGSJ3sMlNEwVcOlzT7OPxjKa3oniE6LnPC8jzyfDBQI0RcFZJj
qkzHw2wXs+n5ikpFoBQzFROlebYkBP/YrtWgQaK90KS/BZhe9+XUnVetsbYde3oB
VRY1mvJGBfpno4heK4OIK33eyDJV1tdfDHXtraGoVSHXeR2abRlEE1vqxF6v3dTH
MgBm/tsLd8rIqEXYd+itR23MBLB1W+5MB9BUXwXft4VVWpeGAIrFq0Zyg8VsXej1
LfMF/sp7XdZtlW7gytb/49bRbveOB3oiddFa5c6rn0/XEG7NV80bLRqWYXbm5BuN
ynPTGrQVLIuq6C2UZtYT538gx7dJntvoksgLk0N/VJcYyo2HEX2o9cSflEojkB6W
6znFGmBvwbiJU4CaUUW+zGbaowPzKi4gmiYSpHJREbLb2xqOJEqXY3jk54Kyxhoo
13DwJePQeppvEb7T9VZAXznLpMl3ZGIIP2MoGqSKXUlN3tYiarFJMC5iDpjVBRSa
k4Bik8kbwuHca8qk/bWz9QmuiFOEgVwHLRofHHyTAg4fm44b0/+XsIST5z8jeQeT
AD2Q7MLZPf+HmH2F7UZM40JtlEvP80brrDw8z/0cwRpEHpC+BRu9ZHCmMw1wxNdT
XkXnl/IcpnppqbBsuQ9Tpu+VcKZeg0X9r5uQkM0IeEw42v+V41MZuSxXSrw1srOO
6T5uX/hexoBCjfeUBsxIZ0mYuzd+F6cRGvXg05i2YTgcX5Iq5JmyD3+vyklCyhE+
5t5Haj3lH5HT6qlIHsqUwtgNJg2y03WyjznWlMP7DSwWLxt/CYuBe7R3KQx+aP8F
htva8rtCIHSuFg60PcAw4K4H3C2uD15KRXDtsA59AgMbT63n7GlY0xoq2PusntDr
YIDnvBd7wNUThH8kCEPdcxr6q+z026OBIst4FKxvY7So7tvta7gimYF+aCnlJvGE
WSDa8oDNNsLPnYFmOIQRMRtmJqaLqo8lw0TOMtPi/UtaQLzJnZ9Y++BazMAU7BCF
LRA9Y2lOR0KWCSIY5UhOgDFov26lKA4L0njEo5nM+fPr1C4dnzWEUQMUKcj8rkAs
LFqsmkakMAKAs7RB/QoNyUpsZiwip9f4ilFfiUS9HndsNX6nV7AdyAW+f4xOgQI1
LY/BpU8jIm6bq+rDtl0NNP86lMaOfd0Bs9mEPzWL3ovLpEQbMqWq+f1m+75QqP52
XSMTlWnoDLU/Sc8dVU22d/J9Xf7qSgMB4tlCpfb02rVIEDqxMYoB/qw+w3NlbXFr
JaE3y3d+zRizfVWdoQA7WeI4ZpwLNwXefmuJ50TpAWskMBVOryyRrmhWskXz0u4Z
t/J08+xxkFbNt3+5lGKkIrhC5hGCE0nOrl4PviuVlA9dpMFC8QoZPGXEsa05QzZB
ODUNBiUOymAt4a1P8EdfYpfHCUYpTBXDQhKq/mNfWUTIfrDK5BOfyrzbj02H7S65
nq5TfvjVKkl0ALeLOiZOOXYQ7R+BJt/gqLq00/3WDMS4fI2Ge4wZko1BDtdLWtpw
aw97ECK9tYuql0/t2XUY5BFFbOOyinEU2Nu9zAIiwW3Ky7+YwW3SvxUyu0gZDcn8
iGg1T4cVC0XQaCChv+Yh5ISBtLUOIeQQMmTAuzutvmEkyRYB1XOXmiRJeV55q3oI
yz1pGmU1F46apUGgFRxVH032uEo8M/0QogG5FVJyn6iydlAuzLZycl267eHxXtQ5
nD5hkH/ocs82DeIzKD/wQhNbTPWOvAoUIEQsGIRZYH23mk8D5Uk1CTCAWImp8P7y
EY3iIim/kv2iNrl51iMIcDe7LNMhZcp7pC1YQnoZYEZ5wa9Uo52qplLVbV2FQQD0
4QNnynv8zY9/oLlqKghvVwwSGm/vE8MrroYqYOhVD0Gz0yYriuqX2rti+FbNbhcV
A5Vk/zaUMAHrU2gJk48rtQn4Ni8uBzGf8OF6kjc7doKy/EiiF4zpjUU5UwzFh+HT
0O1hujZL8A20HEjIx5fQSYfiRubjmzu2M2H/wGEYvstI0tfraAD38fAHlSiWvgQJ
2kgyjRcxbWlcKpJ3kx5tCMWZTjUWqGO2SxcIajtZ+nr0nYmmuaYmjjIZmCnvHq/G
EO98E4QXQEkUOQNarRHQKwTvLMqlE1qaqBha0ZuCHq8NMQXTT4ugaJQTk4/MMWSt
OMlU/K4yRyN0zA86A6OhLOwrbc5uvYLjByv300em+aVDrs4UASp4PSAztuTdDrQh
RdnAdrtfYAGuE5ab5HS+dubVueJfJLFxFFrK7XOzSWYBUVEDRoAwyfy4xPaPo7R/
9K4caNhRAf51vhgHkQsPtGImzcOZ+2yo2H57Z3NSWGb0KHlUzSrfNYUQxXWgwFkD
HcwbtbXU9ZLup6UtOgC0BgYLAlf7+cQxEfYoP0kwKBncn1gITXny2mcwjCcXOQOa
axIwJNMZp0pH6XPe01LGKNH9wAwLgV16cuUAayV7n7uCo+2zFUTy3nT9hDuRMs9k
s6XIdYAZN8k1ViZXxyd7rwa3arqMYtDorRrDBRHp/172tcNCZ6D7cLrLfG5KdwbR
p8S6Ew89cr1GoSHCJC+kBeU73a+VxCUz+wO+Pgq4yNWh+rq58TEj89uYhtEkC0dU
8pobNaCaDOQ4VVHuTYWE4q2Zf25jABcNcZ2PG7Lcn0s4dottE5VJ3GT1TyIax0YZ
lFkJrl3tq5KevlvYhD7Rzy3ejeXPRPcTdrXsgG6/EEd+4EYNDZwjcV+ifUuVMoBS
EIyf5jbGSYwG2bFD3PSWtTFmMucJyM8HRAulbLtqOlELnXH/F4QEjdbaPxuzs5aV
FGYG/4NSvAupiGN/xgx61a/+zu93BZP7HBdp+P7UqLNukRmPL9B0dKfKNQd0vhuE
TU1tanxWAWyWQhQtYeR8RwVPg8l/mylsp3UJj/5jAGKU5iv6H58mjrpG3TZ1++8u
/9+TdfxWais67g3s6yE0E7t2LZrONt1wBekCKhOjWOAX+6lslvr4s+Fxt/lvqhFA
qo84WQCWB70HChRR3u0wT13K07xtIkjLyhj+QQe3Yau60VGF5WvDsqqeLKoaQb4m
5N11asBRyVlTQpT1HYVTeSkBXPKwErpJ+ufKYi/u1WeDc5zc5k0nLUgO7WwYHmcu
Jiwcl6YL6jtG6FJtmj3k6GU7xPjsTJCNh/8HwYcI40lNaxSsDHQgDCMyNQKS/kRS
/8Sy+2StZd965BrwgkWsv9hbCWiDI4trImMYbW4nhkja/bvre+oBLtSgjs87aoOU
HLjngkAlILMl0gt0KbPmOxERtz9+F0LWZ22m40EljzTt6zLr0dWlw8bo1/qQpDdu
g+4IkNLjjMccELxWUc5WVpNJUh/D8NNt/HNfbZnTeYv80ivZG8d2BrmcDEN9ylp1
ss3Vb47WLlU90MrAWaMm6OHRGgT+YyI15Yb8ieygIAnZlEObMaHcEzCPpPN0lmPQ
Idj59cZLQbPmnS1E6fG1UseYWHOj4gSYZP2Zb7q9H7CTcDh6Vo9q+xVYx/5cYyNh
aEwJpZd4VD1NnChQB+vJhOkzzJl6OYoXnSRCYVwo4rTM+cHaMaPBmzKYovAzw7JJ
2gDfcmm2nhn2WuIXgnk/s9aQoitcxIv1uyB0c6NPasb9UJGrIWpockTglYE1q1Tk
9Hr64k/TltMHqb04AMlvxT0NtVvOMXpamPRXajAdc4asou9Pmm16/DU4zN2ncjl3
qNbsOnQK9xww+tr8an9+YxWd+u9z8qK43QNQXk6Tho0z0VdhXdkyToGEqwD0+E+8
w3OYgPQ1vVGGxzWnwjvQkmD4mwnkOyYJfZyVJQRBvVMKd/wkE/OwGAXS27ACzSnX
7QRN4BPxFII8wPfao/pfNGvMqOpusrInGNUb0zXAxGK+/ioSjccA+2NWtDE3q/G2
3OGTDNDZ6NIaeFk4IQOCNs8LPYP2A4phwU3j1t2ejbjg7c7DsQBDfFJ3p6UnSWdY
Dp0qVf1lhvRlQUC9R8ZFJAHc4N0K9Jqw4OVPNqea+SDmVJqVy/MOxRidQ8BKwE/1
uyL2sc1HACtMVhyPNqlDxPXqM5izllgShZIe2SjmwUB5NI49nWdCGsBLahXW1c53
/mUcVnh+IcmAolsszdKoQaLiQKFoX21KluNYNkU+BhtE+cwEziK4HtZVF277O78p
6xHN7GIwJy7kc2XsQvcwWk1sXFpd5G+BLlbd992iJMsCaH98bLmXRutOElN0iudn
RGXatPYfJFP3EUeZ/vdKIovsuOm7wQtOFCMPA+z7Wd9ShEAqPc94IbD2VrUNKKq3
POg+aV2X+N5WG4C4la8gNunzvcBtq7qIKDI54RuJ4OqlL8gp37Fo9qGBRp11Q0JR
2BI5xBxzyP+ObueLFJmCG3VniKr+4iwCse7CgcGiAn8n1NpFO5kL5oHAzBUdJV5p
TLHk07O4Qu/W4OYjTCkcqakWNXCJSZbKrWfUS2BbxsE8GOdaeQ6K2Kdjq/roL6U0
g04ZgYQAlPLDSLTApiL8os2pm4wFPTA1CG5C2m6tKQZy4EE6Te3FD0UpIx9Reo3i
Vgl7zPspc1BIwEHGR5j53j8App8gcYGaZRlwtAgwxgtU3QlHmshw4gpxJ8gHGMmF
1SXtnnybVK62A8PmTjqMvyRGDweHluxN8A7jTTyNtzwdsUIsv8mGecIo3YnfL1AO
eTBDvRg4sAoJ3ojEP9iecwJljiv57MFhwOdvVJqBR+tXr3E+/FB6IoeQ7PdBR+UX
0FEML7r5MCcZl/27demkNx7OxDTTpPRq9tOOsBOIr1qynucxKuRchFHfryYn+yoP
gFdyY/E4BUceKKJ5fn6PNEBkSc/Xjp0IzxYnemQoPi/Wh6bdi1tgJI5/p9GWISRY
kNn/Cbl9GWD/7rxStvKE9S942y5cdKrnnZ7/KCq7DPQnTC+zR5YJ9bIB24t+Jw2c
uaEyRZAhzgoStfEagZUXX69Hha98wpLAPW9Gj0e6ThMaJGM8KOtJ1pvLZ5+NKrhD
DMiN+3w0jPwti5BWALF+kChYTTHVrNpWjg/uIjUrN2IiWUvtvSjSfSJG/oltYdHI
0pNZubusnly/uRUWnnvyRekmaLRkVI4hJU0Tmdv0fun0ZcN7nohWWEvnBb3O+B60
kpjBdx2YTX2ZlPF7dX4FjlqWSmeARK14uea+MQLfM3PLO72C3CZY4+uh4TnoQXBG
JUJSdaA4NDw5NCKIEr7OThpn+/IaUaSs1j4/LN/Ut9n7/zNeRqGzeOwfjDy3O9rd
rp2JXE8ZJzXqi+MSgMkOGy3YBMzqn2fHsrI2wF8NycxpJeozEebj5VA61kB65zkt
Zvu9VGG/KTjWnoKKm8dzfF4pehyQNuuNBOAIqRtRJu+P39mz3npQ79Yf2A3aNY2a
kn6G28BmE0Bw7QrETrPTs5ZmZOnj35tST43JPzRoEOm0haE/4LSwzF5IvmLchNFV
YHQXacENgDq6SmzYoqdjDt6KDdfs/mULf4eUwhOq6eqOQqFw5FmUPM4JeHX0oAqK
sJ69xdOSvySOqZimmn7ciivSFieGfBrxjfpVVMzFz/VlOZmQ4U9JVHNEPlGh5Tj+
XzHstvOR0tECZnoYbMnVx7oJBTAwMOverQDMXgKIsgynzUqK0StwsuZcV2ViceZU
h77vT6DTuVFUQN6XkuXkXS/plRtPh8AO/eW3PWiQ3Y5PR5D8+BKngunHGEabricd
cuswKIt3i68IsHZfK+xLIjr1qk8maHqJRST/hucduWvop9MRMUCPhEmUMJdpWY13
7Ga8w7qwVT8UpIYbHgg4JIper/PQ0hSDfpm4zmKykV7d7euaQLhFW7ywxhPv9OQX
xBpFjTYgZLNNnXQv0JVN6XgNPYdv7pbe/U5f3O1NQWAowXzAyVxUHFBPo8cxnsYd
6axVeJKqE763hnzJb/ssMkBoYaLnaxOM4ouwT5WWStToXdu4JR04eNbEqN4Vynls
BWT8Cw9TmgInZp6RKjKctYD44Io4fC7zP4qH3NQ7b0S5qAXIDllzy1pYlSDpJeiC
vVZVZ22/3kTyRIDIwKkgVzakYGBWV8+Zu23q8mpOUVXYPD2dTKVV/YAhZWl7VazB
yShSS2CopIqA4MMDvu1X8131fWxrQW7aWxQ1zDsPSMOCjFkZwGX5s+vEdGkPCkJW
aKvmQWk7itnTWS1HaKplH25iA8keqXnxCpBrytwLX1EG+TVdyems4NPG0M+XDej7
FqPm/lTHwubb5QkqgOWTZIV0zKEEDUh/+OVDOgCQOeYDDs5wYLgKuCrA2dT2gR26
dBteY4Fu+QNzNQ02JQFfeud8004p74JPgVpZxB2dIjmip4qUKK7A0gA4hHQSj4B7
hOwbIyBJDXXfg9umzYQPvgL718zOO515jDD8nJ8DJ23jnq8xhUws56g0mwQw/v2k
73d5Zw1NeTT8WdgMnExgz6C5R2Yxt/h+H55Bh68f2BdzZjREU3j8J2WAKDFWfjGD
ZOMH2LjVirDnWePyH2oX+YQ5gC+f9Pf0ZmRkUJZQYma0WVEf+f0JJYHCMz22wedX
AgsNeFSCjfXK0Xa4vG8OV+QaaSHM/13Z9zs5YRDF5sJ2aBVUrZiacDnxjbUgng1n
O5joMlKGsZGEyci1pU+eV+I/OPW3Xh2ErIFtuXJgG1wJOG7X5hyW1FEFCMCP8SiZ
tH8XgrZaVhfiUcWyAyh6tv2qp+oH5gL8nxCEuUxFsVhZp1QzRK0RBSF7i81+o0g0
R09/818/3/d/GAtVPSh9e/yMxpigTjNPaTMJVpeRZ7FeyjPFE8QzXLl8RK/kQRo3
8k0h6IJ73Mq41tex9o80WtwuH5jmGoKCKfv9CC2zN5KUwGQRuRRT2LH7j99y1kfG
Jsk9dAp5wPjofAiGSHoe/1KWLCKMYQ8B7+5dmcm26pLVDs4AoTVqNHUqTuMA3dIJ
MPxFxBwZMA8FSacrfYHzUGdkTUcJSSBigGfBXTG4KHdy1nLXqmYKdVC5ykr1VBl4
Zcnxk6tRIrzRZYpzpFY4Km7oQG8tmLBycqls9XFXcPat4XmmyAvTbmQSq77OYpqY
yrqRJZ8Bg3cyNkNbQ5iVKjbqReVYxprHYj0I0llVQ3W3qXUg/0sJ6wMyJaLGS03R
oJkR6iE9L8Lo3OHPY44L4feDzNiCznzyAV6JsCTxO8F+gBnEehjeet9ZMkst10JL
sHSssfKUdNbakNP9VLkXmqgNyciCTAB2kGBnUP7zy022BXH+gQdPxTO9aYfm+WFF
439rjQztBd1FVKOh7QWlr7rFMHcvHpm2XPnRKSJHOehFnXkg86iX2yTDYFzLW1Uq
FV9w1BjoZ11kLOOdehVvxXTLGS7p2yzyylGYBJvh5QC8/Cv1mkO+m4ztZFIFFm27
6dKFSu81K7GoiWAjQ0wDmoFaOahUh21fzq1m5yzBYpU0hlV7AqM2eUEJ26JmnWTp
+azTspXtuswVSDc/cX9jB84IxwgjUOUXA2pd6jafiOeMMmzkF5KiIZ6aCsrzEOK0
rPWtyXFOxFAcjr9QBXBew6gsox/3P7E2D+hm6dSFkiGqZHi1WQ4WsPZGWW01z6wT
mFIFQy/6L6+mJgFdopYX/OJ13codMz3Z1qD1q+wsT/c7442mBpMtK/8y8u6KzNMO
CXVs4ctLABqj1OB2nFGTenlwwFHpOclXGN6L+L5h+WYbC+NcYTJi35e735VjDFag
7eymo1a/4cRj2jhxEn1vp5CCQcjW+pj5ymr6UzZMYoZRAS/R3oXjQjcNCUzEc3gD
aK3e95EjIkq1LuOEO9FqaQPfI898vW4HZOywIUk2MGW1S2nZFBZSqLj38O4+Hr4Y
pTcKm6bA0+58wTccnjzD6Wu1dM9MWJc/o4cEZzWmluCX7jYTuPN3KGb9eqmU7Mry
nzdKVJDGPPzAksGj0SfvJOiO2cfK7ySKgNdnRV7yWSIIFeMIosuvG0erBASIhIF+
kjn8Jj6nPIxJmgil8dozrF/fTk2hUweTxbXFcNgHhEAuzxjBKEC/w/cmagoUsM2E
sjGeyHFPCYF2GnzQcf5MgEpGSvxkj9M74y+Yx+Vjpi7VSPAEhqEgTEtQZ6vSBMI4
DBGTvbghyzhOHMy9vxhbu4ctot7IGErP0KgVX8ikaL3RbYqZlg/++iiNNKZ6tOJb
qPXulnPyBZhRhJlnnw8ky7J/tHB84V8ib4bLl3eM2PDV31l9luAwO6TMY9I/2Xns
p5JyB20qWhvSqi94CYECWqfII46JDLKWXEG9Evd7bMdofon6ESgQvakWLvU1v9kp
4rq9B08ybnYTG1nzBqADF/GgqXab5hz6dN2SaskamTOKW8Geur5w7qmf8noN2aXf
gRzbKF5gXlaFNkMFsWR6JzpHKPFvajymSCuBp1/zkCdgybJE8M9wyHEieS+gvBYb
wXh+3Iy2pli0XDw59BESlkQbYUG38/KfJWpIfdhWx7A68Dvc5Kkn3t1wO1pdGTo8
Mxubab3LqPWtoPxEh9jR3nun4HtT8fRxCNnxPllladCv3aMjU/sku6aquN0PcDY5
YMvDEqeGo5V3+4l6vb6PVo7PCc+1vufAw/XgEHafteveJRAwB/7FOpnYfs74KN81
hS5cYcnsQXsTfwo3bSg63LBuh7iON9x5EKIzANq3le8RP0vM4FCJ+3Anexn2sEAA
rB3gFxptgAbsG2+Sa6NRlIzbNjDqhALKJZoThYYBumyM5805ZjeUoQbkgUMP4lPe
fAHvhYkuXSsjCjeN+7Hd7Tx+NMpVidumbh2X0ng5lT7n2ONbpNHAUkmDv6D4f/LE
Yc980PHLedcqKBBJMjxeTqyBfdNBXmyj6sJhCzTNM9jV22swNkzWhdpf9VnTs12G
Aj4P7/sFldVJBftFC4NWKYS71TC6XOv65AfEjHRnmC+xYRnL1mNil8zVpmqBfLaX
CtgxbPuziPme17YBy15q7IyLF9XBGYnseznGAJshei1OeDrRofutPK+iA4FaEo+f
Gdtjd76FjUMfynRpyIpwR6QFM0+uSZESqhxIxXWzzmXx3p8MlU8ncH/4N5nCeC5G
Y4udb/RRF3//45NbI0idnbr3VqB+sSo77rEbrIuKFgwyChaGQnvglSlqPo1K8zD/
Sr0lhj42zdjce7cl+5DNcJAmZE5xJHbyJDyGuBE1uUa1ujUtAdc0Iwk905KTlFs5
YYAJSTXVQ3EZm1AcwJFou1g8vm4RA7UNzRA/yGiNtmrmTmEjc+/T0eJREd2oQC3x
/lWs1YNzsgyW7FqpVX541B5LDnhPjMu8sASnlJCyWttbfOT5PZURDEjGLrPkrqtS
/492eLe8SL66cGXvSoEhjylQSRncV8LSHsQxuRqdEkg=
`protect end_protected
