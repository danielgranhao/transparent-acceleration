-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
L+f/T3zqCrSHWamoifBE1ZtN5SKZtdrKXjnsY8LtmjoYwdBSxFxpd0fnOlvl6NH9urc7NWk1SmeL
dgeD3vV7Tllcp72yj/gqMx1n8ic52pxZaS0DyWH0qRoFSwUh+P7HhntocwDCZK259uV+5H2UzV94
C/IOhnjCxM3pJprAOmnDYQxC/K8xkCfG9HYCgDJuSkO77xco0rFpaqwDR+1a9mSfrJ/3DxWz7rdE
hgEftt6CjsE7Eb+Fr5iyfRhPn/xRHq3PnKFcVpSbHn4b42diappoZFUap1QE2CWY1YpFQ5mqzJ5b
j+gvHje7rNy/1BfACRtTQDqior88LP2rBgDWxA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 49792)
`protect data_block
cX9ADhzcQtwhO8mVGMOPFF2ioVw1+KQ2xKJDv32rggV1E8gm3QDWvSVvEFpX2+6GVC5FGIlWfFNm
PpkVLa9QPXrqkMmKXAX5scZVUBetrQ66Ikw7TgI0ciYDywOhUVkanN7nXqKJP9RfIvV2T6GfdILx
3FPLRWwW1FTfHZUGUZI2Zu/F3k52+/neOQ6EeTEx0EZrP/0R+DanVXB6gyORKIqGeV74dDbyX5GM
iiBM1m4MhZHDX46s3bWZkmfb6jWw2jaIKXuwXoABz0pDHdVIwKO7a4m7/0+NgfQfEfm2qg+kpNwF
LMbCW0fZmbor/xw7H7HVHtkFpxvDHkd9YHS/m59A0HVYoce/EI+Mv9Ucq7RncDqhDIlhD2kWI9jh
su4EnA6D0hAlLgk2YTbpyd8aPivDMkgoIJ8xksTr9oBKFxBG1BDw1k93wdazExwimZi1e479W6gC
Ox5ToCKBOQygfkoPFsFazJzmyQdTQlM77RzW1oHZPN3JLyzxQJisUeKm/TpCzP/T3fhzJFytsg2B
Bpx86iYuet3KmavYsrdyOsOCNfJXCZ7/Qpi7w04367io1TITHsVJMNXWfd6c/DnaBNl+bdYisDBz
fZSTAh5pbiwnjmlyH83mfsOU9j7pe8JA3+0My/HHZcFWBqhTvYGuLRP29nK/JcZZ/4TXX7GidZMR
Mk8KkJkn4buqM9wbTV/gshfNQr1ofgB8PBa8Ublwg5obddQkK91lxPXFk9rACvUWRXavY8JKtHD/
oC4Q+9kgdM6WYvMtwD4yixlGVZa4OIQOaK2djZvRLa5bQIAZRRwCX1aGRfw3fa/+VV+oX4cCfFNe
D5rKw2Cg6xt7SuSBKaC8LWypKdZEMlcVOGk8hoCYnXpGGh+9YmPZGfPqC6BWTi9SbMgYOst1sbbV
JrU4R+9P6DOn8S7qTB6nNw4kwPg6OZ0Sy/21MINZ6TFVcNVvpc0qbsBrd1Q7HhPlFlOCs0upguOt
cy0TocmpHtg75Co7gm/lZzQCGOTUD/jDLIvNVUzN6jlVcKpK5wpcuLEUVz2EJ1Ls0pjQGH9wyFzg
Ps0JycWzGcHg/wADPszKCFEZ10NbXVYtyjDwtYMFcJT8T9h92QPwQJzTVwwAn4wsFR+hgJih5/bc
gMd6EzfvfP2F3fY/BtgI0U0/BRwz3msNNAnBGbcdkzmIJrc1UhkZ6y9uBQPoKN++f0fv27qsLaQu
/9bqMnyqd+akSGz1Uj1kXzzR9RCaPaujaIpJBSE3Kzo590JlYbfBAht8pdNe8aXooZvjjnBBLwKW
j2d7uSKaXrmFZ4o+kE6ROHaFYzfa9mW49j0ke7VPbVHPNVod+IhrrzE7Dp9N4s6sn7KOPpRrYCKX
3Gl2kpy3jZUtJct2ZFqzCnvybLcdo+phNUjeeDWdZRXg7calmH367/ibnW/+yRePW4+gBHVJH25q
5pQ8C2x9pX73tTDvPEdMZWBFM5I9+3vwq04d3ECjoxiZ8FtCvRxrjmVHFCJrOQkMBETnvxfa2GdT
fIEx7QmLw3vk6ttOSJZZHP+5nN41Dq2KpInMkQBMADgAMv939y9oj34YwBy8TuIhRuMhPXLubW1L
L+GtHtU12pKt9nqj5aou2Z8KwftIcz9FGxz2onDKzdsjTw/Wu37u7WdqfyTL5ZdhhIrOVWovyDpP
PUI5O7iDCN7WHkC2o16JjI7y03kIbfGs5wQ8T7Nt1GLvGyy6FXG9LukKzhjyB4hD03Zh8yk3QdM/
z8zyb98uelpdVIc+kL0/EoMNvigjuvd43JXCD0SGdAgF3ZZjXn1cC9xcBB6OxUR54a5Km8Dc0xwL
jtU6aY8PeEfbcXNo/fVmThEvzDa+kEI7ldJIFZ/bI2qbQRJYk4nYJB7XyNBlcOEGDDaKmmO5hm7t
VKp56eZ7J9DAVgR1LkdiqQPIfz2YJguShlNKP0brH+IftqbAcee5ETnblpFgNcrZ5mn0RPgpLNpJ
EJR8YS7cZzGXZMKHRMGRTtkSPMq30ktyKoL92bkT6aJryoSQMhCPKzOyO4GX6IKl0ufqchrC+ztX
QGdL2Jt8PpRtyU0ZbMe+wgJTTplE/e7mIqtsZC1I1kqaN06TYXTI89mIqfzANU7oFSLdCf54pnJa
FXYeEuZPc9qSXYGEn+pkHH/U1Fsh+jzraUZDRxPsN9D3fWifg7PlNugrfQAyih+jMalf/1rW2vRm
d7ZmLLbs0wOi8JL0CCrx+frh4wIUearjBUUWx2WW+uWXwc4xqSzZxUtKxObPeRuKgy54dyAHvBVU
UUis6aF4KELuC1MM3Nh7o/Q6N/uybTlSP6LywGqiqpvRNUlVBkgcfAwUyUBM8MQjvtTd9fpLR9Q1
Yt/9Mo1eTHkr05P6gF62BT3OKNS+2XkEGeL5GFGR9E3G6axSWPvVB+T1j4B++lQ4WNbjXLoMc9iD
5VdWmUvqjd/xyZsmMVFptz/Gr6lKOxTq/kqxkL0UGpTCTf621hWErGl2cf9Hl9je7HQ3HaUQrUh4
04Eyt3Ir3TxOY8OrB2qFYal/R4Fx1JkuaXaqtLTN/yLOX5spnSM48Z5hDCu/812G+dyALcRSgx0s
fMHngFu9jWAeLtbX7jOGt2+IVT2s6jXOnuP10uro9oa1ZQkYy9wEGmDpURYI3IyO4rGVJB2T0Mts
LSHHTRRQil4vLMYL/rengb574eZstQ+epZaDkqxGbM+FZjNiA+1OsBeMnEe1iAVGw49Zlth29Ua1
tt8OkGhEL7OGbrIlt+X4LIHCy6zn1CsSMvWdI9M6wExUO5F7GfjgtrAkkVK/udwxxhQ6Qc88FuA3
/kdfcC6XUPzTHVIJcL3H2hCu4vg1EPHzYKo37TZpC5Pkfml38RJqbhlJtAmzNNxTHV/PvvSe9Hyp
Fu9zKPtkk3vYrLFF5nfeXrmp4Wglzc2bBx03ZrlXKs9Djc2OkHYrXz3awWGqs2OyvllPOhVLwM2A
9FQIQtEUkee46G0BThyniJrXWNFqP8T3sgqJzIDCnKpc0v7uPpgg8IjcqcFa/cwQCEBfGmxy0UBx
ZwTOzRQMB7jEm+mfdFxl3F0+XUfmvkAPCtW0+MWfn/M9XFzFl4MRPJgDRNW+evTLOVui7AgQN/ay
YpwmuSCGNZm1X/IznXqFwRyXCqQ4wjd/3v6aTqN6WrN8qen7SBKwMNdOp752xi5goCg2oeQFU4Tf
3NjXjQ+W//na1dY5gODnKie9NEtb1tvtMkYSDYzTsd49NzJ9kHVwT06vtCwGBYY6SakJP/HWQqVG
ElC9A4/hlE0UdLMOXIk/lQ7pWLxJPiUEwqrzonXuq0Ie7LTpN/mCKhVrj0v4YXUJNSdFtFsqGYXE
2fL5K3zSV6vnHm96pMcl7DFuqVen8M27TEJi7aLouJ/JzlD4p+S4Q41nYi3aEuPlsvCl89XXNvMk
9xAa0NbtMRBpA2FxBSW7lFhk3IZXAPZNagrmGSnZbl7cUIL4eFlOb9nuCYPGnqPuLpxHfmGZwdpF
FrBKZEyOqvqqNJKSlZ0pg9ilWTMYFPiJrYsLRF/YVaQvQUEicCUnGxuRt7WegN085yimp2zcgPKd
VnMM8lLAoaQymrgvfH894o0+CNZ1Eq7e5+OeJIunwFDBi5l7uUzSA4XNV9Cy4WYaq80T7Pb3Ymg5
Pm0T5KZciXtKh+evRlv2izo4SpiIc3sw4JUwpFJlyoYnoQNAHKnrTVA6RZCgrIV8KRbOeTyZfk/R
H77oVWRa3d39q8b851gHex/iC7qNuj1VSMal27QI+YRIOIItuQtsiE2jM3YATvID+V2qr4n6mtcA
f7qoBOpGwv79le7Lf9pvNoochu0+r+hNwDCNThhiQbCAdClGShPGNb0S4sMoBbPa7rgfc9Hz88uN
tNgntRN+MGAddiBAmv6I8W/33RiMEInkBZUW3kE9pJlv/u4TPF02JVcBK5luirMcAkBRn6OFc9MD
hPU+m8Z7ovcsRbrbpUNxMft/VJ9MkIOGH2uBCzfkpC6dzldor1cpXcgiRPRsx3jQPa19RUAWdkKp
qaqo51d5LVLTSFLHPkBQ7PCzAznt57zNnzwkXIDen2Z0GjIZZVfNt43soSScOobCzLw2/ut67nU4
yHCrT8scdy88a7eFjUd/HXrdRJiUc9mu6aeodlkRq+LfuGC+VmXCurr0I1y0XO8GGrz81XdrgZ6B
6n2Eys1Bg66WDQ2krb3f3QSIudjoMiw4HM6U8gYv86IBIUDdsbOtkgwfrG718x2MybXvw+GReqnz
rQZV41mYSugym8hYhF5Lo4cZvOWJcAcqKrLRE2IXzKzHhNnR47+9IWL7me/otUX98vbbbdJQeyhL
cBoVNe/zDZEZ9Gi0bqCxiES0B98zGJF1/6nUCzsQ5mVYPNPrHSTL1kYvEg0l43zNZ4KrmJWxSgqH
xnUijy4NcUD8AH2LGP7CBKeyX3k2JRlB9e1/SfELe5uJIGMkoUzXdQ85L8PfbUHZInE0iDpRq3Np
8ZCvt3gjHrzJBuZ/RBY9bMyWEKX/Rdy5kBCHWbE/rClS6OkUoiWz9fJ7A3Akh4YhW5CpuhsSGP42
IUG112PkwtMZTcMIMUXbIbaA861i3P7LizhTpOdKWBXamKuHqELN7q2yMukBu1A6GhIfx6lNH2ty
3bRTNaiA/3MOKSUtmAUaaESUPAUHkbCs+nxkRxPN4lC4j+xF7fwhQL5lDoXQZj6lEizzANBWC9B0
2TzFqXEQeCDKYuGfNDDFZziRmQV2BXyBmrm3V68JYY4Z6W/jo9spU8cJX1NadFUo1dqG1hSwNwl3
2spXGOtiHY4uBkPMN5JR81hYRnrYbnXyTY7TccEGCXunkWy2pFZiOt5qv3MkqLK1hsd1FKHu7P8c
FHOke45Gxuvzx+YsmwsJn/AZLS6ReUhuRUxbC+2CzN4peDzSWyCA/PMQwqz9oi1K+A70SW7DdaIX
4NK2x5/XwYQmuUNT0LF9TB6iikRFv40QVuKzjoTsQPdCH+jPYnnk35hkR2fBPtPHtWSowtARHRl1
T69UWNqPVaSwLgV0EL8di6tNXS8tlNzqTwKWp1RRh4McxmiYNuHtK0AWYZUdxSMTVcPbjF/Bfqfa
FCGlbJGMQiSmVfNKkjj495w43EhgSD7ifNkPA6BqIqzA91ISQIs8Vp5li6lrbQRVwgfwQ+kHgIbM
u36IA0qVKxhWe4CPY2TJIs/ZP11jrIvIWVmNZiF0koSzTAw3BoYUCY7LVgj9z3wlha1QVE2YwTGE
A0qORYnog511OrUeP8/O3MMzgweXgYZy8FU6rP+0ltKhQQXkSOJfOdffzRh+s3yLYk0sAk+7p+xZ
vClIXJB+NGtct9M6pyX1HJFQ59jy3Wwsyr07aYCL0oFgy6lGhWkq3txiPArBxE3cYXXp9MAhmQuP
ibrB10QXpaOCIjNUmACBnhArOZ1ZGKXP2dgDyCK1jsZBT50pUSotzgAlX9tEfAlOo4SGCjxUC030
THsJkEelFhbfp4+isPXWz4r7DBvgnExp+u4rLfvKSfCnQlJBVGOF7qm1kuAN/W8+4iJlLq4A9ytG
3EfYn7tfT4oWVkiCqfQtRBW5dgezecoZzgeOJg4eB46aN7XCAQUctlKyGjtYUqRdBC4qRBPS+p8+
3U5siNDZtwM9H2C5uL2n+krZ6pmanQzkX4rLq1tDB/W3SNzoM5GiUb4AUKP31aXYYG0QJfFbKNXa
9BQNQvByLrhg//MUC5CMWDA0K14OEvXrozxzu8fPXpJsolyfyiMWU5Y47Nnr4fRq+s0AKpWqWI6P
knCmRs6seJRd+Ruk4DsDLCVslrWDusd05TutOCB+nPRrrVW5ILksMuNC6lfXqvHeE9HRJSqvgmu5
TFYYB3kkrNFrGGIKROrJeDBdgF1iBRDuZqn+XATpBBNJLW4F+c6TsvWiKEdGLcaDYq17mhajAAdR
nBIt65FdnKquVi3ypGkwT6H5jmyevNUzM+tesNNSAVS6i/rwFgzVRzxN8XljOViohX6U/T8EWE0e
rlkd5GZjhGLxO66fcAswA+wayRnpoI9hIXQxupIY2qQLC0vdi+RoSto5Q5Rk0uo1pvGqG1MLFTu9
XwFgLQpKotBGtV3U6dTIvIuJJ4CEpZx4VGdPBcixJYXurNZjgc3FIn2JelsUJZeVMIFdZQ8K9xto
b6nHGn6KfJHnscMRfVdCittrCvRFcWFqXhTnnMclm5jt+UzPzysx873aV0YRLyjXOJ1vmo+JesPC
/YyVwb01UojevNb2ThfauvsP3Z6vADvEhc5arn5Jr3MPSBXn+iDBhIzvl5j6o0ojpCv5GGK4luQo
s4M6sDr2SbzXMOsYAGcMxYealn5fjEK+L4yg/YXLJKHi5vFzXHmbKHmXMqED6+VHpLgMJl+uHh9j
oCQmvog6jIivtY/bnljxkeeWdBzbzMAOmGbrqeLdWIGAvlzU2IUVbGJnYjjLcZPf0OqGnvCCcJM3
R2mCShCdYJgBII7vBupvsaE5+jt1tZpMpGdWuGK5eo+B2Ur0dr3PsiarZTbdK9gIUkT1NUuWp6zQ
iwpKMeDN1R+JanUfnhyDTj0+8AGEClWqw8yPR3eEH08cNLI9LR9ms/fCGgjdfgBXKfRwbRLwXulN
C24v5dBK7jPa7nW0pwp3aVgmplIX8O8Bq78VpLmry1Z8qABz1dZ+2vsNgYbW/+BWGO3ADbGjzT/k
Cpfrpjl/KMPuetqI7mWEJ/aG9RCQwIItE4cOQiAeO5AUwGMuFx9KoTcix5VTQ0VT7qVFZYRoSwqG
5t/xGbzLR37ZgtMc2HFUw7kB8aRQrnkdiajiVDQ4iM9W9f9iFvSE3XuhnyXp1ZdrM8BPcdg3Ahru
FeP2DuDW2gL2qSwQA08CJI+i/nasF2h3d/wJG2TxITohFOz36ydrUcmLAKmbID8VTThcnK15Rrxx
qbGzCltxHK498lcRqARGmr5bJT0ef+FSi9XECXN1UoHUq/zlSUqb9mSZdmHCr0IgrW6SJ2TjSG7J
fdL3qU/zusEmp+9YtZg6K37xhtTRy1KYqpKbkf21pq57S8F7j+Mk/GSKJt7c+sd8Arx7tvc/fRfV
Eg2xhyMTZjQ3HlG3UOlNcmHluoGOv4VYkpiDT1ZTTC0LqHd54TXf7ssqk43PpPIYJeBseldWwwkP
cPTG780ora5A5YKZsZRlsW3EaICTwH0sE29py94F5N3+d4aKkWjXWuhECpSjBSQ9BxvRoRydOse0
0e2p6IAfXB1nGhf3ZUss00qmenHOIrL4ZQrwBrabAeFL3zMSUE43FAa6vXrMdUy7FX/BR5VZxXy7
H2o7yTprBwp3HOtU/OaNGoy7Nq09tLoSt7vAz9sJwM5AlWEjreU2CLqXZ31jSma4xI6M9m+tfM5q
0Q8Z5czECeOhnVsSK670oz6eyJ2cZs61MxlK6Md5zl0Vd8/Pf9DkK+dZt1VOiTFLWCjbO/tWVJyn
BtCwuPxdDrWA50lmHNzV75NHMiABM+agbosIRJxTcTrVEbHQzD/JJo1A9ruWfQqR6UBrrnY78YJ8
CpyVWOT/Ja/NxQfp83TiX40l1Yn/LfYL4LzG/6P49g7XYIHvi3iozx1p7LtJTp8wV7AadWqDqfEC
1InZuGge47Nj28tc4NnL+xHNbiurxv6k9ha3u3MWFO0DmLd7czz19+rsJ6cZAdg2JuyunDHP3yvs
vsu73vnV96bIzlSXFaoI/rWb+beZydW16CLhP3E6e7Wx638F2NIZ7E1ij+Wpp9PgeUoy9AdqpCUw
/woxUaT72B4j32MEw/Or7ytQtTQHZv2VrAe71zH9ddwdpKRq/usQBYqIhUW35HxDQnQztIq4zqaN
hvDBCaoQ0iqAMx31vyJUwcLJG4pHl6E1cs5Af1J3THF+HklR62mzkQHirJhIRskBz3nwkTR+Qivb
bZns8HkYsbFfw9RvyCzNydFYuPnuiBSKIsjoZ3apE44Le5nTkBREUJ8gfc444Nd46QlL12idO52p
QViTipENXt/TInE4/XSwKUvHnihSkpsEYF9mveBj4dR+dMSBKwTyv78OP7afwBPS2CsNoXLV/ZQp
GmwoeL+FAccj3KqBXWddmJRHHGF2MDbO44w9sguFh8a1iLY13TOO1HdPVqvc+BBR/adW4C8dklcB
0yrt/iN/k0yiCvDP2UGGZSJxt5rF8zKJW7vr63dyeFLl56+E1790vz2dPnVxEx0aGd7s6p17Ai0R
sDlN+Xssc+vOpmUya+fAOMStOUPaFAP6IQJ1oZrmCbS4/N2HOAGnCIktBoUc43WI0q3pi79h2om6
iaghRizOdxML7vgSjnHMbOV61fDYsPjhfxm8D7mG8vf3TJhP8QTYgnqOVPJL9lq+l8EzgpN3fM3U
giqVwEK/O02pKv3gAtAwaM8gAq9ZNHkIafuruCKhhDQN4kf5CUZri8LMtPDO0LGtYjiD6aG5t0tX
RIfgrn8zYBy/n+7+4PHufd0bC8pJztkJrthQth0CKa0MdCOP5PzIQ95Awbv1pVhmgCo9M/4GMTjL
Vdblb9djCvc2bp22IypnkM1ez/hV4zM9LtuiQ4DSZiDq+8LgeaWjd4sNt89cOZxig0Omw0jMWnLa
njo4awRqnjBsIZEW4DT3LU8N56jyZoQuWLeIMPrc22osusEmwJzAjXwiJWO52YZL7mgDFk7t77rO
eu23YqKMX4SCJQNrFk+d7/5CNFw33HCvEt6I3I+AHeiQ7HUT3SEFA5KM2deXHNsa7Fqbx9Zg3Jvs
rRGGfMIjKexLwmHlzF0kWsrZU/5UVRlkYGc/J7chWf/+00yZzf9OFCPQYf53Lg2UdT3rDaqWtOZZ
4CsgBxDDjYHT8M6qqdFiT4cCKAm4V6gPd/k0K2WtCwMULUmowleDQdliTwnh4Vze5QT3Z7gkIXL8
NRrZDNZ6sVWFlpvQIwQOn+YcXSCEPoqx7aG6wrjizZrxW/JI4OGb3erpuKo6HQGUnNjFXlkTj7IV
PHsm/zNK0r49apRAc1WLffjazd82AhYci5WIZwIcBKLu/MEoWK+rRi6hLNIR1Xc9zpcak07nZcTy
Y9uH24L8hVu/gnwfXBuSk8Bk+TrTDzBLs1gxnbeHaMgkpa5Vrt8pqS7WN0gidA8xO83GPBVO/90G
ZBUwnf48KcPHoVq9hEjye5MSdYZW+v//FrJItFy/biN7iS4ZgNPRdmyTNeZaETuc08BgFBiNXUnU
K2eZ5XIHb6XpHiZtjpoOt7zb2EupgD2GQ16EUyu06o8ON9I3q5UQQ2ce1rRocPCI/HfwCxCu4n56
V0dx0vFZL+DBcTfe+lKXa4OKgYfVjtZYpC7iHoT7VSHHVLUG0UCYQix21//gCXIipv3FyQRyu06c
TTZTBVbJXNT0C5XSH3dv1zuL6Qq2f04DldHKwVifDmh/v3BQ86lxouHpJV/8buQW4FO+RCHrjdpz
cYtTSHfaEMNvLEuopGhCFYfHQ2cj/J4/ZMjd5LfJMjvUY58PmPbZTvJJaYWvhI5wjeFswtd5eWnx
L79k8EYIGxQcgJG1oK8hqJrwcQumxi+zmhdeFQnV00C3ZS4OBNdoDQcSGkWwnjDnD89D56d6csPt
6gDD5PPJ9xAvlEw89ls5/7KLuihmH9q//iAUks9s1u2UKComWTKYke+RAvZHcE7JgkippyrxW3qP
+qTpPx0guxBRCAkxiLEf5UBiVfPVHg+QaBv3e6mYf6TjPN3tERz5zoVto7Atc1JGQ6YAawyj3xqK
uuXcqM/iEjC7Gn4ZLvJaokkz+AdgzoTQ7QGnwazT+JKKsh7JLaqywspLg+vj8k1h2LBDlbFslHyY
kRLJKtTJElERRjm4dtIuiklw0+bNMiPXQQVtyeQ/rohJu4EM14178OizD8Vsx0NFzKUJ1TZ+01hr
f1BSV+mek0Q97GqiWrzMgMhltZibrxoXEPKqWwhlbHOIy8IMq2XCVeP3UnFM6PoZaMWplXoplIt6
HVIhjBB4B+E+YsNEVAZ5hl1BxL2mvDMj+weSiAhaucp1d2UN7LT7vx+yF95WUNCx5TYfaC2sOES9
0Nw+0CCbhuVGHWm6HVLh0OpeAbIGqujCniF/sQ1ME+I6EB3pYD1YWrl/5AvzngDcsWJLfxneAe+F
mvJ5E6B1JqD9muqD4UF1Cywl3l0sTUlTJZPqi86gNqALGndUS3JKvIuoVnvUiii6siYne9Fx7Fgd
nkBy5Hftou9gBe1XYthVDtl9rzvJyldbMjPwrSaa0o9PfxD3rvbW01DTodBJ81fii+Rw/NoxOCrN
ANpQFocQ8JVrTYNGJncGzHAs6AVm1djMWh8BXUeS2/C6BmFYHu0aC7oe4X48getwYq7oIaBsvTkM
8k2UT6Sb1mLcnusnt8JdrIYMzO9zicB8PXgsDRYpqbhqBUq5G5mz2fywRTu++RZF3o0ThYFdemMb
AiIM+EROJEAWRJxonTZ3pU0erab0v3dmRj1f+2GMKIW8PAwC7H0uXJg2f1ZEFyFjkvxrPWTZxlp4
2Zsk2+P9LEv7ghjpoEzCzZp+80KUn2G5fG0wr4c1Bz79GJRf0dUf3aexmY8W6D49hbFRvlkgSujV
aeEUcUQqssN8LdGNv0Q+PvKKMZlq0ytxoH6EEea7tlCIX1dB+ckYqjDhlf3lYk13hS0L04bdPCjI
YtUHkSrpJ/tnKxtdb6J9YHBsygSu2sPXhVhfKtFqlEfpbu1kQUHdM1KjiVBlnfoq3eL9mbRyN+mc
qISnuvsnsGeq4oATVaMzmvXjnukcGvIQt4giZS5yi5rKTGjur2WNR7qlh6v3VrOoRunVmv6tKYQp
Wop482ErYvkoouTkax8vhPVBmdqsbFfT41VEWtEhK5eGeWX7iyaIBniHMKN5ef1q+h7OynEbFuD9
av1zVq+Ddj/ZjAItMi0n9xKp6+RUXYj2CgmCVpwLNbeYoDk3nXh1cMFJfiLOVzZjJveQTGZH4//K
iY5KcG0UhpWPmai0NS1V0QuxlH5SXNBdrfs61+nsSOT1hTy/bdb5xVf+oXSHbWlVdeR68E/Kq3mf
XGQlcwtkgUUeV83ojl78i9ZzNzILnj+viYqcInbR0hbr+68p1hEO0Rzyb69ck96kswXPJ5LByCWG
XUpONj+Lf3qXYG8IJ7kzp874VT1Dic/tjIM9ZlDQqOaFYI1ugvqVWGjHtm8LF9KdoEKCW8UftahS
J6tVyYdLc2fsisvllyVWowUSZEAY6lFIiW1BJa+8UBptjweMmbJkHquTwB1Q4Pbml2E5uffte2c0
f03LV3KXWXc0UirpvEU2Ny/ZvNU31G+QvEHTEd4raeBBNxtUpS99G/5i0y2oN30WH0XN8QrMfFUe
7JiuYOV/mB1sHKVdTgXjEaEmjuRLrEZFQaYJfLuEDRyFJwiEDyjNVkFTLOlewJikdI8l/VBmOGZP
icn5J9ACBchazIqxOdpYMC7oGSBFXsTUwxE6i807Mhs/UsownP1YE9KhvVCZ/TQDAP5uewU4VcoD
F31A6Mok7l/0iW2Fzi9MP3ctbskv7gr6owQ1L0XhMy/b5TsETi8rguBtFL6TGRGcqkay7UjNfmr7
O1Qc1RxaapVmQPKzIOPtkSTHI17u2Hbn3LaaOG+FCanqt8Wj6laTgG8u6uBIxLdTXQYTnxvyGeex
maD5r7AvFwF5gWGT0rA2kqWksUTF6G0DjMatGKujT94oO3L+txFelyrbveoZgedI57ulRWbrRLsZ
RcABv8HpRh1dr6rNE9TRTgtLCrdD9zQRwFgdy1uneHBPe/Wuxs4RrRUQGSYE3fxcIXFWO6Pa9qpA
wpcR2NjTT/J4WiuMUNJMyBe7863n93PzBntHf5VD6XTa9j6Uj1oVKaK9YuoBuFnWl2gaImSGkrcy
WvXx+qC+glps1OlFBqucF0h1zIex+vOKLZIQiDtGzXDM5fnMfaCbvVGs/rGYl+DxW8h5jtqt0IiB
7ttKhY2EnwY5GwShSCw9MBX9+4guwBiD/MiKXjoANaZsiogypO4fV2ddafXFchTh36LBKEwhOeK9
jA+qgfFvtbOqmHGHHyTLuxSPedkp5vKsu0x7S6Gt6tZltwL4jDTO0wJyzqTUGhEQW7CWscPJupMH
6OfZEh41Pz7X4k/sdGrI+7yfm0tJ1/NNgmy2MyMdhYWxyeAJEQURHl7Wj+fgDYh3bLLBqTPNJw5i
/mmIx8FRsqgAVPt1N8SUSJ+iaGbuEFILfvEPnxsyC3O5LHCdccxKcDblSKBFTJINA0iVHN/tcVTg
RCtiGBBflo/Ir8bcWWlmIyMzOq/AWtEmcfJwW6zGtujJQgW2aqNo6lNczYUpu6SQGggztDbZrzOa
GaqCWw+ZX/Csk2LwpcegA6WP9YGzX+bSYSDqtkBdx2gP1D0OjIPIHArvOqbdiD5r/9Kp/oaQWU4d
g7bMDVUW8GXb3aysBfAz7n3ZQJgOlBNnrcWCQ0SsfFCY5LMZ//IDk3HCFCz9H4ezHOixdgp7G4ar
vJVvFYboYv7EDtiFWbo/plCrh5gGQVNQz9zL8/hDThC5EPkUljXR1xt3ZVVBOLCC5r/xfLrNLitW
V+dikWM+QLIEgkghXKFP6nWTSNbmaDq7TBO0lOw2U914Di/6rAZAdaDKIfr1NcexWfVSwm3rX9vb
8eRw2/m7l351h75H3uiOn4rCoDm0pQXXyTzkPw4a4neUHFj1paWRBCW873he/kioWRVNQARPUCZ5
BE2Hmj/u1KsD4COpFEn6eDLk1AEgAGwmyQlEyg3YalaUEoUqW/tewZ3G7OMGf+m0xGzVjHHmXnji
O5xltDO0CGKXAGAWi1bVQKVF84eLr0lhlaU1j8QXPGGa9OCrn+UqsA1/8r2bkySN0IebIPztw5dW
XYloxtNcG7+fiBNCYWAogsmlYh/0n7uDYTySrFcYG3uHFE6pxYsJIfcklYRvGZL8kiMiCHwSSt16
47nWndamnvZuZChRd/leC1dv8jfPOAucBXvSYzbAHOgizEEcm107snF422nyQY+j4JVa0yt/pH7o
jMMIL/QMZHSiy6N5wcCghZx3LUxvOrIRkkhTwGLSiEjyVsZuEWt4IgocATl5eFYmYThAxjXB/SSG
eL/cn35rtpUcPyUkpIzU0MYcp+T3ZpntYyCoPaV/Gk8F7DL1gBWJHatZPpdZYe1v9HkBKNJyUWgT
EWBMtP1VwULdHRPF8gal1+QD7PCI2MLSS9n1YQBvDjcqLawWI2bJ7R1oxqcNnt272WyQW6fEnT8K
d9AdTIc6dZwbd5z5XbiBsDqlfR1NjRXM8EgVFbJCSZ89bD34xwMFIzz86pbgSna97oV3pHga9GBx
JTAMlwdtd5+sxoywfkwOdD9MfUaB4VFNBhuZWvf72Mnnxj6RjnzC3Pf/t5/bJoiifkUXE5lPNF6t
yIJ0VLpjye1Upe0ccVqkcmRAsRuKo6HMBL+MCYv+erCBF1LOCTju/z84eGuWqG5RYhO5P+CKnkDV
8k9gxdpBKVeJDPAqS/VfNvhwHuxR8D6q2sghL/ITbC06oG0H0GT40rBeU6ATIdXiG6c776iTLTeW
jks63qzC8ql5dp/kvG2JriXAWqsbZ5KxZgaoNb4MNfg4eLp3pjbCKngMEcwDX1cd7shzkV9K41SX
/gTmWe+b/zrfvmXvhmALTUP1zxYKoVgzKDisDSipVd2zN3QT2naaOuBQn7DMbcmftyPPXk9a7UG7
ibULJQWKG0NRUHHlTzq2cH5YPM3Vdr977TBu19q7/8J8Bc8lFFbLDTvdIkrjSNNP4MsI5O/HXT8H
OjAPlCf/x7RwqZMXMuy/KKTv1c6M6ISzSRzv7qpFwHwehshfWxhS0a7AEvMDPPzBX4a/uLINhA71
N7lUo9sgjQaDWHWWXPvgLITerBg+zuXl0lZuRdTbX20dN8Xa0rF7kdmmmIvdGJ5C6I1SVxvpauk1
Ndqg7mLKW6h+6dUjDnmzi67xN5km+eloQZYlhdkeBipRy4BtMz+muxbs3eT+FgSvXpfF2Jew9YIN
eHTGlm60XhwPkBUhNbw0PPT3Ia5gf78n6cKkJcaBATeeyNjSXriixb8nEYC2nOHghbiObFC1POHg
uYIrREUis/7cJreke1gCKhWVVmx84s3cNV0cKpASvq1bI1geoPm3EBRcl8Et/Qcv/zo/Hmk8BZ94
kiZPS/cJ3gKBecmRWrtmtNbNc/SE7NDVnE0Z6Diq8pWS0M8aJMuLc5RC2EPO1RNZ8/j6Pbof5ZgP
/Eu0mWaIQAuQqXtYz26o3Wa15/gLKg83U1CNdNZHD8FFrUbBjaHjzTn3v9SLCn7ikKEWjKcbBtCf
P2pyN06BpsAOPBTOqotGkcJblFfKLp5qkSvRHC+91wZ3VHVgpSzMVWuhZcPvaTr3dAv+Ps8vQgdM
jow+WZHWeDqncvuNBUreAgYiq0DnSAmXw9pyoAUSNNmeZDYZyagvk4voIeWZXBKx7cjfaHZbvs8L
JHYS42SQt1FK8Ya1KNeeOxHkPXRgq8Qp/jiTDGn1IBArbNJt+iPmpO58phZvNFVeaIay8d78rJsf
KL8F104qm7kIcqtmNYuCDGvETNd3Xv9yq6qNUac4PDOhcRL36TfohdxGjC3nbCN726UbZf642L9L
+4s4Kyuua8gQma1VcXj7o0KI9pQfcR5rMQXnwcF9whAeyGatWQOJPKi4irDAhF6bhykgeDfazkwa
Gm9EjC6oQeqwP5zyvA74C0cLGcs/7bnSBg63wvbRwSvFqUY/iTmeXJ3anrcufZOI+XAOc2ui+HbZ
3fR1L2vGooXZFHYZtWyV65gw5bGIbKNmo4BBJQwFpknWsf1yM7pAofpUevvYc1nJ8kMwKOT6HZwe
//lKRW5MCjkSmFky3owjH1E0n0gDFy1HdL70dwIQpZcHnUCjWH0f0XORsQ/vNqfTtZUTZmWFaarB
dCptIvAuOtIlvQ6wcQ0FBeTCmbmBLA5GGuV5A4Xc2VtbMyIuh4bwYXDtVuGtItJqUmjp/T6X59bV
+IQWSA0hOxp3YOR1Co4pheYaFXNZkkM8zbTVWEvR03h6YH91USNmH1bknugFz/nTWCj0q4vji60B
VndBZyxAR12xE4NxmtpY0Sc4SnoRuBNPaZ+HqF92n+/5rg63tgCRXf8AqVrJfMO5+Tjia3c3n18V
YW8w1Pb+ac9MOpgWdaWH1U2zcOGjlkhrVlzf8JI7IUgqtoIcmSpThQjm7Hu8AIW1zc1tSL8IVWbK
oUaScrNoObcMCjDzaizNKs6eILYN1EEFtyYV3+QfZGVqb2Rjd5H64x1I43oVXtmXERg0i/Yc+NVs
fJqL+c77C1IvetcZOvbgc52KyUyXNEk91FSUvHGNm4os/TVDsclqJ4A6NwVgRDUirhfZtoXFWAp0
n/f2DROBtFbIu4HL/LYe9/fIF3u4UUrPEf/NieCfj7sFkf3SHH7s3ANMSp3K5amEzFTltQezqafZ
x4dmwqP5b078jNy1CvpKKX8MouOoryHRI0ZRTa3YOyKxt6vFHrzhlAhAb75nIlIzT3iX0fAO88mV
703xPKBep1Pe7IPzS+r+cEu6c3YhigauD+DFrZ6bS1+JR8auCpAfqCv8no6K8H4Zws+2t2yscSxZ
qjrG1WtTTyTJLtIq0thsp0uE2Uhhn2KxbnK0E6KF3L9TfY3NWk5TyRus/WQF17fCnKs/QlBnzN7A
L0VkgPSRaKfhMrZ1A9sq23Szl45AYLh2go+U4F+vdfZB5j9TjQQygHDfyWbrZ9F84+wB+jxD/O7z
sb6zMim5AQ7xIylsc64ot3l4MKRYkwBu1tmJB1X5eJPg5EVdg9kuk6LmTj48mUj0l8Pi76N79PEm
/DJnOAJwL0dM6Li6ft9EvdU+MozHkEs7WYJ0t6jnFM5f31xAA2cCFshQLMvRS/OsZnzKmBu6XIOv
QhlHxl8Da18s0arDm2fZZD0QfuoiHhAvN+TLaYXSB/6yoh8GqsvinJV1JkeRebGh9IGS181BieW0
A+oClP5VVbmQ3Yirhtwnl9fKXrsKlzmh/73+HzpQ+znDmDaff+k0pZ9h4Jel/A1mfSSXIS+vKbJQ
GGNAbAFnM/6M1z+9JoHQ7y83M81n4PH/8eOywW9y6qbqY62t9cmByRCyZhDDN0SjTkQoWhLMKnpt
SD6wdqzVPzAnibfv9udME+auInc25S+m4oJ+CrWoJLY8+I7P3aNTbnS4laPHemfHh5Ch1udeBgz9
b87SDTkKjO+bWSHdCa8zrWlLu9wnQwW+QzcJh6h2Lgow0Vk+c28iWKWF/LpdBHfQmfWOK9Zz7v4E
a3/E/2m82nWICxIY9XplpIi+fzRNjH+ihwZXmV2+mqXeEcLl30t01u4wIfqmuM7Sc6RFLMaE7Igf
xNrN/40gd4tRXsX9eDRwOOx/eYJU5CBqNUB+1avmylo0TUaj5Wpz9AWmrR7IHbz6/NKDsTVZq/M+
xKHtXxrZP0PeL6tL65uVg+vHdRMeHoaP7xz9SUjcysjY7+OBoEfk08m5F2aKgOVU4CAB6bGr0Zsh
7LWwiguNpMFOd3UM3DP/iP4xPK5C/xDil2Gt63k11pu4342PwAgLTBd6DyOeUpfSdD9OayPPO7lL
Q23CD5b/VPnXr+nz/Gj4ON1OyUo/VQVv7EoiqUW+ZUxdNKHADXmbrVMCBAwYgPjmDr8lgQR2IYAo
x/yhTix7xYSPzCQD2GStXy8cTgH8uy5FsRpl2/jnvzXsMcrL3+hL6loi/+0myRscHu9z67bEpaey
H9Ihm1661FirqaheSSzoqkj5NbmDYj9runU6++qAFThtsgyW+gHjPR/09cPere4nGTBNVbGAEcaa
js9nk0KhGE5YVQsW4+xdtcKYsabDF2M0tgmqnLxHMa6gVRWf3FV6b2oWKbO+mM8VungilNwEh7na
TNNLShgPYv7j3eIirc645NDlVc1tQbzFBpztOThNbbNPm0rNZPD+s6AdegxWIz6kwFdcnkygprQl
fAqA/jMSywHFd/md9Fn/nJr1+w32vs0gkVhIOC1JLJcUfk2J8DkiAFVbJfCTyFqxld5tunEW9yaQ
8ifVxlJ/lcL+73le34PIR1374P9iJCItbc/O1BSbJOargSdiRBqyzvHN36swB1PX10ptNUf2g2MW
hMSdko3Pds86JeeZE0cEY14Nwv4g9sMRiNE8w6iOsQcU6pNKfNCM6Jbnj68JQcNqXtu7GBMpl0Di
+keKEd+P1r6omDZHGBi6sBwYBy8MYVhcvL8mEZAWzw5nH8zQNG5KxQliWUp8fJzgoH4mJna/UYzK
wvA0Xu/HoN7EhfkE2F7LTHth64RIOEkCHxm9cto+wfdX2mCcI+1Hkvx3CrMOMovUk8tjOfd05Z+d
W7AhB+i/lLxUDCuK9xcbEvekjypZIZD4pgyy/Pkerjfww6/qs14YPhr3hcwcmF7tS4at8AnHgayU
XWyTeXC2kSAJfjAYTQEH7ipU0tzjwc6qfgVB0Gft6YssXu5Ai0OUX2XZk9LN4NmJF94zOAJv4z+j
Wv5U/p4asAWgYXIRYJ3EyNVzr1HqQbAhW5oaLK2BvT9+1SfxoUcbaHPSO0N3GaE2/Sh9BH99HvTe
pssmwEkwMDh6yyJ5Alcnv5AlKX+sY6/cyesSye5ONJQFl/xwlqsKekD2V0Ji8dy/SFXsvmwbWBVL
cTjzkTSPj63rmOVhJTusWIDfXUcDMsJi61CqjIPVR7KxxlZs5JF5nx/7AG4+mplv0dfPh1r2EEPa
O0VNFcRGDaf4v1aiDTRKbvbby6uFblV/AnvTf8zya4RZOYtk2welJ1T/qDXKqFq482rctIgCTSLV
FToTEZLQ72fRtKwjyWHlvQRidius6L68bCeOYQGFAwhx5cf37ZmfUYzzLBGYCfnMhOtNdmKfzSib
sMMMieejfvlzmrg8KxSSOxfMq/ssucXSPG8W8glfvLqvN7juderqk/zZQ91NN2IHGc14amwwWqZF
qW6gH4050NKMsD/yfo/AqC/pOonDNER/RSpzUiXZ9cR2f9fzVMoX2Y2VeQDGmtxPYldRuZTEJ4f3
so57JtVmDbl+I15Rm3LJbAy8aWkctXg0HGkDbTWwjBv67sEP/Der1MQDxzu+wkyC0/y2rINra0cq
nzy6x6dvv4UOTYtcurxgA8lWgxlTkdJvXV7joYTw7ibGVnN8isp4SH18UbEEwoRgiP82+P4hLvgy
HDxBNN95UIJv3AXklFpyb8AY9LOSlBI7OpXlanZ8UMqqCBzTTyFzFeQevwJ9YN3SO6nvCn7yVDD3
efdHzj+0dcfX+R286CSN3obynhGhN7GS4/JkurZTvS3jqs/jhmPjOZFQmWLoF7Mttp32k+wV61Ih
5KYTuqaISqyGclA4veTnSFsdxOXTDv9rFo166QhsVjtuGbPcsQAGk2HY7cfbK/cLKrs34KuM5DU9
ISFy/XooXeZSKFqXK/u+wwUzMViLWuDGj/SXPUwrfbr4CBWzyXBVfhNY9k9UAsFl3w/3ADsfLbZs
NBwB9EQRFdROuUqQEh9yTR+Ugweuk1RiF0SdME17b/FufyA0+uVHpL/LJzo1kQ9X8ZKH+AD2RGey
bL4nvv2afNxDC9qe0/jlWfi6VogPsc/FMYLhxkNoCf8NBM488Q0IeTd1F5gTfYnvjtxAZh+Ub9yx
uWNNKS2fz82dOhLGqsebmSwxGuxMQDgZrTZ4jzMuGBrUHqaD+oaGoH2lPNWSZnFECEF4RBNHw34G
T3aeMiAxRtsomjPXgLPMYiDtX+y90CNDOe+C5YiRmJoyN0fgnQI+jt9Ha12vWT1n4Sr8bK8vNWy3
GGnsa3QFcDpP3WIXV8rgkPWNQQYYe4Dnc0zzkU7f0vCp4/36KSK4b2IRcQ/6lxUEltVfO7QV7hn2
DgINDMtJ13uYhLoj3oYGR0LgYBFecojKWP4/2BB+BqfQwsvjwJBMD3WdX7JNO3Nq0NVYxeBnqY70
wuGwvhu/IJHXVysUZ6NXhhSDbmiON399jvYTbNuHGLT9Kxx3veQ05J+MxfEwK9uxkIljbZj+bIL6
WZwrxxUZOkGtb1f3GXBVHgFa1WbciEgntmE1SjVKEOS6wDtPlwmWF1/831dgsGrUM/5MOGupMYB7
RthsBUyv5W62CD923zqqAzywcdmVA+mW1/xK1XeQHh8vtq+3/z3cJelIxJSW1pSojLG+H6n5NGrI
1e10SkiUGMKBOKUBiZH/U31fcDpiJM/r0SSx9TGip7B9Crhoy3XzOg35tjZNxDD+9TKylraKHRjo
ORkoA5IivZImwIJ99zYoene/U5Ll2NjRpTqnTnJDI5xG+puBrhxqNiiSbfB6bzcAqKssfJNJNsa1
TG8Lj5+9esAUqDYO7i/JBlIXRl0NE8+V8pyNYyVA/BE7SVof/U058EebEd9MDKopPLGzL4JF5g3U
wAV6jVYAFRWokwSFGoe56kqcUJR1XFzzSxe1RAXEtTz88vnhiOR0FjY8WyN9tAuEIEIu37iweEP5
dh7Fso5Hagn7t05tSCloMJpoTUlv+mnbUq1FIeap+Y5vkoDz2t77nt6cu39qhA7wEpJclK8RaSmy
aoKV+nqU6abXjrpXwDu260/Kp6x3+p4Xcg4Dy2Jfe9++4wvWaWaqTescd8ZkSpbklWhRhtHkzgeN
mRhf/j//wXzy1+QrloQ2K4dzFcbKJma8Myd1Dh6C/KpvzSq6JnFkkJm6yuCKWbWQ/yvt7dJGS57C
b6L3g74B7xALOD1CDV6RwaOKXR+zq+o4sENyXt/ghneOMspCe0qxm1MID+IOcs2z3SQWUYwGoTtK
D0TJsHriBHCykUEhKDtCQ7i5cz/RVOVny+YR0r+xWoTg1Y2iT29Gu5zaDHas9Lvl6+0GtBMyuZ3T
2gkNzdodJGxUu7vbtNuVwB2PrIESNMisZS0IKJnDsnBovgrBE4zP2gufX/6zCyH3koCYkfdsJBft
LFenNdP4xJXd3AQVuTp+UmUh6dhOGnOTonQBTMuGxn4hd/QlJXGvd6T1/z97YEHSWda1GAylOSQD
EB7WBJtfnTdCRHzzO2eyFB4ZLmC49DD8CxLRlGqHVveRFClEXOghSZ1Ec8/9y44USnQoeJJX/h++
/5/1W8NlvA5gb5Gu/khFXbduiEpsv9XnF2e8jB/RuwZszGytP3rO3z7xFFKMlOZOh0qd28hiSYel
TmBGTCbbZ5yq3rtCTaYLppqN/ZojlBI2wZ/kUCWho1c0OtOqB8BML2gipQluB0dcRTpZOGe0oYiP
PtLedakwUNQCv9TQ3jCnipUJIklt+ZG98bTtO3DpZ5j7msfBKlz5wgLx23M/dbHgXx/KjzwzYaE4
7/yJ7saSUVR0Lr1x5maaeJ3L82mQ6JQY/OZw6bh+fYdfkGebTAfZX1f4KIOc+aGd5Ywt2vw+mcPX
5WWo1k7Rfm3MLMuzfb14h7mYVPj5smFuzARThn5WMl2NP6D4cU6FVqTpqNLkXwtTvWWLNu1TtbL7
hZyBJq7WaxILWA66V9GMRdQgV8YKJVePxThmdLUL+qbbffPQi5fLWnoSlN/obFX3zhH7qF1mIaRI
g6u7SHFlROoCBvzNAF7HOB2Waak3xvU/XmcHXUZtQC5mk79W/2fKx9tbUIzdpqZnklawGKutpzX4
Jk5VEbpkQSuRZP2czn4ufkzwfAMqc2knmVc5NYBuaV+/C9tW2CipHQlLzfoRkAgOG2gcTL5YKhen
JQfOzmCe8R9XmYN0XaLIA3ZxcSRcf18S0LBM6wi+6FmRIkPgM3XdSZ1p+KwgGoERyeiA73hKZ1ES
d+5zumnI9qc9/L6WEi/HlNqPJaZt/L99aK0zfpo9TCP0wJQdrOZ8yU28KEZPuZx1Dy5uPvixYDFe
Lv85RdgRMaEhG+zPoyybVhvqmTBSRKJ5qyfshjTTbwExim9H3wejJFTtVoz9YuV8Crpw+23+hCEw
Cc5BOiu3UpkSWYTwA1EEireRA08Jp7+4F6SJ8v2Hl3BPvA85LQNCFTh8qX/xrxTiHTDb/o+C5ZHp
QskZwJIiIO2T/buuMQG3cavFOoKaJX9309cQiNptcT1OYxYui5njs76hzLEUaW0sMBky7d9/D6Xa
9feldcROuJxPDJH+tRQI1Z0ypjqvwInMi8ILQozBv0NzROgklDx8XUpJEHtBljE1zIzWC+eK197u
qb4nK9n8jsl5sg4u5IWml/sQgCKf+tHAreb+ljJ7HNuunyAaBiQEtrJr2cP12/Xr+Drt9dMwUMab
jTen+D2g6RRHjEGT0BIaUrc4SWFYeaEmRUeSdwIg7Zs8q712g66C7mFHrpvwKmdP9FT+RK9sjkD6
yXRnm4CpOuEfKo1UOZo2hl5StcbPHpqxdSONI4qNDJE2QBlYAM2XRaV0wIahKub9A48ISMMUT5nT
hRNSv2xd3RDzXYD7vNB69iqEGXQ9jrMxrdpKiaRPwcsiqOLUUbBGuuf6BPx8GO7S0YVhueTcvF8o
uxQOWimFdDyuf0DFTI9LRIAvPBLLbCwc0l7sakD1NSrX4TXqyLgwwda1NI80hjn8qowFlo84Z0ZH
F83XH/b+GaYQQ+Vmu8vfvDWeipDXHWoML9jm3w3nXa80gAAj4nttKAckqR7xLj5RlJ6PcqHAF4rH
+2EaqiyywEk9tNSoHrX8PZE1hPuMivAM4gyUpp0wOXbzu9gfgg4UMzEQW74IA4h03t+Hhh9v7sN2
xUb4+rWK7h8Sr/xo08Etq8qlXIjHhxqr/IN64ez2NhVgO9fV8SmRYsTa197NAabJf+sA7AdGPcNm
qAINOwJ6+06ET8k9KpIysJff1HPi+K+UKh+P974BDaJZ4bLF7u1EMUZEmUp6SEPABcZYiSZpwEuS
DZd9wSLmA5ErN6YS0ndAHLIUJvXuMx3sz15E6ksasSbCglHvN2kgiXnv1Uv75IyMVquzUFtoxYM0
TfRuA7M89dgNsh6hGBWq7oFBNQv6pdogdMZDWzHv50aEab+IS3MnzaLQRTVgbzrpx3D/GItDoL54
BxhNfT41Hmk4mXszu6wuLIFgXhMM/NmYAlZi+zZyfvy4tj/JHpVHNedX2NyX7yaHDakYJHwm1i3L
6geJW+nDC5dB4s3uEU9AQF7gcjJbvhhvtVjCY+9PsWU8LgUnhADY95iJavK7M+A2Z6bprqdzGdXM
QUaUWVDliTPb4nzeArxckJTC1iyW3EfVK93+uguq7Uxa02kJLi6G1VjKQ4qY4DNZ9nHAVGTJ6R2w
7lOd4f6rSAhKqSrQWMA3xx1YkoxbsDu/Ax4PvruVofKwM7W+Bgou1TyiljpFpPFSnjEdhV72dIHY
mcOqLc7TZk9dbaRj1rUbbEwpf6xwiK6KrR+xro8e/5l7kqbceUxROUNKTnq8a+u84SI+JWyVTU6K
4UHnd38UrVSOAN/KXqbUQ04TsIuhEHump0gbsre3nDziNbjGH9rGO8ovF7J4ZJbjZU+ZxTb4Zxqk
ESRSwtE+vngpkxqR2JVWEAVkODssAYsyBbOE4UCoyKIlbKz+vdfpSdGD8bk/kSw5Pju/jX/xbVhz
8MUkgcVozikt8MxRy6UJeiDWcRaY4EnmyTljyXNUCJfap9ZLSP+LXd20onnf/axtKugQe3Ie3sGc
644fnIGWgN+BV/chxxt+wqnKzpQ3OV9QFJChBRm7gsKMOfGeskQQe9tZA+oEEKCGdWNrPliAqd0+
zawbtllIQhQ8fsioImUM5ALVbVEtzSPiz6JrOZiz7oCMw2golbrp0XHkMAeQSPhLz/CoGLF9EpeF
S01DBYCiFj2bYqLqbLJAqA9d4wUZahCMhwMefe6nKXmkzXIXKC2afrIckNIQs2Amn2/Ev324OEaM
brOvqYuJ9lFguatqourG+DI4ENsezs0GjmFinM6ZyvrAQgvLo89bAUQqzt8/is/pL4VnMsoUVUpD
C+jhgevhHidY89Fx22Ri1B495Ld83WKnz1m+WYOZFfRuBhE0hxSuSWDBKZrMLxLCnsQjxuxlCIBK
eMmtnsLE4l3U63jzji7j74bz5bVR+OBuYKid5RbfOpBOF/biCAu5r2QXRBaKMu+QotyKQCkCJlxT
S7XDIFKSRchL/j7UUEEDxdV88q59zkqF5fMv7q2d/bwTLZwd3vvE70koqs5JX/g64tUttAlHu5q/
QGa77N+YT4gw0NPntsRhs9yp6wDRBwiiMAX10Km7FHRYpgiJtLG9RE3Dew5obx7b4qPCmj3OomwH
ajVfMhxddHFnfCdjokhIfAtTHXUC28KuAFrQ6m+MR8dYYkmwK9UR1FiUj5OZ9vbu6M56KdvoV2AK
VcNkwoxXhxzo/nixMsdFRzsC9BggOxxEs7E6cMY9DnJQQcpAfTBBh2tPhm168Xmkktdv6XHxkGMZ
12OERpT9fqJXMPdPJasRGpymtF4MBs6tJTanbOyGi+HfyTyDuxzr8LoBNb6sI92FmHpEnYReEHez
4L7texGGizGByQIUcskkLoNbhjFheFJLTS/mEQnL59u1xh4a3TnB+461oq63oSImQLZE3fSs6zhS
qT1ilYhihw5zl14e1BKHdHgAef0RimSoUm0i1evHNvADhqOeOjr7hrBR0t6CT6zPZTIflUMy/erW
yl5hMovs8HhGMBnG7q9hrtKTWX9l7fWrIZ3sRtZwClXOnDbgdoY5gAj+0/C8p3b7bhi3SbWwS/sI
YbliTXtWDW/LXilo7HkUWa1bBiDmC+ScYaRzzat36/dUTMvk6ZkOlgFfpv8R4a/2hUED8K4EoneG
ODBmujq9pPmGbJUJWvul+/c8oUye/0FMlddhjrYbo4xhlsZW14gtJqYgjKmy4f+N3aexI4mzwOkH
8QYdi8tOMbWXSSS4flGvARmohzeaJ5WQPTRejGYW6fwOj6+RF4c6uyjno23TtDQqe/riC3rQEhQn
CD53muleRPbT2YPv+ugazgF9cQERvUViaNKNsLzNLJtGmzxF3empbWPp7Z0zfr8XlilPkL6/uup/
848PJ+GKR+RJuUy7T3+ki5jO//+rNWysvGzUdtzXl1tXhf0jRrka6q9LpdeaJK83u1BONW7p9ARC
fmp1yUFwUg07RaXTJqJleQdB4Im6mKCd4VTLoQjgpqw7MiCLj/T6HilN/+58aR49Xrq0CzpUJzuT
ZtXgeC21KPJAX18bTjB1cEONGil3VSXMuWbNHRSIigtT1IN8FLphBcflN/bDeX0TyVryDuSLP9C8
Eq+KnV9HJ/8u9q8kvO2TJqESiIBM6vCdPjUhs9eMRBUz8qb+1zP+85ByrxrJDI8/k4i4pDv9oSe4
YRyZqYefVxtXNbVBWe7GzVM5K/SGid810o2zJbRsCHrBg0PAwZ+PzbfJkDhf7cp44M/31CPLKkmJ
8zwLr/rAuaCTs6gtv/zl6FFOd9Srs1NdQJd1fRGEzxNMwzNOONRxptZIk7tjn4qlvc00pVkm8JRq
S/+cQ0KH2d2MmKcaExbb/wt7DcG+1nzsH1rUojdloITa+/PeImuVYGgriMSq5YVKewe+2s3662HF
bSmOXsY6MeLa12cPeu7GcQkyEmV1iwatoKEUTmBjVZrfO/BZsgIY72HhqAoTj9ABWKVwnI3Dw/T4
wuTsE4XgeB/spfANORhjGAhbqmpAIf8ZShp0uH1VJd/gCtYPMbhMz6PI7SOpqyXxodXkJ7oJU33X
OPp3pP8iGiCRxw80eSeiam7UVMuHBPU8O4PpyjCGaWCW+JyfmlfJN2NG/TiGH++sClJ5DQItLBMQ
1OvhOQW+gJQYDLhAkdzIoMPFHLtZwn5YttVCG2Xq0D4L28gaipBw3CHdrs4rl7fCqX9LA/QQ6SoN
/oU1wFY/OOJ8ARsPkcfjTQBlCv+ZtP4+zSxgL+Ul2VQEm7YL7NzYs5U0jAXq91YlPtbk6592Xp/J
oCY7VKHAW5DjEkVxamb34mhcqLZ/jZtKUoslSQwWoFDkUys2viOZQNgKbznG5XZYIDw3ycicu7S4
HGBBBmX1qatkIMMm703nxIWaXG/F3KGBzu2kLSUJQnRzqjOlvJfZr1NjLwNaL0yBZCCZ+ZWCARTO
lJXAJgjikqVs7pPewgzDKfgYjhQGhIxODAUZaeAZUlhqCk+8ujo0w8wy35wJjt5oqgVzOQXNFqQW
58U5Uz32whtMQ4aoL5aOFi/fyvIGDsR/emsbVqtKN+1sOkS0AZKoz6hB3dGe1eflCAwDUdh6kBWM
FRy0epdJsJPWWZaEzqG6aTm6o/5p+HwOhuSvCDRQxouyypiLEj/nYK0cx7SAWCVz6FS2oTL4O+vh
ZzoHMgqE9NDaEswJ0eVzVhQxZSTB7DJaXUpt0MyWlmsQ2d/1Ge2AbURgZRU34ICD16VqoaaC53lq
aYqfFTRXAJXAKNEV75F1mvXjK8loz/8t5qSyB7jwbT9Y7DcHi3Pw+M/XJ9DO+9QHzAhwDEtffPVE
7p47DCw93tGvKkx3Jx7W2BfgdYnV5Ex0+nEcHlvyZvcY8qGZCcZRrW8XbBh216hQcNJgBSiwFPxO
GWaHp/VDvUftUPiW0Xu4EZ7s15EUx602hFpMCoYupnk0TswV68FRphTW9DI3O9HcycTqnzHCXvRi
UhkCXwEhzSMXyFn1rgkzIXLNCqXVSxB9aSJkEz5LL5y23KCQG4JA2gS0XxNn1+HLQ3Y0QCY7TRq+
FKqa0iJtGi3jDkYhTtttfwd7BmoGqoTd7l6NZfLehoPmAFwzknJ/V+lAEuMyr7fpg6ZPKGdA0bcI
oTtUujoWXBEyyxxv+BEwGUs8G1TbDvM2wl+2ov76na++XwZgxAYMV/7sdNKd5yoTQWcgjei8aweC
FKtnlBAv6Yh6Y5FfzqPq52zziH+qdXoAxXVs3gPZWahnNtwp3iWOp4fc2MDSFBvseGJ57BaONxvR
F6d4VKr/pMtAnjWMcOBLcMbwGxLVyItbWobEDXAe+ffDiNaaFSN03r7q7VBQW9Q0cThDZ0O8dHBZ
gj6TQkSc6meAmDWd309uMQC0ctwL6KcZgJJ5Yk4u7ma5V7IS4ADu0wDYIuV2efeRVc/IAbFLsTrl
dgwKPGCed9YsCcghc/DLgOQBER3CAdjUDO21JiAW7X5VTWbNt6fAU8x6M54Y3JwDTWicEmG60YTZ
lnHNZWCI4NpNiucdrBLNrFkvjJKS10BpOsrEpxAZ/SS/+LPj9d/NJaZzvUovJyns8KOS/3MwgYYL
WxG0RC2nFD1Zfm+gENTq2aNeHUfwnYjv5g9ME3y1iYeDoROLWxwBl4GalIdG6QdrRdCpQXi41ssy
9VytlK1sr07lwfBFX5D/ONMPXJz1VurxkVtTIf+odrXCBPll/I7M2FY15fIpUpTH4X0LXYnqL8WG
aBTwVVhVeUX7QPMUlrxtnU7p694JuHrpf75ZZgmqu0cEncCMyYs6owt/CHl+SIniUoB5wqHh3xmT
P12HfZMOnb38AJIXTwYm+8nwMYJKL8sHNDoWtIe1r31f8OFHuZo3WJ1zmBrJB8ZTVmT+NPkdZpJl
6yX9HkDxIbqxFz/gLHvZ5uC9bH/e5ptoxeRgIuw3Xwt+WFQDVq/xVGvpWRpduQ9N3yU3PfbFz8x7
I5oO2d+LGqTYDcJDB4O67wWesJ1La4+LOefMw1cYGbfcIHkzeU+hiaqGjQaA7jzFKs3gImkq1g13
FKfC7D7rP/3bGi0EOlmKwTCi26129XufSsYywzFchP6SeqWGEp8EkpuTMy7r4cz4GepcmWwNPs1z
peicqkSoEz4auy0eaFJDkzM/pD4Ugsr4CglI+gsZ7yVCQHBdtJCaH1YQJRwzHeJ0pmEusZPdQ+GV
P756ErNFknSSGV3kYwMRX8qyz+yXbKxSEwGlYNFf6lCpnEYty51NSXnin0QdnE2WYeEEGG+Qih9X
otdhxw6XD6bUOfQIVBJOOVr+JM0agMK0Pm+/AOSmhsc3lz/7UEbgse10pyz29ypkHxvjgLC5bbVU
ONDM3ZM7Fqt1cQ3gbPNpZ24IuDWpzuwBFArqdI6QxG/zz3V6SEdw5j3Wcv5yZOQEtXkNu5hLXyBw
n2xrZqCViYqwFqKGJBo1X3z0yfvxV6msKBVIL6HkGFsCtzDwGAlFHUEUsc7X33tnOnP8gREQX6/x
DnaKMVj0i9Ki/5rD8L7zqMaCQ2DOSBwWdsD9e8n2Un8NAzF4KTCpOV37qEjX6+AZQD/C0hXPwXLg
W7WaoROByhpCXNiQsS7epR07j6I5HXdn+zk3nXOUok0t1ONdS5/2UOCaTsCFEYA4ryPZXbeE54aa
5sRHX//sIbrVfHV3UM0qnYx+iY3wnANC0jZDTYrO0pHT70PVjEbx24oWXBgZ+j5PksvGSvAjylsT
IT/ZMgzElxpeUnNaFqMKC8X4HDHJuw+plivG0EJ6d+0L+vuo+AadYU+Xxr46foFJsCh5xnw6981D
bPn+9iRXB4bAnUyVLbWtBdHfxp7n/U5tjYTEwB2su9U2poVWNkVSPy6M9ha7h+8QLqa5FyQ7T+cG
m/BwFOpE65YAbPoLTdSpPvzkp4OJBPT/uP6RuoVSmHq/QxtrBxKt0ywpDgzMKWRR0ndWAWsOIo3u
+6o3DqrHLPfRZR9gHBV19kG7VU6i8PVuGi575ehLCNh0Qm5M/HhPLbIsYNKTXGOndwqPYdT326ij
eYwjxZUtf5rgw7iiiJaCQW7T14rf7pLCvhTGqU5l7afD+14Q06m1jNceiQLgDwuYL1Tc//YN39lK
6xR4HBwIzeMPMv/k7NEH/JZyBkLDa8q0IQdAsK3op87HSBJnoPodlQ8UKVYdHPy5xYo/wHEyiZa4
dgkXJeJUohz3GwcmCJ4QzROiJOLeV0xZ9rj+bT6rxwA/MLqvTxZ45X3g7Tu2GuKcpIPK4rXakhPX
MIVFis2N7lrw34OUErNVHukz5rSxBn94E7QB5Iip+M4zNATMALXAtWSyMIL38aAT+YmFTrGfRFT6
YdY5vpz9dXk5qpCEcSAJQPb/LX5ug6TZ0kQ/Ddq3CDv7PmxUyYo5B6msIVAW+cymyCtiZP7zbqZq
ZnsY2xEGssibs5eNA3wzL3IpHF0u5ifkAHSo0YxBoqTSPTKfMlC2bCbPutC5zUFPIHHn22TwFOHg
atclVsPiU817R8qhk56jrGpRYB78m1J0i34ILkOnIJsgqXtcTou6yuwLjWznmmO3xciUGUVZQ4b4
ZKde38OFlBAxJ5k2GzXkDbDam/3D6BdE01QCU203VDsBZ4ckMLQK6AEMhM2M6kw0Bm9+9hzfXIKt
vk0504P4bAkW/AjLWNlJ3jK97QAQHS4itHIWqveaxXuX0Hyq2PeVg5w0uDyJULzb7qa0J6fKTJxZ
u/Qtvk/QajUEyc/Ozvm8cdtDvEbf/EzISbUjeOMRkPf9bK7gXR9jNI06h9MfHmqXxnGm3jrU9+ht
9qZIpOBxD61qyVVieWqbykBWDtvXl40YLZoZ318ZW1b1qNOhUz4QB0KhQeWRS93jYhc9w29G0OD2
DK+t6udLhf4yIhNv5L3tvr5tzg8thGDRzX71Jxb/5C9FWxFDfnxS/LgI+jCHemq678sxoasiWvW0
U8a9y5TRIL7/cXOaCP8Gm1XVevpZVO0Jvu/m4EiiCa0gbonjb0pvylQuxqvZnHkzo71DKgbiusw1
8mod+cRHPTSzZR1tuA9laUUOyoLKvPK4+knCgcx4g+htL2WwhFcuW18vUnihYWVMe5Z/AsQpvxPY
ouPuK+HQD+jnyqECU6T1d4GuhqEmO+/VV/rtpCcCKy3yI1Ad+/xs20x7rxVIwj2BsGlWcXZcZO88
l+C3w50iyRKW8iVOCnCllYDYCxvsYY8Qz4pIzUjGrsFuU9Ag5xJhdNr+HTDRVJefF26GOmV0jtyb
Rr/Ko+yxFQocjUs+VVMnRM4SsyN32Gta7l1321m8FVGDu56fxV7N1ZDmbELx0Hj93jho+Cpo+lx/
9XRp3xAeGZWxD8fjTzK+l865sZ85VdSQ4sdp3+5P5vrSGpdlo5DNtkIW8tqEzCJ1izxLOPAHa40U
9rrT8oIwTpwHRd5YDsFIF0yYBcPp+qB6AwOvXKQfXI8DQC8fKeeq96rBkyZCbcgBvm9+/6qA24nI
C/+CVd0Xs60FRMeFbOX26RJUvsNQcFzLvAtj4m1YV+KXtQ0sMxNZDVlrTFPe0RdUQBQobU53V7B1
k2KMmTGaC/wR3IZX4LZmXWrpIDj/zqQRrm3F6s5Lvl9QfP117UNhBUeJez8cFgkF4DKhDtrwKUNY
H+jZuJnned0Ff/gOPaL21WLKoSaDBO7kiI0c1t9aoF347ekwmRSRLLH5E5Lk10dc126VcmlbWa1T
gBMEp2j6TTAg3AzEPjDgbsAHc5U803lKx3tSyst5If9C+KjpHnEHZD9k06U0wV55iEC7yBTCxvCg
V5m5GLmuxGncoMC83S8UD0W7/ZmngeTsPWyHDdu2pUoLQvpV4MmYoqKZhIMnbBF/jSMI8hP85o++
RwhepK44kClE+AfvqBZuFJ4cMvnPz1cRExw4q1YxM4OoruqD/H+YCVZUsYY7mTNFGc4rb7yrMmOp
VRablZ09TEKe+J7M5Vsu2r3iYJXZiiL7JWYu/6qkPGH7WhVPoZSQ+/q/by0jTSQZuawr8Y0IH/Mb
PqLGswc+IIYfqt5plTs8TXnVw/ZiUgl8B0sfPBl1d4OhrRcA5voGDofJqq9Ts3ZpsjxfRT5vAICr
Ie8skVO+JUrjVGT+5yN5jWSaQV4oIJ2i08aR4VtxvCAh/52bkixFl0EgYmULWGLlepDXgr+a27zh
OxMg6jpjapGb2iBN1E+t87kaGt8GMwe+evBCiZIAsDwW7KhNQYq4u3UV1eJzhrP6brugNeiyouyA
ofiDYuJG9vTC4q9pjXNCqST3n2JBakQK0QTEvwHfhyqTnFMUu1vXO8BG/jbESxvFT5Q70QakVtbX
MzqrMA/c9EjloKWjYuQEaDfppyMhKD9OyahRT5TiYAtxrYeptwHOnxAAiC+VCh59F4QQ5L/ZMNMU
j/Yj5eXaKz2iWSRaE9Yu9QjgAYuF2Fic84BVp9QKdc8WZCMphr/HfNFIj4Q7SN+sEC3bsnsPIgvS
mM+3lFYgBKIbeq3b7odohkVJ1rPLmbp1TvA/DRBKCi7wy8VMv9JKpCLsYYoW0MGJhSsQ05EulhAM
ezDlfUl4b2Z+q/Z8MeUTGL69l1hcPz2/hCg41dZipr/L0yrXh9hTO5Ej7+IgF3bhQiVSWxMuYAjR
XP4SC/9rlewsxycZ+PCqUXNgJflEnMFXs36uKLbOTaX9nbOlG9nLKHx3jOKBPdme/FZVDOyrR0kR
JMxqY/7nRahmh/tSOv06lQ/0Enb+jHuV9wzU5LnDoDL3ir/tU/cngttLpiLfmi2OiP0FFUw4Mssr
NMn3wNRZ6M9THf6D0m2f+qe4dCBg/H4oue9xTDxgowtjvVawF743ragz0iKpEkhPQ5g6d2wchZ3Z
ZypFwwqhKBGyE50VdiWQHjmga2r33Q95We/zFvQCHvjrRXekHYq+wFDBoAjOUMb60MI65WWxdPKg
APkc3oLofGxvQoac4AUiH2Dn6Gr8bEmZZoYCilWMcSDrbyjotwo4Ow+maDHGgVPQ8aVMYBfVe+LJ
B2ylYPl26KwYz1kfU9oczgfBd2zEYSS6jqwrpW/5MRedyZjH6Hz/EdJoNXUSkbl+xcGg+cEvohkH
Ko7SFb7599r1jm7qdVepQ5gbeACO7+AyfB9N27tbBKuzXHEFNMMuF05sgadFBqU1b+ia3zGSHGhP
o8R8tOUUR8VED0WTWEvY8O6x2Ky+aXxjnEWIZyyKuXytoT0pY0mci6cYcNKj8Cm6F4SGcQ9tak/9
/eGRrVv+hqu/WxDJZPvVSgtutK+pGvDz1VWT+NW26+3JWoSOEZswMtdab9dAS2f6j5t2UFao5uAg
e1Z/0Dnlux2txL3r9pUi0e02aen/e/pysk6FbxILk62f+DYLrurm7U4xhREV5vUW7OQEUqj5nLMr
ZzXOB14dZgILRu0HLBsGNFlZoLRWEF6TUuJqcNslNg+KUy7L0zGHpKN4qbauZPvp8t6Z+jsyvmw+
ZPlrGuQ5BMK8cpJi3B6jLKuCfxmEwQB2np/6eZhiGDurUT7WlFiO5SSO38wPYznfyYyxYNk2A6vF
3kI6XYl9j94s9DMCg6jWwumAcAEAAYjwyxuzZG8c0F9GxyYx1AG5pL20tBPCJMPBLboN0+vlGKF2
UirHklP9AfErnWe6wVnwmSmAe/8yaOEl6/rBmntQwdVeJBdB5iuNy0Lke8LymG9ZJfZQJ7Hodkn7
NpWBmHYB082IusXhmoZ1tWq4Djyvhsb2Uooq3XoYvbInFzfe8bC8pZnDJGt/N2EHW3VnYPJjSTIO
m2wYagNWVBmHWh0CpDAu5vJr1+5P6hE9zVahLK6/9LysdeJYfilKV4OlAKLxgqvpOJWkGBYrW4KT
iREzFzwrwpEw0REyAXmTtIgiZZb9OxoripBBecPqFook7c1JimBzkFEYD8PMIBaWtZCQuftc+iiC
FbzPOiadgZrRFxl87F2tUrlXiWG2LStE6P0+Xbj+nag9T4Z76oQ6Nq5TbxzGM+cBUNfgbP8q02zF
djg/RFZsJv/CDWZT15U6nzq8OD3vyVkZchq7YO7dFPiMEq6XbLORJDyUZcD7P+Uf8Yty/dkYkBu1
UIOm5WgVCSlHtgQZcatHv1pEv3UfeDQC7l5TxgmM2iBO90IJR6xdYqrOoXTpg8B2oDG0fDGTLLXq
M3x197DR2csevoHzTqoxFtznAXscvyT42FnbxgMIpIifq7Nba5Z8GvaPkTZ5/5MPLQUyFJgGqWrT
DciMMWsOTrOQ9D7miRjrYzHRp5GuUdBamF1Ow/Zg9iT4mirN5hxMOPuyMp0adxjaYpxaUfWd7ebA
xTXOsxKLTrHy/Z/wFo+1MrazBuFuPLECv1sUUljD6CXwnqD2rW4RjrBR+kluB/K4GMMFwzfx7DJF
kfo7Jm8OUwu+fo3vjKyGPl4pzLrHHzriNjPcZEiwAWXqpk+HZICJWWYpXXz79hyxBIJiLpgCUsh8
HUKxLxQbKVxqXn2TFkH6YbDi8/A6eZd1syUrL3NDBxw57AwMA96ozkd6T2W6kc6v8EUKnG2C20bO
U5N/0V57eQxfwYQL4evDLHGWcIvBwyoFQUhWosLknrOoCYAjOoQzBBCSe8ZEn+BaW+Ir9jvtB4zt
zLoIKnmCCzAxzeh3Y060NwdpvdeJEC3HihE5cAK7d8mMvPePO63rv+Se3BkLkavfw793MpTQpTWI
YLvnylyB+lGsr7f9936Ea/x9W4OmPKzH0ZZz8phqN3NjDn58SsORr6AH0qI8Rsahysz+rVF5AOxA
OdxE2YO6YtVWGD+pCrc+bU3ox1FBDbrA8RwvmZb2oL+p45wBsLVunEnTy+3LraQDNc+m3RLLvyxg
RVrIB3ToYmAWGMMKAqD6CH+v0HifCRy29CXa59iLb7PKmKB7/eWQNVEeAf5t9NMLKut/g/lVroIG
P8P72MAfRAbKsncJ2w+10lwJNX/cZUm13PKV2P/jKxQ8Qm2tUbbLXn88RzX3r+tfPdsJhVENxI1w
2RDK1AZKIbk6leVk4SwMGrZmR9R41AxGXewZgGIH76rbu0AgtKpXwlS4xLw+og8d36xaNREOsD1m
Oj6wauWNhNEn0yasHbGb5BvVtbiafMmk+s9eoz0cqFihZNMefdoljmGMYCiXmd2HeM7g5iihUMQN
s4gp0LktFDJYTRzo9F99Kp4o7dEaZUL7oEnSTtAOIUAOyEtkYiRToEkxh4CuXBrVxVxzivFANlOI
Fnao9FPQjUjIM5QIic3R+99KB0IfZnVi2awyJkSXQmcPH+75/+bZ0DRNgsGxFMUuT638cD1fvgMt
IKDOXkDIbA5DHNQF0pZRt30wbYc8R10tGu312yhTt8RqSRaUq1pkBye932rL8voamL6p3O6+VlYZ
CP/IfU2InVrqamCobngOCryL44KsgBopNvI5Zw6iPZkGgbhjdVcTQn2/ez6Zm0Ns/dXedFbZs+Fv
Ssj7GVuwDN6hPi3K58SQWdBHpTkeeWXrDkkldD1eOj71AXwMa7VubaXFI94fNE/fRAHhcmbA9Lzt
fmP451JqHGe51a5JjHFBBgEVeRyltL2sq0afKNIVByD6fDHPT96rLkgZ5TQ8RVom1B0kbTYu56xN
UKybJVEBMfpbPOC/wznzER7eE0iPBqfl/ug/GoAqh1u8pcnjJg26hsHxij+KvTe8RJUfc+s/2Gfv
ovwlasFlLlKqS8zHj+OjRj7kTlg9WZqydlZCX6F3UH9cAOz1Y25DIB9XGwEOceGSaQRKdoAB+zF2
gu3ebrrnvVuRlEnhDHetZ+KvgUq1YVPx18cJaZSa4ZVKfrHraAxKjr6pdL9YGJzvmperpHmcnfqW
BO9qRNVLE0NsXBWkjj5pccS5mkXObsBs/cw7KgbuWjubUI+4+n2SW/Uy5yOZwzBtrmj5ByLsM54Z
RVcbcZ4e5McpI9ZQjhZ+bGysx4Ox8YrIzpD8XHzrE0PcOCxZTv9U0oK0dqgrxLng/tIQc130bP6t
1993i5cHGX6idrTzASon44xxoGECzQgJxrf3FFOBsDG23UZNnLY7D8AZwB6OHm9TEx3QVUG0nQsZ
SvBrKTe2bLI4bhKOmi5qYynDtfvLaeVEoXxiHi+tfHopgHfE7aycyQ6mDcQfuqJbapSVmvJhsiAr
9/SxPWEvDCdR3hAqU9CsoJTeXQDQ4E13Lld5gxjx/59FhKkT9VLp3+oP8tU05nHouwYInoy9Y5RE
ALYlrw+Ud3OqAuFs+KG6ttt6gvoihmvu2JGoQOddcOJIC7o6Sa8C9rQlbKgEHXU9OdgDMnI2lpmw
Ea1lXyNJdPuYQbeMA3iPWj8daNc6TXQTri++ugXSBhfy+8WR41BMGwKhKUq+2aRhmqPMCKfgtRie
5sems0HhwRTftXnlu4/e6YgEHXnvbSk45Bm6hVicD8EVysqUHnoGGZzTQS444qlHpR1VgpBi6dEt
nTfc0+epSc14pCJqOI54qEeGDXUs3yikKCRm2PLawVRL5NGve/zKRgEquTnj7BXrHnw2z6qZu3qQ
SDQ5loyv3TCrPYkC1whsrw1QfODruRYKgp/evk2HUwHPZJ7iVQB7S9Gq3Zgr8fvfBPxN0fdqznJA
fcjz/iutSvBaMidnmEDfFTG25ZLNQJx2T7deG5I7AVB4TMFmLVCjOV5Y1sMf9e6xGJzxeiCnmMMN
iMnBpo1oCNBxX5ufAay+2hvAfB6UhzuySE4De9ibHuD8izBYeFIEglkp0eYUVBohc8iQKBvmuT1e
vr8zWI1jgvcfwrX/UnRv17GAX/xUXvP63Uc2IFT9LTDrWmB5bjW0SsNFtdByNi+H7jvsPwXZKcnP
X1SqKrJtgphAGSkjbzG6KvHA6uXPKuvIbEn52EUuwzl78ZVV5gKXGr+kbT+isvO0nvD9qI76AArO
yF48oJtZGIkbxNBLGsP6cJhcMrq61V4VqCr078MlqsXfpLTg8M2YGhiVZSjU2ms1WorYLHY6K1pS
yeFrt5Au8zdRzb+3IaXjnzle6o5OOtJseK56ZaTqCMjiUddc+PRAmWwp6MHVkwdPz8NOYdYMCFTR
ofWCu3YeczIezDgAkOiqSM6lu9s9U5vh3ilohHVfmFnIXquIQZskczOVjGqaibbU4KIj/vfq6IE+
DvBdioVJJ7mWYcFmKLusRf2+gZJqRQjyi91OC10Uw54FDc5vzagQ2ghPjlTeJ8w4vhAqWPUSfl0G
A02mLOJOAydfWvfpnvXgrMip8+ktVxl36tOj3U9dkhO83opSHX6g38OJgAsSIW0f48HtbAEnEz5v
2WZhvuKJAH1OrxDppSAwSV/xA+8O6Q0tYA53rNbfiMhZTffbtn8KoU0NJ4agk2wuYpNkvpy7BwR6
OS+uD89n/RZDPby/oMRHDDv40AFG/wFBhDWnO2+B6DarAUCdoN0VCy5rKbYkmD2cEqI4O2F9mEle
1F62VaR9T/rNJNjBdpNN5CNSRNME03A7dd0caJQRF5v7iG2ujAzcQ4PEKmw0D7RVraq2fURiIJw7
KPURy4Q8Lhruc31lkyFymWy8MaovSMwUch/YWHuqGJheRfGVXtFyZ9KGRqsqfRoNAfNU+RZ+Wfkk
5XkZq+U9ndHU4q0I+zcMgf5UE7VXnF8yO3+2y3hlT85RRHpx1Il4gx6giXGOirZLCXhWwsZjh525
oVEeh0F5InC5A7rJh2Gt2k0YvS37RAyK49Wyx2nemLThp4SKroblFLKeqbu1IQHBmpg1/gbwKpvZ
GEZGlUUx2kA7NRBTs40b2e6Eddtf/aJ3Aq/Hk6bcJi31K7p2s+4XdYTCystISs6izrX9/AQKtOTu
SU+OR5DFJoiFH3Klz3xtIpRJ6WCfaDXuZ3CvDmBTiUm63RVeZs9i3P1vGf40mHaRiuhixH8O+x2d
Fu133DUu4+WRGn20qYAPlHaRBepn8GBcY7GF9BP3SDEqgzkiu2t9HazbndUlGwk9DKqFAG43AnaD
ybvnk+pk/Cv5QxLQeYvn7QYXMTjakgUtlGsH26It6UmfLV19IUkPMVOCReIU7mvuAajodsJU5QkD
tq6liVWUP4NkfkdK+3IHIMYi+bvPDAhvBr6OtHbSFmsVPesg4AKZR2B2ei7aAGWoukRhkAdg8CBi
I7KV6ew6yXeywVra91EDW2Uz56/1VPtB4Okogww+Cfr/88bZ47JgxN8ca9C24QU3pxhXjAwypGYh
41Ohw48tLXKUB+FdvXjK+CbGt3pkVKpWmVUudYsq8c3SgL5XXmmesH8aWDQ/royc6pxVnbhfKytH
jEGCVfWBeCdYEJN/m35ub59rZNdCJgumyUAyA0ZWlS22mm4v301qwWInmpUjBv2EtfDHhz7GPwCq
NLqdpAst52cp+h4CmH4qX81uQY3h8NIBWkXhh9/LVev8khBoPExhVuGLEAFBofO4MbjISGYVNiZ8
wN/9RYWPS4E8L7FNQ/Db8v3/dsJK8l9pGkoxF9voy4AZiGTypsy6Twuk7hPULfv9KWZ1hhhY3HWj
qViXcALwzYe3vpaX2DFpHL/0Njj5UMqUv8MlTbt1dHSbmfkNPoQ5jtwd4/5x44qy5blgVcUg9EtH
KV2cAE1ophZbRudMNcMMwp/jXMn9yX8WcyBdAmqK9trAJ19eNA3wCPuAZOmwZ0H2fF/8OSsITPoP
6bOnyYvFN6SCYT7BFXUOitjExexCWOEvDYOWo4dqijLAHtQPXcqBqf7vcA9pvs+siCCj5hScFGUK
afOFJgUrBYjJaLUYDiDuuHSkCESK7Xi9mERseL9rD9pS2ZtPDaRRZ6puabc0z5SCBVLPUD11egNT
imCnQ7UPjGAtq6vVE+Z+9kpmlwZTIMfAEDjuucMDYVKW/ilstD57iRqLvRWri5raEUk6WjngFCyk
dbRUKEs/1IrL0Yd09hQMtrcuy+303nUyPUD+GcVk0gkosz02OyvkgCTmx9DUiQNoaM1JU562QOah
dWNUZd34kLXuExQrtljO4gGFftmdrFj0yXCeiWq8v7EhNey8E5mttB6COc8JbYJtJFzDcXwifv9y
fK/wixco4CCOFESbn/rMlOJ9929yl6gfchD3BEYSK8+ETEKEkj0JGkJV9NBhcQk51MfmFBUCemLe
CtAH8b/Us4i39RuR+nUmRT2b1jwkNLW+p0S0hl5yte8uV9L+7sC5UtvcAX6bETIwet6aYJkA+SBs
+nGzTuuy8B4pH1W2sWAh0rrGwbhiCCBu4JxFpq8hJOplDqzcRnb9srSKpTQv8qdwLfZ8tnr3FnSP
tsaNS7g9E+hqjbjVrBMakhzNMYdXLMIWGoJ6Ah3VPNmLmdGXouqusbPPx+yZIVFI6AN8r5Y+ZRjy
/e/8A+WUCOjfGJP7Ozg7YZ6dBbcvhMbw/ROunwL2v/zMW0f2KsRTmGxk6BjIFEFe3LEqP+681tRt
i9oqtkWT5vkl7/oWIXnKMVqX8b+IZos0fWpuZB05IKa8qjfBdELZNRMtW8sntP6rmlyxfaev1b/w
KizoGUrNtiln97SU4ixQktxCTngue7USjT/fXoocrdKxaP8TpidJz0X8LB36RWNwtvk6Xn2x/7DE
JbDg3jbh9gpq6R6g0DwNYZ82in6FDQE/mXWqegAp538zAzYfUf1qoayyLxiUkmMxxVO5Oo0JtYV2
oj08H1FsBQuTC8vPl2bh4iXsxOV3ivyBgpPPeGxBuVwmXoQ9r62MgqeU1bvxkMZ+BsJOP5U0qCUi
CHNDIjl3uB0pCoHOrdAl59x3PviWsGRoy4CK8j2S1ruPwkC2dsS0AfDWgPQZAynewNg8mzNka0lK
oqAXeDpp+6/KO9RSlNdFAPZrNF5C1RrjrmxKNqLFoyHZ/YHEhqBdcM4ol8AQBd09XBS1vnkwuHy4
JYZY7FLSiZ7uvH5xELC90uG4Io9GFZXiZXE6lhxmOWPp3H9/3uFHSYQvihlelkOWGMEX55ySrJF4
9C2vLLqz6qtSabqBf1xOWxHNdQh1hYK9lIbIbLXk6kjl54gfdjeOSzPqIUzWf5gBA87c2rNrBVcL
QW8SjrE9427pPyvrhj73dgusyH8GQ4FQw9ec6cBXDqTLmuneXRVjfv3q4NeGhhR51hJmUiQ028t7
Psv1vE0lpWKEVa78SRA3Ih2aLF6+9/NnlBJcnxyYMCk6bbTXPWIVkT8bBXPBFhDeT1SSCjoXNX5h
e+TzUR+8TKNxKnw7/fyN2rJiodI2wX9YsTttSu3Wrg5oRi9vBy49LeC2kvcpf70F79M3mSgwx5b/
UZEQQjQDhFHrCrDZEKFJB0ROl5SwbaAlsTHup6shnxZ2KCg2/WqaONjH50fLiQffupzL63UrxTBt
BqDmmQZbfNRCz4CjWDmKunQ/dZZNJM1xSqaoIE7A2FbMilkovdZui7yysxKSXOINLghE0UNoNVme
EZUrrLIYFXzIYCk4MSJybNhb/4Osn0LVZh6I6wpiJTV76im+ZKBtGvPzu0EhWrv6iVlIf293OjFz
UAKhEorQMHLRNzpG8pPWq3YA+FPkwR/j5QDHNd8mYqXNULuRjJCpfzXQgTVMnY0BWfxxyzRfLfcm
Ys9XzRmOzjtOQRhCr7XIPlUTkfYr0mcSxqs9vL5p1znDase/LhjSuUJWMJlQsY4rW12znNb9G19T
9eNCXPUFWlAXHuLOER3DDLeLNwwzgFFfce+7oGg7msqvqu2X2xCaK5WMlo+QhMr1vTcMH+TbkPbk
4WV+/bS5c2Fd+5iYzftWal7kbYpDJ8hphg2L1NLFW3Fh1RpIRZjFFu0naHnOSlYZgHH1jQqL0toM
8UxLJZyTq6m1qBkX28qVEZHuawu9oIaRmhueF6bPlWBa6FkzZQ4trjxVpFvevRwPjLpEBn0UDAcM
1LZv85ZK8cixV7CsF1OxFHck12mYnJsrOky8uELBoah6cEoJ3VmRWINCsdQb4pcmMVLqWwaDo6UX
2C39AMj97qdbHiWz/vqlbbi6WqH4HCyj0sQx1ZefEZZdSFHWN5epbqL3DJ4GAyD3l2XBaIdZ3Xch
11O69hkupjKuCxFz5CIdPMuxLOB8l+k4FnE0eL/MOnqFbY38BH+2eWw/E3vQooRp9FnsOLi8g8ot
ZbbSP+aInATAcJFJ2sbKSZeXv/rA22YbjdYVd8hhlZ1i9qt7w/SYSh+qYM4CvGTksWJevYN/zDeZ
CwFkGqq60W3K6NxaUc5gDQ1+FcV6Oeg5M85DQbyd51Btkg+0FnANSyooFhZ6R5YQcpBBdmi2BdtL
7TJlGqrih+KB+z2vOrQmkemMuT2Kie7E+1PrQO80+MdpqSjcBezgJyizcOLU0imgyTn0PSSU4hBo
+YAY6eNIvv9W8V+5N/ZQPlL39bvbYzs7vxWnlmpLTxWtMr5Av7/DZcRz+7oK5KhFArzg+5zVNG/T
A+IyjxnkasAVdlcVG79KeY+Wk+P76LKDeEsGTjTLrbLZ+iwbUkWzSerXYXcwTvRKzzxJZj5eiHzb
t0IRXObuahstoUSdgbR2ZYA1nyAy+onPejBMUj//i1IE5up/M4XnHnmNnDFclUWE4RxGKvEnWbDB
LwdjzXuN9ijDQCRM8YSu2Hth6Y49Q5TCn8oc2cCuIcurrgkIJXn7Matd/fH9h7CGMA4zG4qRBZ7o
KHO4QrnqNNwq4ezN71NwUDzexnOy7QwsJjIrTvKuj0/zBq8rYp5ctRtb6ZxmM8ZbJ1xwl1BnaaSr
kEXmHj/5zR/cY5bEMxH/VeA2u4QBFfmG+OET3OVivNuSpesTPi8xOQ4aNsu1D9PEWNeF9BQQuIce
CaW88eEHrWCutC+dagtrkPMzQDWm8oKMoQx/0A09a7lsyaxN9ffSXKoX3R8S3eil2QOaJQ6EOO+s
8cxVRPl2TveflTU1u2ZdLUgwpgwB7R/z7554uLPA1mG7Eb+cmpL+urxd9KC0PCIBdtPfHgIIe+BD
o4Ur9gE7kP7GxJsTU+cuZ4B1lYe7U7WZP/ePKpfuwD5c0DemoOYrMknaXUzc1Ph6NFd6NGcPgRAJ
1IoFqsq0Bu6Petb4QElEVII0+sfu7gCGR9j6M6g1MtlTla7Ujiz76UEbEThNDHuhkpTYZ8mkbCvD
KNM2c5XPdxuEKrLBCig+T2AYhyriwN59HztwEZZU0jXTIGTAld+9xvl+ty9ExbOrCMdq7nZqGus2
pEcDuvF/b4Ye4U7IYjoqIAbMD+kZTylhobz/WDlZVbIHAAgH7x77P4NNTSKkPWRWohvSY8xqV2I1
azMzdXVZuC8ifZPg9BmLWnyV2O6ezmidxXdxNSmMkG7aSA1v9HIR74GIbQYoOkt6qTSfrNGa5M6f
K/xvf/91b4E4h6+lYZrXlT8add8eXPSBMS+DuRvBjDLdptiJ2ap3DjK8TqnMxUnKFfzph4C9lM1Q
vAxvi8s0e0tR+YwuShVFyzNmCtZeMdDBi0ZUQCc+PxcIXqgZ48x4tfSJO7cHfqbK5tOPKoe7U5ri
yjg7GYK1r6kMXapib2U1/4muA9+zZ7OQ3G5YC3Hyh412FLNI73S8H7mcoXnJA9PxP51lQ3T9m9yX
aF6Ly46N3beClFikSkqSUZW4fNc3QAZe/JVUAJmRS3K7GI+2fReULYWSU3sveU22GKC7o7W5Pbv3
kYLoxLdW6fbPuCqpyCEDHftS6Q27vE1HtmaykYrq2shXL8zcTwWB1kP+tDoDkv7NA/4D9FsxDlgQ
J1DU2FZZYA2J7jhwdM5DBm/9OaEHVnFhiHXjBF265SHt7FyREoMq7fN5SYupv4lM/TiJMcf9H2mI
MQfIj/FH2dcmYuObCwNOBcl+e9dTSGzr/ZI3VEbu11auxzOP4IcvFOnPCbWD9eJC1qPmIVHSkTcI
VkdWDIV6zJYcwSVKhflbfd1N4kQx1oB6pYMxpwS+aQQiYgDYPNrl+/NLN+g3v7PJ15Yx2tABgTgu
0jtfN/mI8Nwi7yatKETzpSfjdSlFAw242SyrYWZwNFaM5jeh3esI0jxmekcA1pVCDa6pmUuXiek4
T/LKNiqOSEMcVqmRV+dzj/CZnNyYWFTdSrC5eB6zDtMQxDchaznGOAtU36gYArqpeMJ2hszIxYFx
i+7BTkGh++ac69ueydJ8Qbv0gTK8b3uoj+MtvNzlulbT+J65AcPeac7kd+uqaL/JfFHOr6Bdpw1m
XBf4I8FI3VMzRFr0zqoEhSpkBtc06u6skkG54h9hVw24Gb1ccoZYvzS81ceJtC+q+tmLK7jtoyBo
6UjHerS8EsOsV1muEVbYuF4tKcYCgKRnU+w0AHQs2HAMwNaKU6Z6ZHLCS2dDnCR1P0OLPpTcBbh1
OrnN4PZjQj2n6CEb9ExX7jlmpngG5LM7XTKeIe5F9BkbLlYVICWXN64C7IB6MF3S/fQDObguXjCL
jhLTyK/ePxbWEp9m7JpG+AX/K+Bd3+tLkLTmKsUL5lpOL3cnAtMi2mPSkt0+FJIDKqCzty3VLVHH
xtdKucZEV2E0lvPbnsKl0aOclCvibaU2vceb535RG89gIFySfF6H7ajW/nVMEFPVggzsWKfmoYvc
njZ82ZfBaTKx+Y38uBXeP7PM3bJanYqnOOgDhs2tAXSTMEkY1BxZVeFNPETGgIFmdjtpHKGaXrGR
OitbQVZlRvqiAQx/XuabzoKKSI+RynKn+WddYxPS6O3U76NGvGTMa2f49xvANMINaDLZJJRHi+zI
yLsG0Y08R2fQrFLkgJR0TioFk/egt7ibKffQQ3mr9uSvlO9AR39V3KtKP46cXN1g5tdLoT3XDHEQ
CyEo94zBv+j0kw0LyUUp8dBgMivVhEOfwi+mAI1dVBJidhu84rVL+2KuboH0eeidbVa2+ezMZj6K
xAxnwRwaN0BLmTWR0JTG8RgQ3NKfi1dD5nvS7vfrUDX3DQzf89klmKMoJTRNhjRYY6bykj8+6VfT
Z6D+Q6a16Ly/gN33eNHHss8GcTj5gMTaTpit2EpPXUyCwT8fdLLZu2gO0OeZpd97bGl1vBLlZtH0
DbQXIIkMw0WMA8UZFZDrJn+HQPEuf5BTc/VU7xyFWYPfkE4cMs5PqOewAdJopYYF7lmJJzHMcoYK
Q6atdb5Bbe49Y5RcjqIqKRaJecIr0ckDzAfmYKyzqSL4kg79eib5/CKnDEld2RlZYUt/TV63MNnh
sp0B89AYYpM2HT9J3Wwm7hOilLzzi1VlcqftOA8K62IqwsqxqBfgjSogw0NRP+GJUtpqJZ5FT0Bh
DtSghLq4gIrUAqfh7+bpYH4UQMEP2+54LS7fT9fygDfgCT7ztu07qNXgASU9cktnFYkIxqx1cc0D
x6affYAR186Y721uC5RaELLuZTbyl0TcqKmnyY+QQnSfWKqTFXsDxxvy48jOBhtqZjJygzhok84b
/Z4mwDbQ8EfBOjfMxwpFAqZgIw06zoRAwrDDRzkiKSEm231CF43+pHeV9sNDtsGHSCWhXlTgnivR
WkGn5tc6Q5AEuqX5gpAgn+6ym2CPNU9vZ8tgqqljou7/c5nALEj435k8mzjT82X02JdK0ma2B3u/
zCfi9TqrzwuN2GvPYPvGs5LuEshuxayEef+m9hJGMf+mWOGo7OOrxmZRy32cl4DYKINWXLJ1gtzj
0kqE2tBEujegL8Y+NK6aZvQL92xJMCSOJBAfB01zwPBFQTX52mnjSKt5rl5XsXUM5QlcggDCdWt/
PfGErVg3BEgtVXhaqnp7JTQYSGKOTHmpGGvt0pMHsaFol2DZIBau0YQlbQc9yv7YcWyXj/PSZ++p
Hw9HrU0bq1LPgFEfsPI3v/OMvHLPuV4k+r+XmnCiZOGkHlOispVW7r4y+Hxd5hnrnhjhu3HKfKcq
vnQhmJtDd9rucnjVYgCChqkyJOFzQnAv0uOrTD8plcC4KiDvYyMJs90Nm5GhxAe7Pyu9i7UzDySM
wIIM5y/Q+j294ObIZdZnZV5zzto0VpUMukFfYJWVfes9HPuD++TPi3njsBLkiBZepY8Fd7teUZBD
NUcSZxdzQKfU3oix0EpBNqLdabuzUptFCl/5ndxRqbHT+H4X6kSxxefn04bnTQ3YXL9rbQoPvmSt
Fe5H93Vrx3u7xdAfRQLiQ753d9ZXUvA22Sn/pqEUT7PLFY8OO6uUPc18eTaTYrWWhICVekl3Nx8V
nOHa7D2MZOEFvHifx2wizwSyq3uCcrAiWkBAlnAbiJMJjYJVOfKCkHSgROF7uPFCYKKz0LKryylT
XFeQ7HjEoJYQVrHsQDK9Gc5VdNMBywji+RGwH4XUwHrxmBmxyfgGVtm7N9DyMFv+6ZerVQI4Wyci
hFmjp3/2/JZ/AJIa6JmTT+mM9vG5f9ybos/nmM1+1CksjUkYdfKx2kw5a1BnG1WnmWQ1FqvpxS5y
xxKjCU0E5c8zOSO06tF8bXk9locqyJglwhloXfSZZygisUWYhDFqDy0AiBFW6tEYBoF1SgErqM3W
ckwGZea2WhtoYBGRzFyUomZ2xhKnxSuJ2pBIUzODQBhmhViT5gjchK3llHOKHAN9PwZ6OJjMOd7C
Hl08vXMBRu+tsDahzXKqiacDa2qUyC4XsGNL2V5vcxghObYcFaRRzLvJ8Eg/Ff+aDCi/JcC+8njx
EV0VRgeY2vpx9fyqQZNq62p8koRR+0iK/FVMlPMhGYxjYv3Rkd0lkGrbRJuyR3RvlckTn8uLewNZ
KK5y60fMTOhwkMq2mdaXT0Hsx31GxCMlmgzuxJM4Fb4SijP9jCEvC0m4wszO2NYeJE2AYbCoEg7N
2/SfWuWgWUjQz+K5FCNPkq0mnynwDm3feR/lqJicZfwwaOVl0XWXRD8CvulwmzE071+x1/tPH22G
EVdMTFxzwzThxe3fgdYzM0LpzGR6UxHmQ51sVVMWcd3c8Fl3SAdlILn1Ee/lZUntWqyW+czqGDrs
sX5xwGHM8I5lTAYTGAdS7L3Dx5RbmcZrVSe9VqcAElNo472b+XeX3l1plGXtkRPwj0E++5FYwKe1
Yiq2qkbT1TF+nuRfVjcjc0sgt9BBG+liNpVUv1sEXpr+5l9/dVN9ztiKhea1GBZ2tQCQgZX/9QU/
5EQ5xgJ+4OkvVtDnRNX6rlosNB6MJcv/mBdmP0p4kmpKX+wSgrbWzVKhGgq9fyDx4BeMO/h7ydFj
DLtZqlhOnYZaeSjo45R0lXfhrz3k7cyffJipAB2ZIa1udVhklV+0+frcJVRPkBmUV18R13twUnQv
BhjLBSM6NxNzPVcervAO/B4JtuORRS0QfLC/ap1YWg4eoNS0jJgTV5SZnqE/v/Py6KQhh+ZI19ef
PPS6qI6yVNnsOhASzwIfBQbK2XdVtarNvAw+INLIsOcZHEp2IVqw+Ekqw9/CbXSr8PfbyAP1BdCP
eRkkksw8Krs110D4/Bcw5ZN6TGJlp24THQPVtjAV3tgbVagvhS+/rfTwYf1NODPXPzRtQA10+Ew4
cL+RcSqZIB0Ta74lxhaJ0F9+0tbuQjRQkynYXtdQK17kx1Cum/1uFtA8mJfTUx1wIYKCne0A786n
i7oZoLcR6G3FYRtcVGOScRpbq4/psgYIitOStbdgyo48wjIbQ+t/Q0l44a1uwsw2kbTH423d/0vk
qOPKVQXViZ7vRse/+GfmYIC7J1f4+XX5PIOY8Tmu7FUH66mxCSVR6lrdBbWICE9ArX3dzQTDx+jx
lyn7Uj06Ssm48LO5W4XZmR30VdXhywI24+w5AICVC8fqpl2Ryj21B7la92WR1YZAFguXhXuDmu0M
bRh4QZASwqxsIPImCoJURYGJSRPbsd2loiNCjty4s/o5ZDsUASR+HJPh4mW50c1dhhGKOU+fFH0+
qbErHs+O6jnrbHYNeEX/OHUAwKy9BT/qwderoFbPOKTg9H0maU1BtSSxDsY1P4dZePufOmETrU4I
dHb6CoH5HboSOamzeQ+ir6xesjRvioxb4AftldL1u3l6D3anWnHhUzxrfHvqhJ0bCOFuaZeJ5Now
uKmt6TRyUe/cOQ/pH5K/6lfqDBYQ0Sm7y5Wpe2QQ2YruBQKGB0AT4X95NMlDpS3bC84Dpbgb8rQk
s3gSFtvAUmm02v41BwqzzMAEUVy+Y8SnRpDpvXN7+cH3jGkYRRwLz3IXNQuDswOZNwqFw877chgH
KO5KFP5VFHtR2lhXHcJrxpMz4MScBrYeZNC33AHv53+5A3m1+DrMgdbSFal2m+pERMOLylyMTO9m
cp+1Y8LhhSqeV56qbD2zKX8s04yuysUCYPWIlxwOxewxS9/3F205NFxLuND7OjnETd/6MxBPJLPI
loJt9A2cqrnZhkrHfz14Hb6pyddsXhW6Bc/dOiCKCMyqfJ8FYnrcR++3PM2+uyMa8fpk9KL2f21V
1wbimPi65FD8//I8qDq3CZZPTs9d7HI28y66zPOhv2fuJRQnP8xX2U580jHk5suMGLKnFsRbWanR
DD04k4vUM3m6bGNU+mLEtPmjGfxNvm2KZGFx3Jam7ol408rojdnYc9UkoqQoJqlxWaGLMkAotc0j
WCsBOebQ+MIzbcXEDFl35D6lcWHa9Ymuh2q314hiTNMMYoQ7VUJTio4jxOOOIGe9Mf7EjNh04DY6
8fLHZCgTaEmkvWJ5Tbh7flSSST0TWwP9gtImZyLdq1wxQxQlRDld00e1dSqRIixHE6mALREz1IbD
Z8/ohPWl9V8gYV0Ofz0ROBjNhy8hfeSL6Rd4zSs1pWI//9H4rRNvY8HG2X4oPrBBubHaBpedGKG4
r5rO2IoV6HvJUxz7mQltFjFz38EWhRDqVGHTKS5nZ0oztDgA/niPU72Hg4LwbRMRLZnLEQHfYBe8
izXBmFpCrwvlgtTSbf0uQKsnyO4NpFueWxLVuW7D4pXZOm40yzuBMDzGHX2/CqyuCf/xMyPmHQ35
rqGVciD41KRJ5AGPLeAIg6PsKuLAwCO0IlAVB0/0KOBCBCrlmGArttsCNVfcQRXVgqwNDjnCCIFj
38aRlOArTnvrqU0J8RKBqr8cCRG1YPBMqGiOcnBYvDf/5TFATLIZR6Z7uue3oE0YQvtrbqAgpbFc
E2rfdpfCU3RKvsqu7qu8CiP//oXzW4I3RDpEC00DFSKCsIkZOPrViBaBdkH9dl8zAAL/MhaFqnRd
gp8S2Y7iisbji0n96ed7WvYB8WDYrmKRwj6KInDrCkdOfEfG8WxpIbMUBpGcMbndnQ511Uq4rlNS
/Kj8vW1kKYqqdUOWeHfccjpHJaWCdFoFFqr8gKf2PL8WAKHVTwo8KQl4mDf3e4kkOlNfsP7QBzkL
60BssovmfAK04rObcazDx3bIN9Je0iTKMVEPzXs2jLeBsujuC5K/ePetNqsisxgaPsXYQEYpOFa6
E64zezWjgTw1fegX1OEaDusw/rnhnZIXcwQnMlZOUsj7JBJdMyk3zntNuyeDtAtlN9vDkuuLXaTs
udBy1tvVGqmoFed461AA+H8uUh5e5DzGha4rOeAo1D1SfpZjpCUePNtwqOmFBTbKHFm1ylkvJu6E
uDdFYKtFLOqNHMSAla9ZC5OdmkNJ6FjyYN2RJaRnLmlRl/oZQn3/Xwo7VjupKeT93yh6BzPAUCiK
dMXPF/1FYDpKM5hippSgcd7ByrTDkrrBcl1QemQsDHN3OCJzoduDbylqOqJB08ioeCQEKo8169hL
fMqA7v4MYRMoun5qQAviuI1yCJsbq9ROkfht1B0ky5OWc6CQuYFxL48KVs4/4vKZOKXqJ12ycAiY
EYxnNP91E9mX8btkZeC54RUD/ZKjQP0kV1Npv17mmO353Gf/+jyZ4BDTUB02/G+/WwqgZv3tRPVc
nFB0mk52aq8/wZCwORWQJCwhqri4pT2P/r65cYu82V3e4nbybD3SPvEgHqAzTE927Tu4fBiKaI71
+hY5zjoHpgbOzNvWdeYP9efqYwMggtiIU4bnWaBDSB66jzTo/Ai6aMsBCE7Ehb7wpQY7mlfjAsKN
J1IXHtlye+wChWnmtAbzJmM2Hm/ITPt7IslGwI67m918V+R0lAWCO0HHyY3/m0QG3fCC4XesQmzJ
sh6B1ANlzDK0UhVw9ES8hE5POhCqwfrNxkJBAyoESCu42GYbjyZcSUvEu3LcoHXZJu02R15lwiXZ
oqNwWDgihbavEmXUTuV4xMIudJLI04JNauDsscK+wmfaC/vkdiTUJrGvF4mpeRmKxBWpvy9Hq2Rp
PfgHYSgS9UScy8w4WvJlAHWr6W+0kyMcoLnlZ//yy/CiDnbDR4sQ2yUlVH6puRuY+L0tXKUzW1ud
FlMirXSLQ3+8ruTFsGYoJb9GQEizFoE3dYZ62nO75YMoJJR8wiIfBk9czILyKAhj0fFpC2MCvhGt
5sP/pLLElNt6YeA3qW2McS8h4mtFQ9YX5xmkQc2ZCBBdOXfMCgmV2kMPUA2Kffb9cboaN5kAR/dn
v9/rD/ULJGX0ZJmkQmaE21Jmd30dnvdUEqIv8yt/0nUx4o3OPkBsRGcSdX6Hf5IwpqKSSYtl4gbr
PSALqy73UmGrGQlp9dmrcx8x/CJGuZhSA4Jj3nr3VWnzRWiVTBXyldDHA+OGTq9TLs5wjOd6Sb2Z
g4M56OhvlrTp2ZI8MMl0sla0Ssnm38PL1pB3CnmcuYWC6Lie403Hl+yJ1lOdftbiC5oUnceFdR2P
N31+olaFlrou5brIK5B1jab1tJPgMEhH+Ycl+bKElxbPo76qzZIvuzpRwXvOqG1VlwjgmBs1M0mL
K01HUQTVXMaya9wDuPtX/Wo+xugJmqtjySKI4syR37KFH8IUtIB/Utsqd7fI0jIHiViHJj3ZGfqo
P7+e/A5UPSAH2FI9l1t9vfqA5wAQQgAukYmdX1jZzpNo8KuzvSpwoiv40HiQrb4+UVh3vmy9iu6V
oMxl0Hf0MkqnDpugbsnvp+mmp1gJO/Nb99Bs/NmJZ9trxHLzdKdstST4RRdyhVvjaCj5ROjEFPXu
pNRZXKVYOBq5Pqo21BcaDHUKUqgbL8Erczbg+XCySqPqx0K7XDfO59Zn7eSaNpkEOBHln65p9eei
1FnLyn1kAqFW+5ZH+UJfWN2ypaz/5VQwRgamXellvvpyHCq/iGE9LVGN0guZopBneosV3qWwin5/
lo7iNMHcQOQy1YZYEp5NzlJs+ogM042hESF8jdDGHaWRfog8P+Alrb42vxTDJk2ebn1amukidHBP
1eqMnnYC1/IV1FVhR0iSZOKPp150nTw/sx3hn1ETg47qyYJnJ+848EPsZwQw03p1sTLpbGV7J9zu
eI+ui77AO10MhQw6aQkN9qzBVaSEqfx9kcTiKSejTYIZPTlF7CqOtCJWGFHCuA4c2rwcLsAPCVEV
NTtgwonJ6R4QE35jiYUz2gnRDIYgWIWZUNwuGtY8Q7a4Z301DM6a9Zyxj/G0FrK5WnXa+ypAgN08
cCn4/iKj0+8QUf3O2CtrpSsUyKlJWDQAtcPp1LRwznl2rRianCNwBGAEljjIIYJ0bvzSeVRMsYXj
qmoMjrqxfp4c4UXPfKxae9m7uCUafUdM8bS/f40pmFWmf1GRty4SuWOr01IoyQqJ0C32QJk4Bgq/
bQtrYTBqfbr25yEJXdFky3T3GFxx97+Ni0yVCqb+Fl/ZE64WW3/ThfIyEqZ1hwa9nkY3ycldDEBE
TF2lAM3fRUNW2bUGPh7+PCRpMrC3uqRbikwcvbp9qEFOsAo5WXzgqtAUFtrzXzvYmlAGaX2b53XY
7Lrspk/c2DG8tU73ohDTz4JuLIdZZ6XT1GX81nnSmsz/E49y8MCU9vZ1axrLolKQnBKalVRlK420
AMMfGdAivyUp+gzGI/jONljWoez7S86wVxJCQYIzhIqoFDQHjseEH6ydTEjv8dhKhmnA0F6C/1QG
7CH00uj7GzWuKOngzzJggPOx2sYEmpCtikE8KvYpE8fnW6e6qNo2CMuWtTyztnFQRxgzJEKyIVoN
/Rj1kqXzukUpFggbY4G/VRT8Tp2wXuKRDNNuId0OYAr3QW+xsgG+cMU3SEmhqzKkQeGLyoxonxry
xmYcovoJT4LthNBRxOgio6JsrvH70HcPtp8NJGrPamYe0AoqGmeO6y27i8uk7L2u+EUNfJ6sLHbt
6ucElSdfwB1xSwXNRb0wZMgSZ6rdJdKsrR5onrAedQxzQaLvC+D8cGUNucrZkcbAWaUNL5UgkWlN
hqGhDl2BwCv6lhbIfrgArWsGMtcJSsrfJ2QgKNMSE4SdQMchCYlfmkl1J6n9Yl4a00lhALfbnByD
PWYOxDFpgc6TPFRInjDn16zYs4SZYGzJfYLzFM7+SUSEB6Ku94cmiEMDl9e+cfpK5kmELeYNux3a
qUxun8xO2VgkJpdQpeNrXlOVRZfv3B9xdVuY9ldneerp3TdPmA7rIkTkqB8gCl+Uc35yRU1M3fdh
X2gPLOp+ZOrRUaf5fkjNvY1P5P5mCCdZ0vKvhv3Go3MiIzvBmzx7XUmYHBN5UM0CsII4lrnF0PW5
UtC/8wB0JWCWuvICduplKX4Nm2H7OeZXlvgWvUbEMI0xsJiwcNMExKD4qHXN/I5B+LH6T2RZMpLV
qazTbecjnJNEE51LH+JIj52FJTygL57ycDs4a7eP4h9QhBTBP9vpot+Kfj+Yoqq4+/k2lIuMF7bV
wh6J0iSKUG2/PGZAcrKZnh4tuNERXS/Z2eu7XEgyC53H3WQaEReQgV9MzcFNqhzBBDexdAfI+8vl
HRDfOZmGdJfyyfe3NzIkzmq4IcDDhDmPOK0AUngciIGlDxNzp2cHw09tr7wDaxV4X7w8CU+5BqaM
0KoKNJyH69h1gSuvTza2gkrbjL9AFDtmnN6uCFIW2VaGtUHA1/wuJ3bIFmU8aL55iKiy+s0zHOOT
lEeKytTvl6FWNKpIZ0GtjkIkTpUnIfihAmNqfUwj3Eqvfp8FhHyrpny4mAMtIygXkXYV6BRiyYPd
qHiS3wnh7FYfvKbZeqWNuNbgrVZWMyBiOuyDyoGjgWGroSclYXYSllN+VpsgE3N4CdETuDFs138r
w+evaRnj98mIXD8kcdydLeMbFERAoBbnFdiQEGuKZCpQH1dMIQ/uN09Bw6VoHIvncjq1PPofRp1i
ixEfb+lrp1dlocZlsqf69ithRpaN/p9jdxSZUhJHcnE5RhZG3KhpuPK8rLZPilRzNK+Us4qvLaNa
KvXKFM9n7gbcBAd0tE6X9SdjROCieTNRj5FACHGdhiW1oyIanVvHmP2HQEiLm5rB2/mFQLSFmcpR
WFkTGEcHy7zHCxlcrtqGbb5p5YtCYCY03wQDxHuLJrLvrDnPsg8OnzXnzek78m+8pU0vtE8c9h7c
ceYFD4khJlES01yS507pIedE23rNOennHI+UoAxmdsyGdTkhCUlHb7D9MTZWWvaHxX55k12A1xIo
4igb6qPeEGbmff8yw7O6+Is4qN4vOlij2k8i1ZwgUXiSj0xYbrxnCL3Jpac12ua64xsivLiK5qPr
ROsv37Mcm9PFExSCvWK2gkhXq3i3tgWJXq2GyfJDcIjAYS8RHNrwzx657vRl+9Do2MYXDDtXasAc
CKeKkR2Lfbt/8ejvgxmrxamVex0JvkQeDLY+IedCAool9YBtkaiJm3B628WVMYxTbifOpf6uPzPi
1uc6lvLCFHYtECNIgbsafLd8s/52IwaE6K3O2DZRmkt0CrVxHHVLa2RNH+Nt0btxhwwCr090dgpH
ShOfebH3ONThAW3OlFq398rZw8BlwEKmiNYpA+NL25w0XaSBqPEL6/tNYGEZijDoBwGBDP3dBuUO
D3Ln6l/W2IgC9PZk+1e1slQgoKLBdT02UEsCrA0S9ln1SajNBqSXbdBRGjHuJ2WnWSmQ25YvK6k6
EmY/sWi9rirw6AdasguRzFRI1/VZ+RAzg9nv846bD/0WhSb4kbgpI3XtRAmJOghlBap8G+4TS7wM
Q54/eWo+y+HQfY3UJDs3BqMljc8nJPQExmJowuq+GdgyAhqulUOQ3uaX1UVIcRA1gUzUYkEKC6DV
/oc2i7tg3wnG08uET2P8P8io1R3LmqwXoJ7aR8FkEQ5aVs7e9O0oZ2kAbaN0/qZfDx6zFQk6MIXN
aoyqCwd9L9PYmUGB8LXzIrXNy17B2HKjPI8LFz+Hgx4vJDzQmtRh2GlpMfmuVLv2SDiFwHYMhnGS
NeVbm13tMECTISBZYGkTppikokeZQAedizZ+M+8SdKLeAEgjfW38kwS5DEfielcJ4yc3KD5fDPZV
4wYDrZu9nPLGFBDifebMTyAjv2w1yS9JMvQoAjC5sQ6RFW+cj53EL8tcTfmMY3lBYV7Bs68SY6R+
H3+DYquap1qFFgSdkSYHD1C8M205cBLE5bcPL+rWiMuG+CGUZZzukbY7eAsq9YjyyJ0hG0fHJ+/A
ibxA7dzuNAyS4sqnO31YwrrTV6YX7g3Xr6POuilx9YS/r3f96jjThyz82711H0DECb8R5MIJWVvB
08cE0epE4jS1+SiEekyOMzLmMUwskalfS+OmZuS95wXivERreiJfw/CgFK7x9xJcS7KxsA4HCq1Z
FQO6EPvsVr0JFwYZxMJZTCPCYWITShnBPu/hxXr9hxzK5Pr1vR6aaHH8CF44AeTWkQtDY5TDmzZG
8oxWOwkFqpnADeooEj8gJ6/Hdg/X5YA6CilZdMHGmTD0ZFrKsdoCKqDdqCftc4eB35/ZrGlLI/i/
PpM4fU/UjzzrPuglT0Aw/2W2ocJ3DNRJIPOHLkDbD3y2VNdqPQw7bbWrZD9h7IpkoZaVf3jiFD5a
fBqZ2c3xwyPeJIYifJFqzlea4YkARaixc2RbFIVR3QV9QXLV1Rrjmx8BU013We46KKS+IqM3v0dY
IhzUockUJddSVYvzfWVE+aYHUXsrlVbnUdtMrZERZBCwI5pVSy46i4Wwwi4HtKkD7xEX7a7AW4uP
YZXy0qqaDYUviDOnfMSBLJGnITxpsQ/R2Pbhh8vT0zGEopEgLfMr9/PD/e0yHKhqIDQDxKs5eC4k
5dF/OjC2p9Vz1g6UTl1SeavSobybnezsHDszOMRvCAvIDz9zC8bjq1d7PFk8VuTS5HXuBJUETBaA
+ZdKpy3hmy8twk7OF91ZZAx57ygeljLPbjYf1OFI4LQlTUPVQrh4p19Cgwivdy2wTf5f1A/j6tPX
ylk6e/FPHS++admI9hbHwHciwMCoZeK0hWnhF5ho1MTkpSUuPgcwxCGRxoDPwx9Kt331Qs+Mtz3E
8nMy3w65Nsx3kPnjpP/lgZTxTX7C4wBbWKRpiS62v5U2s5dX0mu6SedqDJBFZEJgfdevX924yCYX
5oYW1TFwM1Ho5n2e1sNFExcTPnJzgNFMKbHTM6SB2W3bXVJJbcUjhVIfXxKrxEzCgOhHV6N3bvYs
cV8Xf0huFcfYIw9WrxrvFtCggvgCltcfBy1gnfxgN6xxAPnfoyrrH5OhKCHHsRhLqxbp0EqaEiX9
yoJT4L67KGBc6gM2XTHy6L+wfvV6OQ9axrnIak4DqyUWEavTDANndcc0kxLpdN8eeSo58Zzj4nu+
/CxntGasGieEsuJAYuCcGVfBiDbnpbKs7j/Ps9QqIhGceX2GQIQYgDMlK94T2rq531BC2Kd81bqD
URu0HVmbEdC5FcJGZFjjIa/TUowiuQUdhvFhR3xsE2JVw5bhaT1KAHfpHIkg0aSGpqV0yK31jzr2
a9e30eLOZFmzxyD0Ub2qV4/fEKWi1oJRHWr7iQya0IqorCgVTzTIXWKc6IfHLnj+f6rHJiZh/hTz
LdM4g3S67RQ9MauEehqRo8XjUjPF2JsjFAO3H5A/Esm7pNWk9UnQGoKTGbuK4tzxCSiqA9dtRTDC
WsEZNSP8Vr+XugIWS0smKY+ac0Ko6xJAJZ39gu26BKpVV/M6cG+hz9PY46zW9sSLaZCkbj7ayVpn
t1hvGXoHpNS+yFmwvdzjXueSEPp8LajSibkjblMtzSDxMnKFbLic4z0Rg3Dm3o10yQqWzQegTK0l
DWJ+FY/jw6gUMWmvNKw01fEAvkc4v6YyD7NIKPY1hMLcoZ5GUjIyq4naHSSaMI0B7sMMaD7IK9WU
MrGeF4eba95bRrqKo04yIYAClTRdq81a5GBrxp903VJe2W7/TO2f0qZ3D5tpcxa2+WTplnPRYiOQ
IV2U16/5uXPOmFw0DS3tju4wjXFV0iZES5IpwUpnmvYWUPnjj0YAERQRb3C1HjB63pay/dYCtInV
831I/LItwcaZYtQ/Iz4dqwmAIPEAe0+VCiWa6hZ6yD3P4pUxglfbdfCyPiwx/YMKkuqg2CK9zGwt
DJ4vsuG2vIbd0tUP5kgaC+DpJ68dfv56OiSqfJ+jYuqfvwKAKwc5qr3z9E42PwCf0/KU8rqjzTRL
tgCVA8JIWbSEUbIjNwNKcWn6vQn03sYOkYNLvRIMn0jpa8XdhBQZcKLgYT8f3Hu1i0XZLykyOXfa
84WnlGMNjh4OkDuLxoaDokq+W8Rl6tM/m0iobybyronunw5qkRJIt0hmh/eFkymxJ7LKKkPKZ6D3
Jj3V4q/3XT2yoMsZTSWZTm5c/tK6CN7hq1h2UghiHdfgoOOZop7UWnINf1RzOAoqAxMtg7AzQyLo
WYBdbhS2Lz60pQzHH4tVZWoH1XTObpAB+1dyeefN2ANy8QcPyIVV6a72pjsxTIAYj1J6MAshLIjn
VSTVJFoBgimxbvV+BfXUj2s7GXpzMoBIrkNxnYRE8M6ihWlLCDpd6+ek77dDv1WI6LA8gO9Y+77M
4F+jKYmLcifPZ4WCanXaOOqsWFungDg8pFDneTI4gg0v/f8i9cWkpl1ZpvzZH8ePtcH0MR+7GTXp
o5OZAcL2/NFtHNaFaRxOMto8yTDlxHFUocDkUucaZ0La+0Q7GQoAuJT/W5DmBQWyix1ij9cMC28O
4ZvXkxPAkAei4/3r9LzgJODv8TFUGtFGG7gRfwqbsUUBc4f7K1YPVTRZWDqRU0rdwS2PVrfPIs6M
oTkxv8AgSuZhThSpjhrPmZG/lRKOsbhzRUz5rFEdkCrIZZUeiaqe1kg2fApd9D4m8G6YaX1Dhz+P
jgsz45U9Jxb8mLpDGRe/t5slZtrpYi1+FGuPa6cCx+RngqsoeSD42jVxqo/MLu4M/6Z6A/zwZwda
TFLZcTZi0SrSl7IHOrFJ4c8SpcjqhhPwkZnJnLROWRu+1JrzVNKs46sI3rBg+kQHMEf22fQYh/Ng
rfJBMQqiYPBYvktpw8tx1mxwQ8xWy60vR4ixG62mw6ailluzjWQYmzCZXUdf6lB1ygQQtlfmOaQS
NOrek1hGaqrXAh0dBwE7j8X5qddDP7RwfZYHOHoaEzcXNAbkOoCCXuw5LxGbC9OqJcTgqaEF1GbN
Iw9A8mcczaVY6Z5fUy9F88fEYy8MBwp92W3pWRQKygUS4WErytDH1PgEsyWod5M36PYAZmNsbfc1
PJZHEEyKxc6hBOR4gg1jULSJ9cdQZHPuaYuD/W26PagC9ta9sAB3LOO1C+aUvHINmDzYMzRKRdTU
QSh9LTz8b0r6Z01QEcfWmT6ChWhJIUetUenfkHjMsuAV4lD2MmuYGOoNVeMqUAMesB+W7CYeKpgj
uXFWF0s5m76fiRM2ey9PYHE1qVMtrpP3g82GPYJYeucLFVcXA3Fg2+nE1ngbDOOxPqucVUEK6paX
4Vnx9jCllMg21UTQ+uUYzLnmJwEDHcYrGswhyFQYEIyp5vEZgJS0K7PeipBhrK949SPmp+Nzw+DI
ibzxj5Ehad4j6m+WM1622rftFGxN8s5QDDJGYHXYKTn/B9HrWX0EI0ZGvP8i02bpZO6ItFt2c+bR
ueiohuWIFb4pFZunZsPaiGnbA1Q7l+mxX4dFh6P4fR9YX1nt9W9I1VYnmVN2hu7bbMcUCiZaU5G3
19FrybZoFVK8kbdWJixO4am+KujQtHXSMHtx2fLmKN/xoss64g1okGidv4KFmOgrTK34PdM+1e/Z
1MGN5Kn0hqlu3Pl1HINx3VPnNMQBwAAUAwmZ0JKzCP3z3zdx941Z1Wtd882o8dGrBvZUFRJhvMPP
63T+Y80ERNpBl4oD4OaDkwqb5UxAtaN006goZxp+MgbsWKx2yA4Guyl0hj9wP0nF/07a1kdE7h2T
kfmuVfZpLhZLyqebU4KHEnDMUZsw6HSpdaFMS2dBBK4rAg//azddD/HQaYXBDiZtC21+r8+Kadw/
oYuvLwa5+2eTqQcpl0ZHVe/tl+N/aBfIr6UVuEMJCQ/iwxcL64rXeeX+JznChZfh0L9yZ67yaHwE
JRY+dItnC/sBvEP4bbwbYxiEvXLhz5gdLVv/mhq27m/dv1IjbriG+RulXouEX6vyA8uSxpOir87i
xsQvMFibtTNU77YJUxa+DkVPFOQJKGwXQXWa+EcGX3G0V/fGC962bjP+GGaCupU4klFIJm+0cOab
AEYlyKJKgdSAhr5zXvi1l7mtrHhBNtHyrqmgsJX8cGiVhHU7vjLMl1+iZ27KKi4h9Fyv1C9LWomx
sN7NCoNLs5W1OlwcLmZcAmH/KcHvw8WeU88VS4nGZcsC0UwiCS/qdiOojlzJdknpTIkKNUivUXSJ
vUkYiMsILstEd+5NIstArCSySBCeiPQd7Aka8ALp3R3tRJG2EfzVBoieyb/g+XYK5Byvz1EYRH1g
BE/UHYCVlWhGR/+YsVxRn/T/Oj8gtgYbzHXeLqCqGw6xZ4PmwAEFqiTi9PqgPnhcedcwe1NTfqI/
m0DAVBijI5KZgIST896aHOTvayIvUj7v7CBBeJduWb47fGVWtEsNGUcg/YfQgxA6ZV1ve6NdF1x0
3k0PadDnHz8Ien6GrtFItjOS09cTGyiDDA4qf7g3jURLeZrT5fPwlamYwKxSRRSMoTfSpT88ivnm
brNz+/ZWPP/CcCFDfj24YoYK8VIO+s9f8zd5FRVqKycjMSmK4G5Z2YnKdic/83OV5eCd01q/9Ihm
q2VC91iBc3XWhVZiQyE5MNkSUj6ZaKJnzdTW4pvRt4lQddEBUnw6PealJMU70wX4LhNodKou2t5/
f8OcWdILoeY43mwqZK+axdSxCqkIvuXran/2fmCVa9PR5EDEewdxTG2ayh6929ZMW4TgsTqSi2vn
WTKZMKKNSbHZsEptNHCHsWflDgo8d5fkRbFQRnb3EBxJrWh+6/v/PGRTYZIJg5gXKDJA/GBacqSA
TThUpDlzqssVBWhRPC5b4N76bKTQRlkXo0nHGUY0/mTA785g+bIGV6oH4GtBcmbA/26HLajjUJBS
ECEj25bavImxc8rESMr1ULsmN91pCOVSpCBuNtHSI7FaYkT3nQKXIs37/wF0vxaUZA9PNZlyYIXl
82d9w1KAMNGKLla7CHbo7TBRQ+T8X59PYMHcOTE8gvy3cTws3bH2O2Mqz6TrLsaIpaao6qfup3AM
pzgqol1S68y78De8P2Cc1eFsmp5yzdORPH5955iY5Msb14+W+oCxC25uf7uN3dLOEBYHec6fUri9
Aqu2X7GlB8x6RzfPe8ien+LC2QYIP+thzX7PeTYNChhP4BNuesAZg28GCevvdH7x66Bo83f5kqyZ
5CMzzTe008GL+k6qftKUpJ3Vytn0M3bvYKCEzBJ1TJLhiVCwsjzwcgvBPWwF3Hk0VyWO9SX0k4KZ
K0LZwpN5MogWoE2FKrcgWq5ErQOm5UrNyGHBBnD8aORSIbP7fRQb5v7PukIaCZ4YpBgk//XEMjk9
zLAWIB2SziDvb5Jk26fyhKFY3Tmivu99Oat7BX7qj27sp1NKoo3neDXiyRNYMyL3zPa44HiAfJ28
brq/pcopz8xI7D1lPM6tYyKuuWMvkMdYYSrUl0jfKUUjggfM2IWeSzwaeCh+wLM5wE6IO5oXHpvX
rr58CQqMM3W9Cm0dFdRoH9OG4ho1jSJqkMRD1ugFssFIhHcj3+S7OG2zP8ArF9JyZS5E1QcnNZW1
5NrM7hqRHwpeJ5Sjb9a08bGiT3o+sbNGTsfYarWWDUnRkDTYdgzF2FmBAc+mzJ82CHnEpBpYEYfH
s2dwTikpaQqjzNv6eqKBkTaMhcUfbGuM3aXSdrqrmDzVMff1a89OZAY500Aggb3QBHM5MFR9Vpsg
4UiU35B5FW7Mrir3kelJi6nWjgHluohOWuNsXcv2FkdAc9hR4sH8WGeMiHDIZ6epwiNtz25tyGTm
sGK94Ea72QM3O3PiJTtP75BG//0JREZ+X0Bn/fF4KWkVOd4XMkD3rj4i+hDJqMClGA1zR/yiI4SJ
Y/9hN5OjrfxFmQzqxIGDo/mE0qy616tSwwIGvdSt2z+AR3WTmIgqWe1VpHGIZe66SAeiYWEhMmCV
wNlpdUntICojQQrBkpf/PQ0l645SXsrMBF/lNcMyHG/gpNFU+pKlW1gk1nSpzrnXgNZ5SXq6hz6e
2g/txzlOkbwdwmHFvXcFOA1zPRPu4NS3Wax6e2/TB3HG/+WfHCKGPrgI7k22q2myIb+cujrH2vSj
mN5ID6Lqj42dAeDRH0RGCGK40Ufc2+cexL+CkJE74WvZ/2NZoIXPc459ITIH9AKRKg+FzAfAvD5b
i777pXpS7SKkznRUKL0hHggFQQrZX0uydBsUtj3Ijhic0J1AojaoA/2pHgRRRQGYfu9DeUQ84nVA
ccD+OcfLLyrZqtRgENFZSvK+Ze8Un1ly6/m5XaupB8AZnn0h+FlpQJZSoWEbBgs3woKIfnPeYmVo
40xlYsSSToZQKyiWVuuwosi5PUagXDC7w0eD0qEUFI8k7PyfPNr1X3ciwGy+kz7Oj4XkZCBE55U4
u0NsbC3c4Fp0zqOqMB6YPuILHyNuIpKLZRKS8dVob5r++X5IiiHABgpws7IGayEZTfHfaphOPKU4
OSC5N6rhu+Kw+SWe5XDg+CaKypb4nImzOqnO/14aFHlmlazv49Bt8A7pWcropZtS9mVbkREMPICV
KNCIkGq1JDsDfhmJrGl2nf70ndzSWqbkScWiyxCYUm9ocEoe0fv8pGr+XKoVDpgB+qF5UeNHj79e
L+wEUzY7ffeOYgbWyFbDy/H6UWBsAD4UEFidK9HQib+WV1AaRh7f898FiG4VtwPSkm+3/ngHcack
62eInLR19PdA7TsSjieIeV4/LZM+o+YB/0fW94hv9A1FvlJIIB5aflv65sdHJ28SIdHZfGkeCxfp
sEu+1tRoOGaSk1Giktso5BgtoU0tcLAHGTeEZ86V1zIeAkaFrrlxYhNAvfI9xdmffYmlfhCRnnLc
SKoOQ/4nEgPmkSF+NUY47uzeWVHGfUT4QDeM13d0w+AhepL6gB1hcvkeSi/Fu5YYwWEhjDsh2oth
nw2xKgLwwR7legOjHDSKiIbmUZ6ikjRyY/fD/8b5NO+IFoaBlKn3gWrUxxixUqcw2dC1V9dzWV2c
+v4wkjRXO9bqeRewvOoxavwAHJsAsGPjkJN/UWz3bHLKCnlF2JdSGESyL+MkzQuuX2Ajxhqrb2s+
Fi/wOrjj65LjkJ10sY4th6Z7F5xm7ykLaRz9h5FYs/XboThPs6nV88wmwBsXv7v7O2Zb5aqKzsKQ
imPlujyEOUXDzhRzT4YgLxAOLheDwEJaqQTPgNHYNQZZ2gy0Zz38jzzjQvnplawWhi/b8UCs0fY1
yQQzNXOYzk5IOhCeLDTzm6iBu6hgrBeW0LtcGC6ynG2baudVF6pGSL1w4VSvmUg+v9I3xxBsJIux
w39UtaZ9QgeNwdBaAKkrRdCkb8g8o2WnfuJ8jJj20UinUY8EVuImoOggWIO7nEPUM/5ApzTEpG5D
bZRMXKH9J6GnZmrfYw6ECJslHz3IOK+cW/fpiHBCrDWoZMyH0EWueXSeJ0lMy+47f7tm3oPinGrx
dGdGgb//L91spF+iWA1JWsuL6y18W4UpRUiokgm+oeOAPIhiY42ibn6DtyrR0xoNTYYBnh+crGev
KqiJQRoz3cm1tCwjhRvtdrSHZIROL0nPfhkKZIV5FFK2RTvnUs2Y0jhluJ6Y4KQAQcxhTr2L5VqT
oae0TqEATRB4aXWijinfY3KC7AqPTkD5ysbcShPU5g1cu7W5QsWaUnOiupuEp1ocH3iZBBZs/XKc
YzBhfcWJEudUA7BH1F0SClEwxf5aKR2Ahe7iUhYBh027ypCbz1ivD+lC1Bf+gPK1i+/8Pzx5Kmwa
hwapD7/C+ohuUoIRr6B2u01+8xEi40yTRD8Yl8/ivbPh1pbvZfaCIIlIdxK2lw6dFO9ua+06azcT
5Zgvq167XfAmLpxzn/mgnrydmkaxnxVdNJMkL8B3LUlWsudWu9b6RqKictDLWHcbjJPcqc+4MFqZ
Tj2aajyhceH27IqtG6aG944WfXDvXs18oeyul/h701A5Jb9TmhOqqDp/noZk453axaUg0xxlpRwW
qx8MFrKWFl2Dt0QZHJtXkwjbwcFikJq7lQ98WKe7h2ZeSO37tZO2SObPUGEP54DrQIvetOyU7Dvo
CnymAiyOQEmtgMM+jLeP1aoGcbDpggi6PgWySzQUKy8S/gq+gzW37U/R1lep0GMI1PNMYCh/lVL9
oRjbHDrADRAAUIiJ84CIRIVpbnYp8QcqnSpCNoQjLMVYGzC9hoDSku8Bs2zoNiJh7S5E6Ff1uiGF
UYy4frZ8CMjqbiVaFkfGueWsNwBbkLyEswg7jW86qWiaBguB0oerpPCWRp3IWZfmaZ25fvC6zVyh
SLsoJvQz1owmAVq+QqBIgLQk/qkSlMNT3JyAt2Ve8D2p4diZ8W97io3cd+QvQPQ0IIL3Q2iUNUor
XFwA8UZTdGCXpbhPfMKwfFjFNa5hdUiBxpMJSByUabbHnxzujcqopI02v8b/3n0UbhSoXGO9iEuT
lNQl1PW5SQ+Us7+zN7M6zW0I+GKC5JNCt82Ij0QA0UP4kHULT7tO5os2F9Q2/+MY5XLr2nSph2+I
pPR37UsIddjK6relKNXTFPYNYNoHA/SyTFDu9SqL2CVAp1vjvG7KgorB00oDvJQzNegrdnHu6d1a
eUa/aFGb7phAW9J4dOq27VTExS6Xy3dbM1HJmWOKl4pIwCC/hJc0Ar02ZirFFp1+1k1QvgjiQlZ8
eGtF10ugPgbaSc8V5OcTVO4DV3rdDDrSdv53Qd9ovslRpJq0Wq/Es4hNsBz1xk1yJm+tYUWFMslZ
42WSz8s4J4JtJTLKsCIZRRbjSDCVDveR0dhfM/UGYlgZTwApCQB4aQcuzeXd2ChXFlXNV5wZkdnT
4jjOPokNdMOKFNupEWD0fsNocfaGqPh+Y06tb/4+lOhAn/BwyDKiDKv70BWMthfBFPzRvioWoyj2
zFp93kdFVnJcKEcD7PIf/o1rpRIQ+1Ha/ODfGz9ZM0adtaiepGkURXeDveNhUZyja4FLtAUi0C+w
cpNqeQWb6WZQfYZ/klaM7H0CJMIpkLmtPiyMnt1frhFLt9udqmmU4itTx8uvCGWPJK5+Z3s46Qwo
j7stJGFs5LTzs0b1KKNUf087ujKbQfrScDRSUWtLn0oqF4RPmWEQx22J3H/QxXzRDyc4FEIICEsf
OP5fitTdFKVCFofNXBERRHy6PsS/7ARjxcco0BK1XJDYVdFiaQUdDGcvE1EqSv+abiQls/IGnf+d
FKzfUNuF3sk1ilVJw9xeDemcEvekCqaoaXLrMwVyLVHw6hNlTIPr+QL0v0401Hs8Bed9/PEYBh8w
Vbol5S/WJr5OBTRI4CW1cA2lcbX4sHK1z0pAqRv8WqHuzcdMVvkcMoNw5MgtwvO7DBsamaZmYOll
erRHJrAvvyj4KgAKQUdSSH3+5wxYzFexorGbkQhKA2GS4Vp6o7we+7HM1fY8vYdhDY4Z7sxX1fLm
bgruP+S0QZqhFzQQWZuwAJ0FVsyJj5MATNRkp8D2JGwZ3xjLtGwi4AhYEtm3smJHAd4/A3YrqVtE
OjFwEWgRbktTJO/Cj4IjhOe1TowHkhUduroYMMd6oEFPnzgKZ+88NMyXuCO5HE07Wizb9D20il87
7L75DdmPnlDMaKOlSThN8t5o+wvM9OADixOPJNgjdwssr285yv+E5SlpJCI48hY/mO5KcQ9E611b
kzh/iH7OmkbBPqJntpZAkbs/rjxf+r0B+Pk20sHSs4i0D7Mfe4iYdT3HM6nNruojKxdvkPd8J3kQ
Yd5coUdcykqxWKBuWGcmZUKY+Z0T1fEUq4El9jozNiVe6Nk76VsX7EcxuDqtevC/5UxJPgUuX7h2
gY4gEQ5HhBY5JWnr1DlEGVJ70d2Hhzs/SGxQN7reudG4vbuG3StxmijaNu6TYXM7pUwWcGsW/nTh
ETDQWwhcj5jkY0pjn9n/B+BVPGRdeLf+z2GWL1UQLbAJcdpmmpUDXyUK2pXCbNDbb7JvX9Rbl5DP
3pyE6WuuAtX2LiJjAAagXnzRGg9mel3UAVkmPPIkSt32s5b2WA3MYppjvCd9Ghoqz1xttBTHwGdF
wJFVOnSMD+qZweviaVwaqtRoT+yu9Vl3D7y8ZzGUiM1+6b6lS9DpiBDDZLOUtcd/G26Me156EBQX
dlwZfwMUAel5JI7FswJO0TIlXDWtSczpbETJ8f3uIxfBC3cGSt+6CJAWdaV1mAuF/9hgfgVSUnLa
2XA8KKLtT8V5LAnGowkULBU1OkKh/wSWUnD3yNJoU4lnPJPp78OlhsEpoKT08chIOtx3B5fh/8fU
CwBaAOKxudw1npCE7tnQB7SYHc473ZdqpFS2+UHjCHhc8Pff0FU75FdVf+NVobS2jiYtSom9ZaMd
Iibge3l9TA931Onr2qAbT+NEjKOXV3PhdspdgsQs66/xJOjwvgte3uoE80qQu2h9pJHX2v6JkmI8
kWDucxnjIcVA23k1uFTuapSqvsXrDDPujivyQGCEk8lrWsDtYMQZQ1QWifkK/pmQu8bbF6rmSHiQ
riGQP6WzjHO2EMewiaaAgr1GuJM4fHybyf10PmJl5AlNyZMQ6n6VK8plxG77TpktDC8xunmGdhQc
D2/sou9vCg+hpnvr+pUpVneEgKDrq74vKS9vDsCMkFvTF78MnMpTyhTyJEJ0jTpc13Cul0ir4S+4
wUbwXdU4ca1P/qFFn0xsIgs8n3Jo47pRPqXpvmwmOwD29bXolQqDJC8WlhxGV8jJGhJUHYfwXJkk
k5Y0aoGMUnzc4DMmey8CmyziBZJDjJ4DmrglScnDvQ+ehURFpZign5ZtNbC/gsZCojI2ByFgxxwc
hmIc4SqgpcrwQ4oM7/2OqzaImkhTIimBCjYFphLKdhN+JE0graB6CFz3zrc4MASrCcuwr9ITZBQK
aHXUm/TQUHXXFt3wY0aWrLLBp8sI6GKm+P3UeVdDgH21mD+mc4MAR3+O15IIg5v/irS4NA/Ro3qq
OxsqDaVkhZEyLFcevSBOdzSoJw0bV07ef9jPKQ+idiCM/G120Xquhj43lPb1gzcnP7DjduF9MsqZ
ggg8Z5NW+GUk4UwxEgM3zgfyFP//pZtF2cYIusS6i5cuSsqLpRAbBjlJgiNzC1GSsjrXMLsYWs4G
s31z1CJ6iIABNN369DDty/Dy8IGuHTtIRU0BpCCQLAqHjBfn2aWTHb4pl5nKONJX5bdaxed1P7N4
6x3Yexgu8GEfpHpjFKXE0ppFbav84wTCtcyqRvuN6ygQczjTn1v6L/FQtYVxiH9tjph+zXpXt6Cg
VgTo5MYiWz111XGawsIBTaVzKKgQQAC0tDbAgSvtCHCUeBlxE5myFzZEVvX3k/d0ZROSybyMUaJ+
B+ProMIFFjh53HTh5Y4TWTtHDnXPSLzTI6KWt5HNMjYvRSPV82C0rdBvgbCbMn5dbRQrJ/JgCaNF
cBAEOnlwE6gGZdNyLOMJIc6AKP662b1nxvE8IMhlevqgW44vaWhBXLiW4BMxxLu+CiTSYJ5PgDW7
SEC/O7l9DIcXvZ3DW2WkPoHEJKs3QarPVjX58ghLAWeMQY0rHwwB/4f7B3j3NWo0tpQro8LzlqaV
z13/Wa+grN2mN6hCfDdpxEtLIDpWLGUpiuYcAp7QaGnrwdoFU0UhqFuhU2eOjCh1j1ZUcqvlKKdX
+uPMb/0AbiXlG6FE/ViJUxp2VLCz2TZckr/oKG0/eKAlGDyP7+RLWRv4RtIQOXG+wL/8yEF3CSr9
7NOnMfYbtn16iwJ+ZKvwarmD3oBTox+moJGIQBiu9Lb59jN6KPg+HhEKEo5foM/aZHxlx19vvsPa
QZsLsq5y7Pa2z6Hr+dZU8e888wY+U8GmIH9HHarb9o9G5V2TC/1sKHYRg8WAa2Ii+o/yXLykdtX8
1lsdfXBlgR3Ivf8Wsz0/4p37tEZmCdw7/FmwkMTRfq4X57KKfeiLjbsgVkRTcj6fgYultb110eJh
7Npm7NMMblEwblnWNb2g6vGyboBUUc2axLto2tv6RuTwcBI7Rx7GHHU2bZ3QaaSezBDP9+LWXBS9
mTZSa3/sDZu6YgEw750YhLgGwFEebo1qj/NAwb2HhCA/dGXkUrOghwfOVK+YHahMV/fsQq6qiCzu
OzdKZJDulsghpurWoV48sZIdUVfVXUOKxKhHWdwFWbuSwGz5BLwWJRM3k7m4cQCGh7Dlfo7ONa62
Q93vel/IfJmZxtyRlLzRTUnVUbV6S69IwpQ1l173bdQrwLrVCxqqbuvxvIKrtBtSWXK1qWnfxEH9
rDCC7aJ2yVRv3IDeyeWNona7wDbXeA+4nleUR6mA/4kFqY8+TGJWqGdFTTlwGy3szPKALoMx/yiL
HDQlBX2Bjqo5ze6JPt/YwAXyMlhRLY6ShId+D9Com4qMoNi/bGwlsgpYrwuScQiJfvHm0tPK8RrC
BMA14TLMtax67mtB6D1pAwU3620exNPryxs8d/i1lB7L9s32Gbgg/UNyMZ50qmz2rC6H8iezdgE2
pL28pKUMhhiJIUt3MTJub31RrYog9MCwiSAzjC1sWcsm4SBzE5NpkEyRoI/C1HOwGre63NlKXzn6
PJbZTS/PZ/NTCht297SQi/E4CKZHLYSP8FFnFtZ2emHoArEevwwUZ+1Q0GG8pBO3IDst8u7P4Yhs
hlVosXP80kKMrv8Qel0N6hGL8Xh+AM0ttRyRAKdFSlTu6iC686DrF4fcr3VAME4Lhw+64v4DAv1r
XIC/AKgTfWFEGG0RQmvTBUEFsnO3RQsiz55HiGaOgsRU0YKEiTzZYmizrPUy/ZVY0hdCQoFL7O/z
jvMQCryfD14mPNQjOm9CCRzueqH91jaXMpci31VtcmQT0oQsP2toZODvsoX+tkO8c5uvxiyGyPnc
50AN0Swt9xbJLORTBfoBgm9F9nsIDXdgXk72J6kNXM6Jrc7V4iL+sGBNRE8phqmni9Xi+kha8cgm
VOPvklYLwiqjRcRdRt+C0LHXfM7S+DsWjFom8vUysjuO2zVhTDtOq4Sadkz1XVsnT/FigBMSuCfT
DJtDaesl/fl4lpoJjcXnKaJ9daK9K+U53R6DGMJ3t9arM3VE3so9kbULuSix1lMbO5xdFrLNtejZ
1VOCRwt09PWBjAPo7SPo/bErWKdqZF6yRbGwIerj2Raji6/CJM25H6prt/7cy4AbOIDlRHeTa/2w
nLNYuGHQZKilW+iexJ6COXrf22tz5nNjW+jpELuRsevKHIEC7UM6ZfvwpRsafDw/7MOYxgI7TtGo
O/iIlhjFawKUWMwikufZ6snvjTMYjdOppsI8DyiCBqVGykDop+0UvEuYhhK8KyJYjEWOFdy6X0uL
CmOCvWMw5HV+T5XbfeoEfuxLiv6/1psLLptNyCExBBTa2VUEMREIRyUizH/i/SMUTVc+EYdF/U6G
uppgHvZy3x025FqGgess6+ZmqOjIY0wp4H+deGekMeFXxiD7StkgRq+u7Ig19l35sieoJZ5Skmuc
w0WYfv6GU7raktr9kBDSC9gQARU+h6wliBaHhUWbMZiFj14osA+RcW9BT8t0FpkWR5VNyALXmzXJ
/+mwyPHV4C0nZmgfu2Q9JIQyl/9heA6OX96+YvK5/tOeUM+dKb0OEmzk70stfdwhAEyiZH08aR+f
vn2dKafr3+d4AkQCoNKJZ3mI7vE+J8dvmMh6s24LlUwuvDbtp2FEGBNQ6ypLGjsFh8TFZIujwOP3
Xnto/J/ZbdwPaXDpb4IXdz/7WqTlS69d+Usl2VnTb3kKwqbe3EVcLitVifqZ28pqbTSt8JiSx8Tb
zwc0Vx6va9RIiR6gkmnaOZJm+wPbeVP5baIXyQixKtBBIPQoPnS5JVANhRtYTHURnoble/PEbGUy
pJnznlTS2a/YFlXW+K8D5vcbfD7KBgIFOoT9NfcZRXJ010EcabQ6cOyF6bNQfzWXobBVxOpam9Qe
RRwPoUOBKp/foGFTegtB28kSf2Ci4+rki+M2kdUCsqnyymLxjPvmgOIgnsOEWbYlTIX4LfnXTXle
7tcvPSMjaxnbTpahaUXZBZwSdEM3qRhDKx3YqlAOWPYfcWgSOtn0Pl9/IHiDLHp8IdIBRlmP6Ok7
N2+0+zh+BX3OO/nQjGMiZw8g7UZdmMr2rSbnJlf5FwpCSqDU7hlLdHQ1LkmXuv2Mw/dqpfpzRI48
ebtu8FSy7CnfK+5qND3Jy69oildoB9zlifVs5S0jYjDQo0xDsL/TIVLh7D7nxYfoGm+KKxvMoedD
cTkyafBM5hGV/GhtmKv+ktG+TruLBC4qAFSdr+LylWbj0bu2dniKKAtQvy9KCvcV/HAx0R67QzqX
A4EJx8uo0vZtR+OrNsFAzfDgY5lYNZCQx83n5axy7Qr11l/LyBiFMfrtVkHgsMA30drI0yzGYkHT
am08R9R/E5Y7tgbfwznfUi0s2ji3Ctb/TW2AKJ1gU120SzsvFoF8in6DWO+BhHqLlLtJw4v4KAx4
GTWgijwTdujsOAIwsW53md5XCXDn5JP8R6OnVFEknyKTpiazEeJEQ4hYeRjCtD/RcSaw4f+c+TYe
Bsm/OeSvfIb8iFg2rDnhcOkiRhpuo8sw0Z8mis/unnFpLhKxD622TYfq2IhW+cBxi8sAwgkV9zRU
7TgX6CawPbDIq2uAdQvt5ERFNkkSkXFQH053ueZ6SUxoNDurVhS5BkcTwSDMI54gSlUl+cRZiATJ
FJUkoEuydwpgzSH4Lrz0dApOfuiigZW4X/y+2zJlwQwynEo4FKLnr0Tq6Vg3CPAsLrEFsbSrPW76
u4EAqjD8z5VwhqJgA/e8PuQsCdx1VeMca8KL045g6hnOkcl02FNj+Og69FPJhSfHWUFOCujU9+Dg
6wwjW/XspFxPdlTaWtdR93ycym20Qogv+MZuvi9a76vywEnvpcczImPpNtOQKI9X6/qBl2kSrxAs
JXeWtA50pZrXkNrcVcCS7XC65Z2+k72nMkAwMQtUK6D4zh4RUbCg4PG/N4s1da+YJVVcWVSKmCvl
WOU/xR4e5Kxz6GRL11prko4Z5xLtuSmb7h/oSGgrmYd3ia2YFjfQ1wEKCLoVBR1Ftgi1SFGPqAtq
I+vZ9mBAEcTcPhBDDTJKrOG7Ey6Hlhdb2c6x5KYY1fpka+ndOwgCh7GJjHHbpKyytRMMaohEiOMR
tuHL6gZnxOa/OGmO1knB8WgRoI6CzJk0H1NNyaBp6Eu7LLBIfqCy6AmxqICL7zp4/D1y86BvZcIp
kIL/hDkixyjepYiKrPqCU3NpWyPxERWQC3oXviIgiu7pRszMXIvGfoBPUghP5JMbpnoO5p5PANCl
gTysjKqXvMSrcVvb4U17IS9Xuhl2Rw5ksg5zoAU01qYs+FTSs/BmZj0LusItz0o1FVs2VA3yGyvs
Y9AkbATcIfwmSDsoWjgpgYd17i9MJhl7JvrR9Y1/v9kveFDGskT4ZVSIrB3Wvg3/Ihxxscr3Rpv8
GVDXaGcFNrVdS3qjHH/b88nCZah7jnO0mjXVy3ItwmEkiZBDMUvwSU5J72t/DNdZL5RwbifQsD8v
jx7EVnx/0xM/XnFhycCaZO1OcgGdUlhK80PkvOK21w==
`protect end_protected
