-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2Uchr95GPkr8JNxQqMnMcGQqbGAUqRts+iRTgh+sqG8aqEYAxj+nEVWhFQgcdLPV
UzDPSOth/TjOe8c0Q6et1RIuvePFVnzcqS3mtZ5MzzddOk4WEbYuiDrui1QuIJUj
LVNneNncZSCM4WfwTO2cXbvMVwh+m5eCkwJDNOxgFDI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 10704)
`protect data_block
6lqveXZP+8vIx0vTgwNMyf/xCF4pRVMi0b1HIxlvioNuNA98njy9+i5oevU6cWTL
IlFztOhr2aGpeHCyiLiQGvLfNyUtFzm8ONmpnCaA5OXQCN0vx77V0PBtyP9Ivdhz
QOr6Cvm1MQXjjixpA94PvE27RLeei8FBCvFa2Ke5eXF/l1Jxx/BEzmUCnZ57HSp4
Rdd+NO1dxwRZA+SUsFsJPMBZl4+4Gzf2yd/wseG/hUzbeBhLEJ0ukd5UHC7V8EvS
OgHHx83pWDDKUG2UsY7PH7+/8XMRdE+pTbDA3Ju6uOzusReamJCY5wKfD8dO7GXD
vPnIXML36syD+l1gRU8FZSLN5XuqAmb6TVg+vfccnAr+VsCIwbwjkQAwmcr7sfpE
PBgu/PfnILxlCWorFQMgfCqPhU+xcwd9pmdht98gM1k6aJxSFXygF1WeHGTtsL1D
WRxAArqkxmoDp3Tk5EE0I0KB2nJTju5fbbq4H/3oaJAdp1DhwpXXmqOVbkCGk1ei
o290Wxh39ZNagiSEQ2+uCLCugpuWQmqTds45JGLsj94rriu1cnVywO46r4f44SLT
9ncjIYxlYw0NadPHtyuxhFQnrgkk3AeefVBWIOO1kV8m14vYycUhUwcrV4YlcLGB
1qKAAw9GH2gxmQou1fQYWUDaW7Zwr2tuhmq3Nr4SZTWvdYQHt6QAGWdhsz50QAk7
zMvSuzeJGTmr3o3qwWsDT1Weg8uvZt+05evUGV4QHT58Lqa2iLY9Jt7GpZo1rgJc
W57m3DhiSx/A7XHcKgUMAne8PMU9peZ+uW1OQHpsfiCJ0YzoXjSghp2hIszs7bik
HkjDoSUQ+dcZdHhe0s1A1QeAeYhi6CvjWpQtnZj0gJ52BN/iMVOtxj6u5+rWPf55
6o9yLg7qt0guNkg+47H+dwXoLanWQA8YFJ6wbuhxShxBpaq98EMkY0mOTx0PAX1T
765xz0KSX6Vd221Ojyiqbn4Y052+4B7vxIbaxAxQl+HcolhMA70+ZLkB23mE2X4x
fcIln0K/DVnaQpG79l/gBY+IIkKOguqHootNFDXHdl/cHDLNIHG1FDnX6tM4BFCZ
lIDqdNRq+ZaTjDIfw/ZYuVcmgijLKEXj52FKEIuXvaD6CxfWvYMXzmFVILNSBHtX
VbvGUHSe/SWR/LmrUtOXCpPOdPye8EM4VIK9TO5PG7QHFpiG9x9Rnserq2dGSKwT
CYad4gyXtN4VrvSLp+4tpU8LHUa/czC2xxWg4LDaz/QUnvkaowGmap+xkyzGyAmg
sHKuzbXKl3Sb33+xIERfhgeIogVztOcboJSgJBGwdmmkzWW7Df/XMdpFACCP00ll
LiONxi+Ib08KmfDfu2WghLAgPIVkTZx3LtXpNIpnmUT4zOKrFSdgbX0FVtNd49kU
uubNos+dJZjc6k9XaE5t82IIXWs/QoM/SMV6SCNwv5M6aixkJVFhpSJuSLltm+BA
yUAjFQzI//I6DWfBOLG6R7EoMGUrT5E1SmKMZbaPW47Zch7r3qgmGg+G09psblOF
gsT5XfoV5F818fLAsAy6PXiKuDn18cWwebGU4Rugct52k8GQFwRq9QMHwITpezF+
ud95TH1l0JjtiyVSsTocwX/ahWz4ThuQ2m37gvq8l1l0h/XaB69s2TlGyW+apyU1
OS7i780Jkdcfx/C03seC7doUBszHdpwbfr2eUjrpC/qPKmHk4rNP4Cenc+w8TXBl
FctUObZarFIQw38ehXQwMqyAEJQ+WJVSU9sdreo2fQdC+KD6A8o19zasudAQCPrH
JEZVHGRhpmz+GEFjOdd64uAGO5Gh2Jqe6VsAJIu/sBNU8h1TSU7JP9fofqz+D9eH
0/b4awBiU2ij9BQkzNvIp0Q7DKCVZ1N0qjNjFhZ/oFHt1jROSfxFwEkC785oOH4a
JyhsKO9JT0m3QsDZ1KeyrmTnLbho6bdvJh65znO8YC3twmoUn7WSdaAIqkFSycj6
icZKU+Jhl8/9Dqa1asMnTNF3HIQLc/DNvVj73UfUEbSwKNQsVNSvTsPYpL5ISHkR
iHxmSe6BL+8uZdOniccGM/rGvMlyjsvIubwYhKrvFLES2WL/E4i2DZtuXvFnME7i
cE1k4ltt5ljHGcDBycPgv+MQelsHGMB8PihCXu67kifd912lprAGhmuaKyqnzjS/
yRVd1ryuMVvtXhRzD07ljt3JsdrCcbs1INXfRB0dn7j0psab5Etfe04oILK8gtvr
p/B9/DJpgA8uVaBHK2F/Tej5gkTE7TZO/iQpu6Zo0AsM2kDgQUKGqoGAa8v3PVER
NLy1dbVUp94gz3wmHOmobkgDfMonJFw3WdxV4oZRqhou7TEXgtRpukYi0gcodsXN
xlUYQu7VRtBcdhEqEqd+8dJ2t5BHPz87OK9P2hNX1IjSYVVnOrhvRKDQbWEjonQM
ZjMlKDW5UHdGV2CBwTkFJz57N95Y4bwq4OV6zW0P6BWe7FaVyTzieGciidYTIE2Q
bexk45xO1gBkHRvYa4Y0hpxW9OjdCx9wRe8WFdY3n5Sib+ESQWLj59vpOZctVv3K
9A0eyQACVNHHZ3e5d8+pMS9LwqztxCfOQJWQlWfe8uc5rTGkNEShPFhMmbNyeIxL
6Wi9N9DbETXlmYVb4miTChZKQBYJURjxCfYaY7ptjeyaI1HNlgSgVyXhGj4oo5eQ
nfdwVqF0aoJbF9HEDqyfU4segzTxLqmijQ7kQeMtbMqw29qr5K1qdD3ztT76Mwnw
1AQ8Mktl9JahCpCl3S7HM9xlDLtm5QsE7In4SCU/2orU/Rgkh1cQeKCK5pOo9wxo
eXe7u2jU/BgFhMg3GteA6HGCSdScL9wDS2lAqLCheajbwVPcG3VudMUZF7B+681q
CHv0q8jMnRYuWnAPLcunH7cILSB7fHcx8bPwULRZZAnfWFdyNWuwlkpfZB9dl4sW
shnu5qS7Z5xQnGAvEZV7sBmVpKubsL13QpvjOBo7VbYkfnyUsUBjb7fj988R9hvn
gLZoit/vxfa9i9QFWFJjdvAy/i+QuT7VTsFwxOaxzag7c8a4QkCcwWMI4EsI77Yp
hLMImGLYy7joGdz1YeTQhtl4YFwPcTVsNAGU6+Nzjl3rEuaSLc1FHS+NitHuSIH3
obz65gWF0AsZX8UpF63zveBNICf3rK+IsT9qPOhvHMOR5Dsc6vZyX8S6IUlSCi8l
YF6Nb/Rrw2HoqYSGiPkRhqpqwu4Q/bFxEhlxMykdeRoPzZGtGkuDQdY4kJdAu4nW
4nHPVJam5uj/QhdzWBWC0QyAKF1fNzm4q5BfdxFrKSHODBOQqhS5/vBDDv89PZyW
YAHvGaTQDUB3QGmrn3oiWG4HYiwhzL9/dzCt0x6hz5ARPYj8FWbXbh3djCTWd3iv
c60KCww8HmYB1BDxKY0OgLs+oClK7rcfOfmND3g9LHiCzbmQSVNCBNJS5yZYe4ne
idiqogO0Rd5eGyIOfNydO+FlzLPbZDzx+KOjUbS+9Xfeerq8yDaodvT1Mv/MycLV
sCeF4t3Bt1Zfy5g2E3T35wZIpiZU59BdQuhhoc6JOSfo5XEXOwSv47OEgxwI59qn
BrqzM3iHV/DBq4f3qByGzR2io0grqlK/4cJVzDFOBy9Gg7vizRH8mQ0lJoyCUhAV
aJQEAlicrwqVZ6odwCAQqaiE5+c+FfPUJ9goTWdHx+WgIorsZkPEpw0msi8K+AIh
/gO52jfggXW10eduJimxKjUIUS+JYduzFpOT/abhd8M51bNLGJtVtmh0du87JaRy
L8M0g6uWrVy7CkaTY688OS3qFmOvvhUcp7ZSWE7Ef5EMMScIvkUNtdhAzWbeoR7Z
3WAIc8DO5lXlXRpNoBjbJb8Gnmxk+qXH6/OEa1EG2BmslyvHsiropnC5vHPSBg0x
VmxDyBFwWv+Ts6GfVjFmGMVzCFhk0bxr8aYoHQ1yVQoVU5orxcTf61D2m2Z017Ep
UpxQ1b3Eg42M26xcXN3ajVV1mEt3o56EsGQ6WF1T4LjeoyGLNQoyvrnPP9Zd40Mc
SfeoRvgwsFHYVIn/QEJtghnW1ybtzbqKBta8cU+29H9y7EV+SpVZt+I5YUm/G2cu
EoHYmQ2lQhE4civPpCZEZBA8sdQbVHOdTfKrG2yFDZL3wkBtGntjjq1i2NgGiOC8
rdCF3+1x+mBqjGVixkMa46eb0NU2IWu85tlLqIPhUhuJl3Jw973eXzdaYlzbjwS/
Z5o6rb+8XAeJu6H1BYnDBu7peZYT0+Fv+VmdzVm0IWlkXeiIKbOfC+Fy8S9W9wPI
KGfuysKOkAGEE4s0BNE5UE6N2BOA9hmK34bKo5mPS24c5W0AR6q+IaCtlx/IklZY
x1iTY19ZgMezSrgBt4q3pJz+ziyC1OI19ZttnKj2rEkRi2c9RgRW3J3nXWxbxMKO
JFHzMCNwTXN0beEPxWWSPNf3fIA+Xle4vTZrWXhoHtrA9otiFndmjEE1OVf5h8+c
pdzvI6QRXcVIXEwfY6V/vZ0oamSHOQ69iLZR+AmCn2pUBkjhO0LT+wcnpsE5QKyr
MCLsMMSSIrxZAyNUCXqekKd5F+up0QOSN0U5uQUPXKiFfFtH5CAQkpYCmQJimvBZ
FMOHlvTN1dLf9w0KGJECrGD+dFCAj2+FZeUXPYqI5Rt445ZGjRwcpcouGcoYX1A7
n+IRg4tNAE9MtJNm18Z/B25vtBwOOKYcGYp32SqjzJEtlMwKj/y2jbzMDAXqu5VR
hLW7g8jkduSQngSZoOH7BBaX0gWK2aRgxhdqDfAcJbGBMZqA7LcjuRrSBuHUqvaG
rqq7jc3lRWkKtenauOFskpCRh+oVe2C1OuOWFMhFUoKnQR/yLJDxQ1VCL6m2cYiW
BDDoXHxlAqGhCxFY2RdvzzlGOXMXMlltgFZF5Z1+4NGVWmadTh4FAI663jYrlJ4K
f1cZfMhcJhkjyXY5eIsbUZqjckIlrbExrNgw5ML44DUHXs/zW9qBOnCi0RPA/76C
2ALARU+HTWJBXHyZC1tZJP/1ofGWEfcHfF1KWtjJuESJIOCcUm3Qa3Fs7G+n0pxi
HPczY2YwqW5+yoEQCuIJCpioZWC0pTxkb+hOCR7aDkLeQ9zYGY1T4Xbs60zVr1Vy
+lZbXSe+vI7QCH/6VaOpNA4fXaltRUP1kqLkMJdqM1W+iQ7Qj6wySU+LxR3NR+yw
1cJMmThi7KjPfTtJezHdtji9BaEWkOhDDD/raNEl7NmJuDOe4Pg9DKTlVuq0FZJR
y8Y5oM5zRHEuZhBfq0Uv3lTiXRudIR1z/I3fmL+mOQNIWRa8MjWJid+Z6VtYELVm
sPX3vVhrKk/tHZCJQJel+RasM/gm2Edl0hHc+jgPz2QC2GH5w1gR/ehmLTcsbksI
5tdTAu2lk13/ua7kYJr/CARfZ7fb6+VEyyEBTd/SXYlvkAQix9OX/YkhZEhViiPd
QPEkUwv0EOVQAcjDoB77xFGQCvZ3rpjvFGYzXrVDqWYVEEdWjdn3V4F1HI+vYymr
YOB7mythRxLTDUVKf32MvsSe2XY7q84bvuRd7q3gZBDlxG8hauktzPuN8hf8fHUZ
cGN8/nwU6YfOskSSLF9GvDgiN8p9fqgr356zITBswl563TVnmJDTX2BkaH4lHIm9
rCKxNHIlJh9AZ77nkYlsFTpie6xVQYbPir8VWIlcUCSwL0NsLPFOUVyuMP4w1fTA
b3jz4RWtQLwod87xvHsObG0FAt4BCZC+xGbiZIQYMairr6Qq5crG/WCOk6WWGxYD
tP4na6ZGHVxchGS8ocDVvTLJHitFMNAlKfOAQKBB1CJLTDU+pzcyvE2n1cDDARXw
UNSOTSmVc7FiI2iTugspFHoSwAn6+KfZ5MvdHlHrGG7rMst6uPcDKNTxVda7KK9d
ePXPUdldCs+NA2yEXX0Vasqf53rP5WNFyyuaUQ350DwQX9szXW9QAf32gTjuw931
n/vEufPJksLWz+fsk/e1rq3hR9h0PbFYsrEHHvyMkBJ3IrqStGPHrOj9uyR+BnhS
nQVnumr49zd/faQgi75IwFJ5xsa+LKxlyBPn6ULE8Fu6tV6NGsn1YULIvz2F+K2w
xOtDhU93d/odWJihlnuoRmi5cfzoQUefDOlg/FCItARofOyK6dcPXJVlZYc96ad7
WXaMHdfDV9LTFtwaEesXWjJrT5Gem/rNntYaKCRWPTkKojiVd77R5DuyaEoxsqNO
9OawAI6UILhVv8P+Hg51MDrn4Q195LApC1942UV9d3sQ2sU9X0LgkY3tfpE81vBD
gVpJdk65J8yhLMai5QO46C8ZKzQWEH6op0oko1EpmgyGb2/xPA7S5oom4VOKv8zl
0if4C+zOLfe2Ke48hvwkMgzi0NJ38dl/zaCdomWIbZc7tU2kB9/j3csAeTi7EQqs
uEDHg3ZxnzWSa6S1i6VfL8i1udhYowxiwVntO+8GBYLk5XoPaH2dN9S0n2Xv26Ds
V39oJ1pC0zOqP3/ISehuTVH6yIs8JZIDMwtW9XsDh2qX6WtZ+ctTjHqzjN+b86nV
nrzqRMZCThMnfAxAwXvEHBBaGvjIOH1r7b3kIAmEMGzwHsKZK/NqPIxE+nRTVSfL
OCj+RcElSl+d1w5j8U1uZonD9h3wNncrESuo+0pEr7dKo1X1TujuEXvMRE7sknk8
hp+Fvl1BFTlI1Zkl3u5Ow9BIQvsLygp3aOkd/5yCD55GMQE13d0+Us1Ocp1Okz38
a+4IFfF5FP41lAzcaVW5MDhBlWe/bRMpFQ2B54brR2cYJRm+bLnqLKehf3pI9lhU
9AAcXMuWLUtliNr1WYlVyECMqCxngear1PrlB9SnHCzj4T5MyaenEjbvVfkJmvgd
2RCCGNv7juQlaR092kzWc46z0o0kM41z2f+BpOIsQO6UqpPyyz6x+AdFiQVpDnLN
TXJmLLWRRBI4fOx9t7x9Zq2wM1Um4waIA+CFljIUnxlS9ug8lanB6RSxmxOJznCG
hjbTMEtoJPJomanOn/eCSUwGwJJIM0/uRiG8lMXoQ6bh/yAicw7awYBLySBxXJwP
/J+BdFbwyqOc5NBBYUnG7vogqIg0aLDnNdP1FxBY84HazOUSc+GWK5k8p4A7cZhQ
l/Yg5MtpDFaxj3HoBzhz8IbxeGIqFDtM21gXY8baLXo89YtUt+D+04vrU6k0jR8o
wrWIMQ19g0Lhbd9ORCieUFly3e/eEP0uZypr4DpodR0Z6kJvXiGuB55CMbEikytx
sMe+SOHgf4ikkOlmRzUOFEoh63CWeC5xx+V+zTnQw+QhVlwbE6sjqJ8KG3IxGY5H
vUCU+jzJnHJqREmvHApc3Nm3k+GmNWfaCkvqx8dlg0pjHFQpQkeflHRKvNB/45aE
1GLPXt/F0KCVb5ZJOUO87OQwZ1t+TcWoMJmnWh8MN1Q6Nl+LdhRrxAnADF8cSkve
biX1CC05mTi72aA5Biror/e8sc+RQk4fiDlKjWmjB3ptj4nqU2aZfHph2o20hiJk
N+5HtOm8CZN99LVPTz5X2ot9rMCioDqYCllBdinEKqfUa36zjvvRebHpEGt5fHhx
2MEqKNlPW40h05s1bToraLyNDTiUC8+7mF8HImrDviutjrjwPGRGWchYc9eo8upD
MKfgQDN3JyyRRPzlG97R9r91kovpGOyHcSiA2e9GptMONKLpvDQcIA4PXqjd3pLF
zuDKWR6Q6rG/tYDHjB3hBZ4IobH99OwcPY7kjQtaHIbEs8172yjjNE0arrOwUTLD
zKfQmt9JDDwYdPW2RJ6NEg4B/P/lQl1InUR7R5v6fcAv5X3XZuDTqmKfHCx0CG0/
jnsHsxUlhBkNyQIoXu9Lu+AsxkD2lp46vZiM/ZKb7fxzqz2N+vCxWWbqNXdGYQ8O
FeoqGbDiMt7nKuEIcTcSDH36XY4HyF/6NNf0lo99q1Vz1WsMN11A+UVBI9XkLJPx
YLeoxXzfafclCFg2xTCp3xs7TbeukgjDe6hMr/eUcRNn/lovoTDFl0E4BF12hg5V
Cqi4goys1dM06qrK1ncbWgR3bZjTrIbwn6vy2GbIQFYdv6+s0a3zRqIniLsDhdhB
21VB8bgb+YF9n4cMdD4alk+oNO+fAG1x4ipIbQg/dO3YaupBjhlhsuYg/SmxSqKa
wHAdvaQU3EiHLwVLe4MgRCNG0kvtYCGQPq8dq0XjU+KmTpEY3etJHCvmGLaRIjlo
Gz6kG+kPmCDioWi7JwVzeCdKALnFU2bicPramTBVt9KyTs9AG6ifLyZ6S+XVwW4G
3TiLjpMIYzLfMUwZDbCXiCDJR64DuGRczJxPGPFNYzU4Ktkumco9fgbjYBt1GrK/
V3hhO7eH1z5x1V8REDDXcog3mstRqIpvESWB5H9bmOw5jDOa1dX575RaowQOU4w7
KCn5nbyzHmJ3zT3FjVjvHs4b3cE631F484aIhFnAx/WI2BCwLXH0VNve3I8pYeXM
S1hmIV2waTwf0DO9GJItTQjGuBcC9RSwP2c7ROCNU1w6cJmgZVRtBLnuxdkuVDrD
LzuzQoHWU2re1e4e30XWjnEkNwVMHsgVdRrj8khHmPldR6RltjpK1b5GSarr+79R
73GEHqiq8xzeas+4UMib324IMV+hjwzNyOBHpj0l2NhmK8vzbqSNtVb2tF8yQgec
R4HURKjlM9XaFGN7jR+XSymSZ04f9rsCrWALSxej2UrGXv0cxIl3oG2QnU417aer
H/YakidBf5zNpj7YUWN6PhT/J6ww0eTi91uxt2+hg8Ndgebk5BSwxLLwVrsb7rmy
5REbC+egaHKsnJLCDiFO7ARIi9R8FGp43Yv4LuCv86VmEvbq4Cp/YJfHtYxiCYSp
QRvZ7FFLuMSmd5yu3GkthRqLku9UmHi0dz3GvpTE5OianS/g2YnfktdPogbv91NR
b8gNO9A3boVnvUe43i/NDZNRGn8ETX5uLdgjc7q8+Ek+FSvHYnfkipcO/z/1m3Yj
0t7lg8YyoOBLdng5DOZdKqqeXV40knChQaBfNQ0qYL3m8PUXWglY0WiBjQupJsVl
BkI6RxxepHj07loBxwRlJvnoYCfrTjmxpkRPDPTR7KaMFjAUuMOF7H5GcRC9oahx
8h0reFzqRfT4qkth8QIp1U2HqSTXkqboU5U4t96K4JkLrXcBxLSEosGa5BFF4mC1
+9Jjks1iRBNdTn5aU8vV3tydFGARqFAmRFSCyxonlkE8gXeWHcNmQlJsgB8hBdwu
FGYO9/Y1PTH/Qkd00cG1xjYsIBrnTyUw3AvhkHQJz4h6xdag7v91TFQkcmHrDOsJ
Ttbs12z7DJ8xo/4eqwmebZHoSydiopJL9GA/a21dhbmUT5SjvIWRuoObOswyk8/X
cNG+05tFtZbMkSOdb50nGdumpYv6l0DqDnKEnt1kFLQlK1ZRcEvwVsov4ZAQYdz5
cztqJCExLm+WbpXdPsinaANMscYMtHC7FeV0sWGeXpRTJm8t/nvq4y3IaQk9/tVg
KNOJOVHLCdpf05gyP4njX5GlKdt1wUEryZdm8m6gVzCWB9+j1iybOz2a4ALXBdSx
i9xiqvoc1qD/L77BbqIIkYfdTTZu3qprvzpmS/VRyVzjxwHZZ6RpXNg3GgORoXDE
tkqFQcOviBOvz1qnDSOmK92yrn6wYjHeyUKEA8yMKoCMseXnnaewsaBqEFBsIV0t
lszHf7yv8fPtkZakgkbYF6ZHwatEvE2QepgI8lbbkDsTUm8QfumibbfhqwIwx0kg
oNaZhJHTD5JjFQVRSiyddxnGA4QOcfkukE3ULs2Eyx7bD32ffziYt59lG9xEpwBZ
5Jg+nu1qoZOTNE+PRNvv6lmt7nOkF99GBUQjntTZKOJRjPHU7dZMatlmj52YgfBV
LF7NG11TlyejYKGyew3J8f1Q0KwyxN+2R2FKft5LOpnjdrcZ+YM6cMa+5S924ThO
pBke3ZzSIh2fUQrdwSZY58r4GIQMsJBzBdVUsx9rg+7oWij6XX8zTEtbfujon+oD
AbavQVNEDosUC8BhO5TTZftvzbEpmmkYqrxwuzj/ixg3Uyr89LNLRsEohFO5eCTL
Oqk56dUWYfpWB+fe/FBwhDTn3P0ryfwJK/sdEINuXV8cnGJGFDiDJZZQPukXeTke
oE20ptkoMvEfj4V8m7TWgKVnk5EKttExlZfFFYkoK7P7ZSday805KxxgrxBSxvHp
YZbHmvgTmiyfKP2O1A0gG+kzz1P2G8cI2kPaqe4YvoETS3ziODvQVR1TzixyuYpZ
XD4yG9xlBK9jXszTNosyWy+nRVzZk5Dr0Ja5hCgkVCDtmko9MJmZR5eqsH68VmQi
Ujj2Y9gciDxAKG1441knZht4j2H7HEJ2BId+2CjE48vmApNJODHg+1Lha6SYwUeo
kiIJCESTZNhuCCJiki3vAs2Sjac5aygXvhg8w/cCADS3CSHYL1ft7i+WSAlMDMed
FVyx65TeKJg7F9Y4GXou/6dlX2wjlgjx3/E5K8fMeoS1QYRA71ghqh5YJK1h9zLo
sjYLNQPFCXWRYle0dB2AG3xFF0I1vXrZDZaBGLj322Th7/lVTYhXz7JeOXI9jxG4
qW0tckLf6ODP/WLK4sLimhZ6AQJHhadILWstlSD+aQEeB7BhguzGkdZ5mFjhosPm
elFxIUZDx1CNKT4nAl5NYkcpPAX1+vaEqhh47rGWdaXoMW8uFFl9QpwdUoMceS2y
BgJeB3mR2/h88nK5jdyhQnlrKhhqsl8aMz1EDliGrBadRmezZQ4tvnoGvl8MT2Uk
+0E72+IyvJBQwToJ+n8e72snszJ5j+ARhxiH5YGFu0CJ7c5FjPRpNhpz5f8Owyrt
d08JuuGb5WCC2iW9CW1sn7FgJwCNG+khnf0zC0wfZiH3WXNcDGShWhj4+ffSvE4i
26YFjfLTcjXXRR6S9c67toOf1Mr73e3y+Qc+j1iAmPunQ3uzqCQNho/0aGc/ylTb
ZISFC+rOc7hSt+8PesksY9M/hV670NB30zJxhcrL1FkFtqCQOqZsoz9jZEQn2RAz
XIewy6xYiRIxo7UgMEF6zdZWgoBVRtjANXrS9GjOV8vc/S81ZXuKl1Ib/PUmFWdR
1EELsFlJWcifvjLkVctXleEn80oFeT13MG2zKkDCRS5Vl2R+evgZnKcZwr0w7DPF
dU8qNm8L943wYAbAOEiXDQGAmBc4C5CXukizHD4DXbVYOc03aS2y2DmNi/D0fRXs
tQ0Y4UoDKUPfyZ5YedxCdeCmJdJiO/fi56Jihq5tZPqmuDVLoGafFbP/fGO0Hjmj
8xUDYDzi8OIPRDkeWxW7PNv4FP9O9jvYaD7WKCnNC9eqRWeRtDzuqFBktk+xUwBD
jCMxLeQPVop/VZlPuxRGZwWEtfT/K8Mq9YL7oARrgXnySXQM/IsyJHUBT7fOFsZg
cjX+XWiSuJJKUXISnc6FkuZvZpfMzk1k11untaUqzK6o5mEKSO1CrBBR1ABqOH9M
uh9dXny2hv8xh0CY9HIanIIufxLLlVSfId5eM2eeQyribYBz4uGHyZL5WqaSgKRo
VUYdiAcmEULLZPGZpAU3RUKIsc/zipqOS90v/OY88nrYe202jOAthvWGfF7hd8It
um9rhCbDA2FVyirBosyhhfRUh8jPiFJXndBMS/ZOC0Xm8T5di4NmHcxlyute6bZj
aFkH9Ks8U6j5BwQ0LNhcKDRzKXGGj4Vh6qk04jnGkr6RWmn1HHxwNFmkupDl1fYG
5Zu//+453lCjJG/jrFyz2PPqFDgObnaTs9VKfYCMODfq1x0AENLs1fcPUqgmef+2
QPM8zAJobzA3ZFMkiCFkdDtBTUT0g7xREpOujsYdRe3jn1QEznKCNaEL9iVj6Ex/
dkI76rL8QO6Tc/VfNy5ocvohyENEFdGeMKuJoRkzBPM8i97UePsaTiupP5IYyb94
L8HrLtCDyBbm4Hl+XAMi6y4kWN0/JGAcMyKVY2hPuUtpodke/lT3CvgZXO12kj/S
UN+z1EumaodIMUCqi9BEiiln17la2miDhMvX44K4Ex9swFGOnLBKIA5uSC59hrbv
CeoFoOiNKF65g3NPZmFyw83PZgI2EwJ5H2f8sey0PSlC0+VxyOFf9Qcj/dqNHgtg
BvUx8IiUEbqqwC6d39B63UhTi9uSCYfWyBykd4eZG2v1yftOjnCfGK6eoQerA/eO
CdT+UUsWM/tCXx5T6pXUN0IxS+E+tYJ6TMuLy0GmUsw9siqv9JNN5FfxWZUWGMKQ
CNYmU8Qw7jwUwFvrDIzZ0pkHpSf28pgByMoDZevIW6wTqg+3wH1oz1hmaTROIsqr
kwAIxW2ckNPt46Xf/TnaGqyCxeifVTWJf3q8q1nHDtLXZB5uTR8VrCkfQLg5wqAu
O9k18KdARBGO8VXQDmvRn/iAna9VCCwgSHhfjcMOiqhIykKuFS5XG8bK2zmNgt/t
JXlUoshTB/sCPMp7PiCncSNL617gORIXP18tuLi0Rz7OCZPej3UFwUGYA0EflAIl
rIylXXF5PWECt2WxCZOSwBgNNK/B46XncW6cLlCDnJ9Vqzln4GVFPQILx5j6h6kD
3Wm8w9XsQAtgCTAUp/A7fti1V1luzsB42+QtFUJnPQ3+czpALwIaV9s2Sog/R+vu
xeHtgvAN/yNr/EPB8gUP+EXLrvUuxqghiHk02RofLFItTbfhKklH4MxkqqP4Dcch
z9K35xFoVKZif15b4Ug4idmFyPnaLjOrGpstNuSeaJBjlbW+Ju/ODvb/xsUGkmxP
9svJLA//r90QY1JYAecTi8QtRs0g0lhzqq5fUVYlM2pq1qFj8sFK2Gfay5Hj2+d8
PPf0pDB2t+vZ9+77p+1yclntdmndGuRbFXj8/p0Q5XOu2+pMvF9OvO9S2rWe0DFL
LDqGQKb8KKgEwKpEPiIBFSExUznX9mAMDg8AMPRSvNDInEZbkRFp+3/J7P57W910
qjYn9bt9CmWtAyrMOUBqpZpopcrGW2/tI35zW7xsPGe5ysdFZZ1uW7wBLjpiVUs8
jOWaCS/7iAdZEVQNVgxV8bo1QLCiqsj41ehdYMOxIDEIJlGyhEekZATF7TQgyRhr
1lfuYS2/n3/qZOHSDP3sApoBxpiR5T8fs6XUm6l+TLk++xp4wFNPtq4fy06QrmwP
65pcDrV29pd8P0R33cDkHfHiLWXayvFFVdhp8v60yN/u0WHMV4GVieg1af6ZvVwZ
Ggb37BJSM8biA9nriedl+37BSTF10u3Kft1/I2pd5n/UEvNluWDdR6i9OMCxL4ky
alJb1Q/5C9ZscyiFFwbAt6LbHCsA3JGnLbkDp/85txzUn2t8AlhBDDzmWEMBHNIv
fHN8LWwxu2Qyrul3esndmVbAesnUoS0sIswbNfndeCH30dK3GyEnmtsyDvfRqqAp
dCyIE9f3FcMvaQUhdsWN0XmLXYCxuQONg0J7hrjMLzdF0ENwhymJLxN2zGBYShRg
ZTL+69OFbuB8lgH4SeeyqbtDwm9SwWB2OaoGH1ye6RDFBP1Rjbblyn3hAErb8A9i
CJt57FHRWKNeNwXGpjEdVCLmkFGumcGODfe0bj3YDAosEZ8ri2h1SiuQKS3fYgIf
TzX9qsVQmCZdXKPGUKh7NrCyba5t17gpkkQu+oSF43eq92g/BEHQ+JmICGz5323i
/r8ayGv01/AhVfZT0JlqFIB2tuA3pOotrgGs1BRIEwTJ2sg/QXN8O6M1l3qDuc0j
LjSLADIxMiRP5BKgi0/dkKgjW0RgTs+qXEppUc5PwsnVwi4R36hU1HqdYRm+YgAO
wlhjo7CHwRYf7ju76Np/x7GEdn1RI4N7JMobL0DtnXBb5i3/KUYWUbz5e2GW17WV
OhSBn537eZvJ5uQpfu8DWTlK3P55UQ5YwxAu5I8l43+XYlQix0w6Wp9IgjqgQ/vR
ctt6xzfm26CPrc1ZzV58YVN1jtTL+Q/IQv/NqKrhcS/G6fM6zucBmdwKU2pO6/8I
e8kJRwAzxTBI//f2Y/13H13HmwdCy7Ym6YTJVRprq2iDKdfNWoXgN+EQbtVNyjzW
C2iD0ZZ3xRFXO+6oK0ULDpeNq4NJzZBt/eLG9ZaI1UPXrxDHvgAzvNc1h0P6tGoM
QuVI4jaEcH6Fp6Qr0FaBpqQxKdBs5w2O44WT+TDuR8+/hAZEBMOLCiqTY8HnYW6b
sCDi5Ogwe2vS9A4ac2xfqsZdO/GQKLvBXn0tCnpq4zcWpCd7j0I8/jGlwR9zuVxn
QWptHrm9V4WwHKZjrqOTxD1L0/dw4Wx0MA3pvfqQQ7m/hjemNoeep8nltwV/Ug3f
`protect end_protected
