-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
UYdS3RR9Ur9+ffsF/6PRFpiuF/EHqju8QU+AzbRxETIIOFAmrOSNPGay0UXhEMF5
7BrOGC2cdIuMcEbPAne0UuvVOud1ScP3HsTJ5DMPmCnA7dhDtjmfSjdEjVFDjmro
tcSk3rMUeTtK1Jt/JIy9/efqfWeCKAmnKDBuuRIkgyw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6411)

`protect DATA_BLOCK
sEOD+nyDIivTq/3By1lpnFc9qnDUYK4tSxpTfPQx5w8fhDcJs/MC0Vqw/+NjQ7zk
t2faf6AEYslfRZN5bZb4CFbs3sLowfs2f55kit1mAa9jwJj7qWhxQrz8pvqaYMSa
frRtmBI/v1yntggpo3I39E2wEr4YMxRmKqskSFPapOaTCwLR0i5hsG5wY8TRPsL0
rfDQJDaDnv6qqsApXdxvunoAXJ8gELbYYyTiJArdQhtO/+B6wS4v9CCfgto4hXhc
OHGd3BXxk+LDBpthYl0wQNLfRt9J3bLMK1saeAW3Asj9DMaXCCQdHaTWxPXrHMuv
mFi/pduFlrOn9PSoRTFE1E1+WdyxUsKUfVWq6mtS/gZ112aPKFlYy/hXgmBoxB5h
BNGYopP5SfCEqgy0qSN0ELkM4k5dEyEVLMVC9RYt4o/YvTN9KGikQvzkURUkKgCk
RkdjIk0TpjclECoO51jly/pYvSzJGSzwHGlRjuqddCQjm9ua5PdIJRqE/XFrxB5E
Thw+3pXCXcipeHqWxBuJhRrmEo+cUljTiUaRE04RpJZtWjlqhtvHrMxf0+J9gpif
99fH1qPwF3Z31/7uwuQC+HRQz7kNguAoHBQG1wdO5kQrNrj1ENkn5dcnIPrHmI6Q
6mmkD+DC132WXd5j/e5Jmzdx91dgEpDuhEm4q3BWqnOvdwQ3d5D36Kj+QPm/x0ze
PvBteEDnR8Xik9zBg4+UbvF0uIzZuUyAM7nExKBMQGlpmBV1saUfW/cS5JWh8Qj2
ThK3Y1DWtKlWiqtZlP5qaIH8i129InZ8HxnUEif1TWqMN8mvnCiYOF5U0LpZ5uGb
vSpTpIILZ/wEyzBJ8IVSKhLuqWfuIvEo4ICv9tFnQ9+9KFlzJ3rkMPa9WLnHLIdf
JLYcKPHLUmwLv5nQ8MJbxaOtQHefYC6SNi3u08MJJ2URXRgNFgFVTACYzVpQbEES
+CrVBT1lKT2v7A9UCW89XZM/LbKQhHkK2C20KR/qEWdfvf7ENFW17HGAc/dXFkRQ
fynkx9ynyUmcCkzoDEIMc4H2rez7AQeEXs93VdQv0E50ffTBey1vIraC6hOYR+ip
MLnX8Ao3YNPbgMDjVmz1n5lNRv+VezQR4dnjCKrAfXo80lxqrvwlCrjI9v0AeDdS
J9lZaBK+0jMZK0sSvgjd9KTssuZOCPEAH1vhI+uKJmx7D9CrmPY+JGY1ursTmf2R
YFJ/qYcZLOpfhLhn2ZtuTa6IDndF94xF0Qze84bihPWI521WaE+46jiGs2tJGrKE
k1psoAnqd+TKs8tAQMCwXy7/EaojF67A4BZ3lM3am7gBEr8QAOVPDhHumKcLwCBT
fyoN1DuF+CX4ALGoW2D1kk4HOiBwUCLi4q2ndnkfDbY09BwYMnVNEM9d9cdoCueM
DWrYu2q6z/4vWcTgiqXgHJWg0Gq29XYM4kNhJmDzOO/v+d2VITIhS8Dm0Z9MxRbe
HrC99XmSbxCAm/ObvsHuWjHEgp44NArf9fmEJ5mmVZT8g9EH5S5arNlbwE73A/Bq
r7Wy+6Edr66vG0QmkXgsd30BvnVrbZvKaP5CYd579lJxRSFEgd0BVF8YZU9fFXqF
8wUv4xFCPK+iF/kt9x53X2k4tXNLftdwsl3hgDypT6QeYWPWYpTjQOQ8P2xlFDLB
pKk85wnaaiYjhPkN1mg6pKfEI4B6fVWCfaaEvZulWyEPIkeJC0146KykDMXzIGyV
YM67YoWkllLrNA3wCI8vKEJmgbN+MrpA4sbpyt6X+yvCq5d35X02Ix+JCfnrSH8W
D9rzhlTqkKYQC2BLOU5VBMvwr/6fL5fVrmtazRfYbBLPrRI4aJHxNrV84gJRQSsX
BcE27vZvPvlRwm8YkHlBUfjzZ495kvg3QbVsZk7bjmFz2BlYK9AEuVrOjFb+plAO
tK96yDukcoRu5GbVD/hgsMtOeYmrP5beh4mgwF5vCSrOgnQB9Xlv5sc7cmmb5uEQ
nJlzBHw8PfyuaPAzQOLvLO6EnKXyLciw5UDODd6gmnTiF9bDs3fdUrS1j7himBvn
2HA3xCYT+gNWjDkGXlh6zqODsKI06vNUmFoUCkmw+yvBarVnWAAtE9zHT6Qk88Zd
mYmH8P8d17mAAmzTa8iGDKTKRJ7Cz2j1C5oAz9/UWVYx0oNqng6t8uWFuBho0NNV
sLByZrpXFuy7wEHEc4mEoaQ2B3fZKY4mktdajYay2HeQ4ElUS1WfvET9ggPA+d0I
bB5QdkHW5obKYGGwUbACoceomu5lOKgR8qQkNwLbnKLOcFU4URVxEMk0NvzvtXJ0
HdXhtVFbiH/iMmcHP/JTBb3/xqB8uj1GB89OBrWts20VuzbRG8uNhEgqUShU470I
WbkJMvJbDZmZ18Rjnxr7xHxa3QCikg4nCZNsqTET+KjU7OkxAEF3wDilDKAQGpWq
VFlZFboIuUdkXVA2AkpTf78rcirLR/55kuU50BbfAmVetH8r280V0RAx83TK/6fn
lj/SgK5jyxATWpVA/yFnBC87mRnx4b1NtqyEvxz3UI0K+QoUoCPMdJXUVqcUt0Rg
UPSy9+AWH3Z7ksJd+PatSsMP40Qdpv/dycxfwlWv7O6inVIXBqe0pIcX2Sl1jDeI
xvV3hlstFBUnEA7miPN9xPkZLUTB4z96Tjx8o54d4I/SXFtU3gF1s+k+XhHTRRXq
6Ah/wIkTL7fAtRVwFCj1JxXWbQFO/fxvivKaGys+t2MJN5lUK9v8K1AFevFLkX/G
WbBD0/HpZg9k5/Bq5ThW2ITqUrKSHwb9BOyhcQGMBE7N4434yGvULYbIfxBUCMVk
1lj/HoWI/WgMi9ov95TbVZH974rYuYxN5jrdaon5MIsO6FHraoqUFB8mLyi6+Ebu
8y+Lfb3SyyDfkLH9t5dW7bXkAcihY5sFXGy2PcnKAZo1kvkJJjoieX/7aIlEZtWC
/Ff5ToHT2D0ZPk+G6vPFoV9ic9qIKrcLXmAZV+RF/9fZrBJlO1Ko1wsqqGx7qEL2
3b8Vvd33wzx9yCBZYmLU5LkBabrRLs6EdKUtG/asYk2EZjanL6kK1L1TeoLlFyHO
+0BbnbY9YUhC0kVvnfAHFjehCEbJjstIpmkjbXWRznO2dTrcrsgsCX9BROHJDAt8
M7AGV0O2sqxoOW1XNGAAXbNSxM8Dfmu2yAPfXkvbSTLKlq8WBIDriWaovkbfuvCy
bE1ZtJL6f/qdFafQJ5NpI6hI54LqptjNFF5P5Cw+66FT1qHNCGuxfklrowIItus5
alzHOQWyJ/IPAXOdpwE4T4qUFo+HxLC/j1eVpLVx3f9OOV3dtXgkb9woCMc0QUQs
Kdv45xfbbfXEKI4VV4fkkqOijGGytNFkoJq3HV23EXsd/x1/ao9L+QEH18PIBRRK
6j7DOGZmnDdOfxIDRfihdJOCoq1OcKvgjxN3IsNuNbwb0Zh+0PBUFV+5RLvWhBkk
Z478UQUl31mY0nA9zJZ93JG4aphXrN6Y4zvTGgAEHp0nYGBn6EaXnmxLEZYTSBEQ
xluo6katRMuIPJqbV43Nen6hhBfff8bc8dJEG92rD7tB2NFV39Cz77jzkiNx2WRa
r1C5KvlbiBTSUvYcG5RSWiT4U55fb9/mXa8+zWG982MPhIy1pDyxZKTJzPKRkY1X
iw06U+ShNhc2j2gYECScLgXe3OPhRkgW1uUM84Wkws6SJ/5YgYSzzmHiQFmDfiVj
Zf9Q2zjfhQL41u99SzzBpmSs/PK2WbDGxVvJ1BSMQ1M7a6E2UiCrNr9yt96WPGNY
UYaDfQh/brpwcw0qoVjtcE0ZTqsXF139PcfEuovXwrX71E5YZXNsviGmO985K4DF
5jxFXn+uSY7JUQOI7vRkM2co4dU9tW5es3nGiZz+o8SacdfGgV17PFabQVoqVWH3
nDkC+YsQcx+s65ygjVY5xFLdt6IMKQsrDtRJPlqWBrOoYxPvBfsPCFl4Z31N/oo3
qtY2Sf0l25Pd5j+vxIbgxL1XL/Cr+plxlI5cN2dsIJp8vgmfh3+CpQw72AsFvvFn
KwoIhj4zX3b5ltsIeQoIocRRQF/DhVM7Hivww848s3VnmfKT+aQxvbh9AsFSl5uY
hcVOsAD76BzMOLAxWh/7U70gf4orghdW1nrqR5i4tdCGwpEuseJLvG7Rqaq3fQbx
iPVy/rrWpA2g7pwd5jOFVkmEuS+GjAxJ8Lm2LX0H877RP6YCWmbFkF8RHbVQjVy/
kwbdjcG0ZVXrMEx99/AUxb2w3lgLyU65o9SzU8bfGV0dRDOcafO1NmX51Fj6aRhp
sW4iq2poSIF/O482AYVXfBPb3QGb2l+SeYg31V8+B1sAVdDcvC/jekYfR6yx+T5H
Kmcd0iuMEm57UdE9Ws6wvJxSjo4fvQgKAhwdMjJ8iDJGXNSHWoWn+LRJ6g6h5kzu
SXXA7YEvldUQxQDgTRlzRUGLA2E1xg1RBioFB9PWcvcF6P7T3KBZ5kHuTobI4Mk8
3+q8e2p+iFQd9lFh1MU8pvmjhDUUdKCQBVXpscyEf4217+62E4+z2wC6Z5tdjKo1
N9YJm+uNnMGeMiYuYD2mifwTJbwq0wAcRklakJOdS24fZ520Gjhm5WzYPVDAiS/3
GsPgPfpFJkDaAvlsWBZ8Rh9E/ldNGTWLu41b5id7HrG7eZeHG843s8QXXACNmEwU
0HSdRzYM9Jpergf8ALqUQ42frA9waVsmwvcSreE+7kAwZZKEt+2BOii5PXaNR8SE
ppjGo3lbXQCmGJU3KttSb2kQ4XmYRZB2xH0+BAnK4h/rqJw3bc+7yb1iL71TVtPr
/ZdF2cM5kFQYAUD2/HmAZ3pwNoQkc87/VqWEtLMNEoLoc+L4sEOn4z/JsQKxPDHO
h171GIqlWasjnIve0kmcUWVFo9S6jqHzhfArCp96Bpa6bpSB0Eg3IxZbKbWHAfPT
ugNPpgBNKaFe8soWTTfCQuNqWRlBukaIS7QijAW0Vu/M002zkAMP4MEc9cb5fdzS
W0g9eAw8fsMesYBlLVE1GbK6zVCB9RLX+a6Ugto407r1w343Okwb7I/lshfqW/oc
8O2w5H/O7pdivwhWGdkQ4UzXjdU2p4vCbHagMpnKM9I/TSkppbT60kG2VTnuxCZZ
evCoiLc27mCf88xUIEem9hE0HgLWgM2e2umYrdnsRbE4sMvjyAibs/cPQdDttskN
sodIX+52X7HuSeZ9DenErTrPTRl6XAJ7FHyZLqGbCd070aGyzZPo52Ta9VEUpsKZ
tVcoomA5/pH2pMALjSE6zCrf6rAdS49xy05mYHxMHnDX3SVQoAnWPBA3zB2ZAZu7
QaarSkYCxhL3YNuQbnKMarxHB32aQAtydKCwcXPiInp6D48b2fhKAIvTV8SS9LDm
3qV+xYXhH/+28mefHQVyG2SonK2lC4DsLC29aaDWEWyl1ujqU74/xcHlE/1r5S1c
NuA6JWRx+A4HdxKXMEnWHihOEug6h5gGk1g+v57QG7okbjtn4FJ9a+VgiqM21VrH
PzVLymYKcAuow+jlVo9YgS+0Y25CuDz0uxxXVmqRDGJlrUaoDIrkBAYG7eHo2+hn
iEU9Ce3CUwcnJujZUz8PwcufLtHFWYQONSadMmxqSUlsPuy77vwLoaVok0FGgv0n
vxYxMpRqBUgvuuqkifyuC8YoMXgMwF4u9tmLZTONv0HzV/w36Wq5o/FLgJkBm26j
sCz5Kg/UAsJSUeHTc5XIM3ksmeMBY6lSwh7+6CZx4YFdWEBpg6D8WtK+iQhJOWHc
7SKp6VCyt1N24Y/owXpJJh1tBVIpeIh2D30+aSA/EDvW7WNuJWf0TodaVo+tgdAg
qC6ESP1MW9B3h4kg/MjcLB7TInSI4eZ2rnsl4SZ4apnLR6VRz7LBwMYD29X7h0c4
w0xVzUOxHEOgrGU5YdCYyIUoCZDIyfpIj7IxjLK4JG2hsKlPdu4/xLNQ+T47LC+B
0+BXfngzx5WDAhfO+s0uAbljYkREmQmmEJ+HZ0MWnVcEcYzKb9Soy+K3JAZPRply
eUMKyIxqQCQv4c3gfswUtESIuMd9hfwtgG3rmg/GJjuCdQzgKhREwQqQVd/th2d/
cSYpgNgmRrT/skLlYvxd77XV3GkLkTVj4OrvYEg/JyxQEiXSSRuvnwkmcW9kP3UT
UXUNj+2SjwPnzOrn1QAbl/q7hIwRhZ3fGPNBe/3uO/vFuNA6xJ355qtkAiQvIQB0
mxImGkuJXUYxrj4gyNXoI9ULMCOGn+Rb5Kkar0H3V0FRLAkQ2AaCfFXP/6gvRDPt
v98kvJVGUqcQlLpMFjkTa8TwwNv7UiNC4Q79uq3Xx1/M0tkxjzhVyEIxHjp1rMX0
BV6dRjk6WapIFwkgIgbXEpYTON7alKu+Gln+iK/GIreHEog6B3PCg6NubvOeY1HP
n9XksFt/ZAQdby6W1oph92tQxlgaHSzAG4oKMewg59rqbm1Yka+LgDXQlex+r/iy
S9fMD/RSlYix1VPqhs0BCvY3f4FxwlHFXrwksLTi7NDSMJTLKLioj1WW8+CutadF
bvPihpAVs6rVr8MBce3Qh2d6feybpW9im2xqGacbfCYhjFo/VboHjOiwyKF7rBGs
8sFfWOMc/eD4bqiCTsHMJ7LmdTEftyLhCBuWqP2b5xPD5U2cVq6rhuKC19ysn21F
hlNLMy62LlJll212IWA5WyWDFf6CBNjeL3M6ghNxBu9WEYlyywI+sXPw0N07iPB/
wzISPEqy9GgW6sIXQtmXsf+WQL+cQnuCNCs63SVTBmrWTEdUwnSK7Pl8/V84rHeS
VRVmlztcpUlhDaAFrjl/LsWysJlenqrSBhOTkmnJ96ehFZr2A7G3NTEXuzZdONNV
8F6Fh6j8Y7EIsg/gGn/G++wrgJLELtn+jEMH+X5HnDteOFBBoX0eEKw0m/0aTTzs
xPKX88iXxRkjSgVRyjcJymmot4W0fjkXfYM+G5gNYx19K/7bJo4QTvG/guKngbY/
eAdmSwL9CTtWvv4P6vt7u3W6CC0tp9DzSuyABG00Vim49x2HCCvLu0cxW+uc4Ftr
iLEd75ZEqaCK2pCQUpCSuMo6PmPPKx766HU5T315FUNglbUrebywwDOR6eIaSkVk
SCyRXjOMftHANbpeS22Zg1bAmuGZ8b3XxCEpXSrLrgTrHjdY2l9Pk2EAxNR8OcBM
bTRBM6CcG3TX87qRSdjRBfk/yYw7zPf9hJK2lTbPfL5se+GSoTPjIz0bd41HNoEm
2XgRV7HqtQ3YYPaBxqJsLf3oQAhiIN2HWVrkh3MCay1E5lPcZ6DrsY0K4k7MbQmP
5xxYvLGhVE/cgOL3bcz26+tD6lt5inuO5lDiApU0qc7HqaYtj16bnzTBb0ZfRINr
rwJabiqOAXQn01ywjruWdeUWuGFbC+wOGWHkABf//q005RM6bYTsVk1qxVZ3yfG7
GDmnr9qEpQ7ciZvA6mEaYJdQY7kmWpzGSTLvSCOc6bM8iZeS8J3eqonByemw7QPh
PgqLRJRgXokwZT7tkupuywKyRQKsNwhrZ3yAGdxkH+8SybfgHzm6sOCZCOpBd4Rk
ddDunqO97N1/jflngn2O7AiuAkX6nuwjQl/NQHROcxylwAloJroG/xtsBvtUbQAh
3YFt0nX3NLmxl6i4dovfps+8a/jxq0JWFG4EQPBESGDbeh+zALNMuZ7+6YbaeK6Y
AUY+tHxxtgQH+EkCkT7bb4wG5P41vOoMqD/Uy6cpD/yudmUM5NQXDvPnbfoxH7fJ
++jHFA/Lwifz58jUH+VLH4f5hOxA2G1Wboyu1ZLgxuhLcrK/CEXX1RHpqJBWx0qc
iMBbMpp8XB54h8LPoajk+aOyr0BMWOyUXIwpnHBRrnZyZtnOu6NOatfFvRW73MSZ
yONQVQCLd6t3q7DX6Uwjj6xOsFu0PebwyDrd0wa0afAO37g5zRvgN0DW6ksKwJDC
TFcOUPuhYmqU1Wcc/tCReOsA7mj5ZZXni6wFI8k0vR7i+mL+wm7kpLeYjKXf9xEQ
zQxcS1bcdKbKIhoczjyfq2eHC7j6drsTNHkRugRqYDQ/Wxmdc97KVPBncCctQ8A6
MwQvRofoMuyNq5HCB1pM9uRsqJER7QaQMrFUojmhaFZvSw06A/IkWgWKxgY/IDoy
s76X8wt5rddlY6sdn8k12/4PMv5lJLgrENN4pPdwN5MHTNEFJL5oUzX4ohaU8nHP
jqGaJSMySArOaN+sLNAo3s55rzTQtNuyPtLCJ/pt1bdtu6HM/iZtTnSpdrkPYL/L
9kz19Fa7kRn5zE2qeX2oLDB/P8P2kcqgMgdsefuF2bxnQEQRzI63dIR1bcvLhSWW
nlkV9T7Bcw6RhuckRqPR7/+apEjdecGnfySMbZdb3YPpk8y34+Oku8OKIEjrxLpC
NZSl3TFymIHHziMdma92jkVUG9gZGm2H/ANGJOR6TCxUj8v3HOfWf+ozH+bT5YkA
xampMsbeHpP1AISWc42W8Mi34JAVRu2nA488ieU5vv5ShGj2p6+C0Zukego+Pixe
HPHQeLsMOdxZQTP+UKO4T3p9Sp56AjQmVUTUR6Y2uVoqpHZo7R6qGKqKU+sL2ETJ
`protect END_PROTECTED