-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
CsZVfcUQEim5fvzcLxf5uZB17yVaxzjSIFAhrn6GeTFbLXae6QTo1kl5fFWvy1C2
zV2wj/7agQRv4i2kPFXiCCKH4ybP9AQruMP3NE6EX69cd9XDN1yJ0vSfqmAQd+so
o6yydlrqJMQs3MtTRYUEUP9Ljde4EAWzAT0jF698gJs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4200)

`protect DATA_BLOCK
rpMsZS+l20ORyLYguPSkV0JSEuIBASDUu6KWzFkDIwgUpFojBqeqrQDNpUeLazXE
ffVQU3ACQ7Ug8Ykkf6xPaGCpoUUFVMFp0+TSg5/lB7MB9q31ZM7x2+6HOoSG/SBs
9Cd65EEM/IP8nUxnPtXJNjB13WZJImsXzzCHq7HsIT+vmWIUjMuFMcN/09wAyvvo
4oq6ZIEXJdJolhdhMjCi+ztJRf1U5CqflvkrJqAerqUSih493+7Jo2VkHeaRlFQA
BDyUvoUmNxSdaDgQUH665+RPAq19aZIJ4jp527KMeueu0p0aIc5yftAgzH1/Zb7O
SNUlq9BAcSXEcrLn0ypehTyiV+Y7vZmOTUmhHZa3uV5ZGbxv5wErZpdiAB/7Shve
Rw/XiJ5eG84nbQoLt3XXTZqVLOh8/2qoNIQHnBXnY1gkLhDNMaABk8VLdHV8MMAf
EC8U5P1C1BXwF7YKcFkgMqH9xxFEIJCN5mex3/6BpMpqLK1S+0pf41QEiAYwIMJk
3AiSvVueZ9U/5SVJEJrCYkBDUC2LxY2GsiO2UGy1q7DGJRrb573rBv80ZiIENgee
n3AyxNir+PvTyAcZOo5VWVt/Piei7K1thfKTH48UY3EQKyzeSn4ZI2/+dJoYLlMU
u1K9miTuzQPb7AY06CBnHHmKVWRRK2G3bwQaE+ptoKULhgw/GP8crsvcb05FwpRP
Ia67kGD2Mtaf/HhuXPv4qce/F4ool17USFozgjjam/0XD8Conqy+Cac8j6Wra4Xs
AVloboSmBnmwZEqWDUaGaSLLlm29R4cpOToWjpx2lREOEEq5v+Fv3qMAT+IlYdvj
ggeQRp4gDWW4M3m62ON1LkkBGiSo86D9KICihqeX2CeW8ORecUgPsDyNcXABuvZE
TYHMJUBhF/n7SXsYpflteNsrq2edHH1IpFhJiS9zyuZVrr3jQbxScvagZeT31q8A
ijijB2YtVkUQDOJOfTdPlYyl9Btl4RS0XVJ8sM6tzOp4agiFMCGCOLEroto4BHJw
qhsiHY3zu+DChXjInc1FxK52bcF/F5vxrNentyvLnX/iepHt5uessUiu41XQM3zw
YERVIlwDBJM18cSgoYNxv2HCw0LmmAAUNj6IjbPjYDRiq0Mp6CCWk+kn54K9Wk5L
mwtCIgH9qz7leAW6GJVcAS6Veijmpa8xI/bSjhHyZFY9n1yaTNKNOuxFFF5UkMZo
XlqYJXcNxD4FhFxGb91Gln9dc+P8X/lY9jXj4wVRAZ+/OTowX3zxWcgshYzJWam5
FnjPhpciqBlM2oAT/yctoAKXChGefNvn34PLY96Tagt0+QVgGByQj3hNaRk+4kzT
H7wujCWS+6SqdHRMbD+ZBOMXS2pTIEWzVBnLRpGPclAOPsb4VLeZnS28mzES/GgJ
BR9Heue6R/BgsXaVBCSj/qOdRaUYgcz2kznCr7yaVgGQrXF1eRZlJ/zW3QyIOF0R
qDq4nh5UlN3IU2CqQRERV1z1w1KZy3VsoPUxceu6tFl0z3frG0Uw88DXdrtU51bO
S/l0q4ZzC7f6xfGIEBCEP3xhjhbJ4UVVQ9kdfR/uCcQlejVxThVSKAQYBDRPGmE4
jps9UNKUf8sDA3YDs/u3NeY7QPMchSXW2pmTifqo825BWI9bex/C+SM1rYABnklc
hsh78ONIkaMblfwsqvdkNvo1Ad4EfvKhIWEpdYs8+32ySXjaVcX66FmPcxlYXnFK
C0PgGmhGbzuMuMLmG7cw3l6uyChIGINKn7bOWpJ9PdNwITFpeTEdNi7uJL5UN9Wr
rtVPX7DZtuhh8Tw6Re1hCnzJVOLfVkyUuXX1vm8lSj6xrOLeBysxQhgTW9QsLNpy
QhL8RLfHUhQl2O+L0fIsDSPC5Nz4aFNYr8KInun5AHsztrLaPhvZEM+qqJAQA0oh
yIv0b39trR9hPJxjf3qPx/JgkmUIea4I15B5T2Mdo3FOIb3sZ4N+l5dzN91lNOCM
dA5qFFZMGHhGZlFZ4swabNs8PaKMFtXNvL6/1yIOijY+VZokcTfxQ45QerYevbVP
FhpHKjhH9ex9hy5+DyyaR/ggHEq3aUo4i0TeBJLpLN15HY1oX6i1XAAMAanW4xUU
HVrygSjaQxQgzsnre0Bh4Ovk/5ZL0h/TRWofWCzcwqyeopBbEO/J2D66sbx3lT3n
/SexGprJNU21EbVFkqWdSwc9z2x0//K7/BByoAT6vhCL35CLfod2/UYcOLEAwtBa
Cx+6tF2deNMHyK8DVf/c9y0WwEL0Ae38AJHMX+qW9Acfa84ZkUotgKW1OSfjEHsc
YhMPQpXpr3ycDwgueN/yoIHP5OxOSJcYg1ByyWPBTmm5W5kNVIlyrmPJ9aXZ5VzZ
8hz/2oyGmJpYa9oOibGU/wkGfL4ZV7yv5HlBwH1hplH0vdEJ4+F10Z4hnTLSNVWi
uBinKrpOmBWRVxL/vuAUoabZ5Hz8Bg/vowlB9fuGJlSzpLEyEecR1pF+7beL+HDs
b/G/MfXWAr1KI9tg1NqXBUWLOG362O7+gKKMNuzhW4zIibOgh/H+F/4kcdo7qeH9
Glu8E8PqCe9pQP6PAw2UR6Pkjc4UlrnMH3/yoBKn8vlimUAaIy3ewo/Q3AF0HgM7
hpVdcit1KnzEpUavv9Ub+JXtBAeaAE8K1fkstliogQr9fbgplFBUhcobFwUgyhd2
9QxQfiTx3v5uDIVV/I1IvoAWakx0jwcdEcVREmOnMeOodKsgoQxIkcwGiSKKH/Yx
zK9LR8hfIW0uLdmAt4xvNTmodPnw9lw88euTXwj5V8K3hhZ1EBiTaPi5jHYAj1Lx
IsLm7mRli35GkA3KgRFuKGklAdUpgHgdpIhfJ0T9XB5bCVlkG4rMh6k7X24aCrL+
gpHDOTsKd+umubVTLUObUIiCzCx6567jUTb+vbv0RNOUacQZWbdIT0HLXiQSNh77
Q5tFwEJWdLPRSCB60Bb1K2ug/Dafp7s1cl+BREBslBG3h+rzkgBQyeIt/30C1x+/
evxrG12Xc3SiOjCkppeTqtSG6309jT620y5eJMBEjq/H3xvhLYJKfLyXa0rg54tr
JQ3u77hXtVqb3YahwCsckSV/TciNWcF5JWsoXWswlWm+2S2vaONefpRbJ/wt5+Xj
TuEjdVgD9xQnN7NTIbT2e7tsWu09BYWdEN9+3c70LpurvmZLeRVQ1DCwNOWyyEvB
v8oIsAReWJTw3aioUiOSrC+Q0FCPaR/9wyZp/s9qs4OzxbHs2dl6kSxleDe6qWif
M2Qq/QuOPfaTQmNfiBFPcIqs+r3xjsYYlyqB5CXbHGqydXYaH+9B4RRHpWW5gER4
rOUQPhKNeDRqds5qpYvjccfTj6ui6IDG7iC56MWmrQ3qKDkqPFTNlkz3E/4+gu/8
jPIoBjV7sOgiZI+K8bwUWoTYGZAuvqeHNXcERsCrIdca1wM8XYwHzKXdgjR9kr0S
8G2za76M7sBcJMoOOS/XlUkQTq5jASgP06PdNEEr0ya9rtMwB+mt5GKAWbgXpY0g
m5kMrbyZku8/fEfVDyt1xEb6IyPCjEwSle7b0hD/I2XAqKecd8JLD2m3PJWuC70y
geMzY+4+5xqSeWswGCrja4r5uAyGoZdDy6VJz+iQzPjpNHOYlVg4qc0yE+Pnxmkn
MtpD6QaPydUmZFeF1Apo4B1yNIwo0AvUukkdaFNAh0X7tp93u0VHa2OBkCDnIPzA
hgKOnFPU4KJ7FavHW27gzOEsObaovF6j60sV42BM0DwKKqQ2MxosF+poE/9bXaeK
j+MjkO9aWDmp7afNfeVMAPFja4fNGZx6wu8/TBwGJtM4d8ytFO8NycFyxzBfkEw/
PhwuPu9azwc6t19kH/Twp+uAFgPmktdYqenqol+50F/ShwLh+DCrYF0QYqLarI2j
17+/DRrtX/ONEBZyywZnI4OBQ6bLdRVPSTfr9NGZvmtaqbve8L+eTM5xmf7tmAS3
+iXNh3R9/vkeoxHpBVL2wbz7yIZzKOfYJzByCtEbkO5nrPxGL5tDFfp1ynLubeEd
W8pr35tcdNfIVXDGrTE/pbXYTc5ng7xSS2mCHDi/FNZk1fuI+46kDGEThmrMvVCh
3XwyHOnROCNfeFCGcXdzhYJeNQwgOdzq4M9bhpHfFQApyxNabTeFlfjs9jVbGCZS
QFg9JIkT7sQ9zDkql0FBXf05DuVuz3CQSFzGhv3jDgkMwSMNg3xmTI2lQX5E3xdp
Hp3TddjbEkEjSh5DQFh+puPTv/nqVjPGEP6LWJYH3PTWhRoxKvBlRbGKX8Ahl0Qv
9MFlX51tR0I5e+qRck8ZIQQJHdnVjoAAEHs9wKU0h/S3GdMMV4HLyIvEAkCBcKPW
bCpp4BttPn0n5jQwv3xW52kRNT4nkQ5Srb6iT8BDgTqVd9N43gjTsnorCQoNqfDD
N3yjNF0AMz7UmSVjNuzfrbsgSqeTAaMjalCWWnOaZR/mm/xhlQF8XLe0E272TOp8
oGvWd0UUvChN6MFXSMU7J4j/Tum2CQ12Rlp9/8Ew2rMkcsQMFVsfLPSdc5FFuF1p
QKNWCHIxwqW4VCPDGcS7DlrggcOROZDFqg64zEZiQSJ0z215/DCBQ9Xjr9GDegHH
0AdJAK+wddnUuwSwHTuvZ8zjcPFqOflNAfxC2bhBena/qKqLZi7FlRseXhG5xcvj
naiUmH+QXij1QBuwFI2ERcYwIjpxjZV2fBYaY6yAW5zKKYuaSWk4npEuMbpJ4fnt
nk/apBgjowGsGTopfp1RAYI86rCWCQLa6jt4trsujiDNCel/FSEuSB3abJgTEDVi
R/mXj3rRKrmgm/amdXaTb5vjiCrGksO8tOMMBR9a2ET+zRcti+4RhUrfJ3bW8xWZ
k8wo7s9Vdx28Ftn2dJZFuOekN3JD2qoY1ifBrNcixo5/uGo9XJh4ZB/49VGqn9Nx
8wtY+rdZh2oG3udVH9mXCp0syB0FWii20+qHW1evcaR8XXXRYbodGSlzSPJDrkDG
//0jKsgs+Xw/pEF6k7VexAGkLxhZj+vYdL5fYolLLsFPtAFp1hEs6TI+Nfr6k0kk
5ijnC+xzTk3fCe64Ch/M+CaQWLF6iWG/I9zEvcpg/9gSqCdB33QDfOD7dUvxmgyM
PfJgstWt45wKqsS4Ub1tHdd0IDb52w4pQ6E8ZfTVNOFEJMNk8okbAf/U26OUj/96
IQpQre/yRIALsCv7T/bGviubEXUJzAHG3Gf/Mgr7iz88G4m2Zc9XNgUWAkwOYUgV
3M/sujFrVFjd/aeI/dLX1WfcbXgDYa2Sea18Lw0n/jZmzGpWLlNIgj0vBXnniNFA
j0fB5xiax6j+gzro3dLabd1mhj4LnoPDNtKdZVDRYVv/ocQ7qJTO7OUfl+OTX+Pj
hCNbWxV5V28+mqBQj2iJYTjyunp5iQwWlcuI09dW5L6uPKVpPEXkfQidYgh50Py1
DAr0Ab1SfPEcDlRPOXxeQ3n4xZP18ccLLeVFg8O+XlidUz19vl58LBGHp6jZWfY9
uMbiqEMiedwUtQCVbn+cKYl7YER8pO5Va4edxPUitpd6XdWwdTgyxm01wj75IZ3X
fSvZx1i5C3tRvv04wBJS6nhLnhmxFjjqI+0idEe/sKtzcFXaGZ9WCkf4/bTvUST7
`protect END_PROTECTED