-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
EfBaMpxX5hs9AAT5/h0yQD9fmcCWyCfvv0OghP2mCZEqBIo7v8QsleVZ8THodzXz
YekIwiqgm6Gk0o7bt4lZBQbk5nnzw1KCJtXy90TQagKJ4btwwxpX2H453qBleT/5
xzV8nrsifIrSSXvudxaFuIdIW6IB9pfpmpso3vNnRC0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5408)
`protect data_block
YG5Dpuh/sz1pYcR3/sxbKdfv4ogfYTlrTe/zoDsdPhaJzx3+nl+ukVZ8haEtPkVc
SlCqNLY355ISW/hM8dAjQNj5fzy0+Y04sUdXXIYAaaOznzqXoJfc1jR3Hb8dQQj4
A9v7HooZedAiCQT7tGdJewSrpFYLoGEtiSUzJh8RSHCZ1SpKHxuYBNuyrCkl8bgE
32O/gycmbWQabWcuBPKOegXLGMEUW4MsN/eOYmmvDmZ6PoslGKlLJqEnmwgP5fhD
f6MWqpYbGU9NPF0+9sb2ennjKn8KamiSbVFgznJ6w33iFi4xvi1xctjIBLx0hitt
nCMkIaWIvqdcjjFTVAjmR0PkSZGcAbWqmEcPpZzizVoGfyI/QNn2LEzsGi/NA2nQ
jaSsFqZD9AZ/4LGppc4uK+SbO92jKkmPKYJ7q14F2r9Afu7epwx3OfbHsnh7zFzd
XJfyWrF4LSsGCkWLzEeES43jkjAyAqaFIx4w37+xIZGCkdXaM62o4yCWmRQK9YzL
+CDYXhqp9qbKGTf8UJ8aqavXldk6UyxWTng91szYGUB42mah1gXZGZdHyRJ0zpzK
GxoYICAxaEFSI81Zsi3WSdMCTznIUiBb/c1dzgwFl00UJXHhBSDlXc1K+F9dH6jP
Kh2eCqIbrTmK8i3t2bBKjsp+bn0cGfh6kyQ3ci+iHpIVYeKy2Ri5ONJDdlHhmlcQ
mIUMF2ECA3ec7tjxXjvlB9tmfHLNADJrhaOBvnaVRdaoyC9SZjfdlhWaeIY/zvYO
JD7XIIPlmLsaRDTtEGJ3FQK5NpO1OwftiIyug26UxIdXGw5KaQJVexYP9ijLNles
dJAzVEzO75DwPQ+WhExF8VhHkze4zyer01XDGBsmK0uDl9Rz88SChLN0on5AkyUY
0i6YR2YE47nYK2cj+DCNQek/tNr50Re5Q5b1JstEbLC6RrmLb7/eicnUF+nyhguB
POUeyFaYGhEuG/r18PVDa/k9e2dw55wjn63smrfgaenemWF43xIUfd9nj7L8hCL7
QF99oEDbt8h0C+6wfK8A3qjpNG+BrkWPkT/DKzrNxX0QS6k4RN1NnjXooxlHIVW0
oHBhC0aUEoAyq0otqt61az61XfMhdbI7LrpyBK1APoFsFe80SYKhzPEY/KL56JsK
N3pbM7a2tXvzv1c0EpDJlMumDlAh5MWkZocBWNJTrysbhDKPbsJ/QvVEJgiSHCff
J7u9XoKsBTiF0YHG7+FR4YcVS2XvPf4mQPnHyd0/J0RoyhTmzXBEk9jX0vKE0A1E
JSnjxlb4rvNQIz+ID5IawOl2BZpBuAaqrfx5lBw+BBh9SYNpcfTUwFsY/t/ywjSb
s9QYaoo1lVKThhe01b2hdVNoYx+zSDdY63hWwpDwPkv5TAVRhR40TV4Vi3a1MbqE
APhbLQuGtCeOcGl5pJTkNySyjotfHjHHW/yQ3XHPWPZy/mVTEXCfJ8FOe8KRJFf0
rrqxUL3ObtFY5zCoRjG1grlLpo3ECGkX9AWPItFHbup+eQySXeean76xRJ+sMNhq
0dKiSXI7lRa69WKCuXt8gnl0Jxq7W4BdnMOe+Bp/QIEOgZzJnR92ox0a1jM2szG5
n+o73Zfkrgfd+OaARu5oih3D+w86mEAaTJVZLu7xDd4K8fgwIlKMohkooAB2RO4O
jDSgTboIY41M/4gv2+86AQsRLyBVGDYcy1m4K3I2adQ238P29b7nBGmp326U7RR0
daygU4P8SDBSIA4UmxGIAdWl5YgN1mJ8bV/mn2DXoTOQleVWftk7uf8HXllSVTjp
2dra7DzalYTr6uGAO/ZUj9mmyfIPUc+6Fpi7nc+mgrS7RRNT5SGAPnvOHRPNMWvu
cmCEsWngNbjiDMyK0mmJ2YvlRTF4b+JeGXFqPdgJB/Q3dgA6DymWa7MY8ZhOq2OH
84fb8A93C1pF7LdKlQdHq60v7xqOf55dESoOWYfLYfKabOUImoB+21DoXmkrhSh9
NWUBb83VHMQnWrAA/f9g7PxT9bYiU2LFLdpJWiWnWpzvKqpprZRyRhr8oLSkfXEY
8khpsjUnEuQt01UFhEpsw3jpoRgBKFKj4icgdIRBavbAzWJxaGSYAQ1SwH1XVcGR
PeMjE7VoFKYHuYPo4sk8eQkjmrs4A/9vNfwBeZ5T8tPgNwgC2jXFu2o76MI5MVQb
O9bZYe0Fr+RknrtOyBFQTZFPf+nMVrcT3g2cGyBSCKZfwyYcg310RvTrvWfe2dq3
JBJue+i0EWIE1JtRhyOvBgxTMXgb3ODbR3hJ7Scf6B7ApgLoXwTcmTKKpF9e//up
YggDaB4774bF58MoaMxpppVWPC70cKNWmWyk6q0Ocg52eOoXYmXsLmYqVNchi5uM
/Mtht/31q2DMkazlz3/AMcLSyOrsQ5PFaZ1Ruhd7cxX8p2d5wm6fHOIsNYNCwsym
G8HhXKMLKm0wjawgXGMuFdnfB1NeDTDT3E2S89WgWcbjcoW7YClYsphUw2rls9Wp
nB+FDgosAsX9Bfr9wRerkJJru2ESZ4jw++4R0RNr2/34Cda8s93722CBL0L8Gvia
SXPamXSMw5gRXz775AObT9+TzJWw8uTRZmeoiqTCrAxR1JC+Okw7Dpq1HzYSrWOV
UwRpqbB52+F7Nk11egmam1keLFTUMFfmltrnTS83lI7xMSTO1hnl3vWLF951l8MV
+2vVQWC9SUBFhElBpiz1H3EpTHeyFeEe0/xMJsMv7RESsKNQXjjH4UOr7/lq13r5
tA5+LV4JYGAj19oqiJjXisA4KkFhXMFJqfvKb3dk4jsR4cfuecIVE8Q4eiMezl+5
1021ppRMSfoyhcr2GJjCeLL9umIsmA/lVahpQSxpKUD0e7ooOcdB7+5NP25Pggzh
91K0cIac3ERiDYcOpCME/49QN01bYVXX24NZ+bhLZCpwy6bSU4a+6WhVlRLka9hk
7ShAWMZQ9fLCxIDHT2sRYm1KT972j3FkFGHdw42KLVWmeUAgdcpkzXvP/QkMrMsj
3+twqBHg+nJFu+hNNmehcrTQ7DfVklYnrRPd033g5FyKqBGPWteZNV/2UGVDnV94
giNg9RQ3hUEH/795gdrf9DH4ZvF9tKSI1AxcXA8LFLQBzHvaEmrrPtk31J73MoQ2
kavUlPGnEpY+VOTsOk2OuM8mCQD4OUNZiABwVh/A0WpTANmatixfeU6i8Ihwe8tV
J+d5EOvAdU41TRutNmdJkiAekuMQ9tOqYaiq2NStZlNBHNQATIXa42WaRfSL2FVF
A1FPCPqNiW02kqLCbIq8G6dSu4pnvdRnMijY86g7r7ul/dvTTCBmDSGRmiLhtpax
CDMNnNjn3MSlEBt0PDBjtrGDQgirCBDhvPVcPm49ahMaEcxxXTSI8Vhb8mpxGHqk
awDDQ4xe8+8W46uELDQ9jcsz7SJXLi59Zjn1nkZaiVFrYpI86Ig2igbZScXWHA+K
h3g4ax+p2n/PermCfCTBgOwkn5As5iTdtw9B+hARrgq++0AIlQ8M4cbMyEZVR1yA
hFzRM0RMeEFm+/hke5tKE4Klw4sF8MYYudxC2LQgdfC+9fw69SwRY+kUy0tXyXrH
syrJrmpA7lw/SqXW99O7YtsZy5DQMb/P5OlHSSdodsKjljmaPNE77/2T6IL2uQKS
MWWDla3ryioKdA46Tjg+W1BrDyr39lAYQ2j5WX6G/L6QLVlVpyrYvXbimMhQlTrX
GhFZ0xX83L6rO30iDybW1kPy28pmYN545/8mt1Twi5M5a4O/8fTbAYnJSXRTn/mv
L+xBRMrEFiRmIszFiiUwELjK9ZCG9GzTkWtVi+ga8q2hD6YSBNO95+bYq3oRaH0d
TKPddK7fw9aTFyrWMyxmOPMf48lPb6GJAEM7laDJOeBrGroYoxH6DIyJGgGeroze
QSwI/1JrKy4nCY6eCfwlY2wXUSs5NTwkvPedBhbyrSBmNvITjOmvq1JloJiXwZQG
6ts3TA9nYALmYR0gRKadqLpE+NnrKs4FeMEPA3p+c0q78l5Krxfs8zbIEQzYddO+
UMGLxFJ7e1ZgxaQRZMxHyqjT9bgqQaG1Fk21uQ3/O7KTSul48ToQ+5CmCWvyPZVK
t7zhLlyoR9DbW/w6KYEOm1A2jUVlJjZVwQd/9th1KAhAkavhK8MDO8N0cCo54NCR
qUdPp0KkoLA7yjysxab0Bx038riTzIaDxaaSGfJ4+dnZqYPOJCKZBq/84vXM5Vh/
fJA9Noit6k2ncUjtemGvqKSPYOH/l9Czbs9DPbg4WEp3vMPhjrfVm2J5lvmZHWUs
4GnpY2iB6xzH3G0b0NiLYD9ubb/hHbPgO9mZTPHdBuJhDf/C4XSEO+grjGuE1kUN
f1tOU5GftbwFniJKe+TK9UAFkhPf1C5ldr6Q+I+3qv8B+AZhjEM/9AEccMKde/oh
7w59fih187GoEm56Do4+GIZyfkxfbZyWn3dez2IRwBm8YBOIn8IU3MOxaP5NF/Nm
eug1fQWvY1L1/4ELDChrortCViu41IpUzNp44Vp7QxIAtxp9mteyCM2HIo9Bkzda
nWWQQVvJjwj5df7gkrjfpLswa1fPZ19k6wmiYebEIGIISbAx/WSasw9cVMRwIRvj
Z8pzNakaHQhgfADT+sZKG7Y+lac3rv2NKWm75M4yHsl8hap3XOFhKwaazetSzLXc
IhLRt66rJTeLB3JXBkgxa9P2GpHM/3x7RItnCsYJnXuGfOtPDM0zrGA5lQmtWVTz
il30qHSUOizziHAdin7A+OHts6ZpUwpjSHAGbRhwZeNnMnS1TUgcBS4YZnfcHyF/
raJ02l2kxHqHfC5LK1SZ/dekZZlwpJZqBC8LUN6DwhNk3tHIsvFt1emmxLzcKy2b
jxoOX265c9PJfUY7OwPruPnUrNBFac6ThDox28/d6BDsiCbpOkm/sQpC14i5jh0K
lFw7qfPG2J4w2LGrAaLJh4r8nnuCJsLNzh2MhD6RwH+I4LKisXjpGep0D4mLLbDF
GpMMDlhpy9sUOFbaHMyI/ZWGhHi39n1NjaFVD01sUOTntzF/a1HE7Zuv5fxolRjO
qIovMd820fiv8SZui3j7ZlJDQsO/MSDcM4XwmlRhcC4RTyjzlayB1P5M2vjJxReP
HZg4HVb2KvRkukhz6n6nMKUcqkDqnABE63vUw3yOV0bXkC6hIqm6EVQsz0OF7TsL
xmCB1n/K9oGcmtSsPKrVyBS3GpjsAyQw3z34h5p09pBQ1D5cu+7DYYL/2l1iahNk
+CKC+ztGYirP4cLuj0hmsd8NofY+UJJDEG4hcUwzuTQrSX2jX1Rvz4anQEf7D+X8
aYqOj0g8ahc8WBGKfDW2ZSGt+YffZO2TDSzy/lglAndJmqRf28kupyj+pWdIa+oA
RkMAVvXAn+xs3o4HI7KPBsQxwszqY/s0WInPOiGsynnt6jGBftuX37SbEDXcNwYV
kdwI3vgiJOxscFby4J1Mbq+ee7ZYy7kp0CjnnYHpxRtYEYxy0d3+WD6DHzna+akz
MDxfGIdDnx6KTNf/8F/LCmFIHXoKvBL9dMFDetRtgw+kLOaGyapijeQBbkHuj/7f
ETgVmaiVFRA4h925U9U/uPVjK1+i9HhspG5+uVPbb9012pKeWQPt67KfEpXLbNAc
7n9nnGp6wqn9Ca3BlAwr+j0OAwxQZmeg6P4CaGciykbD5UNsBetq8wFf3Wbun/dR
+aaSxLzTrMDVrWiWaJFmA0kb3t28gQA2CpAYS743FHL+rJ7+2RlWjFNsLyRR3dh6
I1g7sc5zqKB//amTDDcozfxIG6Cnrvxi/zhTYn1bAWYbWd3jpw3xlbNWoMuZRzS3
qc0fWInxi+e79vVovyP6YtbVUmSgOyQXE6wUIJ7FHPkO6M3JkS2p0xhtVKRXfFc5
5QnQIhPkzJB5E3CWVbcQRIkKWOuzY8sWh/wv6pCm07m73TxaqxvG5WJgL/++zFW7
uxhiAEGPUuSWmnL6GzbfPcAhRfia6PUF14Eh2ljU1YXaiikvFZWsbvT5TK2iaRd4
0gBmRISmhnTqjGo76+9m4gZh7JTkif7Md8NlnoeyXk28+9pOmNBPOzWkBJw0RfWW
dmqNX9cdZFiJC/r6KuU5zgdgvzrQ1AKUoihO/ADr4IiND8qGMX0IoD/iO6BhLnlK
lRmig0wBFlqfL45b2PQF/D0xdqQt9lwSKuZo44bl569sopmDjvtOO7kc6Df2+HVf
imQs6X2IPF+XlqWFUUkuUcrxubWJLdjRME9ilr2IPOtVgjohsUge/u8hi3tVtMok
kLdeHgoW7hJTQmW3GIO7u2UivY88eU2YGFAdRcx7OZML9Lq3KewmsLDyBnagw2em
YK6KHCxfXrF3Jz7olptAbpHNlX4XQH8ZduuG2CYqq8riNwgOCnIabYqmjpVpz8tA
8rtg3qxkqLXKtMxRO9bZ1/WwehY2qpbYwInY7h4m6aTfII2dQYIwb0QQzNV3nWQu
IThXypZ9Ky5LPoVoyCzY14Yu/7cF4eBBM1pakXk6f7uB24AKTnmNTZ9IwfQKP6DB
MvClK5mWS/N5MKWEC0GXa9amnJZCr2JDvTpZj1zNaH6SbjiHhHJn3a6T62RIVP63
hV6chaISy7pZUkYol8AJDzUThvzSScfSFqr25xGVucwwzTfT8l/yAvpGLXzbcpS3
ZF2cgif8z+BySeB79MXw+8E6YQGJSzjnEPxgF6VPllqej26udv1ZHKz2kRngu5ij
6orBbTpUHFx81Kw4h4SIxynA/+7CjVJ+TFcRAOR+lKp7G0EbOl+tJm8meF6tVfNX
vJ789fz3ZckPWtNsGi3IULxuBKOwMZudc53r+pUq9YrxT6Lq2VHpk4pGfeHnV6Nl
T59CbXmMbWYcyAPEogKgCg8Dzle8ZVRVERV2HozSEdMCi3yE/XBnVHPKvUS2dotj
PfhBUNX7FKuwhLBwKeoXgZ/3A1NMQH4Nc3V8r6+DOJ0QZV562KaQCsg7RzG2kA1p
Fjw50v43ZhhsDibbEpjzBdBj/iU7Q4EuvjZcE/mgMEFId6Ohm8Qocj/Y0acoQVP6
DY/q8vbW90uPM8tYA/yhB7A1lvIKG3t/hXrVUE1iwpnV0Wi/6kH+YbXDTKP/Y0tH
VT/NKCAeiC+wT+tfQ5jE5z4wvUYAZFfQrbspVC8WX2tgI2JEhPUHBcTeanlwx4cy
fAwIy23i6RWhgN2wp20P32OUPyVlIN50ItDwhbrFT8E=
`protect end_protected
