-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
YTOsOFPT8F12vOVipgLeESqOjdZsJSRvOCm4kti7s/aqy7oyRNDvZ+zMDcLKjFqH
LLV+M1c7z7AbnUbpMeIN9b6nuNHqEIPFxv062z+9D/q/BdKfBMmv/Gx8dCfT50yP
tCyKRcrsD0/i5fQeT+dhtJvT6FbVvBz51SIw7PTxKrNz7JVpTDLpJg==
--pragma protect end_key_block
--pragma protect digest_block
JKYKRENTeKthu89tIUTCsp4KkBw=
--pragma protect end_digest_block
--pragma protect data_block
FYFmTFB1O862aPTHtRuOUuV3AMWaQg7rrpjY2/BenZ3w0HbG3+aq22oBaKIO35eP
zGAy2y5mnJ6O7ux5x/DzDs5kItTBKGj3lx1nmLlKz7LXhr6l0+EozJr4LDnlqma8
KsZRHgpfkkk4yWBJrMljxcbNqSfTTVVF1v1Qnk3mwXhoA2uTTa8pdXOmuaqQ/ZSO
OV4qFWGvOCGYNOkuSNFZUfb++NWF3XkQOpZ0C0ATBj314MNlPVgKnEgOkYE69Jbj
DhV2oJOsDf5abDXfL59ki931pSuLB2fRJT9B+beUDUJzQcyb2tLYyKGaHOimPDyc
ZouaoW8DvImMPudEF9hS1OAaiZ5wFC1cWyzJiOn2WoIREh9Qs3Y1/c3JvmkEPdBG
b98h4VqWgZTCGqedFmm9g2Aj+5djrTuOn+fraU2VM3SPoKUbiTOQ726jzxBpGweG
5ph/nHcILEpzEiXG2feYEUsVd7S0AsZMuIjA3hR7mi3w2W/g9IjWinNn+xzuxy5n
5LwK/vME432ARBnHFP+d+xpeWi7jm9mMKW3yMKZx74zFlwX4Ys70qlJZYvofmUAX
5RTOCn/U7ejUk1L4X8yH3P10EUtWZek8g3bJflihcdhVgqRPQzuuN7jHvOKJxB+t
ZbEmGhNMzB7f/x2oPox8qcRh3j/dcAUAoAXl1xs2XcxdakWXn6kTYrXKLNVmq24l
nhZv5mPo20F84hNFmpxk6ClI2S58MNIDVCT35bBmkNAQBGC76NCMagJ+gCCGZJJS
eqMzFWDS1fFSOyFHpdOLGE0p/JLx4MIekFOzAk3Cbq3HdKB9DCkwb2FaoUnBxH4A
et/ykcmfnJ6/s9TPBSsMwZ8/Xf8I+yxhVCdy/wrdm3wrQKmVqD5lLJGwzX83le5b
Gkc88hGTYHkFQEyz9XQ0wToZlp6A0LXiUY9wv8i+Fp+DnvafLet4S9sd4qJfVdoi
cBRgR+rxPD6r4z7Wtr4+Hma58vcVy494XO+/jcTgctcwmptjh66xLh7YDYvOJ5wT
K6/kmcymyDlqLv4ukCZzkP7EbWzzgV1Gv1tBe5FxnImV8FKeeiqtQJ+Jyobl3Lox
54awzbYLyobk+M5a99jre5AYoFPmKG85CoG1KPUJupMGn3zttnRRXUDM0rELlK6q
11rkuHiJoMfxMJF18Hy3+EHHrydmCFUOMmFF6JglbuauRPOkpgrnW1mKl6DXSa8E
DoEW/r94iCHDpz4AHfZTVq1ovCH82nfvwTnDyedfF1ySC6pcevdqAvy+Yv0QMFM+
gL5X2NcGPy7czIYRy4dr6TNjzKeEUjfiAfBgu0jy2r5Zn4TI5haNjlkEgnou5XUL
v4Cpzv7lG0lmX4YYTyRZJ9d4TdReWyMuI6IPsLJMEMlgZWd8NvX7Z0fabl6aF25f
ecbdLZxbFFi/3TSUubyeO95EwJToztmesNpB8eQiZTj9a7N5dbQQx3CWhqUfZyHW
p3D7q7Z/ZM9liER+JK/+KIZ/051/x6shgRsjW7aD3opM15se5GLp64lDTdcSotrm
K7SL6zC6AalyhGNij8lOoeJu/TbQR5MwjKSJbftYKkx0VfnvDMHXpU7VsJbXiQev
3xvf0//6oD/MBDzzKl8GS7QL1DW73EbApHc/wRw/yH3LVl02GU3CEG+o4ZtJ41y6
R7d+TeIiUtuG08kV5UxEGxVtzIaf1WhO7nvi/v7/8O+TflGTU/5oaqFIFUvscHoo
uCVXcY6LDNeyL/TrulGfMyuWDUsyk7b3QhpfRBfKBt9nAOvGxjvMOI0auSBeyTLg
H9MRBkq2LNFZdnkYaEljqsFmG0KyamnJ0oluj1f6uNB0edcTrc70fuoeswySVJwB
iVG9N+cbzLCOP530UWVZ0pKTVRaAHcPPdPI0udzFdAEG0zVjmEM1eRthpP4uNehd
eZ90vzgO6/vF7gGb8+8XfVNmxIRvpqkf/9Po496l/Et7i9s8kuHZzezZW0ldzGtP
CbOC6BgYvftltBBbS/JaAQwkJxloXdEIQpBvJM248vt8szvcbzcu7V2eAprBIzKa
MSaBStA3PgyLQd20mxVNtIvFCuAmhvJdmj3JlUeHzo31VpSyNlaF36C4OhkxtYyp
0VmF1HU1ECzQfSXoskNyEoWfh8DMruOVm5FEahDfGbRD+6eIgWaL1U/7TCwkRF88
V/XQJFLVjbALW7VWpfhgj5s3G/Mmcjkkhm5zlksJyP/LF9+zcXt5riOvwO3kAhMf
myIdSLDrgrlUd0r70i6ulu8NMzdwcZ9o+YdmUU58+gs+VHSdbb3x+lfGpuWltJxy
xD52UCeFBZSfvxtZm8W1r1EbcRRX5Rrew/LI0W5C9I1gJRZBopYvCQVIlOz2F/XR
T1GGiwgUFn6gQq6/PkyGliiI1NyqfDY4fjR15rDHlQJ1Wg47XcIqeEpkMMIIRS30
kJguzllYr0FM9vlqRrHbEW+r1DdtNNYk1X2+BxO4tItXvqfKrGZwq49t38UOJiBp
WbwmlRptiC1FWHUs2veeKX+HP44t+K1SNWfw0CO0W7ANKQ27IZ0ZEZfL9bhLV1rj
6pqokyBT/+Np9swTqvhc8gXPGCKacV7xozMQ3QUTXjDuqCBzo27XPsq6fl/uQFZE
FP+FhianV7E80VWaHWHSKZAoPrvYvkI37QL7jAESf9Jj43r205X/lzjFE+uy62lc
fDOebqDBEjKpD6DFm9vPUJjLMtJ0wHLF8tV5Lt6gKCE+ldlKGl8XffObV+EDR1gi
8yjnmfzEOYAC0VV7ISZ14EeK4ptfA6q7i9zp3ZgLYaNiFlRLhCHjW7kbiZ3pBIqV
G7R402DWWYGFVvjDfwglTzKnpVrVoSh+94yIfq/P9kBA8DXLizwrpdk25Au7LdMw
Ulpsd2bY4HhXi0vfyJq24c3Cz6mh1Wc7ujP+V1G/YREqtXTsxpRbxczKqsy1VaSw
U9SzG29kAOMYzh4TtKt5uZbSMPKAwhF3bvxQaMyIrzTKFpWXBQ55+a2p1Y2HJiYw
WiPLHLY3M4vFayggkXlvI8w5PZHpQVW4S4Nfe1bO001DalEb4bJF83uF4uL1+a9Z
h1EYDsL9NachWFk28o3wmcbHLl4e/AG6bkd3Idhe/gL+8IAK+vw8hIhuIe0NqpLz
BprjDAQdgH1y7Pr1ER6SAOpf6MJvGtfJK6x+uEVqAZL/6Rub/Wytdhr7ETL2ZL9J
cQRoZJLCh3MVl5gnWtAchJuFRBC5sXcqHG81p1DlgIKmBvuRaIzJF/6VNSaopnPh
BguE4sMlPUXkwOA4FoI/KohsxJ3oRee4PlmSYDTOOghrAUOgipshJXF+60twEwCF
V1LePAVvqnrsx7SZua31ZC2sfW0cX4L29rY6tDv4hqgjzL6sMHHznVHhKLZyTcYw
sQdqZNVNFR3lTqThizRSq1MJqMfEndp59YdE3h81P9nNpVh6yCsUAIhDi/tFRZXC
O4Zrsh58S6u+6dqiEa5NWgBUYNwnNgzGR8P3fOGAqLopftKkrGuwET08wiLv5Pe5
3mvN6ceQY8RhURtweTb1sNAWythfnOXkwFW9uoEnu4vxBlGkr198+VAO5mx3tx0M
okpW0OgSEMr27gi/YvZHnRgIc4lSfj4MMIMmlj0sMO4nHs/Geyttqo9Yv58VabRO
wpF/XT6SC+o4qQx6N+vrP3cdEUQ7hp19kxDePWa8zLa4LQHvmHe2J/VFOZ86cn4L
9/nyNZouo+jvLHvxw5x+kkVQQuVOvrREly4k6xs2dC2fGtqbxEuJCACRrlWsGNZ4
jkjX2rPBIVpPyNSrAJEw8SbFAIPsZh8Y+4ntwNt4zyF1fCOV8PF7R9VyRzsnZJiM
HvopdoWypESkZu4fKENEyn2SLYDCESWxdX6wR5LAJfNdhGviPLRo6tJEa6vFqSns
AjPuLU3gWwj9CX3lqLnrzAnv5IYQtnsfpS4Jdno19nmB9NgchdC95FxddE0W+/x8
gNJ2mHAtKwto1W4sk8P1rTCYdVNFVsPzZkPc/8yyJHAFTIURFAdirXdXS0X6wXg6
VsZwWdKS5u0zhCQmYNH4ZvlNS51oZt+0+FpKHpIIpTsjtlNkOSWHptZjfsqWLPuD
snxnw4cJHwSAp5LdG7CMNS/wePH0zcScvETDTHVGDJ5yXAGys70i2JORgYuVVnsA
fj4yLfzKBr+juisnsIc+QlCSYfrvyaKRenj/Qsq5QGd4Th98JN/uYVWpTfzmLbfh
xLvHK9JkeOdKZU6A42G1L/RcUeAK04QuazLCuYlwqG/4QrVl4OH+2bFuWo4Hg6TG
R9MlCT5EEupHPX4jHNiEmcAtK0sFXebTVG5de9BfpP0udI6bQwnM8GsLxDocBvjd
OJOM+/K99VsMTuhB263Xp7Lve7gLFaWdSZdFG/qTAykElnDfDms/5xwgb97Irek8
murkeW90HSithppc5Su2jHnBm5bF/zTGjhfRjK33WuBPv1DAO/CwBnscFT0kG6eL
0E1mXGWgax6ebfDQQwNO6xc5tD7EQ60lOMo7V//kNBi25xrlnFsy/QDbm3TawyZj
8hopQ9UUsvHP37/JwQMCcBlFpUFBBWfb8ay9d04ObOrGE0DdM4limpvnkvryPtug
ml2ztAxUq2z7PNIcEo4OWlvI/sczwp22BBkV3rFXY7HXhnxHCAJcSZ/RlA31MkIO
R5/sp2+g6j7L+5uowNrPkc/zeSDAAvQzTFrHBQQR5d9BcrfTPJG3YN0Nk8QdmQ5r
46PzM79z+X/rq/uH3Z+Js8T1yyn/Zjo4aF3GIeNT95jrlgX6jRB/uX975JEy2Oh+
YLTgMaHUHxXbaxwoG1sx/hmhnp2+XAitZBfhIBoR2F2ccr6ALs2+mH/llaurcdWn
2sWzwI4wiOYtS5DmKjnSnBCVHmCcjn5Iwv1dGFftpkrsRfqlWmIoySxWSvK3hbx9
IgYqf+IOJt6ogfvVUUsewyF2b0OEpLXzzmqGgLVl1Brfe8qV5sNZvipHR/r9oFi0
jbH1+GMzAZe8mxy/N9ndOo4SoZreYXzhiASw2ue0vfVtwZstijHzX8NzX9jxFpb6
zjdpSzUhDGtRorlHjEBys0VIYtgqTbUl9YUAEGSkFj7DQkk5nN5IuOan2nAIlj2e
soE4In2mu3axEfKOO+4a/Ur7qawm8PxADxpRX/H6+BTui4qbdcZh25lnTUcXUfs0
mxOPBxiXToAmh9DvWdL7yDuOY8YlZAuFddOB7siDxr7H5KjT9G3KXlWgTkge1Y1P
3pLsdJUmAXoiFkxVPr2fkwIWibPhmF7pJDLsIJbfbUAlxc7JCemRzOeeKBteE/cp
H74BKi0akMswOWuyj9jZLNgQGzEU+1HcU1ryK2rFophQERS9EiiWem+DHuh7M3uV
33KDu5vvnyP3vgSl8fbllWwb1Yx5pY8U6T+3TKVu96w9eDJMzio+6OAG2qa+5bDP
fVKDf5jseYUzbIgzRWK/fQY0spfqI6jjdGr3Qm2yA1k36chag8N1xNkmPOa1Mc1x
yGW1OLY/GozHU0/S2HZDQYcQWc3bIuH5Q7d9a7vYB8uQ5lUrVvmgKqk3/Pm1uybZ
9+p9a0MazRK47BEMGKw7kMVPIj3A64tDceTOYlFdl5SE5K+C5PSJTkisu0ItCGWo
3j4H+PAry50pFenuUV6SAuOGF/ZxSqLOAPyryhSUZ94xmUIVMXt1WBo5B+633YUV
Z0yRiPFV+8G7Z0S+BpGHqv9k4SSiC0bBFzdfviOVTm3MqE77O5MMoqxdtU7Mbfi9
AQdQU+WQNlFErgPtU4tUD0EJ1lPulN7fZ8w2G0J5sfyfW5lwd38ZY1is8+ew1i2q
68W4F42n0Bc/IxjdysRo693r6Uhx05e/osdqtxk1pRgtpZ52gIQwTlSXNUKScBSN
ajQLEkyTlqx6Ckoyha6E2effTr5EVYeUKxMT0oY7hCIU/xr+wCKXSe4Jx1jWmXYm
7mjO1RAs+HYGkRYfGesTBxgSHEIyuC16LlXxTad4O8bwWq+Ik3ObXYK8vtD+2nzL
mW6bEWLp5g2qxN5DwltpiRYUO61lVubw+QXQvzIAZQ7rSvVhnRPW6AScelyC7sae
RBeBhhFQElZiluuWb5+8VggJH2/ey2IWom1H4adB/OYkIOXFo186DbwdIuOG+7Ol
kUZQ3NM5YBuOpmGg4SnRQ1h4WSksMApxiek0WCqTmGoA4nbkP7y9uS3bSe49/o0L
/fhm8l+bUkT0hv5e+gMfR0OhSAv9VxvGwAfut51Sc3Ry9tWFSV4tfhg1QNG45g49
2eKA85j3Y0VZu2TSjcLI99kC+2H5e4Xxy/9H0SXecnmhFabuaAsEiyxUFzEvFuf8
45jEOlTo7NUfcpXIVGIKoEGvn0kMfgi5Y77HnoLYSTckuZDGGAOqscfLtprapIKe
klsa7unLDIat1QLQv8OFzN+WMfMtSKS/bOe+ivJzFQlzhZWUPDd2Xi7X5vR7dEMj
/ZwkYJfC8+ap6C1tpl96pFaj5BxbQ+Ok8CSBFi+lsfKmCktD3g7r5OjDhzCyNYTA
TQuPJ3zbHhZpYhfPfsyfYImvkIxUsLizgX2N6jC2X9yeUSEVMUlAmaYL/dpOypFH
PxtPR3/JXit4BJNLawkQb7eNklYoI4MywQ9nqk2ETYRCG1vCaIhV9iaTmNJdFnek
bqrXvOHdNJKmi6ng5g5T+/b0KAYlhtKWuqVyz/G7ySeMFZkPbAbKTCo6pmt5mHm/
eCQS6zB7sFjocdKTlxvpkrvFyEb6OlWDo6kpfCdK0Rk=
--pragma protect end_data_block
--pragma protect digest_block
NseU1EWFkaSVjdKiAJ/EbTTEQAg=
--pragma protect end_digest_block
--pragma protect end_protected
