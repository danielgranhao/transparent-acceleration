-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
MesWv6hdP1yza39VVppsM+hZi16oyW0+gz21ersGDjqvgFZrJj+wQfPIVOFzsf2Z
VwJT2BP+0lbsbBC6y6yMkldA1igsZEiTp08qt6fUSSJPqugkKQ61xE4SmbdEXgRh
ewlsnmuGauEL+mptXkpiQTyjBqKv5JEIvW7kledl8e0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7232)
`protect data_block
ZOWSeG1DPmoKUkGM9obAaG8dtXoxtRSxvcISAfY7tSCz6Z94wnnO3bO8fgCxG26s
b0Eevj77AUzjOA5TH6Pa0k7VRL5EnqNNRcc+9VV7TyDInMGTokZL8pPysAjc2iTx
tcLXPIXLwc5e7m1NYE9f7F4moOWOJdgvn9tjmZKm0R9La7x+tfdByO0UOV9zHoXY
Kz0QCk773/yegvLf2y3WigbBOpzuSbtoZ1FaeRJXm2Wx0jqpi7l1fkBRfmABtD3m
jxiHLh0bTF9kzJ2tJE8ufR1RoUukP8+o3pyaZw1UtMAHHWfQVTtrgEI2kok7MDvl
5KGNfLqkzQbm78/OMBLAozw3aJYg60V+8njGP8gUVSlXbfxYp+ESEk7Gjd5Z73o+
K8At9YLnjes3w2aNJdnFmCeLLVZW6AJzAc4MCgdv3FdpeSGzze99YkI2vJmkaWCE
mURA01+NJDEQJJrWlyBprZWMw5zdCcDBKU5J285NXQJkO5IMzDaWNhv9duXtHH0y
tkwOTJGZLyDhiisKIfftM/js2GNuS3aBJwmOMUYeupqedTJjtWsmVqZPC+2rdlR4
UwPQSSBT+rj1R6e7dyVvjEXZHr5aJ9e/TiYNQTBoqO6kBPvszL8BRkD1ErYkN5Ef
H8L0bW69Kzksx/Gi/W6SPaIqQyhWXKFJJocPiXjyy73h2EnEg0X3Yhk1OGfyUJbu
lVFlzgbWLwfbNoI13tExOYHOnO4qsqKVE3KTUG94L0G8txSogrilab91ORBjgItd
7i/LsqpuvfswH58JIe5HD8MjZKLV3NsiI96pEntcEUwGagYH1iQaHMsl2v9h7R+/
G3hH+sBqry0hsvx7Lynj3tsPI1n2iGiyrD4+rdkq7i6cfvl41MRpotWQcmuONbtA
zLdJqUnYV+WzM84+xkfu+BsIFMmDonZxsC5THLE2B8GO384tHkplfkQ7fIWKdm4o
ZY/l85+OowdYwRM33DdL1r0DjitxAkIvi/9cPbSUVqv9GXBX2TojF38vmnYUe3iH
xoQ2/+yxioZFvlkw7y3Lu4TvA9SZ9CJ0v/0fr41i3qdsIdMEOLXKMXREwvi9NQys
StJpPhUrZm7cgNzF8s9RtYlxHK82xFk8o5NyFbh3NAtyamzgZxvsZOS8AerGvm67
570gTQmENizholQ5w2ERF9VgtYTSsCm+HoByo0cLSLWzFqfQaSWTKxv4QM71rkIN
/z2XFvw6zc0yr2gE9XYChn8rQad1KfzwHcHe6A6+0CwPgZjBVbHYzbZi7Kt5u0Ci
yoFJf6LugMrajfJEHMv+CnaFQYWPJdylScJgXHkzsUHAoqEMZyTs7qGlAmTPHOnY
GUZedtFctSEWxZrOX5vj+LtZZYIi3ZLPJWY1FCsmflR3ffPExZMocga+NzIYQsTs
P26V60zLXC7MSbzJ7Z2J7LJRXQE650gP6BIeCNFhDENaQpgpwmD57YpIl6HFYzOH
XizxkJ4+c1iAWOXbYSutF1TsJtcyN9jMsjpjm9JPkZFh4RiN4bC1rVjoh9A04scf
j1WyhxH2R9eGVlJHYmINe4yqE7q8ghs34UMa1oW80r/0Ru+uAV6MEqhZtFopGs7W
AteBHi4ggFGO9P0YXVxrmPeZKq5M/cM8lCZxDiFJlE8zw7MyGAJn5++54oo0aJaY
z8CbSUYv5UUlm5RBUlTnNUjscJjK08tZVKpzLM3d8GPIP0kt7b5x25flOFgV+1sE
uH5l2fUkKA8yd/98bfWnp1pdtTC1K9VmmnjZzosBbKQzkrsnx3OOc+TkYjORaz2/
b6p9Kqb0bPyd7ND4iIyDzFkpb34PbMqPMmC+eZ9qIp95TR5xGipXFzS290Zb2qmi
g+Dk1eWBLDf/vmMLOPct/aJkm5r+nmlWwlls6gMYsXpFbY5ExM42g1hGk8J4i7r3
GtTEOi0KU8u58qJ6YEW9xyL6wAZIbzpj5mjWGeQ3MAQLCFWWBlUipCjCaRihle9y
12hXXeMUeHh3MtBdjbe3wyr6uBLPkA79EKjnAZCVcjtyXbXLudRfbbQVoBVGBs1g
qqtjBZ8nYwnOVE+/0Zwt8MrNw0UhdGy24e4g0N8PQ4lv5iJ05Isw+iLM/sXBmTR8
GVhanatEeMTFKj0Gq147hwOWnvy/F5HcaLvf/0XZXtUwXcIjHl4fIW353Ow7D+V5
XRkQdV/ijriiFka5fSktkJNu+GSWZMUn6DvqGJ99/Ta8lFstic3HcDihyyKTdEUz
aH6P7k5j09DqioC5CrZXYopFJvOMsAMHZxvceq+MYSsdBDCGXBGapLpREtBr6N2y
TTHoDMBXvjU3K6B6dmyTuNgMgMc25/DphdX5/BNTM5n45OmxtDpCfRsxE/hbbmWN
PfIypr336KzCTOmxFutiVBofsMsG3IHUsWiGH0wWNdV+f/Uc2AnqcEutxePheySZ
jZN9OTCLbUPFj56oQ7xC/ZDeaFXu35bB3XR7CAddAFcuoEqUXRaqTNIga7lkKjgy
29iInaTWIu15cxjC5kJTS9qDVNqDk38n0dkjuhGbJ7+MAz4c/DV16FF/ADlpmMKI
A68p5fYVQxPGu1umIaXBewyrcsBn1n+O4Xmy9dLL+YGE8VMDb34ujKEPQDd5FC9z
+veaLLWfhWrdmy73OhyxEUX53blwaUycpsoFYY1XngQxj1Ci76o2S5zdcDke2VVt
Tsl0DfjZUTRawOVOOGRgOPq2OKp5v+yVpSgBrUXlMMRUzWQuV2wNNVVD58aa5zLx
8rZYoX26qMJJR6GxSrwYUrV71HIajm9Dk1e0wvt9H/Mn08uorHRHmKDNY8fe8CP9
qRTgR2ofy4xHnQOb8y7ATxwfcp1gL+Z8xuWo7CyqHpXZYkEMJOFeY/87z6NwK/Cd
PNe9dFroVEMQu9bT4XhVQ5PGYCeUHAAeniOvs6IAsG8wVLFBnZkG5q7/q+Zi75oh
lJ2s2/303BNkYEBaLejBQk5Gy4llt3ZF8RXEhEAC7Vx6/mAb/MsmMoOpuhcTrS/j
y4Z+3FzDwdB6OmMbx33rL6AOvjO8GMejZZTDbzUKjzZKaEog7mg24neHYLYIU3kj
/8Xh0gGZcvxACXkAGG4xsDwJwLqizkxg9kYL7QpTu3m3aVg3HYefXzNd0wIJQBGI
M/Wl0nMdr6J1L4ZiDcQkH87RVxVYfrYIomhftOdZIhy5uv3cXBOOSkzLEBJiUFmM
G+Mq31hHdvQrnzIpdtk4ljBNaRSYEH14JexGYdraNM728IVObjcgUFxP3mxNTBSk
5OIjVTJH2+5eUoYXDe/XryKdtNE+f5nyRoOfXX92aQfUcAKBTbk/iGK4HKTtd/q7
25sqcu3rTzixvE24JLUxZpbAQC9XgvqhH4To2CcWaWa7yWCOa+Ikx/0BzhUYYgNN
gRS93h6rTGNb3e+ngpe4xOFRLBnf3BJZ1GMTfGyASgilN5qCHbPaCf8D58PaLnWg
lm9duNepm87zCG3lI35nIm4aeBDu5t2s7iFl2Y8etvS0M21Y56irF6jThg6RjevV
mdVCXX9GWV96vmuWQFKay3/i1LUwEFSyet1LuVuRnvZd01Hsa8+C5/LexECMpOHr
gnycAdlzuHE4okiyLHlf5McWnQAz8JwxMpCyXGaXy5zg7XgGIydu8BniwEDbm812
eLRt2SAK1M1jFef0vPDQk5t+9inTI9qOMzMkYJoFpM4vFQlVkJFA29tNOGQL2FJg
EIFPfB23SEjsZHdMcbNdIbFNqtK/N95ssvAXmFhiQ57GxlKVoHkTBXCo3gE58lbI
/AohusMySDGJhp/rHMNxIaFReqG2AE1dA7KvhU7R6RNgIZs2souZ3Jv/fMt/oDhx
RfG1ql0XGBlwxHANtBtaDyBMOfhxt/9VLY3f+ZOGf4OLQ/2c7MuawuZpO0/M8jvi
X2ruubaiRYvU9Ol/x41v8Q7x0pLSLTpPU2VySCSNsWx/C8ks5NjSR5lwz/COq7r7
dqWJlOJveYOrnRB5+y8gFmgP+2TalN/3vAvJy2eiKp/DW/rwudx6odXoacqOXNWZ
dP5Lj9rLJ43DqZVAqprfry53u/T8pNNdM8eScjDJD45GAsOf/M4mHjG2/ZK1yo3j
Xve2oje+OOFxoedCWCmjWjY49PYDsrTJNIk/8boR9aYTqiu75MfIhOMasCDYMTvl
9lR4lvpxr6Uv2qctTzccvcDSjSAVRwXU4pg7BXSyeL257xZuWj3GlDcBPyixe98M
NvPEc4L89ZDiTal3hUnxIBn2jRI+29E1orJMnM8l9dDZexokAbe5sTAZhqZ+Z6Pc
ucjHDKtz1f2Or1JPxwlbPJhZu7CsnxdyzwULhXtRuqb1/HPiMYR2PD3hw0bfB6Y6
cci9+ghfis3dA2PyA6DpP8Rui+kCPJNejU63tu+t6kIamC6GfWPHUKAx5uLfeK0G
pTujhwCQGp3jffNby64NM30HuQKOfKUcPPSiqqJbWXsY3GBDx6ebYuwePvdsTx83
ZHzlCWtKW1Ug+URflc+4nlZf6J2jcpW5CgnNDnRp78h/U4Gl5zpJIgs8sFWqajbP
peSb9bEEo5tJ9YvRhMn98lQ1UxbXZ1Y2m8sqpRcsw+lF6HtLrcLk2y4KFKXCIV9P
bGPX6Y0Zlip0Mqy6+uPLsRTz3pPA+ZYihetQVHtPUWJZ6l1Y3v9Mk8oO48PYaCw2
F/dttDusUvmlxUOYWjPlXxM4AehVQK4omybUn35jiakxJRctMDyzrgVun/RFVDzS
fI6url9JSXiqCPsKNXV59Ks57u5m/liWkbe1Vx11ioV3UvdKzcUvgaVtexnZM4TN
XnFkSsaXELSl2CJrwvx7T8CXgQo86CHfP+vO5d5KA/lxpS95iuAgW5HD5N/ZVA7U
iFrW+LGopGfp2b6E+MnNU3XjcWg8BYsoIZLnI/FGxmFP2MpFyPbdEzxj5cBWkNXe
AIbbYjg+ft65fauek/5QodcJls2Jy8GUD3NNhysfR94z2RtZwZJlCfhp0A76U19O
r2xzO/WRnPQFqhJAvBzPUOvPegCXswtSEJCkfATzWe9stgpYJdGz6Rpnm5vFq5bk
PFS1rVkWqDucXPcPGrJggxbDDpas7+EgDkklNm3u2FS5EDtqOtWwjltgo7fm5oFt
78bqOJKMtg82FecoxfynV6+zm+m1f87jVBNMSG2EP40n3noQAziOvmUfhf8xRjzR
oJ3PAvMTuJNIlBpsC2nvyMKBNIyfRtVPiT1HIUPeNrnbmozgVfcm9T9jPxizR+Gq
yl/dJdyXAq18gmkAlFCvaeEX8cwcM5MTZas5RFoPisZRjSDq+Q9F2uliLHvNn3fp
oYjdjO3zLpItjgBWaHf77jRhI8QUyY2+o0hP77IPCfmziuRMPB6Qi27UURtBAjn6
o/sQ0RYM3S0V/MJmjJPYK1uqDS2oNQ8pU3hYRSeS/Euw1BnZ7rKJL8lOzwXhwRHk
BvGGkZHbhW7Ros7vEEsEiWK52Iqiyr8c9dxe/sC983lhUe1hlfX4JhBpyMS8Ou5B
dX/IjVqfDtKMwGgrIH/GNkbQNfoJbwIxoZLQM/vgXojyLMJAvFRbFQgd4/7ro7Xs
3wUhhaHNjflCWeGVwnh0xyo1EHMPKRuYl8GnZNfjBrpWWRPl1r9Wi7w9RwxJahVT
/hNhq5zTIfi6Vom881L0KVUlLn29VcCZmLAd8Ui4/YkB5M6rvW342K3oM9UtvzEV
zNWo3Ic1RmrgPzawc6Lz2oB4MioCEe0POvXpf+0QwntU6tDYkFF6d7I+YBIuWwuT
pphZ1Je5aT1Xe9SzOgAGIuBp4RhmANlRscXpxJK0jCvw+xpbzy101YbN9I7cOtop
zdd4C907s/xj2bX+HytOYRq3CGMoyN5D7k+2+4N4fDIv2v0RnoyqIkfngpAzujaT
weYgY0CYNe0nTpJotkdWzB5sPdFxVgxkscKvayLkWcBCxBqh0+47BKJwD54MMwMf
Xj84Y4tXrvisE7r6fxLD13mQGGpobjsngk19bW32GKkPMsbbB+rBBPosZ8jJA45o
WeI7fxyWYk31ZXi/fe2dVcajA+dKKxl2RolnjSR73zPKMLQJ48bM3MNmoVpx54Rf
Gn5Dqoo0ZSa896f1de+YhiRnxNOaqgGiCsuZNmu1Y85qoueHe2ol42HSTw/sFCMs
kIPIwvsGv3OfRKAEbgicPJCfGIMBm4eGtWjE2m+6i+fKLlfW08VRilEFJG47HPh/
bDiDWXskIGaAvVkwbP4ARllDbQKia0KS2lTYZ0yM+RnSI8CMg0Mv8R9jx1Y7gQJd
jZCPDcEK4JjJ8bNExZIzXjN42khwOFoK3f/s26+2cPze7SC6zjadfBq1V+S60TYz
+nVcG5/+kVGoy0lsZcwQa0XZfLLTa/F8DD4YVuP02WDZKlvTVBn/HwbMUIWLyqyU
hv81ZPWalyUncGzpJ6h320uvTGm7h+j2ntnQnPWmzPoNYlQYEwPXa2ixx47dd0wB
+TFRH+BCUdtQjoavii2/xafT68nCgHYIwBQuVyWslZA4THbjPxXNNjP5XA+Kr/hI
b6eFMwYsTORFFhpfjt3zDnzkr2jCLUeaqlTtvFgyMrG7aQEn5BN4iiuGbgHcUqa4
O4nz2no+RbstkKcAIcKNIGg8Kork+rV2qQX8a0KUPFCZ/DAVF6PM7tljA0RoPEO6
cFbvN7v1VQ4RSC65ElsIbqHj8EoQZNTbLjCgELQyFDAOcGgWbUuUES2/tN/EejkI
dFDG3c/autQClXZpn1KpVi5pYN0b8qIRuqt1nGruV+m3YlkXs8XlqQ2dyP3sCLFr
McCbU2Yyfjn/VnoXwhbSpYiJd+vgespNP5Jz1EicoOWl497vf5tYitJzc53tPpNg
xtHGjlVNq+vOFXiSFb+t3XrsGqLbbQWvquWLdvkscjpx3PpXc/agsW3o8UsrLGkA
R2aeqdmJdUVNaetcdPN3VPuYFV94LTC/dwiak98A4SHOrXdg16LHEGVS+g5nCDFZ
5oTef8RBRcAuFJ8UB5k3dGhqWBwsPO1dI0805h9DcnacsFNwaGt82KCiMpDbqJe5
UJzBqYibu8JB2+cMUF9GMsG9YmGbu7xfT4kpp2uCVbLNRbj9jK3QQuv2Fh+ImFZw
XXoyHG8VY6xxFae4mOKczg44jK0dKRc0qduZYnjpJMRiys9NeVngAqsrGNfX4txl
kx+orkZ9xWaixsG4R5qKWY7YOS4ANHtvc/IbsWJH4S2/4reBlSd45XcRVJyBdcLz
hF1i3MXZgBBRCVWSxLQTucHKicvn7DlKzX+YY61svAIDz9cB3b0DeE/366v1o79t
fSEZY9lQYJC06o1ZmxAe5ij4utY1qryts0QzHpDnVTwYEKux0XSUamrNNMaXZVju
ryAfJK+RawrGvaVJdSpe5s5NtSjBpTD9dyN+oi4RWAUs9siN9JutgB36OScmdW7u
w15T2bg0jMZaeHx/WjlAIMa2tHlZs3IYkGLiA3ZDJMPpzBAs1Pk0yEUANwiaZAAZ
6H8AdxAFRNFKHc9EijZs9b/q+inuU6mcY3ZHWL7uSCNTl+mQk3SGjOSL2R7aTi+t
tfZmzumvN6OTFO4yhGoHR/GNmg1xqs2QmGsM91XJYUUh/oDD37Yq5IGcYu61O6pb
BtAyqhS9MXnAloPMHa90L5+5IirhMBEqKlT+CDkvK8l/BlUL0gPmiSc52R9f740t
xaTeId/0wLscbJcmmp8BtmOlhzSwqXaGZ2dliN2D7U2pwymQ+xV45w0cyZI9YAeZ
207hvMwhFLK8QV9c3rc9LofdJTpyYISdt7vemqhG5KyFO7eh2YIaeCk8PQwUI+5x
+EYxi++5vtCKt3RqwZt7KPMEx+4Syi9nyiQ3oAPCHMIfFz1dqjF6JyS84FwoebcS
/UGGzHzwfgnVAFdKQWOVll9IZHCaIjrhS9dWOF2PV+EHi1s0lWRW39HZaUPFbOEL
mBJmVSVLw+0/f/Q/DVy+awzPa5KK+aSbfM7xZxQJ7HmsDNnjPe+iuF4xUpDbxKBo
nSezMOdeH+FJYZDojYt9mOy8X6G8kIBnGzWCqJ1T+S2Jer8/RbPliOTdpzX+GA+E
X9NMZ9xTDPz1uYkLDEatkTLHTQc1f5nOIQqFvgBX9wposp5a25tg1mMZEaeEiz3y
ehS98cUfsdf5yhPCUPSGqqdw0KU5przWqgLZ34rIrfvbl8NP+SNZ1N1GxKKkjF9F
2mYXcmBmIF3HQf/yRkrTqNksovQFwwdPiLu6S5ehHbaiSuatyVj0NwzsvIg5EJQK
WmmoA3icXFEkncxni4APLfq0VWXIjMbwstmD/+uD6igggrSb7fWLraZi4HcTDOeO
PhxjBsUeCpCxO5NQUt0v9g3mZzUCS8zllfCvkgWJBUeEMAVcipmDDoqxNfAfo7Ja
CFodjo78cpBSNVV9iQDqjT6u3d+Qpwdx9g/2rqSexvS/cqq0dgiSsNMf3EaKTjxE
7j2MqeQBMX97PqbM8JoVhRs45HYFC4TY1vhHXKq0KTedGgiYa41cjmQDc6NqM6vh
dZNDtuB1kQIziVT9uT+OE87ghA2BCBGSal/YsAKsRa2xOMrhiTXBhVxm6B8OdwAz
ewcuJ4504EdUFY7I8ikc6d8KIPhyj/y+2Q79s2n6H82lEXQq24cqC2sYUQcxyFlK
mBzGJHr+UtMzoweVxOP0MVL7gKnDzc3VDZQfePROvvPQ/RBzXIx1cmduSovKBvxq
IiIYF6YvThyNhmadQcVY9AuhC4Bkw7CN9IZ5CCZyfWA9viuAcyXnQG13nBwTKTTV
WXOev79wGFarVXl/Gql6hb4UpfMahT5HvBtWR7NxSFbavR6cymlamjJMdWDmI0PG
qwj+88/ebNYPOJdecdTcFJ8Hso/m763B3Xl/CfYV953xn4HlgsvYbMzYqkPRNFTn
6Zj28FuqQ/YGLQiRAkt82HarsP8Jpz5P6p75i/vZrcxkdkyzx+DArb5g5pNkNAEU
vQ+eCSnIVhz9Xsj9VGLexmv4wme5llP5HhSGBgVgPoKW9RGWQxJl5Y7mqHmjOilG
AhevwWUMBdkiHPd7wJ9eKrolLvQ86KVsw9Y9IHM5HgoF1SYx/CDSNhNzvBoXzu0j
iHR/4Bmpem7sdutIAOrtrWom/w/Thi8l8QVXfavLqURobqlzhVVnaFx0EvAttD8M
G7mGL/6ACGoUWMxvATBMZdzOho4M2KQau04Hqyx2iBBO6VltM/CARijHIqDeloI4
qhT7tNPRO0ahHwqdB9sRzzj9Ul1QENyI+5PKTUnDPeCenQLylyJqNV02U+KTlY6x
YbSG0u6Mw9Jglf1LM+q+Jodjd5KLztaG7oSqxVWbW5FH/qL+j1xr+qMWoPqeqoqp
JrPW9ja9HlJ3p8gpbThctPcoa+1xldvuQw2Lh7kjoYONejdzq0absKLBDCb9uKjT
ivMsK42l8qoG8Wg0WzceJOI7/AQFb4nIXk49dFwl4RPI+3sdi6bjh1FuBOk7IqQO
7PjEJNuBfmejKFwv90k4k8+2JxHHjOk/FyEPVbXGnzQJM7JFeemt40Av9UwEpaxH
y2mcMpwBO5tjLP+BKm+Rdv8RuFlDYeOIKPmtgmQ8vTdC59BKCWhJXwLusNHNOJ+2
1Jyy2+NRAr+xDy7zUPRald/4ui5T+P1IQzPcAPMYlvU=
`protect end_protected
