-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iG5GkLkcmOY9rXeNyu7c7aj/NzXTYr8gbxCQ+6K+MxOWqS09mB0DlhrK7mQEO+b5Ajn/oH2TfDUo
4lQVE4PCeyDZySoaYHwM9NzfCyjjuo53e5DGnTawZiUIxoFM/2vAMsbCSSzIVbfMcNWNUGlBvspE
5ufCfPuh135BkS+64OMpENRX2tKix4kEtcNQXMYS22Pc9BxAu/MHgodS0u20yjHbflwMrafpRbka
9jTCvTNWM4wSGy8CZLoUeg3ieapG1ZojDR2CT+WE2szSxI61O3J2nhVRaPdu8vDfXVEYFfZ+q+1X
K5fSElGtO+AgrOY0W+Yv+pDzms7bfUsKKZ3jKg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6848)
`protect data_block
aJ7ngNhejEVRzWiVONouYmxWeJtUCoCFwzO4k+nTrDkUC3LrGjoUmj/nzVf84Xv9BAMJDc2m1x92
jx2o488L3xu7Oce/P5V7Ua2miYHHhEQip2PorGb+So2j2MPt6XJB4zINfO+KQ58Amhb2VMApoTkS
RRx4qszgzJkA8vGChGS1o6+F3apmwrzUyYeUnlfxxZAZDdDJn9utzgT9fW7N/H9FOaM0JCJM6Q77
VAgFvBXWzKs1p/7a5KmHkSSXdzEJ8Y5PLkkAlbVkjbHWkAzBaaPeR/o5su1qmdf5QDj2bLtQWRP4
T952V+gORZe7j35XEoIdB3rZc1qGGe9CIRrWF6OQh6TQRmRc+hzNp5EQ7LbpAsQNfYwsgRh+7gKs
fYMcNlyxg9F9rDdaUI/G02Qk14puxyZiuge7YpuX0Iy+8Zh9FVOdmGGz4U+FzoWnfLk9elXd5lFh
Qs461IUeuHaVg4QdqCK6t4POvgaxMHBQgpLwLwNFZXe7wLetnesGC96ODgOJBJrYY1zaaotulNzV
NxSy0eVYKwyilHxZ5yd67ejr6U1DfL7HDgfdV8QmFcUrc0WpVrNyiqVSkmGKCjqRe8RVkljE+lzg
182//SzOl2q6NAXTJiWbuIsHIxKwouxQwGjGbI8Gvl4b5DI2sDQ72ZrmMSb0KHWlep9EAMI4Lobf
A5q6TtQKEbs8ygLRDt5g5g6QaFMy/M+KDWjKw9qG2jT6AyBg9mDE6R202RxURiSrHvB5LmrWqKde
yU5orVI5xrINt8b6CQjmYyqa/p8GWv0opvJm0ZuCSOFNATP9XxfOwXhMo6b4/wppnPEuYmUWWo1A
dqK+eIhZoufRBbnAcIYusMNOlva/QZvFY3oWUy8igMOQEhVy53TjGCL3pV3E9nORQnFfvhOEOIrd
y8x9Bk+Ek5fip++lKNwtMp6WiYGebOKvIqAURKyCEi2LDU74LCwuUA5ldF+BPKcnYUyu1lcrXcmJ
mrBcaiJEAm41lHzSgUq9dvPDwvz+ZpJo+eMScvM9A6c2JT6OJWEZeCSKpjb34Rb976nlK55oD2Jq
9iE/zJu47cf1TEBOQ7Sm3GKkEhaL7Z+iBv0qdTrFAKUj3cRIQ+Xf1BhmDAkbrYfo+jIs17YxR6wh
truAl8709fsmz4Joz5QHKYYOvqAV6ZM4tgQXT7pfjmWjtKBXHC6Tre9zS+4KQmyjN/AmQ8s7/PIF
9jXNlk8ufJaIkDNafqYpuML87EM4GRVyx7pFq/ffTR+nhh/h7VndLF3rfpr6qHpByO8CqG4t8iTg
bX612DiQP3w3kbwTMvd/KcKsQM2DoSuwr2gkTraLW6H+YgAeFDPi/W/yuRBddMHXhXLrAfJZgJG/
Dsj8t1S4uv+Myri4UXMbdASfFLmGfH6z5fR8R4vVDHD5Aowo0W1Xr3cEsvii1TJ1Zbp6Orp8ivYr
fsS+5gRpkmFEg5tEdDoL6/vs8LVoK43OFHBRw86U5cOS9iHKgrm6dz8drSNg3095uXfmRfQMKyzT
1tQAMB+88X/XXJ3evWwVVG5Uokew13q5JmyjM0/8xhfBS8ExrnMwiPFmmefyeYtb73b77t7ll2fu
GIjTZtN9pvMViI6xejG104pA1nhiFjvKX2DmQRcMtVS4iYU5oXz7iBO2ZB7rD9bNRR1amPyRvPxB
M2FPcOh2mnMk4ncDqkuao18+AsdK6yps82iS6Xpn1ZdrAusgWrZoHejTiLyVQL0uRTsQqRtOwPj5
EOS2fIhZfNHPAbAQH+jd1a3rlwFVqWJbylZWlprvGDdVEuLUEMtbhV6OPq/NvOnmH0ohqmFWFRz7
dOnFHkBShI4gVjft+rFmyItFd3gYYimtr7pMHyQL1NYdI4F84JyznZ8hugGyKKEMyfho2TTqMIEt
15HQDmnvcGr8CtTimk2gQ1y+URFQ0gPzEYIG1zUPhgkvebDjoIwsbYP3fCTPwnxrPSXgVNwODrio
i3+gMAx2gVCv0+u+DbiYFfzRpXDsMvgXqqecjEy1oodfFv+PhUbe21E4siqR3pvzIqDq3+aJ2Vtd
pLmeJS15LBUviKxNHEtDmymqOjojdZg2QNWwoCaOmk/DxLekr9mMeaJ2eEA2eINQK3l3dIplip7c
ZleRkBoxVLe2Z213pHEnZ7lFFA56yooW/TZyqpXwy0DCrx5p/2Pw7sVvaQ5IeYzY5kparGuBm72K
utAShklkkCvwtwfQJSQrdiQ9Kmn0D4WZqfkfxAH4zfZ2MzboxVzvxrDEaZ5ZzwMLxID+m9rG61yn
Y7TIoeXjD35fub69weJGGHbjIXIVkgA8ygk/k6OC/g/dPuHluTP8dq9Itwrq97A0/y33iQVZkoUh
FR1p3ajgj9FcMCN8oG9Zwlzhe2AiyZ7YxxrD2PRkpu8iA7CYzFK0iBqODI6PR9r6v6xdIRBnjajL
UgbEXfFNnrhwKiZQU08KwWwSWZQ8zUfr+UvJLKvvXR/ga8W+jH6GuJ2nqXcgehWnj7i0So2oizh1
65acPfU7+bhLANkPFl6yk+bkPK2WQLjv5zUUgbBR1il5wgG3akrQQa8tQeRQrQkxCvKCOebAbYT+
mwGeUVN6rmWAuMSyWE2ub1mvdLDrrZTxJtjCc0aAK3kUCVOp8Cx5sGdsTjK4oMqGWPBz46xU7uPU
pCyT4LKFRoHl+47v66UiGfnth8lelX6T933wTDkHFFPhJdFZVy7pL3ChTW6Lpj1od/LtjEE6jJ2/
h+WRxMaicSLRuWDZD1+/0XvtpsCPViRKmzJBtOwaZl1Ds1AtACILhxTdMaGK9Giz9mBJ4V9N29gx
f8JWLRs62UogU/NgBpnyDosE7JMgpqyDdaclftEYgdVZ/jDm86VRq8ixLP0kwJs0CckrsQHA8COA
sndD3PqyfMh9lGYuf4TykvjEmyJmncwG+u+FcX/paLx29MVp/+1Wttw4Q4onLOJoaLiBSYp82rCz
b0yNslBDcVpT3Hx/eKadpP5ACxuRub8k93YrhkwRSMpWUJR9Vyfh+IorS2Jw9uCAwynNDzAOSiR7
O/LOughqQS0xkYkvAyK73/94yn3hCB81K0pgcE65KlMvCFVD5hgJ1kfRygXc20yHizYnIwrSAvoU
57tA7xhna0MFleKmsnFGmPKtgiZiOTKSbywMoQvUSRrh753OENjF/oBF0QEkZB8qp01dRDNV9L9X
usvbMPXfTcei7V48cDEF7WSZZUc0tq2fivZeNQX5QHyOaguh5jZyc4MJcHVUtjNfGG6W8ih2Q3/H
eXQ2DaYXUwVEPr9cD+vBi7jnHzxoC0TT/YNRrIPXCs8YqfwJ3f56dWld8Ei/+DBCEzEld2lnoEYB
4sUSrRInXym61Kcn7ucNGaa2EfxAo1FohDxNzYeEpdUEnG5ERo9QP8jRisT5/lJs+Y05poFCNUST
XqugqdCNpn3aBdhp38GMDEC40eEwvwTFlSAjGQzxt8uMGeaen3ZkruKWRg/FQudPGzu35MKjOsrq
J2iCuq8riX4vT2QykTUkSzSiB6B/9L7zu0FJxbOW/Uxbr7rtcEbJj1sYfEYnR0z4R7BZM7O10w5w
hrlJf1tOHOBI89o//1tUXzyQzSl/QymnbjuVmrNOIvp2StyQaOTNL2EwhXVnc8ErrhojcAZicOna
2nzfxxwF9nWUypWiQdJi4/Yok4WoWT65oYidXp7CBqG79jojcapLSACwTKmXoGlnvWe9PZDJYzgl
oSENDRokN5vppT74K/erELz3NbjoYzmMpksHKqkMUFIJuyQYPaJ6pDu+jX75JpfjyAyfoITJfMwm
B5B9Iw5kiNR4zoxV11uiXAVK79eAJSa20VGz83TVr3wWFM2/KxFC4X7RvJ0yks1tdyxtNP6Tphsg
mWSOEFm7iMjD/14v5yKOmcqd7kAZzB/iURg7onyfOmCgUGTe9ngM/AA3gbarPObxQ2F8/PA0Li7A
UOt6jnrZNGHr+qskyuGkGKqdBG8MIAFncQKcBHoCNwUqQx8CqPr4bU40KZVjqQaPvLOCV6TS6eOY
/ggBoC+lmUsOlR9dDGVFiN+fPeHPArzRt64L9C5MAjBbvcnytnRTWGxYdzTUTZc95JFaXoeVQTn3
UlBFpNeVt0wMTIQqk3+5D3WOzhRWDc3GWH6WSvltUinsvnA7Qg6wTQEu2TP9H2q9Un2O84XNZPhq
Xr2FwR0yRTe3FdmotFaEAFa/OPJLTMalFPES9p1EdJ0I6B94rCZN3yWAW5r9cyWCdwao7nqSXfko
u8OLecR7UbMAbid9+BKnHpqy6cPXm9szcgtWRztLUs7r2xTYrE3dnEDdOAkqYK88b6aGZw+JB/ee
ab0LTEvK9YfRXZ2qeHAZJiTjKOyInrXeuK41cI9NnlKMERPlx0ugoUIViZPFh5PU9FRoBgvVJ3zZ
QhaR8o8N8v/W6pvE/6Ac3nVtl0ogsaQk2JLzc6+SG13YT61NjR0mQCyM21MHHx8ktKCiIvLpTTlX
jxV+2gfmkS6x67uV4JTYjE6KH+Qfo+Vb+xMg581DEW2PXF0yG5XBJUzU8ZKr2T55J2AU/61CmOCg
mOJzvE637wbXOZyEZ6u3vsLiosnLowqAOrr6pCsFjzC4Fp9+9OWiSNaeSuQ3QQB+s+JsVAvvwJXi
5WKkId9Wp6f2uzKpwmGGlhLfgexZyqrAv30+UH1oQ5wEZL58v/n7FF8fVOnK/wQJJLTldVmGFJ7t
sm5pZRiHglAM4G5onsKzApNVoXYkRk70GRdz7XTubtnxhdnh3NEYP2iEpUagEAcSKIrqyF5BopbG
Svqz/s0VkoSZZVwObIKp1anho5OLBF44ccitBoHSvUv2V4E5IynF3hK+Uqthfi6QW+/EIUFTwi14
/Q7i8KFnw9kGPudRV/SMnMv0kgg5DxI68CUsZqxnM4goe8+Ci77tKlM2M5ZOb0mKO4hWG8yOLC8g
E//O9fBHKwBMpgIgoLQ6AWkNO2oDwqjR0EKEbNuYF4EFzNH5vEYcKhmQ9cGhpp0ussoMUFi8UgLM
WotpKKRzikl3kVHRdSy9F7t2xIYvxaFiXVl8dvR/O42VaqmXezW554XGgKdok6D+Z53u4YQYW4LP
wbHQ+I024BbKaNA4FYX57uFbQ6JZOAZ9LqICF5803ucNZjiIH0XqtdSFRv2iDakWNyjPHg+v7nJ2
jrkaDy+N5eTG5f+NvY1gK8YedkaU5hVMjRKNqf2Hg9ZZefWfScnbIVWDDpv9HQcuuP4sjiFvz00P
CuRWPimzsNh0Y2EyzvTOt2WhPcaOiOaEPYIYveC3eFSnyO7fRL1JHgYYcz2HLi2IjbPCsY1lrowR
o6RpAqH2fAZdOR+cXtZ+5uc5ULxmLa9u1zBWzldGhkUcHQ4iTiBfxGdYFn/zlLOD7dfUmY0RHVOe
nTPq0Jc3jfu7cHhxk0gV7Y8sC9ZoHggtHd+e8xJQJ/qAiqRFvCbEmZhhxqt6n87XhSeP0PCV9GNr
NWeA9LWP+01QZQUc/QYCbxu22mYoHMHPHCEfaVfXcFZDMsuMZQxagn8ZCtHI8IdXHOT2W1IBSM5V
xzmWyQdHxTbiUNdvF5P90rUiH2gOT44b8ozFREc9Zl/AerY3oKRbvj8lgXZZYaKLfukuZZURF6OU
fFC9HbyK45QJnMN2afej0OccasQG7DEF8aGlL771M1hbQx0RnafuVJSfLHTd3kqPIVSH9uh6FcPr
GrSLPKXhjyXFw4QZ/hZaKOoe5Lo7WHD3fVs26shmd3g4c3Hovx4L8QZsutUNAC1cT8Mc4PX/a/24
ENuadvGP58kh59uvY3/Zlmworot4q2ms9ei9fE1/FvAQsS+iQUdYBg8MaSUmDtpNYKf1+HW1GvmD
nLrP4Wa5j/DD/brf9zWiPl+JLNOT2vYM8RZqVp/tylCBkdWrbyES+Gtz/zZW5QJtojPgCmhWa22F
RAWwhSlyFRYiklLJUTXCGlTZSuF4Gy25pM4b9GlMo9inNprGFxNWuVT+DuWo2iCW6dlWsmLmBI8+
gt/ypFyaJCwjwe1EtXQJbXgxyBYYCqXIUUk4L9vc84zBuCjoLkM3tbm3QQsjSj0FgeWxxe07KbS0
eWYDAGpPUoicpnku8X1Gthqp7BCIKHEEafQKDgYDVfRFuRVHjhfyo0kfurwXkjzWSU+7wAs1Y7Sf
1UrPwttCjd2dxPuwedOlsH+ZCDwhM70VqqBh0QMeNvU6JRVAn7mu6Bil/LS4Ai2hTm7Ns6VZhitW
ZYksP9I/Jn9TAOsPOQEnUoC3w27emj1Z+PFMxM2e4OJelv1MPJIFUShItYmBZ2Wyr0Uw83ue8p7Y
AVK+YMxsN4g67vs/xPeyACprw120MRgq0N+PrX/3xaxCRBCgWyNeuw1Sw9Yd4xpvxsXHDT8iatKq
qb81OiAhx7oEVQaY+V/UGeW3UnAZItFm7AEfD7FP3wuNKJNs3Kt62EVcHSx+ncdZZmeA2Y5Y4EZf
39aeNM325LUFoDkOniF3H1yy0NzAMpO5o38TxUYPQXxvRmb41F4azIwsW4YFZqTww0nv/9D8xqjj
IL7wx5RDo26vppM3EoDRwGbNoASEfRGZZ3LCUctlBfwFaG6w792r2Rw3q8HiPq5wTFf3NkzsRGvk
HELTCey265IgEWWrXXnCBrMwXVtWFPaq1CtwuUKs3NJ7+fDPzkDSBm054Muyk3PfWxdOIcH1swoa
HSI8b5TB1gzmP3fTzm8wLYe/wxFa17p1AWQDnyok9AzeBTqsrGiJOhQg1eKruHurFMEO/na+1Q1T
gO3n0FuMfbSqJ8pUuWYTlLVNgB2Co9YhpAkc+2Yut2EkC/zRSO1flgcooPA5JB8K+BWTozdMtgjz
gPwYu5IGfol/lEAUrojd7fI8Wt2Gq8ZXaUviedL1ALXwdQsl8b19nX4DVGjEfk6+b2IzD2JWyUPi
VSLx2HTkoFNt70CKmRthohbcDzqFl1Je2lqWk0ug5TPCyW2qGFww2G3xIibYYqdCzPInYLEWikL5
S6TREkAapiBFElDz0z1se1Gw5l/9IGoiemIfDuL1RGHsI6lwrRM5W4rGaFtPfj2S0q8dslBTGvFw
GzM4aRpMwNe8VCXfzcCaXFjLyrJiJb71zFMuiDECcrgKx4x+hbUpw58n8oROwcBZ+ihytIdXpWU6
z5Zl0CXch2q6zPVQr0Qy0nUjRu42v/ncTZdv02XvJ6GtIiSA47fXlnEhA6lKvZUi7IallYbqhRdM
x35Cj+CURRGZYQuINIFM93Y9wNsQMDcF9IkBfZpbqggw9hYSdHSvORMFOsC3KYWHT3VAxzoZApka
ViHvpaLwNmq9cSXPlOMxB4cRS++Pow04Gdu8indHRr+YzDoixwgRShp7kMC8YxQDmXCFqNXse4NF
FlXv939vPJwc0eMBlGiKQJgZwWo80Wmk83+Id5A7bZICyXeQaIqp/8UHyMFiuAysW5yRhQnLAK3a
x3j9fBy0wz9v0ntaiW0DQxdPpqo6hAal79nuMJnuFTP8T/orFSOI26vAM8049J9mzNK3jHWieZUr
p9qhLLizuBc5hWVlwdgJy6JqWsBr0aMg9QHIJ39dTryTGFtNfwtmnbkuC8alEp4lymcT5EdIRMDl
PrbXKecdd5ndPmsWQrysFgwfkXaFUNrWma+FB+SaiwgpeuJsGnvmrqjv/C77z0HLWUR64ZeyEYsV
JKQpVY86sijlusK9u3GY4nL4NoiqJrhPHOkmvPlc730UnHKn4C34q8/UEv3iU1epAh4keVKK83lu
pbKCqv7FFMi0+QLE+nOUNO/N5eidbciawxVC4sf/+hgyNZocs+ef01I6lyUBah4NlRaSVdXcFu4r
i+wYPCh5rxteI/+BWWXJuRNB/foBOMb7qPGn8a2J+85VhZ7eJS/q3CjMwLWjoiNUBlI4ifPtgvCf
f2wnd6N/tHAcNEepoK3h5mTmwMUEzrxTSRd1b7YS1hZHXGelBbsxs6S87M10r1sLowrUjvt1ZAI0
PMXv2nCAttWJ9cwwXQ0qaWBcbTDfAHCwt4DV+aCV6QUo9s3z8heQipiV1YoKrA6BW3IGIAttS9Fu
OJC0JMmRltU0u2pzLuudc42A3mfi76iRSvc6MEMqelokNZng4jV/sXInN1dFh2Ioc8B3Wz1zXv5I
66JeiHfgXz5iY0nZV0qH7fDB9wWT4CQH1uTdzrEHP0yINkeO7SS4MX2L2gGRsTzhMmv1ELScV7rQ
fpitoyn/EqmOtvAIDerVVBbQ0UySMfEbq+nSc9bOAMWIVQyFo0Z92V5sHE6UdrSJXrrJemAZFfYl
g+jMKhpBMUQRcW4L3iDvUfuY9VFSnaSD4HeYMhwfY3NvtZbKBu7dx/CUEBKlx5fiM65ez0VfSQDY
H2sjZ+mSnk6/zX2l3N386LH4NrknNfZlHmzH/nnNUKMb+fA+eBJekE8SHamxczld9zwfbTbicXTd
y8NU3OQIcI4gWxGfMmQLsy0Aq3Mmwk8I0vHENWrb6J7VvF5PK3SWgFd2UefmvCro+fXBTm1yOsKM
DaC+7dGbXCSKJHfWyOJaJklvd8qw+zg3ia+j6Sh0keMBFk8lozTAvBf9Bumpycpd2BBACHCflhDr
rbUlIbNihcHfZmiPCPdYrRzqiS9qcgx7lvBpjA8mKPjwS8ZWRs+2u5n6iUlIG19xWfU/9mulf9MY
ksyIu0oYl4B6RdGWVTPNvsO1JotY0cwrezRHxjxjTtwGmZqhUUmGlRu+Lc3tHtFLTSz+Jt3rxyVi
czxRcCgwq+/w2lVKt8E/EN0fk8KedYZRQHW9+/52pRSVLvFKDsoTthZOV646y4e/EBjiGGyvosFi
sCctITy1kmir2IAAcWlwlsfhEU3HsHKS88DoLRIjpCgoqA1q8cccvXxd/3vufXD7HrUzUf8oQ4Sh
qmDSPeey97gQ0HtTwiQvrHHeZ95+KvG9ni006vYZT2/Bmvec0ubF1dSUUwTGZwkcpikRmZaaO8H9
NfV222QuHkVEzwctmypvleQRgaHoEUHDVLdebOGgZdktTg3hmuyinIPWQefcFmfB+lBKG507bRtm
n5bgXvVYuPCdGOZdw7t06h2Ert4IAaZvHW0N+9Ngc+kpacHTSG9xD9vuyxrWiJ2CNHEPcXBYBCMF
kQd3ljI07d0=
`protect end_protected
