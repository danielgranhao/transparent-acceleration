-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
3/CBj6Bzyq5Ad0A8rYpMz2v9rnG+tHyWRQXQgn+GZNapuHUpXItvOSVHgtBnGWan
nNZXPJFOzPRdiLt6J1n3aK+FhdO5yZ7EgNBljRHTspFabHTddMqEgzsD04MFV5C5
kXqO7WYydhu6eVgCZ61abUTRDNn+ROfKJPABcL44y1OBWmvCJhSTDg==
--pragma protect end_key_block
--pragma protect digest_block
W2xwyWnqzEKKapv5+NKRSaEOjO4=
--pragma protect end_digest_block
--pragma protect data_block
BgbKxAHO/JI9UrT3CbO7fUbvnFQ+eE62L3Ez90whPrrsHPacqlny+5uLh5N1HXx9
HEuWlXJT3eh/7P/3kIj1lX5p0jaHF0iGD8DsEuS2d5gXPtu/9pr3Ql3eyZsGdRPP
AwURuWrRvFsUcAaVGyTLzwc9M87I0h9E2akith9oZavPdP5o4T3v0u3109wIBfj3
pkXuDkVPBelpEY10PYC/74CamD/gWQJ/+AhfcDqwEHTW2fdhaa77Bpa/P5fQE8sO
rhqGNlRyjkQZAVdrqq3Ab59HXlw2c264bjkL5q5GPHHwaA3A3JoLqdAFKI4Qt7sQ
tYoE8+VZkxA2UW01C43fd3CutKsf4mh4PB6Ze2WGwXUMYf+oT60Oa1jfNfTaRz7z
ao9JQvEIuy2UzQth25JqSf0rJSN4BSwnCTuD/Yi0VL/GFg6e7hSLODE/BitP9Xab
OOsFX/GxQm43fNijmRYZgbWGpFkWSb7i3dM9G+JvyodA0PRANmTw6bWjY89kHDGy
2ncqitx07/ZIK0hW5AcgANr3awZf1BqcQNrSiZNccxEZrT10di6iVzrQMuME++yk
+wr710EO0HUjCK7jd0ed4VdHHQcTkGb3Ie34x7qI1zEKCF3S3HYKacXmZIf0QIQN
MpyPnukS+LKd6B/b/z5QHgzXF4Soq475P7QroRfy4LIza9/61cC0IWycNRjV+d9p
Pa6VKHcR0f879GeeHj8+c0AjaSk90FPwRer0biqH81+uKaO5c4Tjc3QkDZ+pHXQm
cAF7B8Udh6rSgSQDM7b8OhRk+8H89LEs7m1S+RMMp3Lrv2iuNjLyzbmOSr77h5Ks
Ie4Vy5ChJ08Pdyeb6heMcJEbkwKFskf3LyFP5eYD6rGnHTm25H9/ocQzPMuWrB8i
Pmj3nI+Ql5soTCPTNbIikjUAA0CcG9YL2H8tSHH0m9LbQ3JUobL1mFYGlCIwRw5X
kyPGcthX3kE7UZaNfzZsoKI99OeXEWQjD6SMlAPAbd3M01s9a+TXfImCLU0ALQQm
rR1DnMwk5wlEOLeYlYxFYJcUv/t3TwvOkHl4PW9l2/rBWpu0BEy3IDXpfPY+nQXD
dHdVFLcB/Fy9CxHdoyo4HfphFvHuo5GJGc2fhM3xPFyERtYr7ZEnKZNqNvc+VMDA
raMr9L8HIIo7Mu4ebTMeLg3EMe42a9uE0JLYuFc9TwqOd59hrvSV7YABmIXtoKiu
Zy9yf5Z0oZKlSTiGYxq6EgV+mYS58uJ7S4LLWaXE41w5nmIlV5saxtWfJSZXZvwS
cAPIMYcrIQLUHYx0k8ZAFYhbnPiZJlNjVM1BgH+kUrXVj9A+zt9eyehVodzyxrul
pwXJxAHdZCM+sX4rxjDwRPsFGKHd2CWUQmAG43sz/pzlk8XP5RyrQeoF3vN/ocVh
PjiUw3HOCZbHwjwmK5gr8aGIAKO0cU12CDZoBsNdA+AjWi60dsmgOXmDmogCpuE/
l2FPtKiS/ZB+gmhOYeWqQ6dkWsaWjEzxsUN7sqIo0C1YrkK/La6pAT2xFeG4is/r
pPv/CguI6SXppluiewUvcTKTM2su/fsFcOvMlh64IzC0GGx6lG8yjjrI7xn13jGa
Se5obed+lTStAFKrtV46nrDfefYnN5K6miCA29si4OQdoQxt8kdhbOb3vO9AuJYQ
o1J9p/BzNIFEezEmDCLFqufRSGIHtuTFIaREUUehE6OVBfiHkGSFc5s7H0tCElIz
RTqHrDmTwF8SL6cyh+FJL+Zz9IhNBrFNojwUMmfuUmPlJ3N8ONBobA+DacdHyh8c
nVnheN1QupzmOyNs+480cVQF8q1z/5DPLPVjVKTDtjjk2hYdaU1RsnGAo2CzLDrJ
f0t0ShnaARXx/mWp9ir4cLI3CgANfBDyUYqyWJASTym9vx6E/IUAmVuscU9pHFx5
gduF6Ow6HhGERT5AG0Juyni0FJSoHaWIDKf0ZUnHDkB1Sg+emW0pG72djmwsF93+
mV64jwykKQu4WUv2awVQzJCP6h862swn3IkgjLYzLaiKNnTnXQJJDVJ3xGjdP6TI
KaYhNKe75K5AE9lMpALVoDd/UmWtinn4T+osgxbfxLUJfppYahy1JgWp7nx8cr+h
F5xZrOogS3RyE0KdNAabvO89Io9kyZbaLZ4odKNwNGr3taGenAu2QyFtn9L5G+es
s+TPZyT6VvxuuJiLqi/bETVMTbmGJApSnMfKxV/Fb9ymaXnzLXzZ1PrHEiktG0gw
GasFBtT18INB1UdVywFd2Xe7PY+WW4g1Tv2lk286Gm2nFmAU4s0WJ8KtWeDmavlx
yadb6W8MmwEt4N8qnFOSrQDTx1qlr1DcKrH7/OwNGNS55cRNuCwENBHoGs6xa1bW
3RGEEw3VgwXreCgaibReDEDyitIwXl8q4MXx9kXMV3ajekjzxGPebLY48GfqaLng
S1CZ737qpD48L0cu6hMeCgR+RYi2mRRT/ESn/5Lz3aP2S/dMIb5HtRNdmvt10Sbh
FC7w8f8nhbs6xhi2e3ZkRRAT1/gEs91EgkaPcN/JSEnhmuTnag3UR3JYaHGRrm7e
e3yzyxdg1+RBCVSuPEX/KmeFqzpuUdgXIMw5IQcHAJHcsksrdb8lQKgZRrvIK0vh
4uz/jpjZMpH2UXfhwPV+rEvLey7Wxy86GGS4Mhl1KHJt5potHDiaWOgaPWOhyFyP
M1kddh56Y18NRKsUVDQmmqHKZTOZpAQAf14u5TqCmNWTTroESGa3b8fQf5t419wE
CSXpcjVvBJ/B4WlVFCMgqaJDuGLkIJ+8KKjyn5DvAdpINECwZz0HW6W6MZ0PYBvx
ihOV00vUiJ7SDWmNPcm7X0qvIpjBcZYos6V58Nt9L8k5uOi6ZHTyBDgGyfxdp5Ef
ydScROSD9XjM3aacCOzts9DEPO6dlDUYMBxWzSKPAa4RnzNvrVY0MnZLF9mjBBj0
rbBBFjDjONSbJvP4aWPLygs/ue7zZwPE/zcdnHHpORsBmLHOoQ0rnfEXtdmZ6ZD8
XQTGg0x/BwGhRi82PDOaXwcujbXgioTuE2qN5mLHxc5k7ZRMtyVy4i5DM9ngtH0c
9qBiz2RicoMV68A3BrU051b+K67IYEeIRXZp4WPGeAarlEKTT4kp8KmhxDcsMKnL
n27riNBM1t+eqWMcmuiFzQ+uoLkIDDy2E7LHcJ4m9biA5YcoVSV2CnFQ3fnWzQKr
eJKlt2dWwoPAQXzXuHAXQFNPhGwbWuCh/X6bRRIFG09RbqHGWcDsH3KVkVpWNqSE
raTrQNobh7WPNCT1ulW1mb/MOHeB8V4xbI/NFP/dKqe7QHK0GArWSA3GhoMe4olz
utrNng9GhZGLW8qNbm2s7IMNWZqVj3e9uEQ5Mpk9lDB78tTMOI1IklPXHyeXjXQu
fyXPCf+/asFz2xxR4EjwGdcBsH0pDRyCKRKR0sebvjd044aPzfoYW8H9E/0atT+l
FBvgODJfeGHPEtBSmHDi//AR6z1pMd7sYZ/bV4/Yu7Q9s5z6FKKqgFZCKEAo7MIA
qOxIJ1SfieJAK2HMTkZyoLv8vHxfMErHmycSavNXFlqG/EjvegajX2okUHtm+cUZ
ctYMoVvj2+h03t/BtEOMiMV/cajzrOdSc7iV6YOeNJ3ebbMjIN58IE+GHPiVei6Y
JgKKIi7ix7DXL7HhzjQGbCwcMXWC/kYSZLCzYLw8fVPeNNoiWjoak3vnWUitK3hN
S+GJLwVmmI4asQYFnGCQ3g1poYNapxCviq4TGaucTlofcW1+CzljmQ4EPRjHe90j
LNFQSIBcfHr7vDnecb58Lb1ZvcLFV0e4q0zxdV3cOg9/p5jDbH3uR0jB6PoM5/rt
y/mhPoS0IjB1ML2aZHwtCTqadOJoylJmrIoWH0AoxJYCZ8bfLrq3ihWp2VMb12bf
q/NAOghgkMmc2mM14v+bdw6jr2ohnU9J8tFRQfzP+JSAcuPgeGYx6beXFhvuQ7fR
0TvVvVFrxLmTkmKPZbEzAgZSCb84JFi0IgPqrXtDMmT6RfokHyAdUdPG30/KieGL
l4MPw4BMQRwhxmVFVnwAcn5LxVLAK2AnYLOwMr7viTWYwkuWmommAx2bjaMLB7iM
9Fko9w40SmwtgJgw/AV5RRKSs4opdYGCWDP0jyBDTi14V4HRTlnXv8fi2c1ybgmv
XWy7Bg0K31erGkvQyWn9PjtjMWDUlV87qTjUe0UDlUNuMMWOso6e2FcrE6034HDz
Iyk5zybB3/kW+CcTYxA6iZf/Cb9PP8KrIvfZ9f11dR6t3Fik4HWyyra6SPHgH/QW
mILMpo1zmz/eumIdhnnNlALY5pBsgIbMc69jkQ26SQ8RDpWXh3S7HBdHKWLD4crE
bns8DnKkGK8+ufucz59HqADVL79xpUhcbRT4D2DY1sePBzGb0ozIczjdf3Mf0ZAT
u6Vl/2Wzt5nWJ9DLkpP7xMuRTUNwCjBUdzATtBouyZbbO/6e2ic4xtV25qFYbdp6
Zdpf58Ip4u2Efz4XWDni9QS+6gNlshY+fqhiIIQC56OBdfFXYoyMvrjjR8r5zHl8
YVkfgaMH6qHF/XiuMRM1jhd3QFC6vPRN/Oqq3e1iKCxBDWq31YdU+B60sv/4f7fa
Me3s8lh5UkIibowAt5MI4YHb9jyMkyL028ebtFveoz44ioujfo5VKu7Znq4mnLVT
Mw7Uirr2tgUdyk0+uBRNrer7R0D+raoTX2bcBaLewntpMFVdWKa7ll2ASUEvwrs2
jn46EGThu5rzoTzk6Xgo/cqrRaV3nj09eFF8mYkLbZl7S8zbdelDERZugZ3BRgep
/2rWJ1DO5bgFA1o4mBJ8X7nIGIqjwC9H6ERw9Cq4SDnXcuIqj/jFEpvq/F51WNuU
tmJUNOYJ6udpnQejFpNUerN+9OSrkMx5Mp/nYap/JLhK6sKQmP527q8P5CQRrNKi
6CvZtPSG/dr3rJu8XVP2xFLIXWDPcusYswT4ZUsoGCqtFUF0JNxqrnTLVKCW3sla
PKzeQ5cSXqgKxGkztb3lC8pZzyT2SvwLZwpxI+osp5/upawxsKKYWM1ipLR377rR
kig1HNSlTYvY45xavppxLK4cwo4/ZJXONQfcwuOQNErln9GnuFPfTHuqaES6XC5C
Y/tHXA+GXe3zC+JUqb9pjtngRa+PWP73y9pPKHLRaJfcFVNUXqHYPW7rDbtlDF+O
nKzmNgO21qXgHFkqCcf+cCBL2gDC2RfJblVY8odjxIq0sdKyUsR8dPqzE9dWOKvq
UTEuwQoHFXgcT6JPVqiIi+1gHl/XfZ0rVZIEiBZtLAAlrNEuCT8vvTLwBU1Ddybt
z4si5nsbpyZ2qsZVb4BMXbfVxl/2iqpgmXD2arTwkvkYQdlKSa9QBaHPTzhhI3pK
57KIsnjPuTdZS6WpcCLT+YR7ofi4lCfmdsydSTPta8FL63rbGERaEsK06tkwXugI
8tRXMLCZmegPlHWOeZshf2UeSTnnkSCPMYTCY9NQC38VX3me023qJiK1TFZ9UwWV
qZ/6GOOg+L3ZFPvuGfehMzW6EXmrkNovyf8CSZFL8zeE/RLTjVv7OEWBDcTJs22W
uYIScGwAnNhXbmCyjlA0hceUuSO3Bl5s2msf1ozF2Wl4zLJc3Ei72ie+f24D/jeE
AdMloto9gOx2nSLd7DUSN4SUNaiTV4v6vuebEM/XsjkNLfev/QVaS464tHLpYZBI
KpxcxpsgRqzwha2oFGAvkx97D0il7IptA4Jxe/oLXJn9cSryAeEGo47qMTltXx96
kAv49RTxZ0OrEQvJwXtgYv3qCci6D35ux+PpV2ApSe1iefq7LkJjuEfCfmhjRnLD
MqSl95b6tFRoLONJA/RnhBZlgPMIUqKDsDnIvmm3AtsujvEfJ+upi1hEfriPw11N
NP0AhCBsVDMRpevIGlH4FDg4eDt9oXhfTa2+XacB6U5EyL9zgtXxC0Figou7GkEF
ASDRzAn6N3hhCBU661kQ1lrdkEtOYORPNLVuxPs5jI16KniojWpIeavGg7F/KTzX
L4jkO7mU7yKD+MXvKEuiViXQtLc7gs3jtVXaOm2nsiJIx/oQTo6SP3Z3g1nBdBXo
oYW635Bwbo34yZEWfDPtPAQjY5o/vGp5JMd4QGGc180Iz0ySIWjL/7BsqyyBTA5E
IJqB6qRNZvDNfwOA9ztTh5oi+/z3xT+qDEO7zp8dBgxU5IE8dJZCQC8JssGuPgx1
TrTuoISjK53sHjgie/qR4H8m53H7WpQV0XYjgyc1Ed+cewQeTkaJYhl1PvfkWb1M
7bVVNRLQGk+XfrLJnJW+RZaKAfHIqXzbvU/e9vbjGxoTAv1/Fab0whJebyV/CuC6
PohyAA1zTctLlSCNz8opCKF3qVBzJeANbX4MCY+X8WEOLW/N3M8aRjbN01odkxmx
fZWURpJ6sqxJh4pqy5vWxtLgLh72fBAkrsxmg9zimqkv4HqfMOSSWe87svvYx0e1
J18MYXR0M4OeOlfVu/36oRCiwIRBYdlyk02rRAWq+tvuU+WFcMxQ8ECwESWGA8Oi
6sRVFs5KF0Jc7pqs6qjOgL7RJGQMU3I2TODXiEPVwyOZZ+KQ/oVisDLpyvsCsrYu
+UoNJBHuS4hMMW0ISyAEokajlbIAw89o0DZm0ckdjTlRUzq/txJ4iq8Ru/XLzf2R
2tmps7vGkMjraHC0hIQYbxU6wPxNVhUdfj4YmLA6xjYej5onYhMxx8wS/QRtoScp
3Swq+H4m8zZQ3Q1TXql6sDEwnRVk2c2Aa5T72reCHLEccDy1lMiCWvb8Z0FnEEmL
vzhDM4+f3YoJbbtCtOvA/IteMUnaXrbUaNutSzKfCCbPgulDsQqAahyD2ApMVsol
ARdhkDaHX47Kzm3jqn/VN56/OY96QJHnkF1JC6encHWafMKWX7VFQjucM4TR2cHM
N9rXsDNSXFh3Wocy4fvZ+lpCYS6FJS9bpMXj6M1kJp76ZiKGQk7OdIuQFsg3Yr7G
HbJ08XIAzihGLmYU6ZXPWfffsd4kaVsdaW5lcNBkM79qolGwO9cfkICH8yfkRSts
g0EyHvyTl+I8FgwgWmdvpBZjmrHNe9hPCv2hrMZHL+PIKlQ7W7N7albqxtTkKmJg
BF4s37ogofc2E+VomncO8k5GcQNo+JycDIqaL5MnnHsKI069WtFHzz0nWiETfFGs
H3iKM57vX8YsQmqJLp0ND39ZZRosG6q2umwGyH/AjAVVou3gIqNFi0U3y/HaREOQ
YkX7zOe6HRJV7+8NeWJWsiuE2cLYI+ta5sTx7zs0BQFLPuYlsuHOOxwdK5BNUzL7
Cy50rc4rYGSjManeEUgy8ntXiG8ePrNPf3L2/GWWKB933XTf19g4z+mA4Nf5QbMF
/Y2J7Izk1SlUFtWgk5n2ezsSs7AKD1H9pbbKgw5hipDAMR4S9iTAG+b5Cs7ZOSxT
Vrmj+hwS8Gh270xF6IsJAhkqnxYczOO12ADmFYqmanbNo1YexrprAAwcet0TrTsv
E13CaD2IeSIw0NI7ZhRFskxh+IKxKsQGJxveUf93achWdp+Q6njlzLt33d1LwxoB
JFZuyNgYPUHnyYmDrnrURrjnWg1R9QETMwhwRHN3VZP76stjC6dsUXQxtqdmPDHs
GxxgmF87xBmETnQEErQ6wQEvvEIBwIZKUQPp3cdUqtrzmGp/WKCiYk0h3LFnmshY
a1XnJZXJ1aZtQQzbCVe5aqtCOOda/rUyDBSlkkbR9Oap5e227YfifwDYncPlWIYv
f3faSLXKB8tCgyX35FTIezEaBt30BIvvV3StiHTJK9LnYD3vcWRoiAOQj5z60s0D
dMlH6OZuS0jZ1wBMongoNgHbCFG6/StUPcWhlot/zOx61rKH1Ae7RpkmC4H21HIv
1Ooti2JXCD/jmIoCt841cnrkdzAIY7LMrBVR/QKjnwyzi9iJaEuK8I8qHvXkoDVw

--pragma protect end_data_block
--pragma protect digest_block
r7FkHdBAKGGoq43eaZ4au6eWCiU=
--pragma protect end_digest_block
--pragma protect end_protected
