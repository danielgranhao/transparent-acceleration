-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
3/v7u7TKvsBw5qcg228A0ivbF2VOHcKP19AGPwnn+pms4Nzn6ffpA3Ts3xutV2MM
HiyYwK13vl+G75I5j5FC6fYXZZVzZrtEahugBBtUxjNhkD1CtTAT9uqlU9K7pkK5
S4F4ZAzyRwx+0aybS0EwmkZ+FzTt4gEsaMv2hyPySPc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5712)
`protect data_block
3aMTWpJzpmWNV1ZknLI64Tixqn+CIHhsfc2KH3F6Lig2RgJ+mst5oXe4iTQM4if4
q9wwuG/rCCpMllw1B3SkvZNsdQLFLFDR+j+COupahdBIGcD77643RuPXA2ibnGXl
v22Ulk3ye+E0mJdDpuWBamY+W3vqqn23u4uJd1/sr3k1YCBXnM//cmCs8aX/+/Tf
2OfN+lF4blYzkhdqqaLCAphcg5AbNN2rzoyy1PHxHOCqYnnJkepYQC5JXCNcbh4T
K/giVkspjkt9XJQcFO6q13cIHnifDYNk0XQQMkd5UhwWI+4TegL6ChfANzpwPWhi
fc/dO0R6xeaGVIdRkz32OJcf5abqV0Yq5ghaRopAvsvuH8p/RmcVjBFQO6YjiXI/
j22ye5gY5jH5F5QRLp2b5S0XuQWbbGsYk5Zmr5Gulqw7vHNPcJ5sGnKo74cYm0GW
MaWCqiaITw146DSlLUUZeE5KLyqNYQPwiE1AyUXiId2PgDPnSuUBIkJJX4VMloCF
n7nSA1GLWRVQ7VN5kvx0Aj3izPF3FIBVmPcF8bRetOXjmulButeNtulUKaaxlAJp
7Kz+5wMVcXaPcciHBBUA5bgIYNFzSCzym9af0VIWwEK7qXg/7WG4hVX+hAkkG58o
dmzK0F7h5HIcZAK70AMcY3BT3s1/Dpcskjg/kzQNxTrumowojDzGH0btJlRYdDLR
1NDIZVjt1dXVe1UI4Ts3Tf9hIc7Lm/6Ng+BcjKZj9RtED1WDvDWbvsgLCuePfDAO
XInT/+C3AMn1+Vt9MBFqsEWvPHFTvzlDZE4u3n7oJhk0noJS6ErYPGs2SkZ8EGZ0
blmgiNhff1iT+F7ex6SEFfiGQgfyCbICNGGBsaJ1SGSRRtHBfWIQVRWO+/tsBFia
u5RZix3YRXKGS0ZN3gFHJ/bBwEfLbHc2jF3Em/ZNF27zxwkSCXWHs6E5GqU9/Wpj
092YBlNw/Q+4KViMt+wffEIgT8jQByZ7xaSfeb/I8EmiuqsSbnE9P+N6ntEbHyG4
3MpnUwtnoLIChBub8kIv4gfNF8C3wZwfqalL6dp/4OzbVR7xEaXffa0waTgwPC3Q
k5ZJCTy6XRsiroDf33psIAQZr84DTKxG2yLtKh4xTnmgxBcjTf5mP/24/RuZ8xF6
eNWG8k7GpU4HFz998anC9hZ1iN3T9ZB2ivGu+hGARCSdxx7sEPqeGvKRzzvdRnK7
ATKx6S4z2M1HqaCv6GZpM0tRRElhK18RoFqaiWXbNR6Mv9B0RM8R5HT7/fXKJzvE
Z2C/qeekTGImNqe+4ilpke7y0J+9tvhkX6InbYKyoS9GNS2hQl8mssNGKn4ADOx5
pxHKDp8YnYayvaT3wikOlEYuCTDOanks3DPjOB9HcN6i4wWxGANzV0/CtrRgac64
86iemX5YlgtiDkjIWWkvdYZJ9VccZRJud6K0UTh9C7ZYoJQkW6QZlCqpXP2ESpd/
Sg20ryRKnEAK17Z12+Yk3bmQYl7TMyhOxLezAdnsP7d67zCz9wvstrN6fOTwOapQ
jcj6f6NMLq57yEatUC2OzsbIkuxfnvba6aDzVg2C3u0f+PN78SFrB939moVB+9gY
Ge86l2ZucdZdYCBeLpIwhUnI2XSUq/i6acVaM4fK4Mq9usFQAPBuxuvWj1ncWkEW
4uOv2tjs+H3yrC2s6gZJ7gh/jtUbS36YReT1h4e9yPDr0S3IJ9p3QLkW5s3BtsxL
s2Qal8/KYW/hN8XkPusgpw2UOrW2LbR820s8D7a1IAmyuEs+zcJmRsNp/IyLyG7C
1nBddTdCqfBebY2kTE+1TlLdaKdsgQgGYgIQa5rwqvL+IrW3abbaEMGmMDoy+Hk+
jr8+hwBY5MNTJOVPyjUZQGeKEg+mqoL6oP9VoAzvWgiokRMN+MjbG+vkPXVUJKbX
oyywr2qPUIBLGz7H0f+ruOO1kOwOJqivGcofcl0CnzIuCtxOqn8I4P6Npc9vUILx
xgOpTlymD/D/gE+idJVlCp7Zz3EZ67DjycGVDW2UAtMuyDiS0EjoFVPj1UelVpUf
yW7tZ7iVaL4ncBYykuUUZO55ziOAyqtP9gYyaLFFq1nIV7yQAwxQTuSPvXktNKnZ
MbonWrPuJskaqT4+GZwT9HwkWjWwIc85h6zlvxaeWrvDB0kxdKpJVueUx+vbtGu1
fcrkU/NDBtUq2LzSsNJ18vyrIjoCiwCBlp8nhnW1aILTqGX8Kc/9xVFHUOGMCdRW
529dfrcG9Cp1EfmB+MwgnpoWjlMblbW5xTRRdfOswskb4BPzl1jUSm3oytIycHkp
JHJpIiSWsrcYWb3iphQW8RV2nONhR1dr8/vVAI0bSYwXeMfIYGNmHdzbjFVWi1ds
8y+vsSWnzIPbl7TqzLQGcf2Xdhvmi13UVMI+pdKzCcBPswwGFrEHwRXhUKQjs6kK
Zky3nUrQRO67ot/MUV+uyfoBfL/BZHXbEFIWT1PEWJvAdICT9ciXT4Z9TToLXPjk
4GKaoumX/10Ypa7oIGx3DL5+uSSUfx5HFKg1vtfyfMHf1+naHWCBFVi5ZOFZbawk
lK+6rAIS5+26/5cbUwDEYVQGBEvZuvxzKwZURPJDVC1qcNSzf2fvS+o+tZLO9RFH
peLjeIZRTXOrkY4KqyNY+rIbVX5VmAW4NO+OLBGtXI980aaej19ecFkGii9JNYpn
3iWx+n6YAiz95FVDRg0vMdwaGoiwh0Yfj7d6RqkocpGGWVT5jqSGEJ2sJh6fUznx
OJPKKKAnYHFbLaFciKXhIp0l8rnkOgMJe5ReFRy966yBXn711RDPR8RcScXtqid5
n0rdaOlajRcqp4RXPgbJNuwdAYqS9OyVXexFUfjwWfrr+RDerhG+x6SNjSJx0vab
7dVik/wqNqOlHWsIHRrO9fuGdyNoMF7nOYeOMwZsZLJbBpjUBqwcU7Dg9iczq+bG
NgXR1FOonDV6fia6hEll+VOOkq5afaiNpxyH0yPt0zUkGBFQRdfZwlR+jGE7jtx9
NbAZPrXAL91S7fEUWVZkqFCcCL6NsGOABAbJ9+tjHUUAAbYiu3GUxvdfKWPWCKNg
iQNR3XUh+KenWRxeghbC63U+WLNbpSozYhL/4/T7yKWVwY5ofeDdx9rL4mPd/SZD
7w+DnKsfoPQ4h6mGMwv2RJCxHrK4C/PIpyMMOiwixHhXrj9ms637EzxjDMA03P9C
lO8WDfCVWFOLJoKx+sx1jPJtjAomxfUuFWrtz6bMPrBhN0+Yp8+ooZQ2P9wJr9IM
dmJby48CNIKCnFEesJmCsI6lFLXO55+YpVrOru2y3UywUrqf4/coUG/+o8KeO1pH
8itd6ug+NofST2oU7yG/PrV4L8PTae8+M/92QTz8rMm1EfMfxpgYHrRK4BWL8u7F
B8fRmnug+AK/0roMqk7SITzvFQ9+CgDXJBykxcEwWvH+xw/xE+OV6cK9d7R70eOo
7JnAIbNIxnJMeNosYwoBbFXhgjcBChFj04HQCLKk5IiDbocuMc1y09pj++o6xuNY
5fSq0oH7BYBTIxYgrN2vrrqk1IXU0tI/JrIgFm0zi+A449J7+vtpb9/8CVBJ+Vzv
26VVDoE0O31MBhiUpIS2lNxws80MdpyvWHNkUxR6Yvtq4BBNR7vEjBDLHOsRyQCL
MCSpf0g7ITrXcy3Li0YFl0uwY8PM7YfFuhwRqgryLEmjK6vFPEzicNy86cFsDxo2
PLUQ16CxLQON24okw8Jq6cGU5wLXEEeAbNCAlAPPK/K8kK5av85twE3LUbQlCZgi
4SUbzE34vgJdVIPUFttTKzjoAuaL72UoKGxT29+X9Om8beQBifF1zY5XoLfLoWvp
fElsM9hIdtelnv72HuGQS3Rc3pmrM8A81BDXpI6+9crrw/8Q2ayO6QiNaIslH8+T
fysL+OHPtgPbXcxUF34Y+gfobKTSjT4tQpCr6BpshkqnnzyOsKfuDJC0Ccl4BcW6
2XwhpUmR5C4TK1HzWWJho7jk4hdxKLwnvM5H+kCBV2rO+ihhbPYIl5BCa9PceysR
5QvAVcuptfyoJlpgH3YZYeczS/ZFhCkLe+v58hbjZQaFP0tSLNn3Xt/uhwoZrNKm
ked21saUnaXnayp3+ldQj5R1BTCmxQB/RIPK3VCuO2LkxmEpeaVfWFBmHezfGOUf
wb9ZZ8swt2sghUEOLyf0fJ0VZmJ1PzHqetCmUHSEOyfEGeO4ErRbBALT11j0uUR4
SLtPg9zKDHj7moAEa5O65Eu387cWI4dYuaHJx8x/f11JcfMsU6Rygf9EDx1q8BhZ
Uvy17dOLAxwSRju6p57NEbYc9es6TGWbP+0DjcqI0y2G1txGSsq/Ky9rUetTabSm
06V5rL7tkCj8sdWgCACElHQWkydxA0U2CUmiqlcZN53dth3gDbt3guXqPNPE89wo
K6duQI19JKRcFHO3Ki/eQN9aG2Qc3PU/KJcQiDfLfkFyb9GMaPQJgR7X0poOfJj5
qluQUeaW9waOTMDd8mhooTbcJA5ts/taKlHLvj6ycguz1TSjWxtw0QoXtiDgChuR
043w+UNqYi6cCCsCqsSABvPo01zqFZupOxjWHYCGXkaX+6r+ZYBzm3FM+pbO6oWU
8ysbU7tUMHV0LoCFbZrquI4K9CvsgxwlLMhsnNujadEBX+e/ebkysD9pAipRJzKq
DVDjA0+j+qhSTxCjuQj88uEvHI+N78lpvgfAnr9I6aswFLAk/rw0CvJNcpcoZwpn
9IpOwFVJDHOPyvVjvcaO6Ir7fek/hQMZfP1kx/fo6t69eNF9qYOhhszoCTQxY6Kh
dHAV3ZCRiIjiPf7SjSl4i11daSkxLHcFw6XDXCYPBF+PXGqlMSR86oyh8aB6L6mm
mbeG3YLNYHXiymQQZQb9SsJSoO5GlUK/TqIbLdU/3huCyGq673gf/rpnkQdiDpgi
plmJhQJgvDQbNESnHzRSusgGe6q+wgTorQOhzlDjDiiJA16aMwXxrUEw9f3ZTeP4
6A4IO1RTE5WeBbGacOFUaubeozI+kdaEwblq/rUaPPH8RMRxOHQz1bHitRb5gIiZ
5ChR19ii4r+P8ELrVGm9+gjMOFCLqW7QXF2+XHOO+GdRNUr3iPw0ZNG9DjvWzzD4
KbIrC3/kKOuQxlVoSXfYHS/SZKAxi95pQn5w6/UJCZMYIYS5Ibuc1ThvzBW7l0K5
+mShJwACbT11Dvl3rDOsGcVkq8nVUYVkibl4mm7YLhVJ1YT00gc42a+2GIsCAR35
dzprJQhEfH+L2hsvYjqZ7xsK3Aq4wVlxexfTVmWtwdIAeEzrquTB0qDNVx5AWX1x
RDllecyS842tC70UAmd3FbpBk+AmDilIiEBit0EDnRNhANdHeXajQylfdwHcKEtR
9VXECyzckVoM0mSOCIwantNG+vztONAlCBH1j6ZvJdi0vInRaTc6VqIMqpeaH+gz
8UXODh4o8jITiLLVOBwZv+eJvukjalmDPubYDNC7sf+XDmC8tdDr930RJHTokUPR
YEbTE+9SD7RszeHIULTfa6WU+1NfET5vv9s6BLYbI/xyiSvMs4kRfuI9FgUbfHzD
HqXly96EpoeBxs4GvIbLa4GHkjivRRXO90AYxVBNoX5KZr2pxcHtGG5UaR6mskON
N5+dB9c2sp++XuveQ4v3PGyZn05X6fcR5+z3QnAJLUoJJZ54EiMJV3ty9NxADHxm
wMf96HHpNkR+oYgr1JXwKTj9s3UuYoVdihKU/0H4SQXVx16YHEGzf3YYDWonnQmG
ZWQJUrAi865+saNWQ9Od1yQeFH95rvMCDYBUfH5L+XrE8qckFSY/RzZuzLu7RTCe
iSYIqATK0DO/sbUR1vG9jMiWqTDCFnXCjFr0UxPOmDkqxwZqvTeGIFpvpgj55TjO
KPVX6hvIjqciIYy3v5yFYjO049V5yuW4II1f64+v+Bn4s1VgG7SEt03pwmBbBL+u
ukazB93f0DaFVNM9+o3rS934Mi8DsYT5WN/ydtyTGQR8bnnSMV0aFGbHAKiSV9Lq
8TJVJ2QxY5oMTS3Y6hDayY2c21hh9DWtcHM9TkAPKsQLZy8LyBKu3hH6L+D9UGyD
ajN1hx1Lc6mrLvoHkNItxQPnIm3C69QFosdjH/GaZrILhh4bFiH8xwvtxxQW2rlK
VCUIha4mAn2TmLAGJolval+J/h+Njqcp2Ntm8Cv1qVOO5qrNWySuGNtqTPT2n2/E
Y40wOO+Ui3vOcuPtkbjigeuJjW+0mjeb2mudbdhh2FBAuEqpQv55aQoU/9OgkLQu
GOoJaFOjaYY/V7QGPxSBQgHEZPCHBAbyuwMqewumAVqrGEOIQ+NHxfe0/XGPKIdU
7PlMoq2xObsc42CGmuIPiHiZ0Eq/lJXzH1GoO7nFk3MEzoyCNQofqi9J8xNkq9k6
Tpsd38zCxIPG0FYvmVZ2DbMedHVJxYwqaHumeGiQgXxl9whf0RF2PA5U+BuRGn1B
SlnnlSXDWlhghg2ljjpf00TPZj1aEFTkzEEqfY0h43rJtlyGiln9kE9l5+PNAeWP
4YBTY9sPPnJFgQ/4fYMzIcpqZt94XEVshIof7iqquJ6Ju3AaugXuX3pSS0jq32W1
imyH4Uri0T1rnTofxWDJoV5Y+bUIoQ5Heyz9rNsunQdjLZIJPj8o080HKFp7L4TB
ig+g567T2mTKJUv+5evGjjTCGqNi81xBK8lnOIc77Gfs7a+Mp1lLfah+t+AvsYCZ
9Y/iJWoQbBnNDD6ZRODLRpzdTlqVnHuYw13iF530qePyAxfJTRfrq99KkcA7G7mG
QoaQQJXofDSzg1L+5Gbqu4c5yTbQrc+psNirZb3aDVcRW1ZLGX1ijXtLbp774E2i
c6XMK8dl60FLDb549tKpOkbTSWUXs02PUYBXy9X9TiCcX5R1u2t6lsfyMv58OwJf
YFFHnxHd7XUyvv1w8waRCvsHgZLfQfxhoq0jQNmY2GSR4Uc8+wghqInsMQCyyURr
tBane7oRMYBxryxlQxn6ouVr3akvQszeJ05ff9u1x39EI8cXZ3bjtp3MBH37lQWE
r9j+Vqo7DCpwnn9XKtA/mwiFa1tMaoQ5l5uktR7KQpGxOKJj6WGC5oUIIEQGzXrP
715zXjLC4nbFpcnvS8ebdlNUiLcDWScmyFetgJLCYKczwadJImhEbEnHAA0VZh1B
ZQtnRbn3Y34P7LBrLySr0m7zJzEyOVKmW8VZprPebINVfe+k5/yE5lMtD5mbSV/n
0/UWQoNxb7Nnmo/Do/7FQvSpANg70xMH6hFQ338/A7j/fwnaoLEAU2NlGQqmE2Se
qjDKfuE+iBLQkJMjLHklJjtF6tkeEN57Kt4COSIzqj0jm2Zu1Rg833wMfsose+7z
kkqi3jq+MFzgwhpsWgTALfQ8geaoNU8JKISZBsaMH9etHIBCaSBZj+nD1QuAElFU
J0w+myPDUiCFxSQ8CkQrUffNBrB4j1Utp5PFltcNp58ysPo0xOXjePrlEWc2Mq77
Xgx2D8xGfFnAY2NWtEcIXROEmASpxmIl8wdszGSWI1m9wNlyUUe8F6VI+QcFnyJV
QvUBtmTjBVwBADsPwa/w80+P35ZvqucRsGYp+E3LVltXrwxjnQgSiROe5NW2ugb4
`protect end_protected
