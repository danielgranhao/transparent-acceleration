-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
mblgYfv8KKBUjd+ha6dPTuszyJZ2Er79pwuDtm4b1HE7UyKyxO2p0DVlTSpedS75
7UKUeuGigcb6o6ooomUz1iBVk8im5uSWfHyIewivFsWaRnwSvdW+6cz809jXu43E
RVPekAsBMToe8Sx6uLBooZXDMI+r0sDX55BAGIcqQs+X0PU7S6WcTg==
--pragma protect end_key_block
--pragma protect digest_block
7BfUr9N44DYqDLGICMTo0/gVkA8=
--pragma protect end_digest_block
--pragma protect data_block
DXXhuT8fJ4LguxfVaeI+cr4Y4G57b/ocm4KJTedXWyjYt9Y3Rc8TlEanRXbW8VAK
6pxLkxFrOqnx1B+o3GT4+Bh1ekobtqMB1UYIR98+M/sExHaGf6ca7Ns/0BvV1SpN
+5fP65Gw5yWOHcZGhS2+IcPRAD1i3Nu+wgi2DQHymJlLxoDZRarI5eiE1LTv4KfN
V77oOvNDcp0U5x/f9lIwbHmuhJ+2Ci5L2RpMAJOjR7TBTBlfEa2gEQUJp1lHsyoI
Or2YhZyOKEBtAM8E3v1wEBW4a7wdQcR5i3ZsrJ11eS4w2wZB2pr5BsMvPogEYfAy
TgMldda7duPAT93XfLIFOKIlw03LJcY5Q0RogpqouAm/hYTdDnvxWCSX2MdXFw0A
juXvwWjsTCAYPiUTO/nBOk3wQ5Y6WMWXf+Lt/f6gfZcXYkggC5CSg502mJyE7XmS
jgwBM3kpIfsck6PgqEWRNOXrumEETeChur5YFQa5G+UeU1lmDJT6WUWyl+R9IshB
kUmHfPif3siAnbn/xHC5bXwLVbralaEr5qv2aADRlbeCp9mM4bTsCgUA7+SvrYOW
A2jt/mJ8i/kxqkYL0+y2iVe2Y6Ip8nILDEjGF6+xxiFickRKcp8mkMiYdnl9RYdS
i4IaNuT9V6EP7gUinJjcZIgHdiZKXeOJhzf3qCQqNO+RSpSvPH0RH4SHjNTx9d3G
XMp++oTM2cpfWdTdMjCfu/YVmZ0U6XP0PrOo7bIfcyyySkTni2GIUygsnvGBu8Qt
fIuBQ450KpEjB4nzAVfTrbAwivEYG/Xp2lXjwe3NMyfL0BEUTZUyShNvF1tU1Vbs
lVqHUxzxhS7RKUHOcR9iaHBI3BnxhMhYlTCjzgItCPGH9BA03Kf8XMxUCeUeCH4z
nbhUeZPB9S2W/48msUvR6GMpY/eiTmoghK8ZrAaT5adsGoWYCCa52Dheba60JR2+
MoWGJiIdJVxAeSTROzns3m7c2lMxkKPeDJNVRx0ZXJs43ueq4OZT1WZxYBZbOewh
q+WOOnkPLMFtF1k7iwxfdWERe8G5Z4ylsEcTSbyJRt/8zfpQfnt9GLs9RRYdTW7m
SHZo3BRsXQC0FMFfUN3dU7pdtmRoppMsaFMzp9ywhLFqAZnm+lAF+3IKNEcUGksI
tmxmHuJ0UzOask/NJOWA1S2B6aL2VNEZZdaR8FW2bRFGVp+G5M9K0RRyeVDhk0m4
pvZO7lWRb5hm7wRl4Q3Spu43ztFUxdIE4cwv6PVH6Mp5EER9VckHYidGiIK8vMHV
mIEj//8XdlK1wal0kICCCyt2DAQmra6oh4IpNT5R8FaQDbOzqkVrnhnkSbEV9bVu
wBqI6h8ivqW0hG7Zw6tpuL7LYIffWBRLVUKZ47MatNPpIml0eEPNM7oceHI1X2lc
tamqNiZh2bkkoooyKTJC6Ad+75Tg86R8vOQ6r9bPR++yG+j18BM/vVluY3L8L+OH
OPQEGLRp7XSvVCerZZxdZShzkQoyGN7YFl4+z5MvLQuNX4Q+mxtBwZ7fa3BpkVnZ
CwmdApAIgDarN7ifVyImLY1A/cCfdqmvWySox2kNrPAZ01xBZCFCCCBiKJaebFsX
gNrJOA1MURvtCz2QNbsnJwR+NJh5jPh86a6quMVz6zKmn4qS6aH+A44f4Iva/Dj8
ZfcGOs92cTqWaXZwHZMpCJY3fhD38NPA2nN59o6sUL1XOof0vwoHEUAvKhjgYTIJ
Y3BdM/g8fHpObletp2FccJQzhjyvqM1wGI25BJLLCLHKkK71SKAzHh40u7QoHxk8
8ALTg6o4evFWVMGbuYYpvgC1rxx2JXu5YhvRbois2i/WU6gIoo+g9UGafQdIoupD
ITIFKPlIbqGLv2BGbCfbuhI7jAJpMYYmrg8VykpTL6NSGj4BDhSPeFg98gr8DGGv
ZKVUhNYLsgA0vTBgwk+/QUsWxCjU1JBmZEtlTBgra2GC2peEDIASg73g7n/WydS2
x06YL9SIhLnIkW9tACldQVNU4KiMbn9jvDCVstRRytHDB3NyP4oXhUDaERflGlbf
8/vZ+TCdJ56pjGwyfyEEzuI0R1s+tx99pNxEOuTfsmQ0q8Qq5qAVX96368r/cXTx
Kbs9oGJ7PnxYeBIoQpIbO25KQPkg6h1qWGQ2HjjzBzCDocuxt+c1wsSbj5YZ5eQb
ojNeYrcnibKkjTS5Q6bXt55UNf6ROpqNgbBJqUeYzSznzviJzLK/ibhDB+5ZXjxi
pFtwop3NJcooMrJEYmtAYIl0AIUw5oQ+yzvAI7Cfa4rSHqbQa9BcubeaUm/VWJ7/
8B7eXLNeS6iP/Dxb2SjlhhG0+5XfRjWbWLdlnl2zyXL4csWPepHI4l1Qgjpc2D0X
e4Y0unfKwbD6ZIS3h3U+nxakGO8I1E5TvXEcQOFyJcZgY3y08arrKNh1rBHKhK86
/SdHKVI2VCq6MKF1VAFJmcblub4XShreUSavj8azcVii8XsE/5o9cS8TRIVhDh//
WhqSsIDrqCFe+BIefIHBBCKaMWkbdOFijWZQauUEPZTwI2B2dTtOH3RNBeSnHoeB
qm2Rh/lSNt3lpsXjqsiNBb8rYlhpwnyPCOH1jcsgH18gnV+uea0FczR9Dt1xZHMY
xEBKnHapNZuDiMT2nhiFsL/uKMu6ErZCWtkeXG1MLW+JrbuYDIbXct1jdn19hTDA
5gHiXhDnFQYCf3aqscTqZYvFYIZsra+lSz2iZD1lkvBwmu9goIcIFIQX7RrqUfo+
d/Dxg5zjyOGScGtN7TECrKaxI2ePRajT5VEKxXJaFBkF4qyDWa/n3606AtT0Mgti
nf0OU8p6imjrYhFzKMVKEOhk2fmjZ7LxV9Ruqslez237mzSUNdV+ro3Rvk81FjK6
p8dy8hinHNV42bqvuHaIpNIgDlJzLlRr07C1C8JsKjv+kzQv5ClBpijsRJFe278W
5xHiF5oLVdDfZzndZMDXiT/v/35Dda10BZyM9THemxP6pOmu1EHIvfxILBZils0K
6SCzTJL/UvEND7NtMb9xNzuu0FZ2632mutFEc54tVTtRAXtXry22U+Q8GJ7InhXD
P6QDifGtRC98HubkTJfGZqSKoo2/paHXNI+y/kcwUe9ZIEwwkQOTaqN3fiMV1YKL
LECvHma3rvweq0bCnDrsI9nVFB3FX0FSPAnDSnRek9P+qpCX4KNDrPXRfMbLpt9j
TIiFTwgcOHkVa0iwTrs3OCKcH/zzMlY0g1YlQsydAZZWKoNvOEiu7aIqIjhb5CS6
hXTpKF8BgpccTTsuKrMzmokA597+1aQdHuT5NbYiG81RHWfJyoZg61xZR8bG0JmE
SmZwafk1cnqcB5iF5ws7huZsE3EHfM1dTZAFNoZbo2FsNP2Y/Q5j52GRiu/zUs7z
1XkZs9QMLrrqLWdjHotASIlqWF7AxUH2Rd9JsvUSp41qTcXRF7x8FPxbwlgIYnqP
zXtaBKvVi7Pn6Upij7glw+bRilrrug3TQIB4mJiBiBj1vwtv1A+TpfB49wB1RW+N
V7WS/DxBK8N6SyyQPFc9C1V0Zdap+TO62m/fFV8tWlVwfdPYLLvhD/2q3Dul3/E8
WkE+YJM/lmbibZj7JyRYavcxqRX06MbWv5SNPWvcDBtLZRckltJES45yrZgPpfqY
uGtW9WZpgBtJu6DHweJI/QQPYfw+Yo7gyqbCfOTqoHIAtEsF8usyMadNkZMprpia
+0pgJmaCFTvTRzDLrTQnoBYxJ7Jtk2bxH/YVaI9UsaFZ0YyPESHFd3UDyWTYNOmD
C3s2VM5vanLyhMngienwWiNbOWblB4VLDUB4ngRNSAqesb6b5pNVY21PHInsMw8D
yMEY4QJ5vj9JCg9F+3wOxa90QeSDt0fCkuj4IoUTZBQH+EkLY6m1xin1u9OfSDcd
25TE22XCt9Ibxed234pZNgOy0do9XnSBrZNVRvLNORIeupOZcZaUc5w0iZ87d5IN
7mIFF7dZ6eMBNWRTlscXFJdZOaccmEjtfV8wC13fm23O8Z8ZwZLck79pg4LAT24E
gARrX0m9Upc4YVvHcn7/G+Gm6q0qlId/greUwm2Ccfj9JEh69piAWHS5ZXcLseJk
9BJFLfgEAL5dNZlPx9XmJwLDVdOZgRAPdo2Hy7L0ZnirThSD7ahlG9PBect+udx7
Ad1TSmNg1SW/ntIF/6zfIHeTk48KI+q9BadmP9QbDOCm00GHzvdeeoi6/XOYTtJI
NqupBOBss1LpcyJeTbKqa+518SphdtUEoY+X1Lcfy/8vtMdO2WP9K23oWg5sdj5s
sV1VbhLiUK+CBYtbitY3Kh9Hx+PGP1uUnBGK2BJtWK74E6gHcVy+g+T+9bDJDaFa
+FoS+Min1B2JWXgCJ4seSBhybBaJaioarEx1WDEAZcryo0CYUO1lEktdH10AGsmD
ifBbGUqTz1c5u/ibGX+VrrXu6NyICul77pZ9tbODis32GnDQH8FjLwHs18+kr7la
YcloTjAd+ZSocBWnDHT9uVrr2w8xwrrj7AjrroGKipgtlMLCO+WuxrZUusxHtJp2
PLOTxt+DTBoVmWLJehTesbuxBWI3LHUq/+QwKVboqkTbzc7Gvr/zvLYObnV3KqpX
7c87YOlny1qO70OwSR95Xj/S7fLZgwSjyQyEsyl7ca3WOwe8/5tkemGnEsjBVawI
2SLdvQYxsg3nwTaLUXZE4+Th1zgSiNiX6uQ7TZSJFZFeDoZtsMq7sYDJJM34pf6a
TSHu6bUG66sH041fdbQQed3kyJ0TQlWl349gp3klEjJ0eGPk6ZoA7GR4NSsburei
My40Mu/hIpNtP0rQ6MKGb0XXRsI5XMgBvMGfLFONnnfqUk5Hj7BIJ/N9L11GnYuG
1IdRG53goH9o+kGBqowsrXr0oPCbqrLppQaYVIYj3JqnH3zlQPMtzKlisUxK8y61
VyeArOIeKusjAEohex25NfRJIwGgvetmsVt7L/BuaQgMrp+EI61cE8qVDfWoPO6e
p2yUbKiAvZ0NJ/3k1w/gzCppQWLG6DYSCjo1AKAnhk4OkhdwkmWiBsQVZrN/+SWf
JE/0/ScaHaPaB7GOf+Lcz6XFIO+y6G/IlAc54Izp2DXFFozzeCECuPCPgnXEOkqB
vcnb3yLCnDxT+F/WfBGpA/2nozO9Ijd3IWo2/ONTqfc3z7NY7Q+dlx9Soovblawh
Xlfb+Gxj2zhF6L77KQn/SfcO2uS9jbYvPkIMMO93KW75qEZsnYOMMuUHor8PslaF
DEojHNaUIr8Q1MsBxmtIfKdYvgxtcY/r/Cy44wHqn2xE0sdmW4AQOXJBDxUIT3SV
C7n3lT2wFEGv3kPAg4ud7LGBdEhCnDqYwEPovyionoK8tdHoG5bvv0H8BWF6hBzU
dsmiuSJZe/ES9bdsbHHtl8IMECr/rt5uzifESX5+vFXuc0Y5HU7GjI4Oileg0ZpO
agBOGRPyTMcFPYjrhexayZDB4Hw+MaXCF3jxP21tdRDL5fiN29BD1kC7REck2SbQ
qf8/O/CdbhW51U5xGtMhiEMj/8Y8FS44qIWxSHexV8kwPKHS7qnKr6lFACJeagtW
xrRN/h/GkEgDwzTV94eSRvmL0fuVN03Nv0HQVNuw+TsqkRO5YvNkNyfDYHZJfifI
wL0hS6lQvZM7qUyXj96tZ464VtfoBxvPkBZRWJuarWEXT9esFaU1N3i+SNo2aCdY
OKkEsbiyBK9LE3nFwcpce4BbUpDalgcUTLTQzS2W+wAfs4FSfmh19Ef3pm1LqUOp
IC1JXdzLHm5z2jrntVYtHzo77KbeNU5ziQOphqy3YcmLL2rWcg9ofyhia/9oOGCB
rhxwhj0LQEjN0cRtpGD1Op7YOoCtpGjRqfnXAW4u6mQB4RezOSQ8/U7K7J3dvzP7
PThUiUU/QOjZERuAY2L8g3oLlu7remj18sR03lpTYt2UynN8bJgVATocQOWOBTDX
8qaroc7LcucH6+HtFMf8G+r8nsk7QhfVpOJhXuYx5Fm74/c0mxNOf8Zsx7lg1nqT
DVU63E8BMzcQzuRKY0WpVQ==
--pragma protect end_data_block
--pragma protect digest_block
agWM9BmVYN6HATfsSoErm+W86Bk=
--pragma protect end_digest_block
--pragma protect end_protected
