// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
//pragma protect begin_protected
//pragma protect key_keyowner=Cadence Design Systems.
//pragma protect key_keyname=CDS_KEY
//pragma protect key_method=RC5
//pragma protect key_block
khDwnwqAoepTTFB9kN9Mx3GF9Sp76alGQ0XGch19G2bPy6m7AaZxShW4+FjYdZtG
OyP2oTpkFpu9b/++szI2/F3xYWS9czqjLZK/EWdnvbb5lY4U2FLCFLSoPv+/7iwM
Q4BLPsbYh53EQed7DYYLFe+2mpYJVwsZy3WqI4bn0v+7IlZ5Usp1RA==
//pragma protect end_key_block
//pragma protect digest_block
777vBLM68sMnVKN5MOCWa/6OH5w=
//pragma protect end_digest_block
//pragma protect data_block
oYoVjF0MlNB4t4pc/b+1468K2Sh7Y/cv2mOBPoVXGAzmESh5n8bIkjzhCuijJYln
+LGzbfzwtWcUUeLGUH8RdhbY/jeBW0Ijna39bf5CXCdTewYpwedyG1ee0x2C5Zy7
b+mFwlsSuwkF19sKj9GUReG95NwEDwjbkNcQ9ttWigzhl4dmYzrFRK69ReVPJ1Du
FuCvI37x2VSX1WWEMABS/vY0nX1d/p1oDEmBUfKS4TXo2r/VeG/HwMhpA16XeYw0
vyjhJ7zw0bjM1lEKG+0fXq4yBAmQOZIxTZc9Nfkcnf10SAqju/cqaRJQuHSopNXD
vMn/CnDTn/kGRT49DQkWHbn8QrhGmJx2ULlFZLDaG6G1FVkrFuT874xCezeAZv2A
F0308w2dATvQvwlnxqVB0T5KEYvOqMUnSZHW+7cpRNKg8HRRg8kH1Yx0QHgOZ2f4
G5plRrHpCixoE3qxaVAjOgla4AZusacPovUC2VY7FlKBQuZp3/3MjiNaim2jZ46f
ivb1LWcgLAVCzjPNwyA90zG92Kii3jLcVXkPELwsI6MWKENZYpIqddsaa55SCHiL
/p1VDNBnYSbYAjQ3F7gn/oXAV2FsfQ3Fks6ZaOeXuyLUcpUH1VPX/66+xeUSDpUG
W0Ri1u2iWsptub1bfH0/hIs2wOKejrmuNH7AYsIWVbvH+i02nb4upKvmXT8OQ12u
GnSnHo0XDN80L1gu18V9sYlc3q11hbBM4zmeuMdeYfRGA3Cu9xfoX/M7elKHOFyF
6y8vaQsAS2Y+UoUgR5VuaLFbZI3cQGHbF+QDYDUredQUQ9DF/FYR8/q+lSLYj8E/
gzYIWYBydOkjBQGzPMa3NtP5FUxtCMLFodiCBzALN61WoX9+hIL9SUT5i5iUpGZX
CdFpedZVh5K6xXbmwHjvJO8v/iJSlIRy/1STtICkmv6gNbScTmqIrKunPowvGpDJ
Yy87oQwjFvu/qlsam+onHhfhC4Z84NzGdP41ZmlHuwMtWb9C8Dkqy48k7WE+MFK6
BsJZCsUfLiRSZLbDy8i2IDrAPuJP82V4mj7v2/tb1cVAmZUWGzhzbmQ/PqgO9djq
QkMiJ4BDbAoeZqvLgOVoed2uXDQ0PW4C9/KBiwrh1xWX4wyqWhywb9T+27fIU4/z
UC93bV1C2H2LfRtkQg6XQSV+Iifj+tIjgsxC5uYFNRX9rsj0cXXjxbqbRkYnfHCw
uYZSzskPYlzqGWYAyNsY1OmS8QERNNOPU0uHr6Vi+NxKBzh3KUmNj0WezURWsaj3
yD2/pclll4dANkHvNd/SX1lEs9LbQRV07EChOy17TI8A7ptEWBV+piEj+g5icVB+
y5sb3bE6tG891I6LisQbBb9eqmUAQqNaD7VIeQl8Zgj87N82/VEC4XS04qm9buIX
JSlzARu4x1NxBhJTirGWhvdx77CBJkggUDQ/IzuDhExDpOpyaCIrZNG/6A71xLBu
yzN2VRUpiRg1Rj06yYbStt0vmuyYwBBfyBjAfJIO63VxCYIjpmQPG+qhQiLSjWVF
fg15DDBFw6DkEl0TtxYoWTah4NuauG8xUEjn8lCo3nyF6yeYgpBSYUMN17naabWE
1OCGYWtihsjJ3a6xoeb6GMEcKTxxltj08cQiQJyCnJj96+OX9QHXCgkPNBSuUvzY
gXqaQkI+jEXYYZJvIESEsg2Y1o34n1/7+9RWAEUKsIbtjduIXs5t7pfXUSxbabcP
zvT/iYoTuorRjYs71xEBKAh3xdyUiMqMAg+n1BRa+hWeNCwhFvVPYtUAeJaJ35d0
0tGrN2JxfNgwmf+95baCt0rLibIHtJzvojA9kirUgU/t6Uzlv5Ali6tL+li2jl9U
RBbsbMLZdk7F1iybdJAYc1t4BLux/jyQPRFva0VQZxXooeUDFKo9cc4Q0x4mh83p
bZk487b29B7ludAdvCfrIhLkjMPmHo7ZHxtpJAeRQ1CPsBFzOed52Te/ZVPjeGxa
6UBPhVPbcA8w7mqLNjwuHDNYHkIawRmb+5dKNsM41EK6wN7RngrueqDfy52/xjQm
+LgXCMz8TO6HXhWuChEzFINtf16Oe3O1mjSE38z7agGr+3rVN4CTRjxirKXvxass
f69w2PX72fG4uD/IL2nSAcPicZzswq33Ik2Un8NV+SPQkjWfrAM8x3PEhs23Eg1d
peXP5maHxgxf6a8OV9iVCztkUXzctTlUFo18NHfAqg7vaUtefIRhES8xoec446nw
i6ChrIlbJDKiz1vhD0wYplYpiFSfNB56pBqHa2FilSw34KFwvfwlFJUeNemMPVhl
8cT3lDdLaWN83yfdHKgnMrJiRVhix+2bGzrOMBQUiSENZWiLlxEwx3Nb9ywJVpaG
B/2qtAsojubjNbKffGhHCF2x4hXJeuNbi1Bukkl9ZYIMJg5aNxYvrk+vACPtekyh
4svQNASy02GWKhZLTk7G+0djz5JKdDCTLNeBiSCHotx9KjGcofFoVQ8I9laI3FYm
EI3um5v/b7jaI5iER66mtPQW9vlKT0MTECIeWsb23niHN9SpMIAuZX4x6ZI7ajj0
2M8MUbqKuQHXPJeIAzqK2CIzhEZutujf8bx2+47p9Fh/bg25xfeudGL8fgLI30NH
EjJ4ORxtpYyf1pZ/4+HL1kZClxtQO/iKfMe1Ti8FdFBxcmsRhsnYgTMdUWdgQdsq
5wb0DekrAvcmS53XWruWuLqe7DV+s2r2hCfY+HMtNQLgdNfPql4lb9kpDSk/IPBx
wwiZo98TVTp0XtMvKrBR69+ehYLw4dB1eBP5gqdNGxJGRd67JaUKjmM0ATyxINfR
lWYpy/enS9aRVz1prV3ocdiAQrUc+hTMXfPnWQeCtx3OEEtMw2xisu4r7wdjjWDS
TORtYKWmwt9NrCo5vBxvk51ZNJ7Sv8SNf3y/DpMmQvDOgA5U6AC8xu9VUuqgd8/E
/BY3WY35DIIuTMEcVExZ/292XJO/fzmYU0NgvlKyIR1/PbkuHiLDuIjawtyBd85Y
q0RGxu1S0L0ZQC0VblIcpZ3UOBl33GzgbvoBTV2rqv7xr99xW5zLUVrXY6PpJa07
XWh5eUMaLjQ2UKJf3kzXxtIuyNxLdBYDiNSuCZTM5MrXPztt8ArfJ/CZWO8dK8aX
TqUXCLwqv9aoV6j7wVbPjHH9nvoSzf9nPfyZu8vbRgvNDKmArKoFvPUAWGLfu4fa
s6GmZrY8GyzFHnr2DaHBQbYal4ctV4KQjdxCp4fogP0AWzUFoxX9GpJ5HrJZ09g0
a+TpXpt15KeIZysAZNCfj8xhOc9ZHKAKxppdSezZqOGFa7pzt3Y6QBIJzZ4FlhNf
RpkFtuC+s71uswYCGuYC81GaIldiTxk9Yfp2kgPiARfdbt858rJt75oqs+COfeQj
I61T5d97vX7Kk69HLkl8qvmV26oSIplExbh4QJtgUk8UkBdKWM6QzqpdX56KqhYW
TdlnJMbkbXdyi8nl8ozWFWdPQ4PD11mt/JmVhaut+WzE2WqTbNh18nljHAaoYemm
bkFQh/BvbRMlIxLn7CSjmP80OakQbJGgK0TNSsvBBHUcDpoOY07r2NtQJky10/eM
0qL7gJQevn1YAePVdz9EUkUid/09MifGv88y1lKrLZaZpftGn1eb1ivZFFgCYaRI
QmmtscJLU5WN2+gzo8rHblV+jAfnmZcYJN/xPMhls4uu2OTKj9FVjYc1t8f0lYsh
OI20NMdf0vKaQFOBAdlut7zrXnv5PPWkcKwrIxxNSbjrfPZnM1qSZ1yKiLrns6wT
uPb89rUnq6cYjZ8EozhVabk69zMw3cktvlZw1LGrW9QuAWYjE7GEf50FYyhxH9PY
G8LwFnA/RMdpL6pa59ZA7SXLGW3Ohk1KWWkRCqn9K4/LpZFWIASFMYdLBaINiZY4
s850luFsGGRHoV3dQT9KPworbhSHPRf0oWeX3gP+lSZsk9jB7THtN8EyFISrkWkH
XGZSGfRLrgTHo9IG82Pa9oHYPdLmi606moQ77bV/lHwXe/qAsBFoyQ6oKjtguzng
3OxM3npKMiJNCqYTE5zLQv7alWs93S5ee32+sRfySwajqM9RWnlCA+cSjVdSg7++
JUzPrrVFqYIZly/LSD83q2ylAylfnWdcqccvxhEnEvuhoEaYaVW4iTqTUOrr6Ikv
ttftuF7bmFMIZlA0KIcF4iBSY7ws748MPKyOjF7uy4SkkWWkyLePRQwoDeV1sPW3
0nl/aj5Ol0VJpTUCnHnawZxXGOzEDxX6+/N9wS2z/kZJnOw1BpvaOYx28bKZq8mG
ynJQSPWW/AzkmCmhih6xSjfghcS1poagS+s4N0x2Y3EvkkrOdu141tE3uAHnGqpg
mOwCwtiGcLbG9HY8exD5lT1IFQ8X9R7MbgDm356pvcmEbztawvLHUURIKRUU3FI3
GMd/BAqkP3jvmYAOySs+MrpClNyOffsozW532HbzjV7OtrcGfHXTc6H9PzoG1BYS
ntEDUABMchGS281D7KdnKGs1cmtLr/EJUI8UYo4xJQLQNdYArj4xRgp41EcBNNd4
dWLjf8SHgHgIW8jXDvaEsvAG4JglB/pL/d1JWJ5AnyoTJlJAYDeC73nrwIyRzHRT
b3klnNBbE3wAUKT14t8uHuSCyfCnj2QG5VSooc6IpuD7fCkktaMhDLL0oDvIypsY
UPjFTh4OvLRGv+Jy9Txnc3wvlb67yFXipxE6Olz4iUQezKWMHg3DZyRMxaYW0lpv
l3Un/F/p5Vp3gGKW5E+4e4ANYNz58XR9wYokpQaFsUWrnC0n8+jN3+N9AXfdX96A
B03awZPYc0dUJi2olnNBeWnRblUp9AWKIq2mkRaKwg37MD5PVWPQj7tY1wECl3jU
2ote5MonPtkuB2Vnc8WtLhTPajyieyk1fa3m9WZvCUbt3L9CUkrkSfb4U+9jrAN2
PKOifoff28qOSU7ai5/rVCfBB+kWfKMkKWa4c5/HorJ228NkgdQD2ZqcLe+haDnc
mN7+rsPWnvDRZ6FotJeY8ixgNS6GFyfr8uQDH8cGXOEaSfuDEy7Yn3GYxBNVgspn
RPosiGLe7F8TQG2hABb9FoHZnjbG6blb+CO1LnbGurr06wUiXPO8FzoCVXkhMFUu
eWeNOkrBqcUTJasHF/J58wn8HF/BgWt9t/JU8U3gWc46lnpFoK+hskCk7ptvs3gw
2DoorhAZsVqfg+KdxYioIQHjsvME6ks3b9/XK/5i5lyoRUdmjX484hZ9BvbciSek
QAUuMKoH522IP+0KAonG6mbqvqpjonIyo7y/Z2qdAI96s4w1PfEXomosDB/R66G4
epWjTfAxDaHkgsFoCZqAVahPy9wVnl4J1CB5ZTX/KP5M0NrYzCwg/eJQI3KCK/fl
qo5ZbCfGGx1tztzKanBEuySa25PI2c/w1ayJzzhEMWEe2EKgY1/dNvt/MaNyxOYY
/UmIcfCtozAZv+mSB7a1jmAR0ao2ofMpnc3xtfbTNPruWWz5hArs0m6pnzCTR88M
AxjqkcU0y9/si5UMYw9qbliMk2qVdi6Dp6JA8QtgiiESBnfa3VR+3uApZ1f+fZBA
SoxymG8aoJilIuhAcWEsgM2LWL8UWAuAF5jtuFOp4OfhEYDqXZifK9JSP9mipW88
ee8ieZkX+QrKHEr1L+2jVo4O+n/CERqujy2cirUs4fNAd4sYbqQPFUMW6vnTN3Rx
J1TPE3Qlq+zycEYoG1ttxJbuKYLA35wVuKXizr/qqBWfbRZljr8nXFRaeRxcp+to
y8oszbaX6g4H+rdEVialPEXJDnJTp/cvVnW5b+D0d+RfhdGhHdzti3hAra74Mw0y
UQ7XBmMxMwsTHcePHTq4mMDKvqJIPzMnO3WLzFep5PzxIMQJHSwjnMAvESfYtwnA
z12PGiqmRTNZECXleXtnTTaBMP4Fdv7gWpnXXSeNq3EFcWjkK8n6xkwZoNxhUuca
K4fxahQffVYOK/xRxd4nT6GA+rceRxiuSTg/Iay1npsdkwBuBqPrNlFWVBtMTxWb
col+1etZtEYIpmnj2Qs0d/Dg34kPyKxKh37XhUrgPxnTLi9owgCrQPly6gGkwu+h
nbSn+vaBFroligKJJqMVBk+6OeewEUAvnZVqdqx2IMOEcv5bO+MMyj7Uko68QW/Q
u95qSsDTsjejSExkMQvIZqa827lzTkj58WQxtGb4NR18QVxOjKCE2HMpxPELqi1D
Kz9xTntDJASeAxK7qeH6XTSO2rzxuMQoGqoUeXCV56Ga/w2EJVY4hL8uf4+aEI4F
XH116Gr5xZIMGBD03kT2frFefXpsnXZ+OaQuqeytaUDAC3qtBjl8gjdV5/2syeS3
xijKSYvh9DyvE6axH25mKM+VklabowanmZHesuoRtMUF6IvL9Q5il5yLSeOmQ1Oz
QkriVXKPHGMqa67Swa2nwPfwHB2meO8fr05IK5grYuTVaR0eFtPwjITR2y6P+Arc
WxIb5aZKDUVVpPiwBvrmaO0K/tkPco/C1G/nQGQ+DkCIXXpfcWnFow6Lpz12lYGf
4Kht1Uyw8yq+f58gMfXX9hQEhyQlN8DxxdLNJs/jTZPhJtCTHokfkyVJwfbHc6Dp
sUI/HgwGD3LYCdXQpl4+17wPmBCeUKTZL9xiU37J7+zobh2BZDGuPL1KD6PDXsUn
PHNK3bgh20IPZOaiY5eSWGURE9V0S7smQCgppxz87vl/TGLDYMh2Fti2fH8inU1r
yQxnGn+1KWrr9q36Yi2PWX9oxhRxX66ZY7aQehEM9FdVJUzOaFCrG47Tg+gGwp5B
HpGd0kaJkV5f94AfmtntsLjs6ZxPbuSjQnIUBMBv4J3dO1ta48x7YNdQMAS959NZ
2ozBRFcIKRQVajTkfZV+jtIV54wqf54cR2YHfQG5Y+9bdDuLbZLOPTbS2s7+Qx9h
a5Jbb3LfHjJkm352KFufBe2v7jAP07xwYZZ1vkh2MFJohypWAbuXenkzMdbLRZfu
1GfhtFFYYjLK9nty4hCBNRrA4n3u/7DhsDATTjK/9paoF7Lg4CO3oXudSLtuyZ3H
TOBFBo9LwRRB77HWzRLtrZS5UtA1kFe7FVqQi7yu4Q/CRykSKEA/yUUcrXCHQtgA
qH34YTNG1eJs5TLmbNOEyLWzFfosqY/nwTbhdofa0p6WEsagUnA+TzBGL59DjAeE
9MecNKzhqW/aoRF1DyYRRLFETihTJ6YryjVecHn8QMPd7u9S3xo3HXLQ/yWFcTcm
O7CvY/fm5O7g1+xVWf+EVI/EwZvTLP6NXIa0tKv8K8FVU5MW98bWBl/iSPhDq/Ab
pYBIR3+WWtQM/+Ty6y3Kyjte1c9+nwtQYxqn3YBzTTVS1DJ8n12TM9J4L4HyUY3H
pkBDZDrs9s37GYrkD0jVdW2MiSxcksB5RALP/gzRn7V+5DyH/lIPSjTA6sfy4aCU
zNfXzPtSB1qBL1JuNRyvUZJzKzbc+OffOFiDl6+6FrG8MJxLFhVt2MFLBp18wwY6
3iAgbt9SDqUo45ppRCKaW47Ge6CELxSdjg3pzpNdSSMHB+YrsCfZLEnpsGWdotpM
Mye+sEzT6VxB+XVIRy+cF0fFFtMYRi4jY7MKeZWBxgPGykkL7D2y+DzkHR5HBDUA
tzry1KPQGFUb08az+6nxHzxvlJRCDVTOmg7jwuhB9XA8sGHT40zUgbzS0XRGa/Y0
l+fnH0wU7z8n7oP51DEZwbWWeZg6RwFoz92dzgv/1/o0pmsM6IUz/3CGFzZDrmew
O8BRa7Weq3yOHzkCWiZMI28k0xGze7uRn2sic/8UpngzJDZW37zQS+Z8VPvX67i9
bp5i1ZfOSQ1w0sLghws8uP+KPJ/EiWQT0TYsCv2JAxJFJLGzSpKeuh40J9+jPnPh
WhCWR+bzzBx2BQ0IdpH71koSA/ezOE/JQQnvk2lZq1aJpmvGyZVNZF1F2zyC5pKg
DV7g2YlFKdN5eb/2Oj/hMUZ8i2UHjpChzFmhUaj1/Fh1EJjB9ZkZMqfOfemGxAnl
3lEQ57C421aKskFmW8CcXCUKwlT9a4b7wfV1k7XGFArc03JhBOKWJpk3CQR2exKS
7LWIQSVlAZmztXDrJKDQAoDLQftORlLTQBodepGjxOjwSR+zuIih8IMoJ+VZitLM
gkXxSwwK99lGNmAkRP2p4LyZMsJrrupE+LzPDjLR7dcra6bqaOsU/4Ha9jcCFFUE
eXtLlIBe9kbGNQzQvG4pfaPkRC6QwmHKdotMwcFYUSiXGyvgEHMS11ticttKHAbN
8S0QYA+9MctQ/CpFbY6ZO9pXkkITHKQMSz6EcS7CrF2JVUqcEw8Gd5eU8dUGrqrS
ncEdHZ6vaGjOnyhpfFIhsr/htYg04q2cdD/Qoe0X+Vg6ZqGsuHMVfjXihJcodaPJ
Ovq+i0lvshgKvueD85gcIR4iekgTIOXP1NYTsMdS0QS4SiJ0dKl/84Z/bw9dE7rw
ApThKfPS7ga1b4OKsrO7xiIzljqqguSnlWjskRwklFCkkK1qOalxKt2586eEWhdK
sloD0wJYuTw1orebzQe5Ni4bnyQhty909AReJs9OvKWPpz4aYsP/wkEMXYKBJ6Hv
54zgmax0qRjN53dOtoXT8bHhqbHPPIYr45t24NxaRvg5kpwlYB17H5wEkeD/324p
GK2C3O56ntlcO+DtVhmpUcd7EFSD6eW/U1Lmai0FPifkqpqGcnDRJVpX9a1qXYTN
s9DZwa84eNhUD/mGxMCuUu4iDy1BMRDvb6WXFfAV3a/k0nDJS8RaB2dcZueXfnPY
V2czuGDcjyn7b94qc7ZvuiQ88VfmLtuHIF0RUvwNnVYWN/v2KOy3dwIXmN8DvYza
qFJ7YUocoMPrNVhLOQ78wXvjrcNCJ+OgIL3Lc4H/Nn0/v+3ojQFpJgRz93ZXzSZQ
kIzM21qLQAbxE5KnHSyO6zHqaGlYCODnVqxTcXYXII9wwg7Rv1kHyJOAviSs6hq5
3TjoZrNqgCPQz6Pr1t08nqDL6YufdvPXZGFYO15wtSfCPLeiaHCl+jTnXHFdonVr
qIU+9XvTvhCSy86jEgh25tA2vr8vbf0pWjMfUJW6J7frYodE8P5X/aYnF2OxqNpd
/lfemaKnElZYpHc3f0RLmSCdHDZGzoKhyTSAaTuXtrf9JvbjK+8yJeZ4itoBtScr
pvfKoZu6qXOPToMOKDR9sqCeLE9fYD/v/qMGxQy0+gaaGB368Cgc+vRkVFBOOia2
h2azCFIx0IhCg+MjmLFan0a46gAZq4RIq5EqspV4nXRoQrkD7feTrYD3G98BbHO+
xlPF/2EFlevs3olzPHcZqonHR4Zxcj2813ikJXw3WUJNrkqjrjyX6afNdPdgbJJv
VlSnIWp9EWRagKLFIUw9O397j/o6eUDyL+QyhqsJ56WofnHX44YpmfrNG8NywCbM
P8UIP7RyneCWQG5BjFIsxuN6Fc6JT1sE7ASF2cJ9udeFlC39aa1DAp/ZOJsyUqox
q1gbAv9I04F2CK/Ju6hr9Y+ZoC9VOIWkcTfw1ULShDi+BPPWndtV1wrBsK/u01wj
uVudvcQKp5esXja5x4pTbkTdy6PfbbeAzShmYC9OMkfVmJpDwoW4Idsrp0AK7ELq
NH0AiiQddAbYgba08EgwRHesxoUHQ7oirAfACKfB1R8bgJ8xhu1Deu05y7EeOx/u
OjwYAPuijPfC2CCOBnHNRdeS7Q1Rc0XoU2YMAPu8/HXoB//fJ86bS0dRP3DJ4sLr
QwZ8J3E4jObWNjN3FzkII8PARoOZ47xUkJsT02KNuEbZDRhqifbSZE1RWvbMouj+
CL3IFha25w5B01yF2EJA19Y8hfEI0uaXUd/u4sYD2hwUZipRbQL50zu+4lsVBwUl
7uPl2klXG6XQ3XWKbZJDugWvChK5MEAW9IIjCDCk4VOSCW06bbox+eXYbwMLzgI5
Hh7olNW7/bWaF0iO1HzoIoeGoIdgUOHSpQAL7FXIzRidZUN4ADFQri6Q9upiglqy
A3+aHo3AEM/bbaXtgdclWh7nyyiV18U+X+eIdEEOLkQeLqJxKEj+Nvc2eEnCl0Fg
94NOiDdeOLLY5nQHwu345E73iSVgyFPITZt5Sj8lWSQdTHhPdXEZSkXUoRX1e5bG
gNQ82RiEhaoaWxiOeD8tmluDUyIDUdE1ElfeWz2O/49aZEpvOpdzV2y8GyX9ZGkr
19Yv7EVeNANFNXEC6MBhNwTcYum+hW4Y2Otrq8Ncutco10NJnJGE3mKtPNYc3FpW
XcSxPM1T9BHwwo2wwgsry6oLD/BIZ7QSIvQ5fu1Y/qNIcSHGTkk2tMuI99ql/GcF
d0frNhewNcUPeuCi4OLvYu0DkfA6RXI1Smc+ku/xXKt+YfhgbAjF0XUpHQuj2gxF
p2/y/qNxcXqImdweIcOqmZnsv5ATJxbmIw9IgloOyxSGWjctu+fmPJXvqNol9ceA
3NeGPIb1Wqlze4r0bSHE8C7QkkowStj2pLBaCKEb2jvU5hYXx+SpGNt8KRo7QLUK
AyFR2VuCb3L97TNEBCvTgtnM5euZUk7Y5CC2t4Y3MzH0wiqgrGPbhP6i95itR2tN
St1KhEInkzdX3A4GeWUt+7FDsptbuumyOlg6l3ifaVBd/ruaXJ6q+9fZ/Opi73rF
H7jhgwgQMDgabm7xRoTl9P0AMrvCWVuGqvJ98BB9ICQAQX2PM8+N5Ef987gHhwdl
K0sPAf7DqOeZ/qG9QcHuYlMpsLlosEiUnyBwjoZpRWvvOKqRfVQpPS2dzBaRh23a
dL7swkMpwTLcygTtGPuPpF7PcmA/3WosdbIxLeG6+ONCv1p2S0RYF3qb+opKMXdG
+BRMZOcGAthjFVWxK6TooI7TNsiqCPeW9mmYBPystunJo7dHVtSjszx24duJmz2Z
Kz9DpJiyPM/oO2MR12sxNPO/bhk98jo5p0JVjytw/Y2vV0eGEce3K9okEJl+cQFi
UgSGbLoWjzo6Utd8tln1Z4imQJEtCou1aeTyl0j6Gwgtjqx2TEX0i8yjtpRjod2m
EGYYid3elpB7pEn/vMAjhw5IKsGfnf3Aa7peCqG72nQdikcxRVcrmq/b0IB6UWMi
wW1Pvy7An1GwKQK/QUwuvpErFImKxRtZFWZSYwCFsQUrGOw0DuwmGrcchrXheX1s
mGHNsxeE2vDlE7caCoy/ww4flOf1gU+iUFLNSMhhi1ACfrT+DSFS4voYtH5837xW
Xv5Sc8zv0aYeHKK0Yo4WfdQyS4Aca1tSK3CkBw+y7OvjAmz/8dpKnHNw+TgchRop
+HkPkDuZFobIDB7WimKeNdZX/YdsMmUIINz2U5w1tMJuYGYdsAOWTgrPfIlcdeoJ
F9w8Z6AANvvS1njmMdoBb8qV+V01NmbB+PjzjZvj4syA6ORnIDPGVDLWAKDJadKv
Bh5X73vABGuRKHX74lyKENsykpTnkKM7KfZFgL5zaGa+8TaJxFBOQ1vq+5cBY0wT
gXMThbhI8fMBtfawG8+tr2sijlr7QN9ctUblagH2zWg7QmYkISBkCK7EGGpUiXtk
wqig+mtSFZ47Ehdo8RgC/1zGhwyzwlqPlFNS+mSx7FqzO5lVqNmaceZ8xNEY4x+e
n3ou5PrBs5acxJ7DKjexPXgX6QNcf1xiSgQjYTEVELBswpMyKwV6YouEcSRK0UR/
Nar0mxhH9+RLdeEPWSDIvGMiZxcL4Pm8/RUm6e8luLdyzvxIiLO0K7mJHCiMdJjF
Rb9wp6dV7sl6glFVmUcFxL+45CtQHnX2Ir2hEtpRMUPyrPqKNEGXMEGbzAMyjIte
amx41TGIqoLlpcPyWsYtS7tmGxdJqsin/6Dvyl5XEuiYlfpq7Kb7iIWdnGODO2GN
rgAVMqZ/ipql5oblgNtBAlXpeVljfQ6T9jrS1ww62Htqe/ItJcZX15HzL/uKUD6I
zZJEcBUF1XhgU5faDOmTEnx81SgxGnPUijX8+Yp/Pu4NErHTSQF0a98c8TiF1y8Y
lnIg49w5TJNdS7kUELqvTXq+DuCNlTSNS53PXn1r9q3Uhb24SWL8IFaQQcfXfrT8
mwH4tGSI4VzWgedbJVF7ARqqAwDQfRRbmlj2BSckhsxUV3Hw8xMJXqnTxkz/2xRh
dvBKHnYoOc3JgC3EQuh6MshIx3ialEztJBj1XIgFG9f72iOtgFgODPvD1Qva2lNp
t78zjdmUau9tT5lSmySeF13maUXpdsfjBMU0ZyUvCQe2zIsU2m7rIzc6rKCYZ8wm
ftit/bOjBvdTjPQmHMCZDyMINGEFAmWZSOht9hTm64ns5CsDJxKn0ubfYcKl00E8
nAdZw1t3AHD3mBf9rcyDTe/tG0MBVOGV6kDEbYK3KBUKxKUd/dmheyr5LvQ4IhVm
AHwRHHzapP5hxI7/3+lRGwPvexLcW/h6fPLvGhm/P6U+xJzjANrpDbmks2rYtFVX
ZEGdPLbo+TvjHb2u80t2NJ8uRh7IEkeo7cvlN73/9Bdxiuo7gs7ObYxcAZPuMwNh
+OfEZcfWqZ3O6tcTQYb0h4ir7mF+4+uxiMp/Y7jA6qVDMMLPJ9z4t2u12AHqh8aP
yvrbEqjRcZmuixxheCEuNAhtpuI7Z0k4rDw3HLFyndI+YXV5v0jo9h3q1JJR7txr
reXyxJY84PwQ0pAF0z1oX58eL2NcluaEjy6uB6hK3a3MTMWrQe9Hh5wrAzsJ0+l6
k0qLRXYA+sxj5RpaYK+Iy5T8+gk/YmK7vYDdcQYqOk4xd7MYARHjnyHJrQjfl5j8
+N/S4/mUwyaZ0xdytWdiHyIvbdw/l7L7I/npv19TP3fOMr/Nw1nuISxNpX1P7eSK
gWPwQ6citamooKciFal4gmbZejwtZR4a4enPs0CoWZj2RSg85i4ujBIp3GxQT8bu
ZSt2Q5SDpGrHPqsCWojGjD5FkjacTdC4FsbnALgkMIBZUgaSplq5avW31BGfE4Ux
WAnWLNWwFciwcbBlpnUmG50qCxQuMlAanWeAAQxOLIFAx/xFmRdkECZ3gf8XjUEr
fRLTdeJhy2NJpmNDwF2GRnHp4Htl60clz1qLZ3j574lUGpkvTb9op1TG/gIUdE3K
62brBIJerNV/M0++jA5Prp+MrlCv7gQ0Y8BLKWRxdePN8GWyT9U8wsCkq9VcPfzE
4IBfO0MDUbogMJ9GFqIjCIDffq86w81/XJj4yMi4/dQ5jE1UoM1FppWZ9fpsni2z
xukATNrpUYM6M2wLuss0+xsGToSzYxX58yXpU21C0ifrzsXyZMhz3/3Hi4V+IoaD
lrMUk1t51cfigBi7iZWyIkJ3qgiwrBc/+mR7kzOaG5aGibS0gzR4Dz7lu8+JeKmn
xOH9RL6aNJJuYIBsvZ8yPe7kbIBhxYepjiOJFHaxOuSlq0iSktV0T/xhT9EH0eqB
MAFxVJOpywm3TFCU+qtdlD5JDoeJO1dz1LAjxq2cEqVDEir0+LiHVW8RMF4Dd0x7
7ChdJvZLfVSp6NHkj2txnVfkkjBJ/hQKQd/sVK8GrGwolu2U8i5gt0PW54mt62Sx
cqqta+yUf+sw8TcTX8SJGF2QdX/i9Beb1UsfL0ocgqnyaJuSlhGEQh4TkKwem7Ei
FK6jeZSW7zsLDpcVnBYSJU1EJy1yuGqKbmnpeMDAJH6hh7jExegxvYj6cCNAXxPW
PZJZXCKWzWVgaz3iFJZrM4rXHURtaFGgeBBIPI2fFi5C4K1+RC4HilBJCf9Tw5nn
JCNlTs/6S16GH8ZGeG0kbUtYo92to5ai7G8YQpuNGSzLeQHPBpUEatdkV7X5R7J3
t0QPvL3bnR896eVpcHTbYe8Akot5a0PiAL+XrBtQRjxa1ZIz9/Z3gidHyUPK4C+p
EB5yA2ApJALZ2d00Dy7lYbi0pud57SNLUq5okW2ranwoglWLOPtahc30dHyC7Eh1
WiE6IbG6km99pOzqCQxwqHFkizGqNAqERJD2sE8KOwOiVV6jmWVVHMqSPWovtuby
tSJ1DNk2XwIn7YgI5CNl7bcb1VqI3J1mciq8EJLH4Zqgw6ImIw+LNoq/hpHhlxqj
nhdnc/Hbr3QpyVNzMar8M4+D01bVXgT9tPcywK2nDHcOsBkVXe6y5Kg796YNT4ic
rYgMGd21Y1IOr1j2+hNqL5UCcyNEq+RdCMDTSRg2j91lcbsH8XhNT7yDtzzf0iLK
ySsiVXRVSEbMDCeyIVcIHQ==
//pragma protect end_data_block
//pragma protect digest_block
ZTyIMLRcHtX9JUj2w7XRFTWP+z8=
//pragma protect end_digest_block
//pragma protect end_protected
