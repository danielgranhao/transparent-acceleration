-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
I518t4Jlzb+Vt1i2tdPzQhr/A95/GMbibCmR/v+5VwwDcqpiJng5HEhewDOYqbF+
NLZrCqfH09RtC6jknDkLvwcbEfoOcZ5AMgmqwBMGmL9M25zwUWK1u7kLHRp9u7FA
KUgHBBLR8dO6y6T/QxKrEQOIRbKClW00mSz/hQJ8Qag=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 42976)
`protect data_block
Qe+y490xSZ74goFpcObLo6qxgzPxuPFSVFvIX1lhzS72yQQHLiVLmBonfleCis87
tAJROzQBTO1cTLF9YXuwxZEHVwF+5PhnhjLFeqqoxUuOwr9SKI3i/NKHg27Oa6le
+JzgG2aLczaoiSXWIEXSQAosRrp4k9//WYAxs7Z53hmGkSV+bAU3Y0eCx3OicarX
BNsqgUMrKIJCFfuAlOCCVMlo1o5mgpMRGg5I/uVdwiKMpPwi8is0wI8XoiFcc2sJ
rGQtKJo5+7jL1ypG1xsloiDs1l0tt5W8jpmqZfXeO/6U/VmWNIJrtu89VdM6clHx
wO8Lu9k9HZSJwXb0nkQs2pbEeqqFAOpPa+FIYyqiVACve3agd+MI6XvNNcJ0Vx0r
JDpiTXRWTEALMjOv3AzQvJVZsEm9qzhudXNmiH9RVVYleY+eCa89gxLkQZTLpOGX
KDd0frH3tB7IKE9opOcVesmuBZTqeHspQsE15+fe20qR26v6pD75i/4f/H1Z1uNu
Cmzzd7/L5X4nlZs87XyTHnIDFHq9/xm726VwsM+Pij5OhwKXUrHxmSPpA9Dz9CLq
fjv1afgi9U9P+220r44lOWFUJS8O2R8EbG4y4O4rLGf4UdwHsGgIYTdrFB3PWaao
qzTOm/wKxIU0x7GX0lFskRgpdegMGftp5Avok1uKjdWcqBbBtj2cq7L/oPp3oI7L
BawS633/KrJxvc6zn2HuqIdEYg6GJfpyFQ9KPdPiz+Evjq1GeoSsp7a/m/TvFCWQ
Ms6Xu/vkrB7x9pn0yapx7/podVtAS4q0Usoxva63W5tIF3cgCsyHbNusY9pnUCk1
f+DdzdDh1Fh+fVZRj4WLSXYWCDkPnprPpyMsSOCQgcYn7s4uVwXnrIXDRExxCgKJ
H56qDHaccYt4jh1YvJR+SfZlaXTcY5ABZyRpJTAzIHybK5Cp1i+rWU4jSzOWuSrN
/KwqYfjvA46TyaGdAOe028IRu28qPztT81ctt7M9hGtCwnUPbY7s3m3glq96udAE
xEt6BLorgEb6OqgO+xy4Iqo+JcsZEMzkkDA/j5lrtrS92JqrttLeGgGI2pEnP5f9
qotJAWC6nswBbdn1M6flb36Z5yAPKxs/sEpNImCsyrBVRJinrMmJjvA4VYRx9OhR
U4w62WJxh4mAeXWHno0Zjc6vSOSTFTQTL2Yr+Q3pMBquzunVL5HgPoPiaHy1cSR3
3AcVXoKicVHDGCrmMTgPjmKP0yurhQ6Wx2Jo3+yl38fG6JjToJvKGUl8eT5/h1ff
/KieV4TyX9tuW2xZzIvGzhc+jTIl/TpXnA/1IRDSpJIjMcwh75Jj4fDmXtQKKZKH
rhLXguQfD+XGj4UvIF76YJGpdbvmBbmoUKPen0jZM/o5YSy9zbES4omUQEJar9jG
CWCU98em3HLNZiViWCPXV1UhbEI8ACHIsO63MxC0T68PqmRA04w4EtpJUu9zK46J
GX01oMOkhNdtglwM+cSLLTyQxBRokUUuart1APCvUqodW8JhC/WdxfFotSRjis10
m31qRP0U01Rw+qY5RoLVt5XEz5oRCm6OY8ZaiD7/fSQneWeY1jeKVlZ1N8ghK1Nh
iFltfwZtl/T25mVybua/jKB0VYptc+HaFCBRxyY1SOpvjNFQycoto8x7t7OlmBhm
baNpMXoxqkj39GUQsTv0K1+L674ZxzFnpyMNONQEmb3EuyMP664/puCXbycUrHhM
OuzZMUBKt/DlmH/mM455bZceHQPHQhrxe51nu3B6/4pvpB8rQH6/RnMWOrvWIjJc
6p4sQN/HQfKeJQelaxAkYXc5Ws7T6mEoGtPYpNOpQ/iGy19+GeIQt3Oocnz8toy5
i/J84enchM3wnRbt0ByRX7reMgfGndsRzQ28L8D+pdQwFKXujS9+hOzCXKch4bDt
0LDMNO9Uq6T8+JL3PEDdNS1HE5LUFDZysFPPYiE6DxGDsjVW8v8LewWCQbrAClJr
QtQiBSjysHkkgRyb82VnlQXVkA37fqNW3qvolFCZn/GkhrVqlRY2i6FDqP8FWqXO
wmA4hA1vd7aSgJmqW63O53IgRKMPEFf07uzyx4LpsB7D5aLnGxnTp6aAa0oIEoSA
Bkuh7W2zYbY7NhYtkJt7CgSuokAZguykzact81Url/5Mlsx5vd4DcWtxyqijnEo5
MuHlZqK5d/16iGoDbE7Z7zXGdqtDUlKEQv5hF/mXYf4Ngmm/ToIy4nr4C35DbhOT
oXSbjYC4KuBTJG4rE9RXEqG8Kfntu7369x4KdofhGtLO6um49gjcCwcNV3zkKiwR
lugJB1K0jwH3rjqsj7Y7NRslWJk3FRYdQzYwjpM91y9Ao36UeKuw6tSCN9eT40oY
mD8WMvV3yN1w6orCNGP/Z0n06cGQuCurQ/rkjw5BcuSTWmGELGYumv89+T+1nF4o
RJdOkomykxF9W3ATJRGC0ZxnOX1DDC++cEVZryK6PmcT+eogxC/rzj+MleSZxvBF
hhDkaXbjM8ppndd14ifhlzulAVCAwjHrAomCktIeAgxYvOW9JeZ7pA9Sd7bsjoYR
3/+bd7F3jE0MnN/gATvodHPoKgQw6tmLQ+2WyvosUGRpwTOUl+509PilifsMhyof
OJcdczIw3NN/BedC84UWrG1T1VZmsFXV+p8nyVDaWHjIxLie+D6EQDw6dQNUXcLk
o0f85aodYTCusz4O9fDhOiNGy0zsQ1U3CqkDY7XkRuukOqgP4vXbP+1vg2ktgQVE
1jSlWSyXad737UdO31WXMVmg+WP9Mz4/eVr51G7B8gNoRXnd/PztatP2Dsz2RHN8
lqbgOZqx9rHWYHIIqxK4D9X71IlcZBSEtfy7rVuizSUZxkRZGn/kfqWov0Q1zDkO
zEp7+eTYRQqq6aCxwjAXlCgcPpR9FG6ZSCjP3v55u+8ghGYCU63PvSZUxepLdkEJ
RFhphDkLgjmj2FUHjY4TEpSHY9M5XZzfylZAw2GVs1aVAt7BhyE76Tg9Jiv3HGuI
GI4TqC+y0DC5xdPiBpm9mjln3h0O7i7GwmWEwc4URUoznbmGlAQ3jdID7Y9LAgzV
wIsgrLqn9y2o9BszSyv1MDNERzmFQ/mtbflQvAiXWFj6zfeoMsu7A6bI1qp9ymWb
9s/HuxtiYfhmaBJja1vybx9BUYyA1naeIl5Hny4AjQNPRjYfBHi/jzn7Jok8XyZ9
eRsZoIB1zF5BVRySCpo9SDlGaXrzwoA5plVQBodHGrkbGT3FCWmuAho6jAHqWhJC
BRhYPFWA4WEB5Bo9xC3jrhmFyInY45InjV6Ob7H9gOqJUSxm6GGa5iEg1hkxqFgW
bz/9hgC8lqTcdspegz0L+RupBv5fFl+TOOL9kG6UFWidP7b4So4ODdxFfxnAyu30
wkPY0T5wQgEklddHI5U7sVixm/enyo0lyoeAuj+N/s0Q0K3LbESRWEJKpq/Oc3kl
5O9iCLqjNd+ZXIU7Setfg8iTX4e7J6lEIbkABPhN6HKvvPwZPUghvLb8LKe+rE4z
EuCK2BqTc3vFxT27YXJYlOip2dbKkz0FTzYAo5SAMG80ifqQriEwU068fftuOpko
tpeiRfWeyJFdjbDJtjHgiOvFkgxVd43NFb1TE4OKo5k5rbAGdgzmdD9EjQ9tB8Qt
bWnLQPN23uPDMeNeho6+CVb9M0QSUatkWhtD5Mfi6kL1mLqR1r5Bg9VxmbWARsfq
qF9FNuexrew8exhw7oTk7NdYZQ5Glu/Tzi+oJFI3gG4EH22fWhEUlDRQQou2r3GB
RNAG5gSfMQmZeCi/g+N4XJr0evkbw0u/w1VhZ3e8/ZzVvAdXiG2TW3wDHeuFb3PB
chDWHrYnaxB2RoP5nt4iN1gbgq7EaWkVNl2Zx00fi2PYz9eIX7LWZDTbbYwpaRmK
W7anGtSD0G8m2mmlR3NExvhaeVNjDR98EkApddqcTaOAC5PYfI/+ZbBK4uGgvRei
5t+nf2ftL4oniVSCbXzVpBz62NJrinqhvWpM+dLrSDAFA7ZFLoOe51UZmC4LCYOj
0VF4y0jg3NPHmB3qT7vz18TxBJGNuAw1HJ6JYOx3CXDEEGgvDERQUCX+plyUq/0r
bJhIOV7hlbfZELe1TN4CHtJa8qy+soWYJzmkVvPFLT2w++OZnr6I8PXSEkJ+4nAT
t6VuXY5LDF/u5TXpjf7j6Zyqb+dac5mJAWvYVe/r5OXoc+1DaAmonbMdP+N5GxKF
A0aAWRXKJyLkymf8DTFmc8J/OGRbhHjhIjKda92JrO0rxrIiGtXzco6qESt0AfO5
cHdFjyEZjm0DcWp7cBXtBz1k8xCUo5O+yxzEHswklApWbYMKoz+loa7Wq9AxZt64
XIyV5jHfSTlW0+Yv0N+ESWK5OdTxdZUt0O+zUEC9y/TTLuxjlkyLtsRd42WkknIr
+tDm9gkLc3GJRWGsg5m+5EW+eTqmixhe79A/Lx08zMIWcDqObiDgofLLrbyhlwap
ZRCO4dYBLQDqt1lqYQb+KAL0QDuNVatwinKVLlPgWoVjXY9mPjCnPxwuls2UnH77
uSCig9ZIMrAEexEOemuTwOnSccC8HYFJqDaDo5BLox9lXhEBmiJjmN3xbdeOc32y
UBxwqJUbyL3cjFHzteTe1bkisDftfE6mtob2pKkfRsMRqnfh0UhGaD+893i3P/hq
5RJBcO0fgCutBdkRIKjeTIw1fetUjSrjwH+SZfrTUYxJRUj2T5vjs+ieHwYXYiqq
jWT2gIaWbGRmWjY0r1atcEgbyuwpIFam0yNVCLVOls3ll947qcQ9rq5D8XKLJE0i
uA0NWPJmuMPWw+AbdoxI/Mfj6F/roPq2T0rhUwseSPzfDCc9dHYa+EUv0L0n+170
ag1EiVJavAqZCmHwPlp8d7veZO1dQA6QPL/58Ar6zPhK7WBXCCxNfFLOmu4aRANJ
5xg35dHVx9O9adbOolunYFohDfgJsYEEGwuzdLSldkLV6eIZSQ/xrTnOG+l/7j04
k209LCG8AYRMzeXYqA145fb3ab57ghX8mfYY03gVtWHXjpfXNjGL/pjYWBnw+mLR
AMbc2xC/a2YTz4r7VbMvUv4UDEH5tKfi1j+JprGoDPsKaezaWOUB/TEINwxy0XqZ
58r2s6tVcBZVN36IqMMkOhQ4UsqOCsu+euKZOKxNWhkGYLnp1oP2YyMjNMp2Yh0Z
G7vtpLZyNrXzR50cBMT2AIWrZ5Fq9c0M7xlWg8FSnhP9obLVc24gKhgm6u1QgAMq
uhqYF7BINj1lBwOpWZhScfKXziZz7op9EFjmphKndxLNkc85J1FY8SgJM2NzLyUA
dAb3/zg2twx3oOz+lml80N9Heq2HN/HnGnLXovFvrB0wdnu9Rqv1/xEQWNpNQUzG
mlqVRmU30hs0XYOqezeo6l1xicWEcSe6Fyz3Mr83DlDmP2hh4OUizfJTYfqdtYR1
t4P9dtHqXc7wovVvU60He8OdPQ5nQn5PwHrOhNL/64HuxAS6I8/SlkED5SvR+MU9
E6IEHYRxaRCKkSIr1E9YT2nt5BIXRRUC7KeNcSpE/yaR2N8Gnj5qwljk52AhRV8X
0k3zkEkb9pGZCMk2ZwnKRGvc4ycdGKe3yBEnG5NWevbnh4vPSizL4FbbYBWRyMHX
kgngxVc1lOfNIAV77t1zX+FlE4p3oWoEIABHM2mXu4l+WpgrwazRef3JI1nAngjQ
y/+LmEHiGhlTdlg4V3mMm+OHvDWM8/06jNvBCIivlijKswvun1AfjVGLzT3XYsyg
KxTRHDh84lqAR4k8OMUC1EIa7Emj1NtDtyiUgJz9Xn4aka4K+bCaDBx661bBZyEb
UUH8MqqaX2MScnp5ope/pWw4t1porN8wsGm2OSMM9bCoxMBAY/zXgujy3ss9GWOy
hHyl3eLULiNDhrgvn+oC4mtdkXELjqc6VtkbkI3fvpHXIJ8Xw5qgOS+/4KGWR1Zr
SVzO0jmQeLE9CjAkavfwIXjGLcSwqG62QrenCPjcXjl/6vyuNmzqw0qs008deKyL
pAUaVR+JQ0ewWjYdru0Rs63tsPi06DDXhb7laR/T+atkdYYMSlnooynzIScFjjxK
Eplbp/DKM43xGwHP2w5fcJGpnsKny6opIfheL/wBORQk4IUdPqtVDZ/dJQQdKGb4
pXgydnBM8ff/raKb7CjpYb9pVI2rklIIZ9n31wqu6Es6aHPFCDg21szGTOGUutPH
NqHyAE5ChJEUNqVCgK4NW9TWNwiOa/OueGMS/QJ6cWEyS41J7AVZmRQrlva6qlJ0
kf4hBlbk9Qmbze+OHWd+W2Ca24fZs4uEn5HVGJGRU18JQ4qFSO8wsyUQlSBLoIAy
uufRA35EiQmEA1Z52iluokbOfv0Y6TxcRGjoqHTnm7lILQAGaUzZEvcARgqP2IMY
diHH5YiSFkJG2mQ+MXtLbfVyzOF3SYs5hciUa0yXK6krVnAyu+JL2hIboqPXkFuq
BI/qD3+CLO8cDCouGQ1HvUvnNzMkTOB4J4cPtMNTJvEweuQ/S87BL1QIlUeGLbDJ
uXSykWZfv+iKTHxQN9QVi8sjUG2/9T023vz1tfbpm6lM5U/MzjUiyADdyv0uz5aX
AwIK34yZ61azhm4fhV7I+gz0GaTAW5ailphkMCWF1MBR+uA9qm9tmI5NJItl01KA
wFfm65f5cOIsRvxqbyT9Azlcy4D1OlpaIzQjq7cWCq0hnHK8eLVYHPsq/osqmluX
T9EiSHvi5VXH6OxndtReP3xZwO0vNQ1DTpxJXLw4RCC6fkkKTn6eKbTuaO/jPNf3
JwarClGVSV51w+Jt54OgV1pM9TW+RNbKJ3DcuW3yDctNdymk/Ef3UZHuFxDtxU67
NwpVO7uMbOKUQWtERL2RnggAqMbsK4BWk+bjZvS5RgwmUxaKH5qgW4sr6j00Zq3o
TiWaud+xpoeJoRBf9LVnHtmsOdDVS3bO3VnYFpW1S2YP4q9EZ0St4HeoeY75McOW
J0CEl+3uv+4CqHGW8IFTs6lZBeRD3jodFcKjP7KIxKdMFS1uH40PQFtIhYgOrYf+
XdvwEAKI65LtBtKfZP/JXROG7crmRf5xUZQWgw/k/JfbeAucAwfvIbBFloAscW2P
CSxcTmgsyCx5AziIqD5XiXMUSwW8JW3F29jXbiKHHtLsEjFmXAoe8Cb8s6VbbPVC
1ygpRa5QkfNvxoAKE/faVrwkA2yu9gKetkPbH7kKbxHW1rKOSXJAKtXm1H9G0XIU
SsnRe5I/LZGSmtTlOlXwHwGR6GfErykmWcrmBr1+/BgFMRwLWllTfvBehLyaNc7i
ULUYEVYeWSAMrTEe6PQ3dJ/0T9VqZnhZgkuoETwbZPK4sqihsbMvK6MeS4SCUpkq
E2+i+O/hlCNrHcimy1JS05zr0bDuA2pwEYtlSI+zLMs2UrhbYE46xEY7or5e57Vm
Ih4CjXG23SwMVwgZ/D2zKmxte89r9tvfMcgZk77PzSGSmUCVpOilO/v+n1E0jcN/
gkkOQLV+dmO5nrxV1ti/JznL9YDdNICVhMwPChoA/j9Z652gPnD2lk6N1jKks0UK
P+yj341ssxluetJzbFZKbSj/Hpqst2sB2NL8FhInpCw6sEyy26FlB9902bUe8XMz
u4QyjrRgcUySpPTCMDf6E+MvS3WfNt0b+MjVZ/mdX2STRVxN+oBtgx0b30Di3jcN
irKf5L6A8qG2V+irBNJx167FhZvnexqAJLO+NG6WALFopUiconMJdwE4C2zYApXE
51cfQMTZGy8adIa7nzQK/vmtDAch9DwwIlxovmwvFvai9M6FWx/fKDbTY4CqDISI
lT79x+wCxLhGRbJa5u1DajnsEMXEc7r3DOaKyuSpRjSEtljjGkU8bYtOaUN/D8i3
nO+pPlechE9yn+oq8fsvzlhvx9k4x2QOq669HzH7+C9fEGtzgeNdtw7q309Gfudg
tzSUhyewjZxrOWKVVoj2BwmHtWa3LVOra6f3Y+Nwk/vT1CJOogNDK+llgi/R+lSN
C+oQbYUXgMyTs/0LpsB70XsWWy8gFUoIcPPcOlVEdmQxBGwrauKgk77VulYFKkRX
6uQPoOo4JX2KpW7TOQFGkIoZwDFailD7DU2Xkd7xyEmFMEV4+lxoCru7QuNAp+cs
9HW/AKW2iCvQbIVfmJOlhE++3JBEl5Gn6qm8o63lXBGpB9/djsBbMgGdk0NReZHb
m4mVvlgBKHKWt3H0HhI1+ZQqNgcJV3ifeti40qngPKEGxt4glOHdK91w7G+yfGpk
BEc1YwtQiW4ah8Y2AVUecG4GaVJAwW68Q2OYLk+RPnMtS09Z0fuB+b8/Y7kG7w1D
sWmDN7w8dM4q11ZubZVVYiPhqS/9DOQXIBn6niQ673S7e4+blAmGiy6PDCt9Xddp
mqMaAngA26bkh661b3euaJgvuu9b3tF6G1jKandKQ0O6u5GGhMAfJqPxWf16pLQ6
cK9Nw9+7jIZ6bzchuDCKaKgr+Jt0zQJ50OR0I7qBQ17Jh4vFew2bkok9j3ylLuEt
AzjJUwi9TIKoF49Trdr1hmRGcgFmEEzLj3smP5sxJrUNGEUA3LJTQEspmjDp1hp7
S5wsny9nB8FAT93YxNqJjaR88Ootoa61UpHZ5r+WWBzZbptECUo4v7pXvMTljz4u
NOkv3J8Ej7TB1jj93q62BVcqtduCz63gk65AMCMlFJdglSM5nLyrwwxVpDEXnxyV
DamuoM/idHJlBNTD9sCeKmMQILnoJjNxCdmEPB7yWLwu9E50P4BQVCx6WgUCH1/K
Kx2vueQMhFMDIYoXAQ3urm1wFFrn7DHip83q0Tl30rQjwPl1d7XM/Q6+Or9SLTww
cF2BxO6wcaYWEvD/w/1EFRW4CDp6fZ28jl4KgHuODQq1/fZzEffmrwkFHEBRumRg
Qrs1kiNR7o74jL2uTmuF8QXPqvKoxJfKRpVXHtoSv0nAxY2cLy9hMiL2M19IGKsG
Ex0JIC2gWKSg9SNiE6txshqNmho7W+n7/EyPoHAqy1eoSOIVzHvJUwdhGvU9jv3j
tM4av+mTpPYbnviqarhYz1qLtt+DKdbtU1x1tGL4h1PHi9cSTv4aWsIs397oLp+0
3Rk9CErbmT21hCwvVAg3qsThT8BSxgaRRd90tqsIIQnDzc/Gm3E07trmeKT8kklZ
fheNcmAVu3kKQuiaawER1zKvgq94e+YJxOk4Dba/bQy/VzpHbxCOJAtvnvG6cpJS
uSZ8SNEnqFB7t3llNbfwiJDo9mCDBsUBHQP6wc7Rjl4Ss+Ruswfr19Ut0mIfUz5b
RmGrsC74NDWyamwRCA8vAhJWCnaIrnfRiy0Nm8LZVz5XDKxRs6ZxmYBdo3lPN5J+
2eL8EzZyuUtRbKrvZRNqUwtr12WeuhDHqkCUiFJcmujKpKy2migveb29JRVy18Y+
H+cT0uokdyb+bCt5JU1Tfjaxx2GfMUtTx3/4cayba+0TOB7MeCwoWOdxSvjPM67M
Q0l0NfsXkZVOQGnoAhxRe1GV4gYj0dNE+jRBokItP+T5aOPQmk06HTGCskDqPbm1
YhdeIYkH7x7nPzE8Pr8zESgvXFCM4sncYN7Ap3wsj+7NowBFpQ/Erzfj2bqjjL/3
LOvl8OAYhO5QuOyHcKPV3EBKIsMo8NTUvpJk7/AQZelV4uHftdRk+9VhvdBASDQj
S12S2PwALWRans+gy6nde7SRwP4oBAGRblCGZr1pfPnsOP999xrExVNO1/6ec1Vh
TAUaSGP4mQ3s4/+SnL70I++xJ7SiSTQwGAI1xTM1r6rUtJ+0t2zSQ55ulAEfTaCd
2xr3p2iYmyBuIIqLtQ9UfHD3T5HkHRB+LwNlShh/y/tZDbv2wPqL/eJ/60r+y0Oo
5V1HbxkMyo+ig6pWzYsbA/+8ZJsG5DvwBbzG84kBIOR7/qlbKJj9uMwvjkQ+RerV
6GgW90IArlLHjIDA3BXiKoVShSZjwBo4wPtbXM7js/aEJaV0go1h0QLJWzDy1opj
AzRQyfG7AQt2YL9dmTdRRSzRUxICqx8zjshguzdSgDQ6N1BfDbDhiyfjWM+tMq7G
acSvAlQQS9Fnb/Bb2UKMuuv2S/32u+SDcQReN4aKIGqeABQeSyqdCUPpl430iJAD
3xV85X4VVeC7arrI3t0si0uJiVY0SGI0BozXLrOK52Xtzp/H+nIzrKwCqBAkIIw8
0UXLgcdVg5ZrKJU1tU9eZiN/kJI8Jdcx2KHFDBJG0ZNZfR+oxZ3kUFtnoKifbcXp
REVJD2gCpdY57AH+cIx6G/xAUnRo6Q5s09pvhqhghk+7KqX/DOXuoVy4MZPdYcC/
I5BaduyvXhB/Ulwx/4sp4gf2JOn1ezT1jKQAr2NSwBKAk4NmQpOAe6F0IelkDD76
WmmXdvr6vm6vdHR6XdoaoXlgdv9jx9a+CoJp4ZSxvfJK215XL3i/6Z5fcfvxrAGw
7sfCupg86dlLtqx29lWUSDY61TFouojvuegvwJWoOtsCpjKKWz+XcUFhPmTkDSok
/SOdhxKxo0GHLtGinjT3WTnrcCD/IuNgHayqxPRSawbV33uRMdDSZSLGmcAaR1KX
uP5EjK0JZmEDsVw3j96U8+VIIBO+tAf12x/fj+nlQgMX9//ZXqkiO7FgIJnS5fmJ
xlMzkOPkxKURR8T6ng+Uvs0T5XgZAcXPHoChdURf7jVQtih2pjcGsTDULRenS/Wc
y2pYHQ4kAqC5mnW28c1YpMevvIsqrLOuBO3I6APnT7E0QuOGONNIwfCEaOi1jZr/
Nao/nH7NGNom0am4OQ8HPjCtMmX0Qtgwv7x0xvjcI9RvOnS9q95RXNV/KgAoC5fR
rAzJeoVo+Oufg6TrU2x/YzWwla2bNaVAw1jJnbaDkGyQPho4oPWma88Hb/keffXs
/32r7IcjdJdURmi6lSU/Tn7p39RlS8WZ3KW5ydAuj68hzRa+HqbGpNGgBF5UCXug
dBxpijOeJYqC2X61zNkxdLbiSlHdqclzxvTfSsJjT7ZyQlrthKACInfgpPtSqjGT
nWX/bfBJyv88BKG1dLwwg63XMS3nwo5C9IDC9L/g0DbilbAF9GjrJiBQDFB+2y2r
vzulqyE8grahW0Ur2fYio4fmidx9Oslo8Q8vho/tw23FciwAGmQ0DHoUr+J+wqFl
uVhl02mTkWh86nCAabvog3g5Jy3/8sx2bp8ynBrvQzksz6m9coVOHD9wL2tsUnHU
uLLSaqvF79roJ9grfs9PEi8wbfDab3E2U97V48IkGTst2zI6mqPANYnNIolIHKPY
aP58o3k2Avv6VPsjYVGomOm8P41bZJCzHUXljsgUXNHgIm1EtauYULpXjUp8+Z6V
Stl0pnuNnQArOwo1ihnxafvGhYSM/m2KwCRPdslMgrJmcU6aXkDNeC9dB0aQnD6F
TXjn8BG52AHHdlC+cZDMjIjn0J/hNj46pQjplgVfBCGsIpu9MWIEoTjEJQNZP6pv
189YZ2clxncs7GBtZLQORe6c6Badgm5+Pbe4mW5UzogMbg4nDw51BhT3CTlNYPMU
/dWnzM2uHdJKZ2vEWbbM8k7IinXMNi65x8/vXDvNxLIFUzeDcIJcuCZbtoLwTdps
BaGjQk57mR5elcC/QPF4frHwWwphdPFj75J512tOnhUf4nAnPckCIc99XaKef0oZ
exlW3Oi6v2jlpng3W/w4sFTDs6ijMgTFFUyutw7ij+rZ/XygJGRV4uH+sXuO5X6T
nsISoGr+Fyq0npaaWJvCffJsOZq4kZw389SYVIQ7RTy3gcuu8Hzog/ZmOUaYpZ1y
Wcn4jBvFQ1jVwE5fdRMFaN5Np3BZbUO0IWm8PcftJLad9aF8dx9Ibk6CQIbQyzO8
mHAvK40byQlojwo4vf0Tlhyz5O6Z5ZcZCYTT4P832gbhInYcidcs/z2sJv0ESYEE
sGV9LT8IxoCjRXUWbbGkerQQ9jdru/c4uyGsdmHcGbDhkmSlAcxnCFFRTsUbFlf5
zOi2/RVwNeNS0DVh8sm/n9rEAGAC0coi0bqdCu6V7ncnFSjFLu1tDW6t+1xw3auS
Lf+54TJJR/36j+OABShp9GCUXbGVz7gCRrk53ITWNIeZC8eVn5A37YP8VCogkqfP
NMXkyC7QqredUFK23YApY7auR1Jtj9R8/Tint77hBJnAhRmEjro2g9MZZWduhTAn
4YQdLEmp3gf8jaUc6JRg9EFict2UvtzeaklMJflSypz6gfJcVDc6ac2GlcwdVLud
PkNA5LtzEV1z9lDrQFaaoBR/6VwSIKAC+fWhK3D0fo2AQVra/Z7ad89wr5ZqpFMG
1FpYq1lCjmuq/+t5LicWaVeLDdc9acIawg+4J2F/q1dgYvoHHCUGqrRPg5t5Ml0m
I8kJe/6BWa5qU6rNV4uB28Hkf00tOzjl0XRchNOWP3B9t63AF7HlyE/nc9ALDiH1
SrkTSfy0BrIpIQsqVfUJyRmeVe2M39SiXkuzXbprSVr4J0DN0mekukPlftDhRTNQ
+EnL7PJg2WIYyBaQscMl9yY+kua5KiB3CjTAlZb+lNFHhBP7Z2zSep7VjBnATGW5
sqzZ1HMA/WJeBUfWRYoslqJL6XMkY1qq3BlvgT8B36dG9JaCGLcHX2IxU3wjvJJy
eL41GVYfRbv04Jx90DsCkdta42eAkZggsAbPZeSKBZEPhQIdUleKnaQhAE3br/A5
ocYqU5l0xsU+4K8O+ZN6vhGzBzekqjvNzwmX0cPikWavPGwu+eFm27Rgshjo6lg4
reF1oBd4D57xHtnJxKf510NRVy+0KHiRM1I6beAa7giVJCnStX/GYDUoQXsQQuHU
Q4QVgvwCjFGUqzSaKW7M/exRfXLtc6QtQ6IK2ByqXbjpWvaxJJLTom/XzzswLcNv
XlV1cSQ4MFiPJLIJSK1pP2rdys+xIhCxfxJphnfslaErJftRm4TzBmzCAc3WS7wI
9Is3WbTLiVHD3uGVOVzyk3dXCdOfA5BgtmSXYwSjE5AHqtB5qeL9pgsmobm9Vqyj
fRYgaMdrdys2uPDe3CDYTvxI98b99R153vc5X1WxzNBmCJOUbanpuotLjBwz0CEU
OIHIQAfI6illn9rFurfHZZmM+yDBsVc1N69ySuTRYFQAbV47acwzhew+IkSx+M/T
oH25TtHJdRlJD34b+tZruMXjUcQh3C6d+UOmxj48ExB/tvlZe85rxaVIHf1PhWN4
vB+qVWUGCqCeWYTvyBfnRftRX1b5GyH0RPwZONPemwgDai0lAJuOacqVEagBYpt+
hTJMj7Cm8Sf4bf5CV9+dG7ZYnoPGSt5fJcCZ1HpM7jzIfTxYBHEsoJ+0GvGEPygS
s74lKJgQjcZzv/Bq/L/TSpVSCgS98h759l7AxJDPgd5ZdTIQHL19ztFfqwPkyrlP
JHt8j82R869PeAzfacEeIhjITPvUVhcHpwNFEFkDaDj7cccYXSc3FwVQ1j265lJj
EY+rvhRnDmB8D7H3qv9UMJztEStLSS1vOCTvR1zNhoQQAbo0Y6QJ/RA0pR6SI5XD
1r78jYWxGRvTleZN9Raq4KmixQdcIemvMeB7DINRdvz0y+HczeXfd729vh03Ryj6
5d5nLpnZ/+Mp3V4kuBhx4SLJkRBXUiVaCwzqu0IXR/veU3MvfSaSD2lak/lbPxLN
0QcTLKFAow0dgehHxSPv5DmGOSLCC+EBrzMQj9do/40MyQwXzhrE/Ee6sk7k1m4g
zhoNor6Zry89IjRKdyoFw8KDor7DU2G4BYcyW5YXWGhu1Ge4rBuMhOetpuzjgpmV
Mbkbvs1r39kNuH/gih3FWvZCNqJ4IPaJX4dfKxg40tZF9p7zqwhIVe2xbpdBj4Cw
Oh6BHRrESiSR+Q9X5d1BGtLZYCwCJTQNi9zjI1SKj30lCAj5d70fhYEjXS1lGZ/T
P0uCIN4LVgbp21OwY0XKXFzPfyKXt08WYEQLKsD/TTIXlHy7FvbPhT3p/w2e7U2E
t9mPbZsf31nnNN5py5z0SKxXbe5MxQGA0smUsBF+80ogb/vHRoi4OAaDFC0kN4c9
HHBvOuDEtGUo43lh31pxLrLAYlA4M3ch4M5qLB1Ts3IHFk6VkReNXxPxRjCAf0ix
i4nb9t7bNAQGgQRNPMmPK2Be4TAfWtTsGep+K9WO0N9WAFtyNVJI99SzNFXyjg9c
9Zh6EFChBlzfs3G0EsUBJodNfsSNnjZREcEeOnem19xFiCivWI5XB1iND16EAAfj
gvcqGPCeBqdsDW1UU3cLVjLyVcTpY3Ey4PE0+YZOm+fNs+mI+7b5kg7ufAlianVY
35w/1v4oESPhx67FUBXS/yK0bbRw3er7NnXz+FtGA+dy8KIKXwbO/g/trEgZYhiA
pAU4I4zRzRWzs+YEa4sDoVjX9S3u60Iu+P3Vjwp51fJm5EQnMNxX/bZM2RHvMslJ
NwuOZ4v5mBLiCXIz535K0tsLbY+JBbvWnUqAL+5b+X+5TXsrSUmrIpfU7aHrSXsG
PfePcQoOkQWibR+5pzLludg7OMGmq1oI7gnVtliqlH6ThE4iov3ZHoNaFeAs0rLO
cEm/N08oYLbOYXnYR/lvvXPZ5sje6rAh29WtfjDu3UNrsdP6qqnyqBQ0bf4hgPRI
lwyTzrXekITAkT8WtR5DekTQ9QILhLns+VMLvyoLuhQIK+4o4KjjjepNBL6GzZsj
U1Jxirtb83PeZZhGrhVRb2CmvH8dLPBTDqqU+W3qzSBm4A2BGpond9gJlGG7fQO7
c7IrF1BctEBH5eTKT7GNOXl39uUE2dUwYdLiEyniDP1UAFgkuQQk1catn/+oz1Xr
VSXg4EbjZ47d3WW1vUgAN23+2Uy17Z19N1KZYN8mzgTZt+Du+BJaOh6XFTk4ofF9
s91L+8bnzD0byC+PZUutn29RuE/5wnpoFznjd9a2YWCRebKCuJdIGYwaoOl7QedM
y8iRmh97TXlN7t+vJUui8HVROQMwMF2inCaVUzMaRp6V3uKoLirLsOGwK8S5P4Du
D0f4y2lBgsoGZnZi1lP9m+YjNiIcHjna9j4YZdScucKWDrPZzRq2Z4HRqNBLx+vf
ciKT1glbtVmF/btxX71fcph6KzSVp7X+ql4UzEfmrDYhkxUqZcV05p1rxTc6tVRK
MIjWz9Qw4FbwwsX5tDoKq1MPmmQYXTeJhDsjY7vK6WTciOaEo0UrU2Z8uYno6ba4
M1N15oCPzkhjLlIIa4qIoVrdZWbvyp8WOMQzsa6cfMVuIPOiqBB9jq/cips9/HBb
o6/K+tKD6jD5DjacOJsAv1KqRsM7RF6AJmDR+HgZJoqJTICYqYx8VfSf2qtgAWz2
yCy4DZKM0ahr6pygaoLXoeDGQv3o9bAYDP2j6ZP6iL048CuinYgLw63+ndPsYY3r
sC3Fo0KqyGA+xAj9PCdyls/kF0zbEAizLZbU+t7mkHGaurzLPcPMQW/Z339KlkJo
vLVkS441OUSZhv3ONl13MfJZsijkkXKzwVZhARNmO+j1uyz1S3uMvueoe3l30mPn
wt3tEzkpFLwIxQRAItsV/g3bpo5RhvwVOFCXa00ThbSvckh1wAgTY1vjQ2RgjLRB
FG9eFRpF8i0eNymV+iGC0W9KZUGyjbInlfrzH/d5gI8rSFQlRgZehsX9MIDWDEzK
FV+P/nT4HXv4abNW9Ud5QqW5ln/zUK6G4V34/bLw8j1opf4W8tXLPFL4RHPzYxom
9JIdE++rRhvVuZEv8xGz85F5qcG5r+nnyyjPSYc21+zBN+QQuxOBiUIzFPJ1vUCt
EFjFQo6hTZAdS+b4z6YZ2SEtH6z0i+lhSzRyfivWDfibMcvSwj62wPs/GIk36/f6
d2DR3f56eyYmzcniUeL97Bh9cTidLB+eJeS4Go3/cja7hTAeVYegpT7KJjdrAKln
Xgki8YKfZG1Wfit4Gvw0rI/bJqFu4/R+fJekczefAYwOg90HD8QMkKYEtR+YHFsV
Y/4u1YOJnV91Vkvu7D6olmPx9Zq3TSUqcX6DfJAis+XEpbitPmXrZNdWcl1fKj8H
2bvwebtAJyK48SCSXqWFLRmcBmQrOqEzbMKr0fQdjupmf++/PPePWbMrvA8ga8Tz
b4+3e8FFMo4MN+lIzeB4GFnQu28hr7wxejndwslf3ujqcQWTiG6laxODMQaomjUL
8EqErpogG4X3IRF+8+AwzE07yjLrQ0xccgKu38Z0vGt5tpIPfry5WDfHwAeimxNW
VC/xB+v2Pgk8fteH5YUmQO6ZtXBzC1qeU7TEPNCmdj08my/Yh7MtYJwrMu1THBYQ
GtmGCceW9NMkoCE2llRO+LXjfMnkLRZRQkI+UxyiBJNwIAuyjRSY0sULgKbMYyaU
lmyDnCabT3LG5NvSGq6f53HIkpQNQsGDNsg/XASKx6eb0an02zVCUFD9Roemuv1t
wezcxktJlN/aRf7dpoVapXQ4mr3p1VsHKMtZoxAJQ4s4tlMbeHmz8GFRCaRCOd0g
84+4JelmYRMHEty9+TQynMsaQnQk+X3vDOn56OonZdSuFT/opdG2HYgG8Nx8Iyw8
mORYs7z0hLH2GA9JfDYvvkDafWC2di54TytQ11Zmj07e+NyYArbAOgULeh7E4b4O
ceUvemU32xdXaKqrZVOV4i074mzm+gUE8NTrtJAZ3HIx7K/fPxhBHwiTpcOuAxdh
nK7bkQ6Lvue6ObRiqR8ZKVu1/yjcSstt4tsAVpK+rPKvf/AJvMAT8ZgKWzDcFags
hV27O9FSHuLEXLgJuGtV+A9JeSuciW8YTOu1mamLy/bB/7EbTSy1p3qTYd4A4UFH
mpmY2JqRF46P40vWWnmuLC0QKO0EqRbrRKew17HN4jG+scDwD5A3b/bR3ZcHzc2o
ppXuRHYYRq1w1hoity4ApBULQ/L++KbABbrvPvMV2xsSLTurspCJ6PwHWvSjI7nz
3oJGFx1KRUti0SiG8A6JFkT3rXKbbKCa6Porj+5eXE4NHaDV0zaBgVVOFcxetVUH
ktqnvVrLXJQNmaKb58au8kZo0VTsd5J8hpBI22wo97JMFnGyFpTACuLp8auoITKW
r3fzHrQmmFlhQZQ4guZmlOfAkkGQ69Dkc0zqKVJmpC+tiIy8dDuDXL1/ing1om7l
84O2xX95r2Z/gUSkKA8L4enb9UsyTgE/xFL0zMIF/SUubDDGHI7dsstzUXnbC72l
+vWB83/QSgrup4SbtD27+D8ddpYf9IsUx0HnUNQ+GaX6bEYTLDFkA4UhPcvNUD/A
kGfZjG/WK54punh3u2UiYAHPf1BqBA6Fo+DXhAf5AF188szk7NhlUoNvjpAoVuYY
tH0+9vfrg6W4jXNt+I+Jmtt7YlJUFE8HiIN8fsvAc3GNFFCf2jqiOTPte3AaeY2O
TQaKwS2zbVdjHVHtjPslpzkQfMoq4kQIZd1QJpP1QgvpLWDiWGsv6LrqmhLgxTON
lWBA1jpjZzvndlxGNIrrdQwacc+vFoMP/xxUj/7gbq0X6zRHvhcnB7ZGGc9H0FLh
B/0CeVLs0S5pcIHKZctd23uvhL2uNiDYlah71CoTL71BE2+3h78DbTEtRhs+U4YK
l0SJJR1f9VRrcowN7gDCWbpt+XW2qPt0C2+ZlQV/AyD/JOIJ1i5tBZy8FSTUOlei
JVAlpZi3uxCEBg4g/CKejY17pxp+h/qU7jKPfkpPi7Qk2Dyg9nIaKukNWdhO5KuQ
6lfqxOnhKkWi9YnYVuOBWaFSieQ/7sdScKYHuWHD4+HRby3vnNzRR+vznnt7qLWi
OK3mDvQlvq9BbKfy4+VPFHNznBC0B1qpsK5roUDzv9obfpqjC6xGiKWnNQlR2XWb
FuFw1HMMdN5E3lyunUmnzOpNcJ3WJH9+CuI8JkdH3p+1Z6Z/mEIjemByYUrFQip8
NrfF7mVQIyN2OTKTGm6Ocv3r/HgehjyB5qzOiLLvLdEqA09SzcJ62zt6q2XJS3wL
Dw/1fyb50aZJjXFJ2fbOncW2Qk5EW2knSVN+ATvXHSB2Az/2lOns1vnx7AooNwzJ
tAXxBp0ad1P9WLe9wCoYBZaIfypHrNKQmO6shYt6EUxVFTbg0cbUFEuz/eoU+vgt
MptPpTx+vLv+Rsv6BjtcJiNkYkUnGqf2/zlysL5JRg5M15hncW0/CEXtctv157/s
FoNGH2p0MDaDrYTMpH0t1Uw6WkR4aJpeg2J5eL9xHoBRqyFmmnreJEg0H5K7L+uN
DXyirYIDbVrYUXrhDxjMLyBpkzXzKr+Z1jzU5Dl71IiSDBeLj97uZ+s7gHwV0Nw2
V1INap81vFNrckWKHPIHMk8jdwVDOds6++w76fgpK7AE2Cv/2yjioj+bB9yuRN9B
/yb4EKl+3vBwEhzXkuiMF0ylrQqEBpikEwqMrITWPOrK7CPlGKfCelJEw90egQ+5
M0bFqYeiwtlQxl0LMSJU4e+Io4QUiqMjM6epD73IpAmeXtp9mp8NvMDlYV7l6TLw
hUXhKcH4jXK84jbm51GK41eAv6gY8KWtkk4dLLX3/ZLnXQsCKVWz5LufihPRLd+w
LqvCStC8+uUt4eNnZf6Z2nD/JI7kDhu22ogmWPkyuiveV/8IvEQKHNB1XkeKeNUx
9M1f2+ihwiEIwakvhUnrZdeSvbjtg9SsSjRQHGXxnzO08YrtBTjXaDNkZ1vntrdh
LrDZ8R4FaDp5Knx8+2ts/WX8jjzY1M25WgYTXGCFX7EuoyJMhiVg2ZsS6qwTTpsS
lQtK83yuISym5S2+QpkqwfPqTBDru7vSs2Ap9Gy1lWZa2FRzTmEwiZ1IWkRXcdxu
WTNfcQgTZCOnHa8F0SIMUafcu7R5WG7ku+J0mJJGBjDehu2gU7zTVhyTxihvuU1/
+2/qFO28x4kAAkkBJElIim5CF3XRkQXzWE/7gxSSBSKygTMiy4uCybwACb76tFro
R73AY4MENuasJnuTBq6nPJKSTmbitJzv+dIorN/bxJY+efQJuRMpzXFIrVN5o28O
uehu2hs4dtwoyhdygfomQXrAg6i0jtu0QxstaOnPEoqwq37qeGhes+Pp6UKI6NSs
L1FQtPVSr0kccg3lS+wFjP9eGKyrpkrTyhswsHFgl+OPKFBXk+IluBsVc81dimYb
DT3cqSOXzLDdzkFniK7uoHSOHOnrClCD+GxliHfPBv24AcnhxtVDYSJftP9Dw9L4
XLlqS7vfgaiG09AHAbaWeOkVD9WjCpDaj5Z8UmB6AtwWZOr5Lt2AqFM9iHdmg/+P
kiYSDdXKdxNllhBwWe2AIpIPY78WIwB6mSjND2kAh/LJ0U3USgslDTwPp01Hr0lV
SeWXGPdgoOtcEm/DrFzM58MwYKb/3q45fh/THWDVrdwrciSS6alATSiYVqHykKNl
CwFpY4AqvYfL6Wpv18PMpycfeahCWNDaBHD1epBv3/KtssAtzHc7+Vry1Fxd7Io3
hSl5eEMZaLWmFG2ONqiiGei2SpaHsvhhjuNfwiW3JYWKV9pdndjVHp3YWe6cIWq7
UTlEn+ESy8HrB5+2oujiQLZUSyLSOB49QjHTyij1i1lSyWYv15uk13S4kATvg0dS
CeHWmKvxyrIdK181bg3xUCDqr5h6iFAjW9sWeSO7Vf7javqcvvhsqKFuzaT4HTiN
g+NELXrpHl8ZQcjU4QhS3iY+FYfA2g9NMYraI62E+cZinM7Hoial8IsDIXF889bb
HS41aBkUJsgFjPy9lszuE1Paikt5fErSPcwJ4ddqOq243rZHvVUPouZa/XVUoFUd
RfYomXKvPx8vzfwIKZLBAsSwTXHiEAo/5+GbrJ6QoW0rBKvuwXvn1v2fiouWl5MD
WmFUhcuAXEB2HcrY6Q8YxlxU7O64sm2S1snewoYHVcXews6fnSAXOY2qE/RcAd+O
Xuxx7WN78UzB0V53yQR8RPq9QI+QI7V34GpwHGkZtw5svzhaG/ZHDIs/8iCyBJyu
glhPv8l/3RzkDaGbKZFAI4c4+6beCfa/PNjONgVNczLYEuPJ2imyY7hq77TVmpAi
wfh97EkNbrwQYik57eaX+zoGF7RfftmHX2FN6cBA+KrFG+ODArtaYQn8RQthg6W4
/BvzIYxpr8Zvrx4P9fJMCFS/6rWuj+X+L21WCLqySqF031wB/F4EZSvakomhcs9L
GcbfJy6y7ySX8+NZTuoKE96DPKCSoqLu+39dS+JcyAz7WWjlbAw3AMjSI1h78FXr
inGHc0dxNyDwxRUyWcB3WDaII2PLNHlJ4UPpnyYnAm2o538BaHbW4a27+bYBbTuv
KkZ3+NJuxLSI3Gjm8rixFCKVlOZakB6MM4U3xNlw/GR8NvBYsUVPrmxQZVBtB9d4
tOFNPtEws8y3cziHLSdtSa54/JJ+abeP2Jz6vyJmXSl+VOxsjx1pEW2+h7oqq9Op
vO4KapvsDloz3cHq6S7oqBKHALihmW6rh8XM/UUb/6/Ps3PJMBmw5tHVU2l4sNLk
OxEkafFA3VXeiRfBw3QaXP07u32YZsRw9+1CfBUT5J3f6byOr++xSPCJXXErNgLp
9F/50bwvv1FFKQaRJgTZQYVC3IqTq+OwQe9NGlNqnt+WLOZtEbF4ove4nbo4J40E
TpLDJkqIW6hZvLYrurDgSMQCeJrKiOPw1ji7dWl6zl2zTfmMeYY4Mv8RryEludNm
Hs24+zbKaEU5srzAPZkq90JvUTX9dLrder6ga+m/pZBjHR/ncx+lTesQIvls/ox1
rVBXKUQmE8jH2jWablSjkaRtpaTvzrNVXp/gWmrtrcRmefzK3e3VVkh/KIqTSWTr
C3CE8I+weVGK50WHvL2IWtiiZDTqeCXhCtlU9ekC6gYJy8l+8aovnkXae1nsTaJ0
qudiLdI5eiNIWukEmPX+nI6Mbae9cLY/1ugmf5Kazybd+6UwbpkcIg5Wwn5KYrRJ
Aq7+oGGUkfwpBLm4Gf18UmWXC4WUk465UsuOGZ4PqY88lmvqpIby43WNvQhijK9T
fvzFRr0evpGhlI5cFmb8paJqEttpNRvTiHbf5vTAP+5YQipQlzu0RcNSE2XhuVg+
/+nSQn7zVU/pNkqDHaYjDY4ucteuMNOOfnWr27JN30pmvsxcleuWMY0pXkAfCMej
sEdHS3mIzoXbLqOcibovosy8bSn7qks8XutwlZXhuWrTgv0ExL57xRdQjLibITII
5J3dXl3BiyrRUKHX2oH1IFiE3MIzYD+2o5qyu3PN10xdFdgYV8kfiYsVBY3m1F3J
kYIoFX7Lqtv0myMsIRg8zsEgCWpsZqBMucb514a+Q3BM4JDofl1zuhGvtYgEV+G/
xUVyc9+AV+jJBGssWn4BuwU9SYwE30RoFfZWCBLgt0zjHRVpHT6I1bn+wAyH0LIc
cw7d5zWzKiaJ+gAjSIUJqSV1FFRes8F90N9Fi3i1Z7CRkrJD6zwLMMO7F337q91A
DsiIxtKMWVPThPzINuCEgA9W7PoYLW30uRapCMAu1aV5E+To8NLF16ypExcnkdPN
bOvlsTdD+n3+uy0RI7MMfQxRkI/vSrkWwvLbxoaiAGicb5ozccSGAZHBH/PFDnQi
ZPRsp9vhVNgsyoyhic8YrCdUTecCf6XXco0omaXJsPwSbzC8X1K8D3e83lJRoNnx
eC5LbTfuOWiGJWBVgnEo9rO63dEH55B5baHO90fpS7O2DFN+HUMQK3AcUEsWqCgJ
Ocgz3hREdNm7M+C4zbm0uXgJAsVMuUimV2AAG29ucnx1yzVXpiVoEbFF6mAHTqdl
lGHOy1F74eV9/7kysUa7oSWlp7LfU0MpN/V2qx1aFOebbHjAXZfdA+TQH7XGRAsb
QIF8DN9uGzHili2FS7CG/FGxcNSCOC+Y0LchB5GFdm5FaYXyDf0+HTwCeqC/AfpE
VnfbWuDn70dqpuHdnCgMqaHG6dn+DHGodGRkLwFR+V5WoZdODKNNQ6GIeQ1r8AwP
AckCz4qertbjRqvPmhW+e156hCvWRdsM0LifIRxWz1FwXS4ctF5PA80i9ICHaXWR
p0lX1a79p05l+jPeoqXc56RnYkDhzuGpy33WaWM9QTueFsW4TjMfuaWr984f+Nyk
W3Se97/wxGSR7sFmlzkNpKMikLkYFo6OMUaSoIZBJ9WK2yjgq46vapCIYWqUUIRE
AEuGJ4GVc3nLTFyEmLhUaNfslrEp+1b4PoNnyg1z+NhJtxZM9e0vQxV1KKEK3SbY
DrNGC5x/3Sw9zdMhGV3RIdYNL1CwuncgY2iBFtmszr88BcKOGGtq2poIlYBoVM/0
Z1ISD8AuPCzBwDJQAZqtRnAq70crx/ndTrdPAiyIKc4iiUgzKyXXAicqeUTk78lM
Rs7c3UfaAtCgS1xoZ5yrEb64R3Q9GZPwRU1nh1Q+UwM7yfq9+Ch8bJc2e1b/m5Eu
snUgie7QuVSMpm36YF9cncGuHws5X03P6ov+6bO14x5CIIz823UVPqNPBuyXDMCo
cBqsOzd0vFjZSquzg/bnANSJUWoNsJicGpkx4wIFx5tUbu3+vHsY36+ePlfmlkpQ
sc22bsQzoWexypzx0/Wy1PTr2e78yUZMGkv4F7BGggs1+R/wTARk5Y9aK7NQYu5U
saBC44Y/U+Pyw0/r8Bp6+3/JkMtNW04ObNSocSQyvSoBMmnyWtTnIQlOP+99cc6N
+ZSq79OzfstPXYkTLXQl0Pw88YxNpKu2QLo1vmMq+d8kwHeyk42dV+K2aotymdqv
jUYwE+WQP3aKjqWsvuwhHt+xtg/wqaXXj9heAIrI/gsjxxNZpUdnPv/odeKaxvQC
FEdXcHJaKAD2ntbnCItLteBBw9fUw88W5yvvV83UlGrwaxyfYdp19+6QLXWJPv9O
giPHiUQ8Z/+ICDLdfBdWG40AZq2QSXEzZWp5rzLJ2ArFdrH4dL6CkUnuWDVK+sJR
bEb/rZ2U773OShKMDuO2Hp1CFHstZAUy+1W9u+oWPDTREkAHIwcBvV3uXZYAM/V+
sCASkywSfYiDSrfvTPXZHR11IC92VIEvmHENc3qJJP32Hh5IxVNim7eisIAcXfCC
MqA+hfxzZkaB/NEcCYG5ARww+aVQtemL6a9Qd9xRDGqoiagwS4yxOSTMdvLhaaiq
tKxSIi6BGcyni46y+ICFPEQ03mgk2I32YNwIE5cHuI1U6xtW4i8mxxRbs8CxyAd2
mDv//G1o2f7AekC6nhJhIsAgg/+UuUErKO1qJnDJ2xtQNbEMJJjho4Nqr5GdYxBe
l1pxOVVPIVNFmm/3ljwEW0uvldduGGmSDEoKmiRmsnyFqCGD8bE07Fo2znNO+fpe
e9QL3Fmx8qjiqEOJfNR0vs1Qsyv9/kbLLBJQGlg4TLJRHGGNofl8bJum+7MRAIwl
YbSWe6JpMKWxS2Da33/xaipWRzhcsCW1nBDgwrsHRUnTxfsQ333ssRnouxda/6KV
dB7UHt6ID8QZkJ3n2zPoE2tMdwTe4sBWyneczneO0LPAhbtTpqG1ZOY6qaJEOmWD
lU68H4PVTe+SeVDNHRz4EbJYMHR5mk7n+f6jKA9mbDQ9QIA5T96O8iv8AqxMTW/0
zKKFYko/y6GAjDgGi6zxqeRV3/iRixTALyugiAJhzHe8XvfOj/yNfkl+ycd2sRKj
UQeMQrcbXmtK5rxBqxh6vSh2Z8EzCYbmz4HiIbIimXLMVIt35KF/q9F+fqpr/i9J
sHzIHQT/4ucxAifyjXJtuO28TjagnJwUBYoHAtNV0WoFUkToHiKJTzw4by7bO/f3
kxxRNZ2EpMQWBIM/b09YLJ3D7YB8qGJdZw7wjfxw0FYW5OB4h0Bb/VgqBQE4asNj
mgoYkR63zh4J1T5v1fPIdU6cRLXuEGg6QgxIJJrg8bxmYD1y3mdCDDxUavXuUV//
Um+HZB1/MOBYHLx9DwQxUS/ltcdnaiJvdEi+tYRqX0HnCx9rrq1eMGL7IgYf/pHn
Kb4eW+XS1iCxAH0q1GcALzmQUQfN7sxrC3/2rDpI3iiZ4KlCo4xdBloiIsyCP9wE
4LVxP4P6OPEYGGtJTx00Gcvk72GLxw/W50tGUKltDnxRhX0L+SQjdc7uyqKDVwqo
l5ThJUKFdol9o1tS/s60/Zt+xGYI9IS65u0lHGHQ40g7dS/v7IlBWT3osMGWGydE
8amjiyhPrLYwYG6iRKzx1WmCPUob8N14pipTD1p1kpXNerogePnYjw3XHfOIZl3o
D7IGN3Kv5DI/IdWgCLdB8WVNPNFGF+chJh27HmSeTvkfmtGVYAx23Pw1AQQyFn3J
diQ99KrzhrFpLlBtayV0grLOdBCMuhsG3bZ5yDBKQNdObAZdsWiq6nUZus+J2mrv
rQdvpPmkPEDaTa+ZU8Qhx8TwwbKsRmlKDWeGER6T3pgThY9f0vEvXVkz1EhhTW8K
4lSj7YUh0b5SWENPFiVM2C3x0qY0ssdV41roM1fmIaArqzSW1N/1H/nuKto4kUnb
ocHELbynURbduFlFBKZZ7PbTc1yguXuQ/gjvVHGXZtFn8Z/wTqJ1o/I7uPZDok0A
hz/9n65oco3HUEJ1rNjf8RP4dZJWNPuwL63FiClT2reXs3traG+tjMKtMXF/yHqB
M9FekczASoxC7q1Oa1b4Bzhv7ned52/QREwkcxa9x2Jc/TfzCa8NBBp80dh2mKen
8vBqLV1V+MJpeivKVCVkWTyU5OWmB5aarTOotwP0qe5iaVSv74pozYjdp2ZfKDvF
c2H0Ej6EMHNfPm8AFRoVpAfVDJTwDkgVXvYkSfCb3uwZC7CQyjvBRg5SEvBIQ+QK
t7IK4bxQhAuXi/g+eAD29LWxUieohQAs4qcDaoQhWWEKhC8aW8/TPmibq3zIAmOK
MokQH1HXyHR1PuE6vu3eGEyRXP10ckOK/1SOggO4ogquPM3sNMxzAg6vBa5f1tnz
FDwLSqZGM1z57kpDoRWdLSCPpUXoQoxKrYNxEWj0HvvIkgUXGoXWB2DWCEPDAr+l
uyGN3BUS0irqZBG19MOShyAngY6GCMngUJIMXH/eSLdxskqgpV6C/n9NtqVFV18u
fDGQwwLOLy/PhToE9GpUTV9ZpuWs+dsCxYW8x+xj1IjA36XVqsJfAG67qFK86WW7
iiUTXO+UXijECsOM27syVLNmyXTU4sqtJxmkctFl1Jc8CED6ZeDHHIbJnte75O3D
GsOIG1fj47sQBkjGY7VsFjP3Ok53rfQYrnE2z0rbcoCSSPLVxsWD9U13y4pV7sbi
t1KWIRGsr/Xxwjx0K3UXTKxNZDdpC7bF1kO2u4cCoXDER9URTz1rtt3AgZCZ32H5
8FFS5T25jBcq/2vP5Cet2aAXfyZpUMrEPs38PYm7I2dAzQinSb2PH+v0H2ILxT25
NSNekOVDvQ63vBnCUpUsSE3W1Y54x7tsvS2zqh5SyEsnqBHm1UGSSShl8VcoXZwJ
joVswXJwHE4+Hkm/jGxc1/LGVRfWZBR82aC4SYTOP/50Pe7Ei3sc/RI5q112LKor
4wCjqH2dtQH79PYAzQOKzW1sVVwUiy15Udyh7Ic+HTqCQ58X/jLPHAQcsosUV0IB
AJUAVTv/izwmRrrOIYQrM2kVUiC/3HQKcC8PiRYTJAE6Wk22ATLQQ3LX9H5zy9+t
kq+vkLzwWn1NaSOQV1yZrcX1Pk94cpfG/GHta77OAwqs+XNnkNyruZ0E5wbTLFZZ
wDaeHuwY2phFXITfWjlnK91wk40XF7DCc2ukqgbBcog3eGVVLgX2JaI8qQAhxYXB
InCFLKn+8vVOhiGOPHZCI507kN8NEBvdZBE9CMl8CesOPhnD8ePsTlWTtoQLdEDM
NhLRj7Pu3wRP5S6o+F2LQc1esrj6J/35a20Nh/I59Xf47VYE4ylki0wZ7WmsyCHh
KoEdTH2AaAqXy2KdBtgvJpQ3qy8i+LGqExDdMLuYKvBF/r+8UZ76YJihMP8ER2ip
h2tQSfbF/udvvtW2NcxHMfrywNWEbtFaKNyB1GQ/cXn1fZjyQOm459dmCDuJcW5X
NJgtZfO6BkUZK9ZE+k/9Rm+GHx/tWQXqWY2iFZj3s04mBcjyAM9iR3a8njDTXkw8
93IdMnTUmiWzOum8jTnAW6XEK0UG+CTe/3a6sxUYLdvgQTtXGl8bX5+puQamQ4PD
FmlqfkrYxJYOgq4gofSG2ypCh1FS/XzpfdQSppS4Kt8IPz7/lysZSoG9paALqAKz
3vHdHSgQtvHXwE+50ge2IBZui1OhYwy/nG5w7tLV+pbTD77PKc92B8FJbSzDDMqK
8cSWKB8R7x5YKQknw9NSTAJUhQSB63mxl3C1ptIwz8ZYdr0DUWiyF3DybggxvyCu
D+/JXZU1ThfGzj7Aoh1KagXc8JIaJ1EFFVCxNRBrVSMXYKH/0lViiv8o8bWyA8aS
L+xH5Vezg7IMpruTc2Rq9yFpNH5UX/3sHMDTJSw0qqJnR1eRwU7vPQGRaAas+pyc
+MxkhJovvm8EMNt5L0A2Tx4lii3bMM9N4OTg6ml05k4+qqqeG6qBCU4Omz89iPWM
r8kNIKHIQa0hnnimiaZBqA8INGtX6MF9oVRVBvxGNnJDJr3PAa7aPfWcG1EqXI3c
FkfuqwNVA4HGjk0fBZF/pUyinLHc6qySDXfB2+g3xfJ2PxuH9Lgp3k8iidnkHxCj
PsS0KAMr9CSsVA4HM5XVxXxLRHqzKSups9qwK8/QdvCp/HR6SXCB9HEbXkTbSlZ4
LkRiZOLBxeNNMzaCmcpoMFp9xXxe03hK97odp0oV1pgss+C8nxWLlDL/lhoDk2nY
V9uhrZYTCKAuzpzszn73REHF9G/OgAfSVnFpYs8ZJHwQV0IoLN/r9Y2kF9ebg1eX
R0PeG2X6+ZxyxncrwHGGpG7etQ/1Ji1EBrfM/vKlZz5LzEWw8Z6cfGlCBQ4hJWwL
syBdQ8epQnrF6t1XOZHYumWHGwAxFNiA1IOcTHZBUF/MM5uypPJ+krX68hKOKsV3
YEZHRVVDBNfvUQiRY2TICc+IanUvyiyKzjg4UuFt/PT4dRRHBeQF2ba97Q+gp5LI
v4QuDknqUN6N0pHBZs61bSDkTth5uHbnXjr5VDqhmr4K1tSHRpakCfT7+K/HsM5T
KBxlOgvwjlxrDQk7GASCv3ReJYJPiLkgJuR/bkeRQLZq52B4FP6J0AlICAn4/DIw
Xd2cHB3lTueLTr2TwO3mp9mRX+zfY+7vMj/xHMMKlQjqZ+xtYSaBIOFTTl/c9y+B
ydRSCpwpy+OZayKHshI+mEjJwhDgf+CKrOM5fmWKygTvd0K7lfpJs+rNS4s0hIJa
U0rCQoyMcnkKN+EzJrNxOsa1+hG9Pc3NuhcfY2XHdn0cCd7fQyd6AgpyXmbY8iF9
VKH7yaYnvWpLN+of8xV9ICkNAo7kjJBxquTgLRDkAXekATZJI0vddGbgXV2HSsti
iUHWGnENiczY4gxj0tg+leQBlVyrPeBCA95X89HXRz5cib2pmHU4RZtyb0G6NjgH
LUI78RcTSCCIq7kaLNFzO87HhffEBIij30OvvGusClCM9x3wdqjHncQVAxYva3Ci
7VXTVdMNBZBd23LToSpZRMgFZB5baN840/+Ij5YMoz8D/cM0pHRnGIy7Rw8prBob
Sszdu8N6/H9avKsbmIzQb/aQgjbBEZ27+NrIBe8050DPqs1NCzVftWDOiclfGjx9
NM+acUHCvmQ+fm0y2Crlodot1AMXQ9qlUQPgBJbTy2weU/yO8NoznRq0897MLg0w
rndyWToPFzE0Gg13vkFoZATRWNAChPk64TGHF1OpF9V1sXFYX2B7QQk90yUbM/WC
hOHQWi7D6Cvwwi1ioR21a/sNb/Cx46RYcBVDnPB+3uJQvmH3KqtkmMzTbUwmwo9D
MLXeQfS4ndzrp1iV5ViM15sK2HlFqkbw8dbWgOOPLC2LJvADSPxLuj/NFt2hlO6N
YeWPEvutxsOXxCPU5pajdEVXvg6AxPPfwYP6wmzyVGynBpY/yWQvje6GMeS0RueG
K1NYIi5gNGzKFey+TX+/iosnsrBV/wxwF9Kd8ycEvA1utwGSCQm5DMT9hKq79/iR
7A0oOmcqrZE+bNPrXHfioA+kjm1BapfYN+ST4qWkmIXrlgeJKf14rUI+i4xe+zbo
qW8xz5YRHXwMIsuZMOZvsdY59cgW3TkYQG2zKYxKIErqCaAf3ut2/CeX2ekY8C/p
ff0+4trgvo+nTg4wsPgtzY9VaTa7civd76oO16OLfgx6gwKJzV0lbJP4MhJFWa7K
KKkcS2moJ1Kbqgk1Jno6//WWIRFzUvJS8gY365IqxqSytWGzsHk3suxepH8xoWRs
QaRSWw6vgOpvw9vEm2MoIkFrp93bFFQQ+RXKRiLCv2bLjSmbFMnmviTOw3kvGl+P
dYXSrasmuQpt1xNobnmduUm/QII45HfgVgTEyHWwd0Ob1BcpacvY6ebJ3TTP1ler
HBL6IjfxQmJxx3uhRlyCfwZiBbB2LF1GIm25VJohmAkbgq4fl0xleTFZwfeKTxMM
nGwf7es+foluoiNGhtfjsXpnrxnZbSRgs3UMg8Oo44vNzf4DzfEthkqDkfAw+w6L
1EdC6HcxfYBnSHh+ST4UloR00Cb0EXjXbz6dESh/LVniCk29eKk6cYr+wxJVrQ7X
FatErD1QpP8SsGsPtDEWECbABseY+nosOU9orU4yEYQylM5ee6a8wcIMEMYJuVTo
sgJbYU06Vcs0WccfFd/0f/lbwnKL1d+jok7SYCggGxMKmG+ngY21e5TwArBY1CJw
5iHjlSvK8NA2B6R0mowiAH+Lq2qsMCkWRWiypW2QgZ+i6pp4vXF1bwPH9Vu1d1z/
KvPSpP6Pz8m22H5FCQ0HL2fCwKGBckNZq1NutQfbwMRG7VQRwWZ+Akv8QDjkpYLp
IagYrGgNNhbCNN1Ehkvqxh7kvauApK0iSBNa3I4XEEcicmgmjUpShSr5yM58DBZa
uiRtCCLsVlzK4fRTlqEkyuvk5ZVgVGvOmppEf2q3DMJblZz1B4DyJWRF1t6BGibE
aj6NsZAz6hrO8rQ02jBUvO0kc1/v+4FeYxAIaHMBTBbkqYcdVa05XATuxPeVjU50
6x5+gY+yJbvfM08IdZ0QQ9fk3FGazv5hGAFZfvX27W0hnQjr/mR0zgza38tTJQnE
MZYBmwRQOfTehmF7wH1gHHfCzQpOEdbYoMZ2ky2mEKaGyowUoZquASb7cn0r8J0l
QuUNU0mg7lFQxhRcClVW8fvELd42yuocgCnh1ZcTE/Wp+h9vnuEfRsXq7Cn6uQny
JUWrM9E2ZuYL8RmM5wDJwxK2sGE6Kd0t06rSp3V813ToLrigRZd4AbAxhmcqxbc3
MqfpdssJhhbBHiJIqqjeXr+5xIOY4B0P4w+ow5N11tBsQs3J+j/vABYa2TO1xLzj
LAiHEuhWQbaJBg+l1ZHKJrhCe5cwLtBD5SzGUxePU9iLo+Vps3wTLTF1g9s9eFcN
puFYwDt1ruVn9XVbyOnZp3aM5yxmqZ3IKmmEOub+qDxEYfgFt/mhgI0c7ITLsTo5
h2U/zsRwbkNLoiphJQkBNGl7O4+WOUOtugl7YHZNvR3crHvH3om5+1sUBDRHtfdb
Tj66SiIr3y8bhr0fvGaI4FuVy8FZT/fxgi7QoRfpjHDnZ97umtAJ0snrKsoVCZu6
U2Qu+qOBg+8LecgXRL8fY2+RbOD1Ua0+/IAf7MIuY+PnKuAtwgbsS3gGEVTecI2T
xwocXbKOD758nC7aWrJtVMxl6XKRgZJWQTQ1ZtzbuajIc9hWWOZMaFc8D/4m+348
kLb7Fgl/TM2FqvTKj6psFDdQDZbIJ81lXiYlily2MtNx4LqNI1dmAhi5ZRmAy/T+
7T8AnT1X8PpwuUhNjSFbjJPjI1kYzQcmkwkXoIsnQKo/7QCVnfjbrAnfC0TmXAi+
b/z+b43GvZ38zjkCBxr83eWE5VWrnea6XB3DrguY+LEma+DIyibn0IDjuCTUcT9U
vaJmJEj1n/xpqdCnz8zG620auOKzhEj0Et2xGlUhv1MpkL8ETPsMJ3HMSzM5CAoB
3uJXwjNMAQYOZRUSwIsP3oep2dHNWY25Um01Qp6nCiPO8pHssviqBIemfITP6IJj
jIQIbIYUuSt0ocvcIaDGDYOpaPrGOF4qZB02jfasTyuwNsuOjD0CeuSEoo26cWn3
x2Hi4/Qgs57mmKC/DRfhfe604qSkAn+67rNQZcn5KbZDmTt/hHWFqwxSzTDmmQer
dr/ddb7KtUXNYNN6qc+eaSHn8N378kFxy/W7v/GUBT9YR/TEdXE3oO+hhVOYeIhH
NXRcrPCDk57U/Js5fZlnWt+bDmSbJRfOX6f+mw1M1E1x4aG5PF3Hyx0pJbmyrPMd
EyJROP9Z5v7Ygc0XmicQdLr1Sz5kbat8YCl7vQlJLYXeqtSr2FF5AOXhAsZxoLs2
pNZ3hutFlZNK/uzQgIKgyWUK9dXBWVGS2ukoZWZMESDhk1CDLZqy4Nrd0FhS6NjL
PmulnfOiUKOnZ6eHGw1B+PCBHZzgTIIyGRsBz/oPOcGZsOXyyM1hi8fbJIt0K3yR
MCaCiBcLp4SJT2SyzGOhmGM8EzseQ0fqkfq3pgDohGmthsQdG/82n/laiNHaBEt/
fP2aHnPTrP2w9rcXCmLkj42MQIaV61QfzjaPPgIsE473sN/UGwvTJdkr1Qrdmq5i
1k8QgM/pt64IIFERfT9Na82VI39u1jUlD/jq8k87fuviXtNrDuG41xS5C0GmIR6D
YWqJm6E2mgkrWoZHmYtsfTwJUlVAZjeV0+9leQ9ODMQDCMWNqVCXzcGaL6bG/u9+
9QsSAcd/PKgwdrz68MsfBUxdjgOIISGkcjN/Z6vfkmRgqgfxbCnUiXbwE+IfKB4a
uZUbabDwOCaiqc6ipxH4iVMP8XPrfRanFO2FQM5LmqtDo487KzjcsO6h6zqiX8sN
6Fbbww4enWxiCeJHjtdKm9CrR+M8wB7src9Fd3lhV1+257/oykdfRDqkBbOxbdCw
IwJwK4KmjwRMzhUWUNMCd5bAm2RP+kbtuRAWVcYVGgusm9fUJ6TwtDtLthF/c9HN
GGetgjozycrS5gNbiQSzNV0pqXBqNMsNgUUHTKXVXLpeDYKhl+efPuo2yaPJ8ZOa
MI/m2i/F+vDqwZFnm9F13KxMfdS0pVnmmqFF+55Z3yFQpFMWC2k8EGmPjhbvSx3U
A8t3vVCuZgu6nA1xsHrjdlhF+mq43Kt9TbsP6YTDHePUAq4WM7drEbmGZdEQ51ep
7r2ieSxQpVhWFGS4Dv8STiDQjKNERQCTiG5AenlkPGXjgaUmJsHRt088l6sIrBFI
h+VGOzO+K2C3x5BKOxJlfWKPZ1QQ6pkmw6DUXzYtMBFGP4Zneri/Yf+0eeME9vqH
tJ+ZgHJtoMhV4x8srCdn20t1Eq4V1JLlOSAnH05xispWurlEtnT58562OPxHqj+U
0Pe4ChxeHmrRJqsPxkFvtjdsCpFiCmjfZBbTzGMKo08jDpIVbHDAt3nDV4oaVQLM
2aZUuap+nUpQmkWb/h5uAQV1+oSTp73oESeQroI8f6jvfxNpp+8T8fD4cHbC+Mw4
ck6GbGxTIzjqLqK8SuKYkbRIRphp7slM8Fs7rPLIehW5a9M9qm2ARkKgK5mgtEa1
rPL0bPR9vKYCi/zRWvUooD2mF1OrVS40Sxjg8UZsGE5Mq700tiB6wmN0dEWFCLHx
u4mBfN4JDkNfxW+717AGKY1JGzh0f3HGTD05rll6YNQQUR/jiZNMkungeIn1/n1z
CdadA+ZrqhEWv4PnqA27NowxYkteSjNQYVDP9HF8xOVB62Qbd5jGVhojw6PBDyRd
kxDRCRi8T9fp6bRX23gls1Sj/6S/FhTKcTWBWw/Qg9GmNSkSFDlr+5731CoPxPzO
t2sc21IadV+bXhuCj3ERwQGYCwBmcIF3Ze2kC8v2F5qd8iwqX2Yq7g8mcPyEtof6
qcBJkUEcoNQIgfpSZsH/sImiwF0FMF2/TyU2WS8MtAsLRfZGOOuW0VnPSf5ezTtq
aKftfM99micehnJL7C0m4EnlLDBoG8XBIvMjxKTrLVdLjMvCHh8NnFhTtOsYQuQ0
r4nXHL9Zgquiostdv4Ua1jThpMRqzXExq746kP3Mfr6v9gVvoByDUPhk5RxNKqoh
3f0au4dzFTpsRp7fEg9lj9yE4tDtK3rrE9Hn0chbrb9g8dLW5fF3/BU3C0GDtpXm
EO0rF7wtQzO1ipIhY7BcT6ziTf+toTFB1nau6db4L77gsfAQzWjIBCzGp/pguPZd
cSU42y5L+BU0RKgtpZKV1UhhaavhYnhFhKgIZHYPuo6JqOwG5p8mEoexYVShxFT0
lTqZofq18FTWx8TcH43gMCSOK/XOEBeRq1kfdwg5WqrytRapRZlrIU6tFkO28WLw
Sez9ajLExjEljOUYk0rR03x6oHI25Lo0DgGCccm1EYglEZg3jSdQyYXFE9LUCOX2
IDwAixrmGh+NWZzJ0GyVRhzQcFQ00km5aBCbgvgUuYS8cXKhhxt3wP28HCDAa5t0
kC8ZpZ1TKOarVoIRb2HgD0/lHiusxoOwuWQ0klck9CXS+4rmV2jqyStNZ0UY6m/j
dwYBjVeIUjMUTsG8XKcL0aQ5oy3cBn+0OtFPkuHEeuCsrcdeTcxBJdCM9JayuEJk
GiM8iCSLbGvIK948zawTuLQ/8TnI3nofWWf+q9RUxwxgKdl4zJaSV/sS/QtMc5qj
eE7wMFc9XtD+f1ANraJLE/t03JJf4obx55DgbFy/FoKGNCEh9e3lx4NbvTBNr1ni
fDFcfDJbNkFQcpK5a7Rafqxb+kPRabsI6Mu8rnv0jVzTjzAtqACoLvvuxwWNNQ+b
WoGq9MDs4/Om/JcE0yLP/f1GXWpOR07/lbmap0lP6ZpVvXRGT4dR6tlybisUbeFg
dEuLlgFC8EljIh9qBVt24rciglrv/95kGAYDXWJFxdXPy7/2+V1d+Ln63757vXIM
zg26NbxoB+xhzD7Wb3Pr1ANa7hrglGbASW0eAI4dwEr03O+gtWDPMQleUtDjpMqK
Rar3nVOxshpOuNoRA4Vquy2gExtmNepLN1zZ6X9Nx/b963fz3h8L4E2ljWZryxVf
WS+ZxRblDkksSH1xJJW8H9qweokUn03o+VFKNUtNqQb8dcDydCxGUabccEadLSWe
kUOpYNwNsgf8/Lmh6jS7t5WQM8zaLIaeNe4rPRUEPZJtF6IjKIdPYd0/b5qJBi36
PuoyBjAJBSh8uOE5ng6Oa88H/r3yma7feyhymgmpdRnL09yo+iF1J/pNYfXj9BPo
8fxUVxpad8hIG0m4/snTXCfcjDNmIntwuRFCl2nwzMeH2ROO3eS12iLM+QiaPuhQ
sHZK8nmnBgbWdU+tq2LncMQVm6blno2CvWbXkbFA1HgWKRie9r7CUvVnQrsignSm
xRWiW3SytyHpK+3C+8fdiUXy7Wljm0Z2MgcYKbKSB64UBnA8TkBbmrxVg1rIQ99R
E4RDMOfPgKWUf+Hi25Zqa6r4yQNi/PW7g+0Hy/XVtdVWAYUmtWg3K6kanU8ddA18
hzCkSzfkruCryuXFm7nk2fVaykH2pbHj3QX2D01sO8T0W+41qdAYtF6jNJmH88Nv
G7tsvPO1aoCChEbcueYXxhx09bxnVlL+8f8HXDkasX6njE3zInIDlsrsRnklILwa
Ee0fO+dtKZEu/TBgUCxa1/dPKDJTvOIDnXiQhAbMZiVD0Ky7TmGwprs2R6Vf1fq5
PeKP4LdewrtWHa9t3PvM1fHYI/eWWAWcja356+Ttg9dmNqoQMq0IahPbVbScEw4q
jBoFQ5NVg//wIeI+Ux0Os5JHrHEvKtAA6fqX4MVppsTeq67IpNERma8NIzpXeZkf
UD3LhsJwU0BpreCjwka61h32t+6QribQxTPh1vTZQ6fuis3wSJR2wGHTvH9aFIFi
Sue1aYRR4mTHkxqtrKBRWJqA3grrIrgByQSMMP9By8lzoqJYw+WWVojnGu6ixz4M
pyJ6qe4Sfktn7hsnr7cH6QMSoAxQTpeOCEvCq8K2XQ0N3Gqd2buMZEC1uuG/wu0L
eegqPD0D5g7asjIYocCM2dE4SYV7p+pKFi40kdAWMBXFqHDXXu5bMiGb7wlLgf2M
ef7XEjKA6YpMnv61+7gYugvu1/Z8VQRjhesN5hk0t05iWWTMCOfFUjWUGp1ASUqV
no4FCnIRWiAWKigGbndohSos6dRyiIaDVsoVWa6ynZL/U9iGXZi7v6RPnijBYAfF
ZhIAaTDXSDfzFsSOQyPLMuOtnDzGGZFpGMLnwLPhNqQR4pSqpRCUDlCFILKxblnC
lkXd9l1hAx0bqV66dmreOu9Wm/bDeRJgxcYplx2zPAUo+nYrWP2mgZu18siFLW+T
53cDShxHrtZAASQPHAnlgb9XCD3cqkNLC2w6a9ZXG5ukxbIDzeGAjYmLTBWDwMXU
JnAQDmx+C/FonP4HbCNUZlr+/ZdQ1hi/4PwfAb3jejSiGEvQfdAKKnf4NN6NrvKy
uRubhm9c4hWN8u5aZayTXQy3MyPGroYkPQ46JixsbyBAjo/S/B0/ziU70vgwv0oM
XBv+zJFt6ot9cVvdtw0QbGznwb6jszmLqYbBeiIK5/O3VA6C2vVyEY8Sd5yk/9a1
VJNK6grTF1klwBsw7OMptM8OnG8//e7ObnS32dL1EWTTp+a2+C/lV+H7/d8Ude9l
As+dgDy/rN2huuOT8azQZdyTMGEDM2XZenxJLV6C6QlN5a9zwy59eCnzNg8/F14q
9h8QSLaZEU83J8D1l+lD/kYSo6gnQf/rj4CWAoMpU8dXqengaLhBgFhKyE7SPa74
tXm4Q2ac2ukwoWwg0rkHL9215cayaSKOSgF2qruDkhVS7e7Z3COi7Nk3wIEHvPDm
se4toqQ/dLAVdV3WZlogpiccYCXJ6NPJhB6abWCghK0L+f+0Akqw0CMC9nVC4qtI
dqTET3RkgR+4zHFLOt6G+mtuUBaFk+/isHO+NBzjvS8MVuCg+M3F/ulqFmupWK4a
WO8Wu39O37q7djQUoQFKfZDPf0PAHc739iELrFznO67M+i1VdytFH1QrEXMXpjzD
tMZu1iiePuMSBinqmmPfh9bnafh/5KPRhZgaE9IKzy5gYkfetC5oTVdsHCJ8tGVA
B1ddexbZ8/S1jrv/hreZoFPjn1pABEGKJnrobWEINzXf17Fsr0QJgnuD+dv2SvoB
KYY4/upODFvzKljCiZyjGD2PfCiujHX5tdaX5j2cCJ18a5conGYEiu9HssXnUIt1
pcxB9brtWw4JfMtHJLvwf9GWSOixHTIpzZao6g/luk0IZyxjV/XlTBe6yGckRTO8
gbUi8qTPVyZfktnuzp7CRSRiznglG5ZgZbErJJdBr3hJ20a2T+jYEaJ7Ox1MI3aI
ZSKe8adpO7YcYCiP1n1mAAejRnTPrPIDvZ2GLNBNnUKw6tVtqATLz1kvBIbANpzN
x9pBwJrfkH1BVIbkXSMtkYhhE7SvOhfzrOMDiIhBtxq1SGWZapTrMyCZj+Z23BOW
7JdxwC7qZmSZ2RAWZfHkTSfIVBt4+7m45D9Vfatj1tW+oRaTHCf0esaYxvU7dO0/
bs9LYsP+VR5eRkNelXdd2+NM1VHmy8QUOFxBizXh1l1Z2oiakYm37p1xCBrf1n1Y
lfqmKSp8JqVxUL6onvKASGobwdeN22TUevASermec4rPyIV5rJfJ1Jc4N61Hl6ji
mnoTjx5gcgZHdVFRBV46MUbhVw8+uYvZkjd33YU89Ya+XnsjPRQePL2348cah5Lr
fo6E6lNRftmesqrlZGKlwN5/cBLRGEcbZtECNOuVemv0UMDg6Y0omWtgfLdF9+aQ
Nwp1YA2NvfN/0NZN7NsOef1fOiuPAOPe1LUAB3+59uycLMPBC+Wvhu/4VK7Pc9oL
R772VlS2gDj+YJpNSA69srpCUCDnXzYHLCyfP9/TmBTJzwDqWPDJHa/UBY051TTI
UxRsLBXTw+wRqOa96HENvNeW+CNrKtTSVS+4WAJejYABNtoBCLE3cV83z5mP7/AM
EUAo3a9Rls3O6yHMcC7Ic6FEx6KdBx0mQlbzllgPUECtkZJ1r9D81+cxF2SGerZU
QDkCsnKcz8+guCJMDQx9VMjkfLb9+LmJ3KP4aoHjtHDgm1roOujQRAdxj8elDnS4
uDen9EZ2ddmrlZTbpgNYgZgmV4J2hBB/sP9H2LWjHRWzqPrIIXMYeEG/75TS8hu1
ZNw4gz3jFvWOJ3K2fxOyAgX//UQ8YduP56O31GaGkHB+znNKLj31puaZjhApzsQk
xMZPqxjzjbc1jqN/VIlLRWAQ7qR3P8RM6hG+KSowUpDLvdx7nHdqBI9a1+xFgoOk
zti/bxxpw9z2+LdrirSi5179osCWS7ACrmt+xjfIeHxtuQ4ITlP9Oqw1V2A0e2O5
nkpHeZMtkWWfTX81IxVWyKRX1PdjbIw1z+p9zAKzb1soYhuRIs6IlAZ0M3mppTxC
vTfZVROCrenGgBzVZHbJ/4YVvwulDvJcm7Qh9oB6NLpntwl17nHfJs5o1zCq+RVo
XAWVwgoW3Id28fLsBTUaGpRFedS8cxEa/Cz00HKYMhGpqOH+ILDRnZPloXVFloO5
H3bUmE/YwZCKlCc3z2WkBJbpR1Aeyit2ZJGBH19cATReUABfzGsGem63E0QMDZKh
bvKILFqeRsb1hoY07p58aBo5RFsJZGTb2i8eoXAjmaBVc+lzed2FaCLljpeY1tBm
3Ep+dc9VGOE2vC/5/CcxRFZO8no8/8HHbeupd/QNENVMjX82zSw3kFO2zqFYVh0s
rqqY4hq2IwmnJfHkiSsADH+EsqZAHCq/3MPkEX/17SjU8JfBtaCdkiK3hDI2uPKO
1UBVFQJ24XRFsn5ZPhGwwljAj9XrUMAsVI/ZQhcDuh8QeFKdxyYImCICVnd7LwTl
d0lrwKc77OZRzRUvEWSUGqqVDzLWZB6sNVopkoVY/ZCq454duA1K0NDozpaUgLt5
3ZXuaZScv02aJa+GjITu0Jnr2SQn+ziWov+lD+Cu9EvCAtb5Q2d8ZDpSxWSSlbWb
bUnttr09kOWTetEuGBNU5bTdjBSi5mGozFxQ4APPCGnyqAdWA6R3P2jI+bznyXa2
jkzBMu74GM3MxIbgrjzc3C0DSiOthnGCmGdWYhLlpNDmMDg3MzOKgFdlAK3FFAVh
txOOL8MeHCgeBlvxs3ixxsoR3rtE4gR+7AWh/knCbXwNrHBX841/iHTmTYIjUz7B
gvqUP31URZoN+TYtaGbIE8+i5+YBMMusFZF88EJe5EBn+ZcsxVlIQOkezX9MFL73
Lae30Dk3AORWLWqU1C1ve3OzU8kFnTD4+sofLOM7XTixS2DtLg7pMNJyK+QA2Du7
9E/yJNsCVtVnKYmgnRMvAjg2lNUq10Q1PhB+JmXUFzB/5zLbXzGIdkXNHXa3LRUC
r5aC37NmLQQZD/L1vvnFPq7+C8xeMjYwAX6xrjOLKVWE74grGxbtLpjQXp/3Z9l5
4ApiXvULVgyrg6c/+vFmE96iXP1GHzGxDTDe0hMPHPpVPrHMLBfZsPVf0vdb/yRX
gHojEZTHNFl2o1XegYF9sfwA/Bbc8ifpRiV222elxRJ/t/SEKjauCU5XYsMbM57W
Mb3y0j1k/5ZzE/52Aw1AVe/ooUqIF9GwlcAbLdDtoIh0CmVO1yfg5W+8KXYE+vUb
GEWuEBbVSxsv0EgmLewTVaDhf3w8EkT+oO3M0Mtn4oJ6T2SlWCOaMc2Q9y2dAoDT
2dhDJ1A9jItjXYJAd2ogo1UkG+Qi/as+hw62WXoQVMiIh3lsu+ZzYtuCpderyhsA
nXmwN7NWih1tgEf+bAzIhOkavI76dV7aR72UMVYSappGUdSmPB9nfCApb2gghzZ5
enDzka/fTUgcyfEzc/jWS7cUK/qU8a8+d3+xhdW/BM2oyLrl9Qvu2tD+2rcS+Pua
Y9AouoApfoHu2j2bLuBYgfBkwM0UhUAZZpG2BiuxbU0cATIKwTvYet+sV995jW45
An5rzre7iQvro2B1jRTLa/5GAolmAR90h5l1TrxUEkOPC+B6pkf0Fdg5QCSQ/BKg
AtM4X/wm+ZC7vTpdUEBmzRcVOuCo2GrWxfOJ2PJpjf4VG9dA3ydXf01kLClHN99I
MgiD/x2FjGj+9yce56gLPt2fMQ5s0aNWJ435iZgjPQvHo/r/5T7JY9D4MOcdFya/
UoUEoxO3S0a1hEGLBN/VCZ23nnG6E7D4jZ3yANHRZNNe3JceoEH+JmYV8SPNGCmm
O7MtqN9zLPgltqHUGO4gXZYYPKEeD6bNpEWalEa7cQ/zE/yDSvNu17btvxrRG7bU
jOLVxeJxpV5W447qcIeG/FS+jsCkbsf4tbxmf/zlXYwtcEFeowa/xgvs7dES2wyk
e0NkUKiaH7vklit296ZtM7rkwVPWosaq2+0iLtNWHhfDPAd/TL57KmoftuFZIBL0
WvP882Cpkjy9LYaUvbIgo1MSBAN+sMkwhI270OeBxVByXnXLGbwVxRvDPbhXUBX8
5X/+2oSNzdAcxKXflRa8X2j5dxsumGKP1/xiKEKgG3bp4TBbHOnw8/N0cjoVHnIu
FrbLKkuji3thxPxgYUKjLQl6RgYw6kWIXrj80C5w+07ItO7D42ItJPGb3T5l3W35
eb0ojSGV+rI6rzP7siVQiPo3Bn/Pv9On+p1PXNo8LTRwbsECLLaTwFwlo7iuBmDb
wSOxEf0pkvR042aUAkpzdKz6mTDRMId9YKe+Qgg0HQkGPu1zG2LCPbbX/f9KIEqn
HrCt5TRbWNKvMDggkRhPcHcxdI7W0mruEPEyYTqMH2PY+uzv34RBSVOfMOxYH6Of
GWb/lSdkq6Lmvjw350JZ9cgIzyfg9MAjj3+NH8qaV9fTt1zLxmisS2NrqYyxAcZB
8oqoOoP8gJO+kANwmXHbN+t5wpUIvKAGbwRZUCwnXbsoBdJ0VYI/E594UtB1g1tC
+RGTyDcJpKEYM1HkvBjDsWUFLfdPFcPMWK3LI6Ns34Xq8pDD/NEdZfqtNAL3cLE5
3lp0YuBi5bNnTeT4BgLjvXshFzlZAk6dOmvTY6h2hpRQGpmm0c0oOmM/Luna+9Oo
sEPIW+AiFFIUBKIsLNxg/BI3GmA2VGr6qEIqPlAUSfhQEg6CotrdkJNB3nSso3io
nVW7lSzy4fcC/XvIuRY2B98MWe1F+S3x/xORUFnehPhTYC3wIPOzTdarKOrqmuS1
PB+Hrv5DK/TzbbNH/Fz5h4jzEQO/5fBOFfhrVX7Nmgr1ZQukKNUhQV897g5EFqmF
Z88tKmiWoupM6ATcp31iCHbbzTCLEqAgKbMJt9B2lfUhTaF3bRJ2Qf6G/3pcMr2F
1dcP+3P7rBCm16UuMBN5y3OKa684Ff/nkeobqnyjAR4EMUpBVZcOsFZ+oJdZbJ9F
roMDoxqgXAoTovVd7OTUnOq91nIwbnzh5EbxNLpq/JRCl8nAkJ9GouhBTT4+kT2P
AuelBvZmvsG9gSCVo6VBNode446zdY2XNFlRIc+GrKpKEKqsSHxa0/ByzFgxJ254
UasGAg4AcroCZqaOvCApbCiRFFt2M88pe7fiXbhulQP7gV/fUUTXJ2oFBGFfNEKU
OmHstJyfzegpeBusnIywVg5n5Kr6tksA4u/rZ4/U4+FVHSF+Eg61TvKEaOcXl+KL
O5o/m6iiCCf7P5azVHNHxU4bqPb6Bh36qOjvvqUbTMWEKyaM10N/PYGAWsbseaq6
nWPNOZKB/OupyAYuZc3m9vwJlAiEb6s0nJewJAEcOT3I1U1eagmMxOM/c7nmaD7o
aLsWRs1YBE+/VZeSXY/2k1qU5AHKZT4ScZPU1pMdANWH92XrIEm5+y7Si2Pjkm6Y
edF4+O4KPlyzVu7uNZi1JUTxfg72SC234sLlNpPrgfi3Mru5ptfJNqqBm43xWQvT
i3dnthvxNFySRHCJ1D07c+MoAk5PX/E3dusACduuKjjg4F6rPunxWQRNO8ALWZlu
NM7MkJFK+oQdL4gx2eA5ZqqZOkTKvDbYPCCPOTziMys/mI1I3rNhUB8d2Kja3QZb
EnfpOxoCiGDuGe6kh2UyZ9zcGf9kco+h+C1qeVS2cJZ6hGhFvKM6zzrMofzTRGyc
uEvENUtRiCzyD1zBWCAC+E8iwqx8FMgDH0zb9XOfeamQEZqxpuypBaM9JRhe5SEx
SLm3f7TjygkMehTzuTphGsijeFMIpM2ZLw/sFqQt1Dpf4wHOEwuXRT7j+SByLiAw
UwOn91SXmoPdv+mzyqIfn8MMfz9CJPbC9QW4TK53I3WMRoFABrGaJfOtwVjMl284
D6hYWPN7CZjrz3KYpbYBxs9A2wP4Zihdk5xLOU+cWSRKjBt4zUSFv3T2imuoCOnM
FmwUCWU+qlYv8sJscbL1V24DFT8xBjhAhBOzbWVBTftNYLOMCLNq4Ct2yNSJR4xt
eSKvn9l8wg41XSLhv1fRUaxl7bTD10Fldp0oJXZTYclR7AfM+ajS7/6yMPVFdJmI
+/dvtgBfWvw+iS1hvmMFl4evptUVx9kjdgZBkMgF1KgmZCWOOm2EUi61wCGlVHw3
o2ntfdhqv88elZZ1srrDXIS729lImkMXZb7QtrASzRxtWb9m2h39CNrp5Xo/xIbr
hR77sMDeMc0vKpD0P5Zb00brg00uTYqNd2WqJAzhsOP/SKtznL2p7EeNXVuFcJtT
kJxa2t5xQe6s5Sq7KdZkpWst80sSv5VbrnZaVVkWEw+RcsPC71vWuo6POMCBXgTT
NTUKTLTfyKkyg7BhMYJZFvzUKOGPB4fpzD9oRMH9bTkszsNT2pSvH3dxDAZEoLxT
kNsfKFe6g/TRW9fRR2aV7xWJurF1N/K5YJ5MgJ1TlAwJgmhFYZiPK882iXhmFZ94
YCDvMuQMehVEEAPkZpR2QJKRO3Bbx3m8VDblZhWa9zCNVBUqinCiNgdgT6UdxFKW
nt7JWj4z8XHGNjUvd0fQalaDvYUWahxpFG3pyjPhp4DZL0dZP6kbAaBcZItG/LcD
G5vRILwyJbxX3LRaQV3jxaHbI0rz1ReY0XBJquRKpGXa4JHGwlOGqEe1KYpLcs8O
sLGdRhO2Ffm80zrYQrda9Lo2oi2zwAh9NtroJ6aDs+yBDVDVv7lI0EP6d8c0/ik2
WL3fSFUbCuocWwGruzA/0rFThYk0hbQh492WYFZvFfkHEP+Cv2OLoAdb+c3qJ+tP
hsstdArER4IgVPvoEK8bXG8gIHipg/QPh6+rCVnxaN8vJyPM8Bp0MT5mbQuPIRf2
eoBDnNy3u8F4Mxn4KiegcjexqLF2qQFce3NupS6yAl6UVCqnRhU+fEgd3h3VNftk
phrYO5ekikhiZaWUMwd3JqnS1dMyV2Ua9TkIZTZ7Hxy9faTOIvvve6qcGWcqWMfT
ZbsLL//ZulSZ6TYn4Ie0N1iIPb8vXM9yT1rKyurhFhDThyBoRphvN+RycBKhAWg5
oaB6oZoeknuxpz+KgbYy4I3puL1hwm4W956aFOvXxXYtx1Mf61CwEbstIwCpVSb5
2W9AkQNVW6bhQgV4LS/qdfFSIMU2ug/H0SlgBolyNpXzV1uy+ASwsephwUXZysxn
oWGgfdS6uodTs2lo+XPuqud76APWa16H0wp9CUzsPTI/V/cCkKgrJfP0YHardhnE
IY2172vfJwvqgZPEhTmJVT+Ydndi0tEGrUOPMtu2UALIuJ6cnnTEFnsiZBRcM5Jh
ehDyGCdJk6nqQqU5LixkmoF3TQnOCPK7XnIFXcB0kePfB/ao7FNCuroW6jb0h5Iu
rzVte8awMOYvp1g18fUgFkqootLFPmtQgvxVHkjP0aRHsZHecdpVfSD/jpVoQjs7
bL6gPIsqeI3FeGiqZvqx2Fm8LeN05yEaYfaCosAaR9hyHIuPt8GQHlE63BUeHpPr
EPfxKDc9S7itNknulH3j839Vw44K+6d94I4AbykBK/n0oyfc1PjdZxgER6TiaOOP
g6bUFIdNOxIOo8xf4wb0gX1Z3uQoFP6x8yzDZHaCEuHvlzPfLGcGD7ws3Jis3bxK
wFb6Pf6KDeXJWKC7PfTGV4stnGTWn3ZQhv8vNgB5NWn/kC6uWPC/15iYuZh/X9yg
OBdFGLfCZVby2lVJ8JLXkDQ5KaaxArPaLph5qKEXdDvy0OyCn/kCdUl5JTRc8nsZ
lWfHLE3vtWggqVK4Px5Ot/kRUqO4k4kosxA7Xx4mccgOsF6UqF3pusuDd8y6U7Cd
d2gQhMpymlt7cuJO2SrdMQp7Hck61fguUeEdsnknWKkzAK4uYf6Qz/fttfvfUQAU
DEUJGGfavgaSQo94ojUnTWVvwPU9oTVE0pAwdUWOObW7249pviYz6XX83JQ9tccm
GhoulMqZhofjDJMYfv2NvGalSOCrRrIR16hIerPNJwADV7od7SopQd/gaIHTjJLB
PyCr66dcbILBthfAiZXlYEp+pbrcUVutMfvjBKS6UhdpRr9gxmIMeQoAgrtvT4QW
lbzM9fEKRek0FFyCt8uZGQK0VNyvh1WuexmkJHGa3EBYQu8xsBN8wbq3TNGSeFP0
N1qtuzLIyjzQMMEzUMdeuaLxLSUzmAN651ncuBQICo9I99FXVnObvvFB8f033rGu
ymt/9XniWT/5d4VuHXf4S3aZ1yIixcXi3MkBZ10lOvdgsEgwf3q8bFvRfgOilrMr
1kSoyluq8R2L0vseQKXxdQTvX+OLaAOrU2zaFIMyl8Y4VXU4Y6XG1uq39V4TWQjS
UjZnMLpuZ10N7w+nlYCHg7TOQGLbwPmWxqNMvlgQqrMZxKzSNCdHWUAdHzSZm7k+
FPf/koWQazZdTsqd69qBXkhJiUToEYEtRM2odFJrmqcvqtPuf0Go8dpFh80Vgg/6
mOYaI8Sn0h07i8z2o0XJf+GOiBBVhEcLgQUukIiYM161AyWELBvUS19xAuePZ55V
J+Ui38cOwpUBH25XjmDr8BYHmFG2SfFMFQnn+YJnUe9AeCs7jMNcn+uUYw5LGcp/
8F0jpOYnIeW6i5cV06H1spakyvrtkQxs8tijn2pz5T14s3ttVK39USl6b2DJGNly
4UEShliyfFsVzj7c5J0uZgIrPDj5dTKfDE1f6SksEzIKG8I10aVuR2HAeEmszmFx
/c7i3pS0SrfqL3utxtLr3S3diRerZLOCsiRSWk+2dIgNZscVyKyoniU4AXwQ+kpx
nPqxFyL0NEQF/lK2Bz59I+Bmo2LfTTtU32wo3WomYvYkWF4iczTf8d9FU1vU6gWs
AMv9GOcEezL5SjL6bLxwi0vvUp6KFOWrRjszp6TdeFFemKtdUZBP6SEJQTkPQmbI
AZRRRISFsb2bCnMstC7ORgCGpEEKGfB/oXSnzWrMNuN0OGQR+2i78m3LejjxegH7
m8tkwB8uDzRStBV1KHb/pAihMSYvyz3gBlpLlP4GGbKJOiVdHhOM7wz+uVdFLSlv
wZ95Dkh9ul+RF3RlerPik3HSLYACB9dNEfCX+AqtfVWaHpLPr6yTve0dD99KMSf0
GZagxZFu+RTRC3kQGPh8B83gssVqE8EY9D91fH5p8XeNwy19Tzi/cuE2sviiSn78
Q6hTt45jcCGTa5w26MuApDsUJL6L/4MRSEcA2n/zl+60JE0mM4rX52/TwIO+XJGA
c03UWQtYZuDZrKhTI4fgQSZjOvCOhobUqh4ZGIewf3T2uEczlYV0BUMvPZwecWP6
0mPcjjcgwH9SytvkNB4WNeupbonTTQe2iv3nTQ3jBMowsSj/saCy0DdiU7aaDx66
v2TBfnibZAvB9ve21nsGcJKkrIsoZfjku6yNUrtKvcJWN5o9esJfpSCRewGhwh9/
E2nKkPjdNS/+/wCENjWB3iZw+AQqn/p6dcVkbGby+G+VhR3iSz9lZ09zLsOY6tIq
5oUtKPsYKl1Xk+JzVI9ujwVjILcLIYaIV9ZxO1jEU7NvVY1Z/oSc3vOCT1UfGUyY
4CLmH0GhUPgVxHxx7z1+2XtUf/bHgOHW8od32h48ZphUgqYGi7De6hKlwyDjCaCN
OhQYHUirFrF8aNrvGkx2yMYX2t2yk6i4MHLOUN0Ke9t9erPqZsgGLZELjkC+CyUg
QHZJBBjFoj/mqaPAHSOhn7ZxtOoJKR+8v2mu/44zkpUZuZQ/Pm/dEcgvt5VwHUyq
KmcTF+k01vOhyq4pXYZhx/L/DlrJvn7znkcd5sOER4Jglm7k4F2S6RKRca+aGqHI
BcUzf/zwdJVWh8RS/P78IjeLi21c9a4OCIXtuzqN16SWgX+GhuWRj+XkY9HEcYSz
hsmRJWAFHyuQpNu5o79mGtz+SMEgpU35TiRZXubQkI9NMHTGH/V3GOM2Hvl7B6bN
yTtOu4lOGNsqa3i1l2iRaBsAGMNW/w/6Jx+YI2Sqe47+mXH62QGtAleaf7ORA4lB
rhF65NiVxTUsetCc1fV45UwasrJqj/IqRaAdEmo14sDo1Ui4/ATlP7VhD6t+nUuP
Cbgrw7RaaI1YaYhaoArL/OsYPlWrWvN4DtGy6jDqEpQQQql3rf5P/MJsPO9SPIXn
UDjI0ktEHYkzs063f1t9WCpLK3IzhuDpSfsorMoD9sWoP5w94eXF7HnY7JiIQnTz
wB1dbLqnMjxzTDJJQ+5M9eDDlrsKii9/7vcjdRPwZz6dyn7hob5M7avKE7AWzaba
j9ji+FbXODUDvd1oeBPZM3nw2HWTOsov3zx2cDdIqEY1aOvVyW3SEqDGEMutboct
tFxFRSNNn9zIjhvANFrRTrNDCCv7YjWZQmpZaByEumK1+ZJvbX0J/nL41P0XyZfL
pxpSkMm5LYcMYBdwDAwooprnh3b86Kn8j2zo07qgu5WL0ag0MBuAgGjvI/dNXL4f
cFBNCCgl05Uqxr3SIywIfYN6Tf1bwumAkQ8nQWoGfbe91LNPAGkAWZ47TCJ2Z8NN
6ZgU8TLzByNbQO6OVo9x7oInmH2d7wG58j0rjsvxKuJguS6k23bANzKyp04hO0Ee
F6Xz1Mbt5HEItJByOoU0oAaQNkU3uilP+OxPz550N9LVCStecTV3luY2gmAh3ht1
CS6nOP28W6NtbOPvWUIrX7kZdptuAmASP8AX75nHisrNSHJyfRKR3h18cBnfIzrT
TiA4q2/3lb9HURrtc6cxwvq7l2rHAZxVTUhxZEHUFCUIWtkcbcdhX5/H+O1iP4K1
L69CHNI2pr90JLbK+0Y/zcrdTTZ0KuxIRfP3CnUCswrb+13X5r1QufxxpvdpfT7S
fu+oOWYF0/6+A4OLOipEd3nWpjfR0i4qv1GOPnv5Q6aaqFcB/nWmfhY1sQTzTpAZ
1JoRg1yZREqdex10Q3icDTTaELt+Rgo6pXri8sUDsbv4q/FHGVWqeepxg1fPQ6kb
6sd8gPMNvqg681DNPO/Bw9TrK7HPcjJu8TZNRkCBfkBXriBL+9Sv2mbn4Fk5GHX2
COXLhYvPWGMgRLgYjf/zfXgQt9p4Jvb5gAXqcQY3sbS1n6PoeTRhdSbOz/wIZmMW
/FqSqV7rJOnd66D/46hB+t91+bNBLwSGIP9QmWULvsCpQF7vMtJiIxzfncVLyxjS
nk9qUV/kc92AOpyyx3Gue1Xs1F9hNuDf1jQLLQc+428j+nLlsoMs+sYUZHBFw+t1
gr5/DtRsEWSIoMISP24GJsPwYhjS+2jhSWSc0ibxbo2tdk1PFgxL7Jo6IS5PNbQ1
SzZZxk7BzRVTiizi1gjfGdDF8vYifdyLwSKCG1kNfVw7hXMhnQNMp7JrdYrHJeyc
DFb7PPy0G/CNAz9Q1KrP4cInTtUNFcRHZxRIRDKytRSebPojpXMHWxhxzrYsn1jd
53mTjPjsAsI8maoCcmkyXR1VSLX8JEt1R/L0cMQscbuMQC7OkR/6mx2M1Q0BD+mr
smA8mGu4CpxXKKB0uA+fYKkVglEnJ4mVEZ1OAs4sSW835DWfbu2JkTjCst+hXEi9
h01myPX5Ajp2gnOFk+BkADfg1D3uUm19ELfCh7zlod85nXI7eStgZMEcedPcl6w5
e55+e3kjAE8YmDPzwqaeU8ppbWMwxWYLc91DDOjYOetHWOilGXw/2/hH+dr9wtea
WnE0DpzLv+znO5lZrL6b6XORncHSVQvxvf+/BMZDqvT2xCWOmdDPot5qLADiJDIN
lCm8jnieH78DcTtm9Vhhm1JfXjzUJJ+AIeFpwo+KPbH/rTGK5MWYXnmhWg0rPw6w
RIgEJpPEtqamyYuiLtG+JDMv6UUuiyUX3d6ab2vPYMhm3VXKaU3fv9KJ59vO2A4L
r+85UoK7TaDLAKO5LdS4KpnIiIWzFPziGuu+yWurDO7Ar/koY4C+ZI3ptHsk5qy6
otedAeRIyka8AEVuCVfSj3ufgRSF5ysJNRTXn1m012NZ0YMudmuhK2C1oxQrTnZC
6AkcgrAwb1+d0pO6nJ0iaBd1czWJZJDdsoUgukszCEb26uSKVazUaDsN5HbpzJES
DU2wKKVSyJCpZN5RAu1Vs7dP03gB2SIJQKcM7ni1uLt/7zAZPqL9F+8cCrWAu3tK
+QGbTTK29C7PCaLrtO4rUwru8Z0TlNWt6YwmFF7N+Nfup9jt4RE+fCziwzMYe8Oi
ao/vB3aKco6Xib33i+wgzgmDjhmjReZOR5obMjDsjw9gbkHEt17eOX9X5AMvN67p
+Lj+WUQkKviodruUNqev22/Ye61Qt0pkMIDMEmsq7phkQdrWsnk+zq1VaKL4Mx1w
5CBaplcKGr5LUpa9dnCmtUGV8ZJSFo5SHM867uuJgZSbiTjp83mGzh76ZPmpj3PM
mgx4LRXvNXOdv9ZTv2GB/pxtSnre5KpnXLLgN2YpvknIKKylQgGN2lYkHosivUCb
H1hMCfFBL8ZBZcY12WVh+fHFxW0wExLVUhv2rJGoa4rVrfIsIOSxqt/2DPoBZoJl
eVHsz5HzzTr3sjVJwxcqB2Ghqk4CaL4OoIIfd4OgluhRdjQ/j2zOT6xuXWGTXdAn
yeHhh/5yVO24KcKSRDLY4j5SzzBK13XHWUObhU47JK0sHF6KcxPA9lrfJ1aMmOw1
KSojWJm418gKN1HvcEdvxOfzp6FiM6J6sXcULjV07HbuabF4yMbNat8LXc42Vriu
ZN8yvHG9w6UdUcBO4u2Hz4252G41oUSfD2XGUnHYxlzqxD2hmjFTN2YgX027xmUr
EFAC29y0LjsCusRW6v/tybS1qMYChIjnvfC6G9W4Zh8r/5V8r7IPmwhoJuVDRvwR
wgXi25BG6OJeKpEvHMf/3KpBOZUrywD1lWOG0HGBKNahKu/esiErNnn1SAA1xP1a
QO+OCDnrQ6nFevak0VUR6csjboM5XfjiMWID+BPzccs4wbaaOoEVDkPIG8DW1v1p
n6cUJz0cSROnTOohnQGrkFgiknn/OJgZSdj8g3UFxL8zuK2haP3Mol6wdeZXWhO1
jaDz0agjkQGNEW9fXNsm4DW9YbQ0Zy/JYH0J6/hMVkLGBf/ahhrzl7AFdejUEO8O
1e6WDygxQ67hL4p43O5OWVNnX9tNHLpj9FKWWSfK728gMGPL03nGkP7pwspc2Xbu
BnCanPCEcqxmB/ibwxr53D+q0+6qI81Y9n56GqI/GG1wFz0YUbBtLrRCUiYDyufK
Z4baPaYmXrhu8bvWqZtgUde9nkYDocxKep9qio3nR8NOWKa0lDd3SaHjHp9n++Kv
z4tbFtGJMMcaF8LfWKny9La7HEbdyI6eEjzsy8F/culncEQoPCr9FO4RngQzL/OW
3EQJHR5dRDj2nk749TaJdJk3HDLSCVX9UhKX2HPn+O1FR9cyJd3Vs5oyyATuWGWt
E0+jBXF/eRPEUmuMT+ChvdtZsLSShkujFC6xIZt6trouOVskGZC9PDhmRBYmwYMh
ODXHfZGpvAAX4GYakz/JPl/pmhBGHxQyMagDbCpaiLXUG6Wpq8AG638UzfBYFduu
kA7RqgjftFqGaV5SXiC3HPMI+30R2F8UH9Gtc4AesVCtRgy6Z5wdWzGYPuNM1K+s
vOLQe0LGJyGhjbYZtCLO+QW2YWOCgrBD+q1V+/jFmlXFMdRaHEjXMjg7Jawy53ky
CWPigRBuRPwYq9ZApbQeMB3Npt74QkUSLa53Ww3xMjtugMi8XR2wbcAze0DAnbF0
BJ2HE+HK8BK/9/u9zr9hjL0gJyXofABHnuVCrBgt0qWgoYUT/AY2C7xPUJzBSfxr
I3fhicta9KSCij3f9LWmkiocKDX4NRc67tKBj8fMi+XBqRdCDDp5raC4m7d+flg3
kBu86XrQEEvrTRz4wwCgD3JkLKsIIrLeAnm53popoPQCzxbUFICcZYfgRmeVaZww
5M76bVL09DxwJULFL/eYHl8hECyTtymiTNd8WLTM7fvFP/8+kWXJoeU8LGIEOfr7
Ks4+aYJdtnuNDbvvKPOyZaQJMdHWSwE+gT4CuLFf4fjU6oFl860+6+qxQt9PWbpq
7vrJeGO2RAnqLn9oEMIhJzX2wIotueFAe+c10WWeshUiXTuFXTgB9E+YXuEuVBMd
g1bSlbE4O3dW92yDoyo/2gBBv6todWu/mOpPjo5mbVXfn6eX6Knl8UXAJ6Da9F0c
5+yQw8s/F0H4kIy+ck1ZyIH5yXavISnwGgjN7RVvSvH80nqg779A3rlLlSCTX1Uy
VKkt0tqxyF4s9wWtV7jSBezaX2IOJCfbZ8fG6iXoIqJHTBJqCMQVau3LdZKogLPW
9PDuTZhhkdQyogKs6wY7cX4fk5k5Oibu0TO5boQxMb/5PcsaKkSwdIAk22YwlwGo
EEduoY8569b2kAbKKU0Mycz1cBPqTzyDDrThnV+3BKxVR4c8eRJZQqC46l0X2K8i
mkEyoJaXXgMXZM8+4T13xuATthFghzc7oj2abG4L1DNVYjD7udjfLva+04wW8WkF
6EqSFSzm6YR5yvjfzs2gW52DWI9e1Krebs+pfwDrXhjy5iDGh+FGkGanvYmn3Cn3
sQFnZlKB6NbXlp4ttENTVOxOdnfgQ/YSmuBpawRxk3uWW/peXDIrzxs8Xcjr3OXo
+rZzw3wkIicnBCDMcTTbxxSMS1+8VhlAhYSU3Jd8/CG9gNaonn38rX/JkWQeRa81
dYxD8hazjbHowv32UzBrwYgtAaefsCvc6vMmzhER0+sJv7bCjELV7NX4T1uSZiKN
9IvX5xbPI27XP8lv3go9UHhAIlR2ApNWvFgvBUFtgF/zD+nW9UoWxgwKdd6GMyZn
0uQ7YnGEO9DCE5IdaW0r468EkNTU4/g8Ku37f0x88vMfaVQ6HDFgq00wenHbbWcE
cTwxWpIDpDnJCb2uklDqi0ewApZXQVsl1B1LcyGhppEk1HSC1i6jNXNFBekW1ZaA
fIje7pki2sHXLu5GoyU9MaGPvsjVz1Z1jjbm1fd4gIbXloRxeus2Tb99tFd8jm+P
71oTpQY8e6eiGvjYa1p0WQDvQKDW3+NH1xEdwQ5lNeRsTWie27YGeLzvyf1xtt2k
yk7GZyFCHVFbC4JJ56mt2xzg4iewWrZHAxvpVfd6m8NU8qIvEktHsQd+LiCsqjfP
mBkzFiyzqeBVJg4Nmd9pYAyCtVn1ZucPYsEGMir/6iZPe1mmckNeBu239eXTV43g
EnvnTipxGdJVFhVm73MXAPcdgAIwKDYITua1UX5TcovvJNUOZXfWE3rkUq2jyGCv
ZW4lgFH7D6IhWYS/yl9m+NAWEw+lGUGZgJifCMRLZpAy/5aoEyBEp/eQDz6Jv3Fg
/+GWv0IvGFQ7kglrhCq18BPFwXQElJi3KqwH32q41Zv+egqiWXfDNRFNCC0WlFl8
wjtOxqok9RrixrUsMggdxFP2E0ITjTONruEF82UFvCdAAaDJSBk8c0fbSCUTeGrF
rLA8c5L8ox+mRWv/p7a+LiR2GznYuVGowscqxOrVl1Qxm6FYe5g10xhPAQEk6q5p
q+LFESh25P1y5McIfw3gPr8DR6KXPIbDqcBGj3gs31SQ7flonW3Gary+j7qtPD4x
fpVJHqK6jL7kWFQWarabLCtU3Ik/Dgsc+L9P96rTjzwIKPeSCPf8xJTsDx9L3Ous
7qieaen5DWPWCbQEzDzwAlhtR3IBs8sP4y2X3f6nfloiRIa6ZErBbhfQAbLLjs0I
BgbcqQBSDAKIU/ZEzTRNxnakkAWbnFid/vHeqSUG3+0K/C7bdyz6aMlgCuUCOaEz
sCxkhAmgkT5squE02OZ1PcjQkcq99rNLQeN1jzynVlqNsI7G2uz82rrN/NM0YPOZ
gICSY4vDUlnFuAMlLod2Dmj1JCX1VkGfdXQB6Co1aadLnvatcBt4wMwbvSBMmq0O
SNfmRtoGLM2So5B7IAczWUcAWJ3gUUlYTL5rX2176e35Vy8edqcucm79R+ucmiwM
q8z4yzeMDhmV2VxGWMd9saxkVNDxiCJdpO8Cgmo54vTh6gOz5CIK/pN/LnqGU7j8
C2UQJLQvTMVHjblQ8ysujcSWH/z6Jm14htFm4i67jO+ACczXsSajUQSjBYjrIQfD
7slhuIqdvdBK4i9rmWaxpJ7qCXUoP8iT1LtYRPjW3tgd0xqd9QF/+C+dPPwy93zu
SBl7xiWXD+0A0e/fDfiaAY3KDxC8ZP6vR35S1OK2zDGIs6q75YU2+FfCkb+1bjbT
iy45+E5c0nme0+v5TFGamP6dSu/OubnHy3M9dwyvHg74+K/wghVB8e5SBxfYxsFq
gFY7kJ4p5cDqCVgiNqcoOMogcV1ItCEBBgW1drZA12yhFQnE5YbeZuG+7HvdFom+
/1ej1uKugl3m9ZXHR1sjPXKNrChQDPT5i/PQy0M6f+EsF0JMLHN0ObRN2d8tGFHt
Sv4Rxm0fA6OyYdwNKqXg3uPUDGjyDc9CLXhw+FIKi/o5CPlY1iUyP9AhnH/DiuJK
aOzeSYNs1+uXYT30jmgsv2eteWxuBUAIEg2UQJu0h9UQi5K14O6xgK3OQhhR54E3
V7Qr+nBTsMzVAC975ZCNGH0jYBg2guvW6wmgEZ4IgoVuT4fVwC4Y0yKnF4fJspBw
CWLIvDn74NI6let4rZDL7ji/sh4cDxN0iCuHGoNFMgv5mNKHIQp11Rbwa/TOKqGa
PmGMAj4e76oT0SxDmdhe4hKxQ7q7xVfREDkgwA2jf8++2Wpaq9c0vTUphCXT5Fwu
WP2tZyYqapcVr3tcac5ga9IBzaVIPD8lvTBbd2WqgdDltifrKvkS2HOA54cccAQP
xjnK0NtBxs6W65ZFqwBTxxErBt/0wGXzL8+HyMpKHQn+7Yn/2xWb+zyOSuiLs513
8AK9GHtrDNyy8HSfgsPmm8v74kpa3n4Pdv7no0CFiTWOSAju6/519CILRnL7dpKy
HzIhAwydnPv29wtpIL7g9uTu4QKYhOL4IXV1QJG75LJ9LaSRpfCR0n69rZduESm4
iaPJy/BxGyfZQPNzAGUHWYHy5jo46TZb8287gAHgQomFTo7QqHIQNjiAwraMeSG8
u13tfkdazdyFnwOx4tmY9UPRSOkouUTZFCRzi1iQ3TDTHwF3csfr3HTYMIO2jkXv
9iGXErbp+9Y/J3nS4m4prH5Aryrc26zjNCNYpg2AFh47UdfU4Kq3tdZLKSPzSg9T
f7j4e7WS48vxL8hxhaVKVyrxyLlxM1ugxBbCltYXO72U9mBUiZroZFtC/585X3sW
3oWrZWeNIT5BViAmO2mEAk9dsi6VsfgjiXIL4TBkqtRqvKLwvsydNlSMWAsBtBF2
A69vmxs08LVAMelqY1k3Rycdms50lHa/4ptG56QfL2O2dpJgaMwBNJzEPQJaDU3q
TSDJ9shyxOm+JjJxEyrlKVkjIF5HgQd5s5yzSFn/eLvkDXEwag5Zy7SmOnaalAW8
vvIuWy0PzJObqY+yqUzHAJ9l+f+pf6si8upQpJhcnlnPdryCDV3fVddv/utjdeW+
x1JMRXYffQt3WgagIL1Ev0t5zvvoIlLsJwsrFNQcSGu3e/98BOWpJG3HK8NaHsTV
sSxCDzh2WA94FaTBYhYWRbzPCEjkgpfbQ7PA2isV/J7tMbg93xUrMlocVpoJHc7x
cZaHwvTmtvltcTdh9lg7Y4rC+i93NNqGDd/8OrDYf3I8UIhAbK3c7koXTJI47t2G
inUz5zFOvv7C33Z2gXTYlFvKJ4Mf+dnNV9pIQVY4ozr72JJAQmjFJwgtNvOhHWbS
eyg43LIihCpIWv9aH/QAmpskCDdAlJYXwC+uxUO6uNvxmMpwLkhAj1Ke1/FNQNs6
WiIjXUDQgxpx6wUGblbfxq3cqmBHa0AdWZE9EfS4USQto0QSdtpoVf+oD1e5j3ds
NxBWlbdzhG1o4Ihfq3jqA430udobsbejsNrVtgxbjh15uYQtEg+V2OrsF5H0MWq+
r+rVVBxquy+sLYClYEioJA/E0Z4rBI3aDuzpu4AUXDJrIUsQxjSFMwxb6CJ3zXmt
WeGNAt8gXy9wjXRwoVSdbkeiWuKU/L+ryThYTcYkmEh+qQm8t35Rs6CN/e9ZCYpm
zqWEMpyPOqqQD+ujwWw7BszgeG3FjtI+myVIcure06w4dcbRtrc8YsMLBd61mhCG
JDMvGIdZ8s8kBJOJuY/el/OZruVURA8MrFkIfELXERncPuZPTxZ7hQZKYs8TJkGa
o7NShNblgLYBa5sxNSsEFLIrjMU/gbv2xA5KbRoKBLDG8buQHkGs33xUqmV0YcGW
gyxvnIOWHeWTfPuAFQciLgR6kI29DhL+R23Ei0A3fWVbk4HxciibTydMDts6szzy
KkhI2vOO748029HngkuPVapskPH3gHoPORoL7pIYRDL9XGZYwSUNmEylIjEZdPTW
IU39T9uz+jxjfHBr8OUA/dbpp7AXwOVDAQFjmqwUDCB5YyYJf2+m3dsf5BMH8cUi
9gyLRL/mGjdchIKYgHQtAAIj8gy2o/WUXANEKUUEXUthV/gXvpvz8hDJipHgn42F
TzI4qN2Mkhdz9ydl8kLQO5lP2wXrUqzopU3NWqDBn8WCvYKoxNqDPfrMLIq5gjgL
ClpJbt5m+M1UaA4KsCZYQOH1ZxmcCJXHZ27XiwC1385B5cZanMhE1Oji/SsuFwv+
5SwcIsdKe49237Udr7Rx0W2vSQ4DhV2tLc3TmMLPjF4eWiEjjJZHzKDKygO+NRCE
SXMZCo6d3WTaJVFFZzISwnrFf+coAd5C/PYApJxXn5Wu6r2Zw7VuclN4SjnspkLV
KCQaRaT5kF2SPSZI9hm6kgNigewF/clfb/9bPgEt1NZ4OxJ6ZYNPZXlsEiDpFa7k
tvlwvApQOsYf5WUxVmuEJ66wNe4XNQGz1uIzQdRxPerHw64fxaDDoqY2KF7GeL7B
PTLO+GafOLA/lHiMhXBW+OT8H5FLVjiox36DpKxmLehpneajB4ecLVyxYeXlS4y4
DfyfOTz1Mn9a8YZRDdSWMEr9i/hxf81zOcRZYmykbgBRI+GT4fL2a9907dUwp8O7
aeohxVOTC45pljwjUnMn/XmMtSuGIQ7xHVXOfZe87RZbyKx9eAq3cHlWHnc4MN4j
EhyUVf+bHwGEO6uLwNONH3D3pFCTs8scFqMraiv9si+6ZwsJHwIbw9j+zbZmjV4f
aeYhvMCI5C/aUsNy8UcHYopmUW6Kclm9Lf8aNrUnKTUMI2zl5c2ADxZDc6nJWyD/
+noW4k0LOVOA6bcS/8AcvfRM5KFlH8OriW37Vy/CS4TkCENQLpFJkJ+MoSiwNrH9
on76QuWYkOAltX9pAF6R1LQ47DiAjnPXaEAa24NF89SP7JqRBjC3LIE0vlHDw5ri
zBr/hjU3dySFC1j+7w8soeFLS7/jiXnOrkIp5bRKJ3r+MCskBKUsL6aQ62BikXO1
JafrA+TT4qcjlJoBVvlL1wQ/bF0Ww/1MRbyZuLpWS3DrV768dUaOxn/h6qcngoQW
BHXTuMiIGfKGb64vwYYnOXvaiTywFyV2lCguPRyL5gBOdO14hs3IOtxDT9jDsIoh
aBFxVWa783l72iGpzsaB9vPWjy9IMQZiSTqU9JjI+gvvaO2IqRqc67u5WdS7ueEb
8aKE7BQQ/S4JGRsAFSoIWfhOH8ejSegFt/D3IuiAzuPO1bLx9gziPkKqSso8wyw7
P4DugUN8rNGb5FGwRFZEtHQ2dQ4qkKbSmT5DO8MGepSBBifpsn1YHZ+pYoDwufcd
WKeATMMkRdkORyX37qeUmUMHohmzQBrwXk1B8Qzl03Ngfbi8uYWWS/tkSGPmSFMe
Y/5+dBUHyPT5S1P4Sv+s8h9erz1HY8BwH3p/5H5yzbB6c/5O9COOpN3E54GCBz9D
r0XfEXGpJ/ggVYrnxTY1PWMZB1V/T6iQj9tUx3C9qxRgndO1f++UsNuQDLuhAKJr
oxMW1aHYd4xyhQ9tfvCpkrkFt+ixBQULqrgJoEc1efAnEfi0+d0UtGTjiL+0OzGg
2uqFpJjoD/chjglBOQGuDAJ+RCrYjlucfHb2q7Q736dMNOUhc6hxSG4Um/FLMcrj
LzEinrrNA9qBbyWMJE6qXnSyXsqqJ6Ov/gdyg0rdHge1cuhW6RFSvAI+jIe6WENO
wABM75SKgKQ4pH2lzbCKhLaASqZ/yQrDjsvzJLcbpApjJL8IORUsiy99bgxoeXx6
JUxbK0bOeyqztB7V+KSajvfmCJDkNjtaL7VxICotpW18v3ta9spF6LmIv2IQlHdy
p8zyhDWHxExuE4FkIqevNmXw+NXTVheA8xvb81DVIDQDL+xg9fl/2NGbdHhr48s5
XrbnSQ7Lg33OXhbqj6kbaIZ3vnJLlCG65HUK+x5DRGPofGCzSl7kNz0yhSQhExni
JdeOlmveqVHnUmO05j65pTOvs4N0q5X3qgaqvD3xHXtf/cI8p32RBK8zQfKRDtuV
95y0l+sYWoEND7tLEeuCszaJXqni+aQy3Qo7U2Go0QllofBfE11GHzfF/jknZpIc
nWB03PVHWEproATc7PrQyW6OvmbQOV7YIEJwDghUwJLeLGtwBFWqaakGeNVJa1Ld
mWJclzzu1CDIjgwg3A4XyfhChejOl/pQJ7iqGs2BxJkMqMKVpCAB38orNpQHheDl
QG98uEtNLUqfn2CFrlSmPlpzzuix5BBpWBgypY8SogwoYfPXO2aWfpPIfEovcf1C
7dWuaZxUfo/WYv3XllCSYBtpxu5RVnDHEKBStJQprXHqkFmVRbZ4e5zq4W6Zn31H
4rrPiFgP793EzkV3r7AdQR/EHfPCW0Zgkf7x7Nnua3BJ6zBXLvGs9EsxEFQ4xsHu
4VZUoOgtQqaORHD7VT6XZYEAg2Bnb1nnI2C0Rm+URILNJzAG/8AvGoYnmOzRBga+
GfrbAr1iqHXd7JKC+DTz275tF6BMI4hmhHr+0njmAn4pvFHJerPajIhbuwlYdTlY
BAJZ1YoSX7MLir5q81SrzxWXbq5XvrYV+PzyULn0ejgtt7+XPhVgk2piz7iXm4wm
tkkML8WT2qRdKd1q3fHktOympkTKzEPnKMKXS4SKOcxJHkEbHxzoDn/Xn/qwL0cx
vpmqHeeVykVttTOaYyykAP7LzRSr6yHTaHUwPdW/KEq6CLYI0WK1AcS7gt/gCrxE
7d1q4jihPrergFiqb3cHA0SA3pslnElnaPwv5EXHCu4jLHYb1k29Inxo1ORKD8tM
Nkn3QGtrFZuN0VnNY+w0q74o82k8OwlkMrquDszgn/aPVJvPvf86VNKg/BnpkMPL
dXKF0TU4QiXkyHozVSsi16KZVEzkCuidp+SHS3HgWPfFkJNVvyjJ4/Z9BqvFeC8A
ouQdL3fTq/NHJRefJcn/oQPHhQHX+L8LN+9kQR4kFS5by7B7dbFSmW4o2s2/taWE
3gnQwVVmNwR/oKGK9mrY1hXuS9ouVU6OO85NKldTIt1GVpwC/A0G/bYpwy+en2xq
OPfol5tp1KdBpeNLPmSMEYMCJXghEwMD/B4FLCOw2DrWvExlF5uLGoQGhNCncYbU
JipNrfBChHi8HXTjGdoQHd5RAoPYvnzGYg9SH19C+SG2m3GOlMZr0VrbUbjLvcwW
95rlV3aK5RZeNOCcCj32/fda6B19XjoiHe/8MVJRRO6sUbAL3r8PRRfvQkLPwz9S
8uNDj6PfWYnhIRiVGoNnIlaZ6mqgshEp6iDpFxA5N4DqNMBD71IKKmDoR+ZzaMpE
+64js54VE7L30BNkqtaTtl1rZ5i9W8thHWC3gx8WMqaiDDSVOJ3mF5d7G7s060kV
UXyvLf5DwjvHJ3uHm67ee0EtYrjqBKyZ+UjNpxOYZ/b7SUO/pelGo6h7CHyUNEJo
sLODvVwzMLktj/WutUVxjQyPSZ1AEWzrjTb4ypnGsuMS4Sju/F/70/5ogJQ3v6xC
oVnYKZm64ECmdDV7QEm9c+v6ftlm+qb40auwi4mLxokJxvVK9cayLK5Ne5JyWkSA
guJ0gZ7A/oRTgd2ffEhKSgc8xvfO/cXD+cJTGoYy+9PkYtlvAvBWWOFvuWzHn+jt
tGv2gt+ccyqWNcXYqtCshEpd/9i1FeKQr0RH5HFRizidjaIqwGHnZMe1cTyxMOnp
mvC9p/mxp8krN0kpW28VT+KMoYi6B19NxSecph08ciA6QkYt1j9w2YvMZPHUZR2m
1LaPlGBSZqyz+d1PVLrQ0E+VO/3nl3PREzc+00igggTNWT9edDmlNMR3rbdL+3nH
0PBEdtFBi0knlrR+nj487lWljY8hItjTedYfhfYTDjfqSvrsVjCRFGewZpI0iBA+
ykJrRrlaPqIy6zHqENVbJ4ifSS3fwgJD3n7EVhKzhzfqc+riK5BJNy+6U1evr95Y
XKVPfSv4Pr+ZSVLwwepnu+AtyvmebyneKDCpkJDaMD1PWRRaGNhdnNhI300F+JJA
MegnSykhlZ2UBG+kXcwnIY3TDrckFeUBQNAQlho3D5jfi6nncmqGk42QrkrJ7XyY
m8ciq9lDCeQwu6bNJf2torZ4/cvJg8kwerVB6JKR/ZLnRO0EKBsoZvy7WN+1HGA9
63h1rUBKDoJ/r2SWyDDveNoEgPRK+jsnTXjP1UuhTpsStlPuSS/DQ7skLnsmOTJ7
6wfgLsZjiMfkQTSikIRfGPRUW4vPC/HMnFdmO2hrcESsrZrhUEb41v2VfiVoG2ns
K6hzXZVP69aWs+RysOB+EyDw15HZPfxL/AQEzZZPq/6SguAIG8MMXnnjITdfVIXS
T+kyrCGXDEVPtXMSbDClPfWaeu32XknBF3V+bgh2ibH5IQHh22CtYDtsnM7bpLAm
+BEoC5BjjuF3GgZ27Xp9i73KWhDyIp7P2sIlNfiTcN1uF/nXTTgtdBTzCcVWHmaC
D+/CA/2I5CbPxDvNRjs54MqrAaTUgj0ODw4Cga9ZlnzrqDesfHkgRDAsftU8sw5T
F4Zqrd2AmSXSqrlYywVPOw==
`protect end_protected
