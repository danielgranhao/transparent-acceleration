-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
dDS7eCs0bO/qf+3oHA+zgJBPmLeFybsVNZtV90J08nuSB/LEq4yOhgRUw4D7BWROTq5apLCfd4J9
Srj8D/WNmFe9/LiE6fAPm209y/xQ2Cku4ZrrR80S9461Hx9wxVpk98I8HcIw/ciLbYEza5TW8mHf
4NrmgpsSlserofsQrRY9KJTPmxik/dN2vS8TKDYO6DPbv1Q8d8BZtU4DAMmlVE/htLS15kllXAiR
PwVsMZ5j/cQUdlnKwjEn9XOL69ngxEx79YSAuqLJ1Zf7B6kju+KkynpvSyaWZ+/EA5RIRffWqrwm
cMfMp8pj99VESZfxjY6hwkZwT6g2odD5m9KN5w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4848)
`protect data_block
yGgo4gk0F5uNtJEFKjp+1kyNwgPtdraIcohEEkb1O6B7C+EUhurrVbkKCNbfpzX3QGnOPIBX7eMy
Z2Bgx97nEwq6usYgWjOQR69BHNMUEjTAiawq9yNUew/ye0HuE2c8f7aLtHSuLgFVLwwc1zclwkyX
vGcmLi7m4yQ7sJIr8V2gq7FZk+UPV6XaQUOM2PeXHOzw6j+lPv3UogdLc+mofl3NeaMpQD1DncKY
2a6cVgXMs2sdKEpB47fRRy6SbuV+puAucHWScftXRnO24MXg63Hu/Hm3kfuN22QBlM4BOJRr0Out
YFb9iHaO178hQyJyZkS3l9PUVP4P4bIqtuECZpv6iL7gwFixsA/DM4NJ13VG5oWBLhSsU8l6tvH/
kY/MvNXMRr6qvU9SV32qCYW5p6DQPwjnG2KQBXEo/FMkMtbZMhE3m9VObVwJp0hUTWdiWAgbeJ+f
j9KuHIv//pk2Qh8zxx+8a8UPVAQdqZe0yQSEsnIuAszxUwle7ljzdUJfwrv+OFx1wQcRI/w97Bkh
kHZ4J5Xlzpow5SpxKFnX+SkF4kwwcFr5VUXZxXxjwsGvoXkDDisLWEyLbz29MPoqb7Qlzb4wuIH6
oUbFDdgksdPN4aqXnn/H/L7VJrKZAigFGoBmSjj3Yu+gj701+MpDLBN217Ej4B8Beo3LXF7BSqhG
n0MqW/mD1OXA+Gn97YiLaTyX7wTjjKvDQnfxdJS+GhvwKYrQ/7OiTK1oqQ4QlmwmS4FCv+y51eNY
6tm8zdT0kHdGYm2aTvh62u/AYZGrZpCasRh5jj3MNdTheXWza9xto30m4RtHD350Yy/ylfCuGxiQ
vLOdvxVs9tJdZ0WYostCmwTu+vSz9xzHOtfqQwwSXIAjqlcaRN7+0tbs2PIvwOXeSD+PMLNl/3Q6
iIwRUDJIN6x1u6jWHrXoGadvZ6+zhjopj/EPgMwCSGvVwmdw4bCuCT5/MJ5DcKwlyvFRC20/SMle
Z/OKKCUqAooQeZ6VYwlPVTml8XpCPkl2GMWx26o3NwqiJECvXAHTHx+9dQbWdWydGcK5DMirrFgc
7NNPCJcGWNd7sfluOOuLff4c/14C6ggvwyW8ByP9J8QRLJiOB0Ukba8oMpdznDBaM6o5f3oQGFty
j4f7hW4g1OGgAdqx7HLp/2EBlFkBMHqbDgmMgrCjKyXVIlDQfjGHrOuSxCaG8bTEAbFaWMCrgpG7
2WfLQDNN91J+9T0js4MQ6fCBdL8riYxPdYJFYRcmOJIJXJHsq+kknniSnvRXZ8+cZmybQN0Ec8jp
CfkINjUMpm54y9uYUpbM1awVdedGPku7e82xdQpv6m6QarhJhH1HZqwOTK2oj8Abp1KgedKGGTx0
xe5I3bK25F4kAurbEpMyqEUSzUahgfQCoqFoHS2KkmnRFGIKy+kcXuqzrbY8wWxGUeYwq6Z+roAc
OeDT6w93iKUOqmOaj7BWQLAI9giwerfJF3iYZZpvfnBaWMV0dP6wH/N9RoOyp7KC21rvHZs458MC
1XAT8WWYkM5szshk65jIZiPPPf3Gq8Z4costaSaxlwwSJI0OCHA/av7v9c8CHUKIkscamUNBsDli
xoGPRSjCVh0V9sUB8e/gfqX4J8gKCtTX1ReP8/drjIT16woXn+n9+51I/6qtzbL1E0zgF2ZSkm2+
WPItKAOu0W/Dh7u1ByINa32x+36ts0yVAMBJ4LLKqew3FXoPiPoeLFN39jJf/dFy9d+82YTYpQW8
1LD6657doPZK4yL43tgF6hxFjQXqeuTPd6M+MqVVSYq/F0RSeWsnfR7kPoSd/xlLvsuvHAbzsLnA
mfJM2RK+pqyieUjSbbewVLMScc0V7CB8e+DyJNMclcL0UyfFCrZK27XYtWGeWOhZIEkNY2RgaACn
mLCV5Ev4vskiclaNOavNjxAb5DyWJGNeG8ctyPiVK1vfRkoUNkroD0gu479y6uBZSmt6OAr7bSJw
MusmEW9vxPT8ihimNNenTRWzEE5nwiKe+YojK7WWBsO8U67vqAMnaSS66jcTgSf9DEJUs9MvMHVS
rkeW26TPlU45LmQhVPo+sdDyZ9uFCtGr/glzfQ98e372TG7OpcsJpwf8TTGQflmWqmjXOCJHJNBz
R8KdAyyg4ndg4+4TENjhD+lNxAzyb5K5K0hiRVEr10r0viJQqmN0cV1rDG2cVsQ7J+XczB2Jw+Rb
FRe0ofd9xT9k1oIA5OA3/VkRK+NzTB4J5H8UmeqvVsU5NFagFDgOm/c5S5Buxi8/8Cb9u8jGqp16
jCU5XoUmitv2NxeF3dyAydGGiQY0bWhP/G4bZ+61RI1jO79+uDSW4YuFnBP+OVNyct15J4LNIeHD
ihjvpQJtc01JCgDWslUDecD6ZpK7J8n0kb51l50L1OmiBQByZmMTFpbh+EMez4jcPg72iEQGNkYV
x1mgD041BX9VIMh8FOPGZaU+ttoWpDiLNWoYItcsar0TZIPItVfL0A9DslixZ4cewigq0VVlhPk3
7vGKntixM+gWKJ8sBnHyd5pvWEd/mE2UALpmKWzL42MmYHqWI3WLdb+sC1ic6E4+7lu2Ofz3024P
LBbRQoDSuEe5RM8n9VWmECXJgbAI0zl2OmflmAsMcDnyxMNIiktTJ0UsG0ST7XT168BxCrv2V4AG
6+boBsFy+i2HSmtfSNbMx5oZCZdtY2oAQxdqravXjYS4K+2Ig9ZuNldTvFO3pZhP53XYQzqeRQPw
V5ZtKIEp6upTVTmOZFKiP1CXuFw12G0c+UQSPyHdU5ZPth9DoFOPNYx+IsloqtKO9O0tQrTp92tt
8d1CSBbJYj13vMowRcyrVEnZrG8HuxlG74u6qr8kaAuLO3RSm0H4q10tlnIuCAolWJ/2hwEpyS9W
ntP1lmsHp2n3DzTLwHvgC8T2bDfwb1J9kIfSfiNuQpzq0gUR0owFTCu+aI0Q0DXnPCfCeJikn5D8
MIVj49e+d/D9WtGNtKuZxJ7FurmF8GoucgnYmoGC7Kg7hzI/bwXKrZYjRsaKk/jR/thS4rj3Utn4
ALz7tfMwl6sxUGKQ0z478ythh4yYj5K61BQAYZcZ9YfHCQOZBTtHD4DE+qtpTvVOm+NdMteHer5r
lhFV7D8rHbDSeUb5XMfqBWHrR5tE8RtQ1gq6wZBBl/7sONch5m3dhFKgvBVyr+JzRAvcVXH4M329
YNeRZf8iqWLwgKHpe8QYzzOj26lhTcp+yfUFxrdrshWV85BKM+ggQqePNaS7OPEgjShPbRGefVIW
DCAYalYknIfIcaRUnyxN3GJy8H72/YZUcO1kMpNcjGjmdhEXgB2qEQx6ApA971Jr7HZN5cmhuyDi
ivp5GHA855pAgFQdDiBnwtp/GunZXKPHsIkUryGvy55O23poNL4YQrOGOhRNOeb9geUt/qAD16he
GcJJ6UaK1GqHZ/ngRIxtrBjvVm1WbMjK4LpHpMiCyLApwrvB3Bb3OZGStWSDygKg4yKdk+7cB5NU
jADIaoWS8QRVQWg0XqL3wamDO87XPflIOfK0F0fYXrfEf1hCPQxcI2m6qN+2q8ivAyBxwoa2JV0I
N1CYmOosUREEsX7tuhJKsn7P/tBjhgwHqFt2lI5gP7+eUpLE9DjTQp8KngjyuSpnQe4nUZBtPq81
c63+uCKWtUeGG2SrCERAtFiPUfw/EHF4RPM3RObc3WTBBjqTRws5Suj+PhQAow6e7+H6i/yMZbON
L8B7ZUU1PgObdwpVRnUThF+g+i77winfw4DwCOzh8vj2BJhhKqqQF6rfzpQ1NEf9svl3AM/3hLFQ
zZFy+4JVvxYb8jHa0EUtc+Y7TXJRzsIv3OV9q1jT59u2pIVD0OOm2Pw9lhYo0RIIwmlyHxne+APJ
5IDl6GVEP0GwvOSSk6hOOv0QqB/PpgfHxN9qz2GAfwpGdseO8WKmhWR52wEwCaoMZYiKpjTo7/LC
sAhQBogBSLBXOAEqGjMZon8nC4QU6NIgDx24rHKZDRSHT7zLC8Xx507Nz7YUV1fK1YqxfykJmSdy
dfdOAorb8sXhM0+7fmMAyAjceXMu0ofG0pmnOJ5xBfl6/xIOECxx93/z15w8dIbawr57TNqAJSb3
NMvswjIdeCWp1mdQfyNQtoQG9XkhCJlJEb3DHrAJr222oU/iV7DuP9Icruw1WjR68I8nU/CyOdH9
ZYaBMdP1xA81FKxrsC2Q8AREfcjZtlUxiPExwRmRABcaw5RIHVouRG8TxWpFslsJAZOKlqZ8o0KT
wA/H6Wwoh8/nprx/SMQS3HRMpK/Ilr453HU0Y/HY5JbaRkSQQjJ6qYXj2ioCAIr1r+a/191LTcih
nm2BD8zxylOJUAhLj9/5f+Zge4s+/J8ID9Oy/qD8tXIGTFwjqB3aGCahcMtdcayVYQ7YQW9lzvy6
1FazEyBiL9EY3V0/MkOn9J0lkoyoxvT3+UbMSO3GyMQjSHyUVAFBOMwDShvqBRWPVXnxGPZXXRrn
GfPZoEpkyyKWpni+JetTKlLCW/kxh8osww8tsok3mjmJhLFHkIao51Qm1TBU1KJk82aGcn4uluvL
+Vh1TrAgW3oWTsRArp+bxNSh6z5CMrxkJqiQs2eqFdCfWSk9uZOiINDS4APzyg3pgpUIbO6afASn
1OHHy1QPTeaWjfqnfmYw9zQJfc4rNsQne0yyT81Tp4lNslIkr2mJ0EcEMXKszNomtJUoDutyWpbG
dM4ZP9zsIIgGmGViRWn7A/3IhiYzx2t7GQcL35K/UyCn5rgHCfuHtk1c7gui13mK5M1s7mCgHeCU
jqxigrCsy/zsN5Oo/4EpJekt0BtXJtK0uGR5AxSHSvTvUxozWwalJMSAgceo6fERTefst0UiTmKv
RuA5BioFPRquKYHSJfvhaDYqvAPp4GVoZtr2sPNX/vCJeXjBifTVxhNP8a6cj+QXS2k6xP5oUZcm
mXzn9Sbabw8g7MVnw8jNJfdm0fhTR2DnOpD/6rYWxzHlGtPXjNnAwi3NYV3SKmsdF4iLDxZHu10g
GE5QucXhR3I9oV/DZ6R8Sn+tAJJK16yRNj62gBK9o3sgBU8DYEQ8ZIYnxrCj6sjUJyysQJUVkK1E
lSXeu/c3eOY1UimwXnR/w+vvdzlJAFZV00T157lwPOyrfJHfB9GjOCL3dzRiuTXkLyOx4mulF9yK
uk/pSoTPR0dkHTkLVxQ0FX+I+B5ucp8FEAmexrnYRzCP73/B47J1LQXUkMyNdzE3AERqakd5XHoZ
B3LB6ftm2kNfhKwee2um1m17rkEWe1WBCk2JUZT/KRCuxidTNFsqOloiicR1l1xAVzDzGkQCp+of
j+HkCZQIokFJMXO2lg9xXXD8A5AqK+Y3d2mMuoo9SyuXTwr+x7wW0RPop3b0NYTcYE5+es7OR29h
92nt7m9CVmcegFhqo5c8azZ+FMRdMvgu7HkRw6wPazHtYIaqD3f5ugZZJNHqUuRzObpivKRngaAw
8eMnC11zzLpMGauXSj/E4rx3dqIQj6yxDFeI5xDFZWOUCFHM/OTSTJ+k5HJ61eGiLTaZR1pjKNh8
o3eJUI9rDyqPcmdWcYS0kSWfuZ/v2+hLD1Z22VnIZKWnk+BkF3C0F9pnMfVL4i71kkco1jc0QRAC
re2+eZKusqAk5dweFJ7LXenVviTdJsQ0fsQfs4LFN6i8YnwJcBragccR0gZYIFfWnKamho4JrkvO
J95HKL8vJnpfhc6nryVCXjJ+qD/owDs7FIhLz9sbVwisRm1Zaa8BApn1ICx2b0tn9IG/PoviphJD
qK1XIp/J9avQ2yR8GZGrqAHkOCA2pdkL2/YbNQ+B9ibP9LGrD+1j0WjKsCfFy+KoxD44EEv0WDcN
K/fJ27osfjAssP3TQN4kwvAEnW0IasokdGdkQmrKaocGRNUwMdHbNILxNVJvx9orWcmWsU7PJDMt
Qi2/8UUkaBgcAIF4gBZQ9EiFBodC9X3VA4PnxXrayJxBd51OR/geIX012AsF1qB155n3I3ndSCmH
FuxJZSkLUZswCiqaKL0gecFW+ide7tLwHh/4+UEVkv9SoEfBFqQzgojfl3aLfvboUuyh2zMd394w
L6WYO4Sz29L6zR+j6m7NgOPIxoSuvvm2sxY6vlODi3RbCInr5R1ZxQLiNlSMjpo70il5mB2qcBan
mhTor+FkZMQwwGCPoA9UFtYSfyJlGgJQvUBZsWN0lutTT3ki1xf4l8otbnlfU4++bKU2zotScpZi
LoFGYMF44syzc4CHsUvLiLyKYaUN1QCiYgHaiIlk4JfcIb/+N9h8yjxRJuhyjeyD0Wl/PD7hQ/9v
uUR0LrKBpSlrHEac9fXUihs8st6hNa2RGdYZ5LxwiMoldSD9ofMQW9Ky1VCC1gyT4QoR+/kAoFnB
lYfkIpPuoMshGORnps1sGh9MCJwe+pjAbIYInCmLBvnKkvffMgTsRc81gsFNHa7VPSwG2YBAcxAU
LK8F
`protect end_protected
