-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tMQfPK85ND2VmrciTaG4S0g/NnHmfjdQDhO/GSMLntFQRLvhYr8xyxcKZVCHKfMM8Z6Sa0CfMtcu
ib+YaxL4+rGWi9xFe2UNy6k64QV/qPVKCYCvWnBdyrSkFDIwqlewT7/05QKIXLYcWrOWj3rt5Ui1
7e7yo2QPVp2b76YxYXssVHiSR1RYa/8Z9LhbTvZXd6/gBRau2npyxclQCiZA0OT/YiPdmlRdu8Yq
zzE7nnrQpLU+obgjEE+2knztke+daibxe4owbDxWQ6AdLS8izbTJu7LdbjiPzEFQQIZHvuZwg7fX
BhIT69nOIRNCm+8NZ9OSgSeWc7twlGosR/nTVw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4176)
`protect data_block
KGuH38MvBMXdORJwS9XbHCLF6a3QN5B1yUz+cZxTEbT8p8zKJaxsymGRfECeByWPN9Go7IMvXAhC
caVD/FWccdoZFs8imp/ZyAp74TnEVOWsHytQQSHyqA4qBu5NP2+r9Ujw1LGZoy4JGrY0JtWSxlGj
lUjb7VcJt79rdqVeCCP0Hfp7XDlfgwpYvfxCSWp28FTCSA/Bh2Bp2sj4bqhsjqm47S5lPvexS4kg
qGSfXM+U3kxpVxDxvIX+H1bIF90PYuYwk+PAVDoJN6Sj2l0T9KRM6HpRKSMGw8vud+lFrvubqDT/
yIFMEOg3skt5PZ26kKGtylgBZMOEnVHFOzY/wleFPss/H7Vj2jjNf2CKJ2DV36mzr9FXhvwO8jMx
Akt2KOkZQMGa0DpResDVK38v34zYq82v9Eo1QWec/rebpuqmG6HdsqNrXlB6yUFmwiTY/TNUKKTL
rgX1uzPCYNvO+HBGSmfjhdUkf/bMUISg5i1NMlsg1vfi9aBWf0/Xvv4tTLtd7ItqnmDX1hV0r4kL
K8SP5LEdP9jDtRydCvPXbE+Yt81jKr9ks8DKV4GsG+f4KwGYi+pbps76I/WAXPHF/mttQZK4mnqT
w7EysKsDgvPhbqsdBVBDaiGDYNuQZBZQK9zQJWXtbLtJbB/cJ9a3SzTsqo9F6HgUGwwQL4qg6dWw
VaPOb4ArcmZHWGgyeivwpzCwhBUmt/JgKC2d+7eLDe1yJEVBldKERw76Wg+qsE17Rtw4eVErBKct
ApDD2P8WYmvldrgHW0zvw2piEhtF8Rak7rbE0UIyJudGW3Wl3wmO7T2WaYWTKNbnUf07WA0c6sRz
SHy+EKWhV32FPxLHolVtnP8WaoHgbgENoFKpWVEsY4t7zJSLY80/Owi6sRANdx3DITEmM6JE0aX+
nJCrPxPHPf4trd7rOML+r3c/bDt/M7an75Jla0ikJ7Nyn6b1akcnJn/6aNbfn81uUA/owF9IZiHR
QxG0iy21r+QXxm+6Zfp5hyy5QZcTXM8LCV0g9kvNrNpaK/a7tDmdcZWXou87k3Gh9leUZgn7yeU+
8cW9RtLj5B+8pNak76i74tKnF/v0U3KekZ84c+kbL4xW/sXZBJgS/aIxDpBMgNrhtTCV+9TifVUu
B/APnMkB/7pJ2Erg++7g4QJNdoI7NBC9/JI7Zs3qIoQewNh1h3PjXfFzqUHqa+rkOq+Z94aM4/q8
JnL2eSUjXsDDLNejDdJdBYoMRd6QuJVr6DsafEClGuULpuesA7iEYKiEt5Tx4sJiZRD6Mmrejgu/
aaVdhonQeHlGsq9XaezrsMCCOnN+r7oCnIUbB8FXId68M8rT9eRCp0pxg/k/ZxFr82zwi69bKCB8
4wexbZN7BfbaQZ6rVZqo4KuHHI+gFMsDlwS/NWH5C5hbANPd5huSO+K+2wOc0vyTbFIK6pkh+Rh5
cid7JatQlw7U3jAXv2f46+q8RYSCuDxo5dJbLo57N9OAnCyxEYFJlxs97NZkfDt+YSRq9rnQNf9v
MgYYzEqNJDVweRMRHIXH30hn6Y1ibuHQYGWvvPOIg5fPkWznAhLFvHzVYOjw/QU+C5AVn4gwPojq
MMa59133jnAkPcKtso/6NFTK5VG7vo3i/0Sc2Nb96Jv5cW/kHlV3vhe1a3UicckJ2Fii654rdcMi
hqrI9XtqfM5nI6fcCsqNWnjf6dFszn9Wk/+gq2QdLes5eg/P9lVW8xZoBOM+okhWUXXYftP3mymR
HotiwsLw3/hUQVB1vXnOb1ZPyMfjTfw+c9awA17tlgtJvJCt7il2ocKBGMsZ+CJLCetvhstOSB5x
dSyr1Ko1pqEhH2oojUu/2hNmI+m3ak5ppaSHCbzJjDuoSZqbMBGU7MptnFZTJKvYZMXpAW81Vm+U
49MSG74C+V73lN+tHtToUyAQ2zrgISuRm3cSxad1VHtxNa1TYl5pekr3mF2N+hZUAYRwKecP8eNC
Z044XF0s7hox4TXhaW/LPAlRwwmh6i1PnYbaXN6lEp+j5WF4Z0rMgFBWvLLVP0Oj7z3eW5Tdwh1X
sK7gKVETXv/La5RkDtOqYWx/M58LdIPvcIrnL8VoVLSRy6/txGzKmSeXc2AcftJkKbwtxD1/ggFj
5/oyMrE9U19zjtNygoUe9QVL7y5rwGoHEeB/j3/6uuwZ24wfP24HCY2jEdMaJwe++3C7/+Cp8NKc
Tg1nxL/qPYjMudTWbmHX15zOnF73CJ+942HhdDlvRO4033nuJVZdjyvm1uyheaYPuCvQ85P3D+wp
FMpxHlO5hogigN64lfCC11mehw6D3hhrGg/3mfEUGh8Z2K3jDhfYtxEZVABlyCH5OQT8kUdmFYyF
mHzGCocJhk6MAw853Li7LFiIQvJGx2Eva/ADYVSEHK961Zw+6ZIhiS0AiX+ZGxEeuvP8Mxvba3ej
QcT9ZWPqnX+i52sWOc11I+2il4P5ucnHHZAEAHV2MnKJdYrC3MQhaeWhjPd2ba3JsV9l//soWDQI
WgF2XTP2FVDBemCgD/IeBreiv9qBIlwK9WA44YIhZTbmQnK+r2OpkT41UwyhBQl1ahmGctY8jzbo
yva1GJZ0eRAl0/Bbmq2SSc7xXt1k5QupVZ9/mzSoYaf1kCHPf4t/ter4mqNjyxqnMP5CPb2BQc1S
aPLxrkA3DQX7zVUQl4E8GO+FUhLwHNKp3PieggovpNhLBCR3eW5IvTngHCiXqSQm90uqY2kwTOsh
1cnyuMTJL4vRkNEL0X6tisIl4Toxx/aHy0crtaV+dREaesGDBchzTnG0CMympSBx5D7VW5uxwzxy
cdHDmoavjophA/Dio4ObCeRicDT1xEIxH2Oe8xY/m3nrgtS4XXTH6XOP7aUvMm7S42VI4b9ILxoB
vZqx1JlQnhDmwfpjjkLqvwPD6ZooDNTsKquDR8hOkbiemGCJOClKdKes3HW6+t2COtcpgV6Lw9sr
cE4JLcNXn9IpR7npRkrK7AjX7fB+8dAJFDPbffxoekXAHtsREOyp5fmNzHLf5+rt6bISFwjZcjHC
9xoc9CcMwPSLOfY4A9WSZRFduNOBV3B5Ur4wB3S/8eJHM8xIlc0gNWNpI/YqmQhyEv2fkiCv6aBr
izzAOcPUbSoWBlyVk7z5YnTI04VYpxZ33nJnwzFiEiea7sIGtLkPv6UsArXojH6VGgnKsvW8gYu5
Nu3XHXVwMxs+/NzJXYhxce2LoulLUynXp5R0dJE9rdCTfNBKU5b9aEXui3+FCkUMzJP0ZO2VP/zb
D/TLgugj9mJ8T8JgVALFjo8gYpXj2Hw2epA7MVu3aldZad4osATGeviaKTOoAA7J1RwQN9NRA8W1
ba1X5etlHSSl8QTx7RmHd9blmkDaUs+1eZiTl1+Gs4vVakHKEgebop9wBSFdHsYyoKeCQusWLfAE
vJkQbBGoOC4YXGuEltAJB21T7Xra2X4y/CRCEVqhxmzX7Gvat3ylPqUXYam8+6QWozN/gXINoVwi
yHJ97ffhOlBBHPexKHkBiQBWpHA673rmpyDDV7ZJRPKy+grf9jQjhZC5sz39CfeW4eMLYanT7COl
zvkrjaL3Cve8oEglSUCP1aoE1uvKiG7rv/wSrl3tk5sdXNKGd5T6BbR17ZZR4TNctjHcBZsQkfbg
IeLon6cDp/672gvri5njni47Q3tSh7es+E2s3hg39tdeKEV1F34P5mj4WWDFNv+9BRfCcvFS/9iu
85LRhvmRHDKgRM01ymcXB+GFlaXY/KQAypVZn2P9bS3oC6FkOMbUGQaBVJ2uG9peft+ejQlUJZWR
I2kvT5PIVqC+ajd1N3ntKMhZZYJhfnq4UySNRfa2ex2j/PrQi17GayeT4HT6GME5LRsBxnAPj9cz
V8v4/rrUO3CL7poOeWqBB0fj3zgdUHvNj5kPVwxB5izzYXwVtHyObfNHYeSeFLCpaf8IVlYXvkwH
1ifU2hTiLB21QLhOVUr7jwzSwxJuvW1c16T+wTCLdnUGuly5rJZIUhsM4QCa7JCsPrOTY3il5iq7
LyJY/Vw8g30qFNmWwHmAXWcOr0sauGXERLaLomWflgIN1ZTSz/IqFZm4evHYYLASaqpMdNYp4Ig3
9HSOiAYM24TYY5emlkIcf7selbUkgkvifBhRe5RlfVwhApJcIjoOtjEPQoyt04Sbfei6A8a+qm3X
jGw+dg+hRIdXAfRcTn9QBmuQ/YVG0K4hMxHTigVdQYKOSZqTwMnJjVh0uj78oWmgRKtvK3kzcjwZ
dNMxd+3oA74T4Ii6OktXK1sVtcvHU+8fredkHuBxefpWBdq3psYWDlU50q8KKDak/votmy36unAC
qu3cnuu90YBoWCNczS8pHBanOAJdM7Tz8E3rna2WVKIlv0DkT4E7saFMc3KyF8uvCIMuINKAuGa3
gwTe2cAqT98cvehaqp3FYfqo0/fClEc9Bi6DXaz/KXPE9FWeYkwCWI3Tx1QLsd6Ks19wJc4k83Ku
bEi1wmYmQRgPWTcqINFThpYtXpfJpzyfqNL3sFfFT4Ts0MLBvdk9IsLUWbeiO7SshvgONVNqZAZv
mvo5cYQV0MpQb9nd7bYVx69nMV8MsfVH+SDfXOeSBn3EdD+VTbARao3jUFTI1c4uwSSAgiRwKMz3
es01+IpQWDFpCA7Nlu4oWt8ZLnXt2ExXk8YOUuAKCuXSNzSwhrq+5HiIkkSclkaaK9+5ulXAIFpL
O66V0865/I8v15BbjT+lzHVpyUcmqkZhDzre1eg7utAxBnadX9SWhTw9kAzDMVpBZ7y1YpiGtvTn
9VZMJ+OuUe0Yqy3lAbRH4Rr5NIRUwMqSGoTHIfFs4dS45RlwBNkOj8C3VRqfr7TeZyQip2GqbWiL
rDWDNeLo+U01ycH+BNBKhZlvKiDQ422UUsDSxyujynN01lZMabq1zJhGJemhUADVfZAJOfEtvg5r
OIfV+79kx/m+rsuIVCm6KFq6POSQyswz7z27MstaoTpR+w2k6XD70f1NunU3XErZ23w7hX9TFhbP
E5ZyCGJwUiBXMDqmeMpgbZlY7Y5pIPLFLzg1HombMhLodiVYvjKrOgPPBZBg6MKRaFBktqlghhit
H9STcfzYgXrfI/Ew9wHNfHtHOdG5orETWJY2nkS30mbmXu/uDj0+asVm1sqBNAAxMKht+qAmpvue
PBlVKwuAcWTSmuGcv/AIsOQH106Hs3DkRaQJMi7QgEQrUO2qOXBe74IhEXKJginmVVlxJc30V0Iy
W2ypfnwJpHf+ntFk1WXmGcNWfMaxg40WNowz1STFqsVJf7zdCeT8onw8z3GHHUm0CvckogN2rzbZ
GcVnYHpksuRVucfNstPKN/R7zCON4pOJRgl+IOVyJBdBU4Qo9qTVogsTnkkqw8Jmexnd7aWGkZbE
TO8mD2jIp+ViLWdAZ3yuOgXy0ETUyeOj5F4EpE2W/VGuoabYqQg0ihVW4dJ+BIogKBU4wyUlGPnd
HPDLl4mz2FB8MdoumY0Zt+Lld2+QAOtEhaxfEF3xTgtpKqSw+087KhyzZPSzYadRLwgVFgppS3yz
9baZW4lHvlmFDJ70JeeL
`protect end_protected
