-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
F1G6VfVYtao2c375ELkzYv4mBBy770duHkm4VxF14LQppUcxm3l3c0fW2a7L4swM
BNhZM82GTfKQh0x16yh/lMKqYFS41aSty5wEtdtPsRTq4G070sqdx1dARlpnaDjO
8KibBNaO5AyGYry0WqHhbdo5jKP+ZfH+J/G6Qo3Itwuradz74s8OFg==
--pragma protect end_key_block
--pragma protect digest_block
Kc1q2KT7wTiZUD18jjiUwoApXSc=
--pragma protect end_digest_block
--pragma protect data_block
swwxjcOJn6pazhuiO1HnW08+iCNfY5oEQ5BQP0Zf6ZEnaYRoSBfETWT0gTgFM6r5
5W9CYkOt9y/A2Hu9Cx5HAI2JARgrxbKNxHBfn1NNKn6v+VLoSHazMIHE7ODvp97k
NcQ3QXVnB82wyzmM9kASZ4FYd2TXUPCi4puxgWxYkoz5AQRrlhp1eNWH3furP6qk
laqFkbb9Ndrd7Bw+i4ciJ6Nf0f2wLL4KCTXVFAJRy6F6yZsnyj6Q5HrJqrx155Ds
TiJkgsaEw6CCSW7lB6c2wcMkTIBgkNqlM0RcMpWp450DT7TWy9MjSHEPm36BfYaK
LUqfXbl3pQJUFcRFeAjE1hCYNnxJf5iJuF/W51PR/bITxFrPvDewsmxhHWQurDio
E/qZqWkULTJR3EWZMY19AV0W6koAxr7+TkJFropONZj34i0lgeijFqSVFe1xKqUi
z1EsJIilF5dKUzw+zIYK9m2W5vprh8cVa1xmtsIcR2lgURemhKU+6KXgSk8nnbFr
zAQi6viCy9ogcUmJuYkaG7b9f5Tpc8kaDkgpXQ905peKmmbc8pzNW8dE3BK58BCE
wljqq8RFc12o0P3BFewVJXy4nhFWjvoAgspaG+OA3YqR1b69TjaVSQsTYwALCwUb
uTOU6Gte4tYrLXBAm/H67DrMAusC9t5erKVmcw1LsrOKx+BltCboTmQLlB/3wcSS
iE/Uk2vefw5Fl742a9DXtsoqDdZweziHIMMRTcd691m8fZmnojd0T4Pp/6t6Btiy
SFQvXR90M1LVYRC8eISi3CCpaHi4Eczhgr/Shv/TeKPc5X+TYNTKReP9BzxYM0vZ
znHmWVO5HUZdikcR4TrO4X++e2R31NCf/jVsdPuj0r/RnyHU9yBkUPlSAIQzwRqG
bkv1O5kE8LkEHnUvQNQgT7eZQSOsLhZUDpp7Y0Q0oAMZHItf/csIa2sryvIQRHW8
fd4mqlzk6SMW4XSbSMEEFEE7cteHWytJhM5jQJolAumb8X/L+zGbbSUWsBSDc94G
EpgWckRZhkmdIUhGoizrzEBECSL5LrDyFf6HzCrOFP61KOD7EUw6as21UA7d3+xH
uQF7BDJ9B8MyfHldCpZRo1wsPNT3pexMjPEbkH0wcx6wnuCPf8IjnLi8bNJI6Jnw
iREGwFRe7GcJrJG+cr5T8v91XK20mlJUv+DEo8Q/i5yAXVgnV9nsEOqdkfb41xU8
85LkYYDoknvIQFjC/sdVNaCAwN2fLNi5zmw8CJT8XUNoGiLmEdOek40J5x5btCEn
AWUetXvN+1SWzwpjn1MFTeIoVVGLwJ0swExd7IpwsYCmhZ4+1Vmt55k56FxLkMmb
iuVUUT/92K0z2wsOWqgdUXsmHvbFXL79bhaqQoEmalOVCH+Pndu+xReJxYd0sTBG
D6lG+l0YRgYOrpvGB+gJKFXEBkEc6E2xOJIXGe3DyQj8pK5hi06DZ7nV8KGN0eaY
eagqth6KTK+wElAtnKHLHlO5Maq2WGfsYiJzPJ7lujK7bR0Qr7srTqApGKigrso3
bpXneE6H1FITlVLjl0iALYvso3UYSELKLCKg+oSvBZA/0YrrhRIhsGRmxksV6c6B
QfucdTQEaMjLsEnFdRfaD7+9DbX+YljDBFsyW25/bQFcE3Smdvtc3PZ5DQFUq1xj
cKcNZN2xHoVkW/fFLBmblnDfAh03IaeeRDuq87aU5MQZ81JHv2y/7Lej4PMQgWno
nni6FNp67SNEXNcULwk9jt0Mc63XqIcSV63ZzYScpvDfmvAuSPqGZ14GGtVEEOpJ
4Gk/cyhYmxB52ZbmSNqyA08xOC7yWKnzPAghaskqVZtT+YMGbY6xBBoZ3S3N91bX
qlAQh3BI24qcks3jSTMLNjttFLgZzRea9EoQXf4F28GXXfrnRWi4F9L/M9PFg96R
PiAp6yrfI2zhfciQWz6ND96PPLV+nj874p59Nw+uj4cMgXL2lKFVpI42J9YjyHjF
M8nz+S84uGVeQiHkX58kI1p3ZDhh2Cmanu+/mhigj12E3+OisARFVDrMDhgP2Ceh
qyB8zL5e7lRCUxqsm4bgdQSKAGBwNGq7SJvaOwveputOoLw3vPFiGm9lc3ctfY3i
YVPjyaF+BJQX2ZqUW/33q3TIjxhPmptnEk2vzVE28aojDVpudTCxCgGylrmMI2qE
xaX39FqAt4Nr5+Wu8K4Sc9+GL6sXhuL+OOJJSeIGJk/LZZc6zkbsjbC8myrB3k4E
3cOZqNQMUhStq7xK+3QAYiouIn5HkSYkg7mOmayYLAs8KW7vMvT+gZHjh/vN6o9C
bdH5MKcpPiF4zKxm/YgiF6QNsibmSV3uINHuFyWqKbR5VhPvGrgYZfeRehTLR2Ue
ebv6/OCqlg+oqv3Hsm+Yh10Dl6SMpPLkaR6Hgu1+Yq40TIYt6cvgPc8KYAXUmkdC
HCYe9wkshvkJIOErut6bugW4rMNCCXaQ/6CZXPYvj4Ryl6CLSMpq4tvMOXyLD2UJ
851g8nC3h8GanWI3soBkX2zRFObFSXM4xJhU/M15p8xsFAhZIEtaZ3fhCrD9Mc1q
olnCKpIWnRM1AaEoc04WFNSNksuUQyp8zGMaPN1Ny4AdJnoz+kbaHCd732ApAgMH
9WbbsmGUJcVtXlbQPSifmc/yHm3V6ep1O8APoiz7tvZXyhmJF323J+3OQwO0D68s
oMjFGnjsugBxZbc6s47L7uzwt4l8TPgMqy7EQjaqjI85DvQOGju07oaM+iLvlIIx
Hq41MuVKYV47eqdQEJx57BLKA9j++pC+J2OGicbmgt37iNAckE+GaJlC1b66JIrH
1RlFquVq42SbpIaTTkHFgXNYyNFCM8iCrPickq7zVLalelfOUZmjK64o/ZofiPE6
A//goSQhZYG8kTPDxA34EOLSuZoWFBG2ZQt1xDPCyEIE8sH3AETzLQu94xpydKtF
5hMLFzrNBTACOMpy8jQ1Zs2KEEf/3aUiIBtZSqBAjdityXVZUTgQ9qMjWK4moESc
UUwJ42zKO85WXi6JcYW1O/3dvga5DnW0cpCL5c04nW58XLslMEZrIm6bm2EDyfyS
DYuaV9Ue4Hw/Y1lgr8c+JGOkncLCrNSqskYWfoiT29tlT7sWsgf9pPYYF6z4jdrM
SENbaE/szfjn99tLwhCUyfnTB7oYQNlo6WxNwkkQl3WcM/GMBpr+R7Pg7lJSosbA
Z1BFoCaxO9T7CKIRlaPsRqyQ22xVdq/DfGrswdUhcdKr4khHkDjQoJLRImsZ1RHr
d0NpOyxKCeyVskhYdvKRIGJj+VW6xFGy+f0t726QKb8E/EOl30nMHMYbPTRwKj9r
EwWkZJ9zs+xB7o136sh81kYoRlKua2J7HHw3xLcRkWzBEJex+UAafwThNliNprzK
noM6npTA4v6/lOgRqy/aUI6xblaxHDKcQ8Xv4oLFZKP2wJPI9C3EAs/wA6yCr2y3
U7a4P/+5AKwl4O0PGkV/HEHpdUvb3C1mnOdeMrWuNw2KZiyOIBQOx5A8ftx4PXHK
zkguxdWFavjNVvDPYwP4qEC9Nz934MiT30tJ3xwawWFey1CRjfvOH3PzanBwf0G/
XiDLhInczKaBxJg4jbpWiodjkBRfJAMAduM7RQJ9w9Cjr/iBDhD0zqMWOaiYT0Ai
n6s+cWvnbEX0gCEhnhzpTOQYYU1grlV9xPHfUgQ34oPjcG4qW+VFu/CZgAyWXi9a
72FoyzgHa1xrnAZ1y0gDaTmVMGINajzrkGacZ0cNsy42jG7RVzdg570p3Lflebb0
kXYv21YqgLYvRj1vsrRHiN6C5di3a+QK3vKgIAEgbbRrrJUgti7UwWYzUJ+1JjY9
/XEDH3XGQBun94ICjxJjPgHc6XH/Xml68J7VQNXcNHV3RVwE6BIxdVbPRGRtelJm
xNJmyjpqKKLxgzcRNR32CUW1esg0M8IwW6IltvO7+0dBrKI8bQhd1W2B3yMM5YXQ
qiLvVY3TStGexaSB+gZ4M6GGCc+LOplPg7yQDyHb38LHK+ogQ1j3y3+fjHNAmouI
RI3Ez538Et/6hujFNevcJCC3CWzTiexzdjd/5lgK2wXtNw6i6/6YaXJ6AAsk2VtO
PKSsAy6YyPkzLiR4rhUWuQ9XFQoEKHJ1FPlaCseszGxSuj8+WKj+bBNiEvp51jo5
G/SzsH0Pmruu0NRvYHvRe5xg83cKwu5O6oEKFOQAVnIvToGs7AR0suQBjY54eJzf
4q1YYn52uNg0A2Hubr+Q7AItnqwZfgFbW6XWUmGEKjb4dOpInHm+yMvK9H/rct2f
6U70NBgyT4ha1yYHMYRHTFHOSt24sMc0LCQ3NOul6iSs9XT5YQs2RBfA5pS/mi7M
zx2Z8MdcKxR/4v+FOZjWcrwe0lQRsKNv8pr1wIC3fJSikGGpTus0RJ5Xu62tPsRu
6Pcyc3MIwZnRzFdcnxGhscdQzUAZcIpRIWM206b2MmSsFhIZV9xPgi+S+xLLuKub
GXTYpGX7wu+iJ0aeyob33BoPRhNbvuGbhSdv4r3F1EB20bQjHnbn59DB1q5FXk7s
VsdzqhLadbxqBlv3hRo2kvWLZO9/o/EtVvEXUPJGY+jm28+xcZXGOo5n8dRlo+qg
IPRjMKYRs8OaFcuj1qlFkoY62TZT83X1D4iw9vds3FYifH36/2GKMxZCjvZpSWWy
cBYnx8+VKykOBlqbmEUDxwQMRaN4lwYWMlXc4UN54j338AmbDruXDf3zZ69CH0Gx
O7yYxiO+8vwDJoWrWD8pLgveStHAfTubCl14ej2aphfjRk7o+7+ROXVm1HX6p8Uu
3sxl4nBoycyvF2mdnTqrFnMx5FEvMMk66TV4GJyYbBi8UaqTYkEg4UZYK25Wdipb
DIgfHNomHVGd9adcWAcAVT0QahO5bCoZlbEwzlRe0RHkqoPkayvrvbggyQcQGuJJ
YZtWlWbekqVyoHG5Po1k+UDoV+KW9ymIljwF1O++/AhAoaCpTCqRd3HQygCvQ9N3
/l096np7BDieDdgvfJ4HmKqV0gozD/lRwbjmDdLpMiDJ+8O9SUx8ev5buZ0gjgJX
Nyg9tK4SpxSMkPSAY7NfX68w5qIvL72Ty/jCxdmHLDorbjm+dgaJ8VpC62WsXC6H
neJzFxs+iNshB6UPfRJqFCSEdNdcexF/Oa5pQPIX/YmlkBsBy+2McreAqthcQAXf
yjRKC1Nu8qfoeJXLO8+7flfLw5Wgox4qOzQmgENDK6bJR2n8tHX7XF7se4thngE0
2YyJYjUIwSfef0MVfH6uwaz7+7qaXJugUe5enr4+qrmQR5sNPneYw94loGplVfl/
fxmCmZKwPawPlTg5eiS+eyWldhZAt6FWBzfofGU9tFP80fxchFvOPyev3lOOsB+S
lZF77Qh2ewC4IrfXL/gwu5Av55Opd6zqeWA+OYwICIjL0fsQa0ubwhutVF6NblmS
URmk49+1QxDnmdBaY1dTXV1vDWFY08Gp+BcqvgONhAoa5mOKqNAeS9W66c1V45fj
o9ndib/T3B4mjxP9lv2cT5HG/f6zCn2jC5lRP4xK9fMV7vzdhatZePXQ2tZ96JzG
gBmKMIrWrMtCwRwWZeps29Mw82PfGRIgYXoZnwE2N6/rNtfF7lNqAs9zl2n/Rfyu
PqKBHUKjTcqtIuiGsJKLc8q6aRiAVYkFuzAIctWvq8FA2mGbMGJeuiRDUBeFbOBL
dpQAilYakTywU0MDY8a9GIxyNAwGuhMD46IJxpbERRZwKF4o8nzNAOLasC8HOFg7
7mxpC1cMyrwcEHqvcqDL2jdtJZDrnVFt/qDBGnOthLCCQexuAC9H7E8qKBPAftF1
5/IF06C/VaXWtefVRIEl2zENM8fjDIJetrukFosvxhNBF/NcbarFxF8wNmwyQ0xa
/XoWOrHGFmr07BmOY16oEVB/n+cVYRsltycqWpFRefzPt3k2tYEhMuDNAE4kC1fE
jY2MTrkZfSgwti4AZlpvnnmBeXZkaG/262aEsbVzIG288T2SlWemKTXa3bm4rRpF
WlKFjaUqscnLGOul7pDPTHPjPc2iVltbDVunUqOaiLv/9WtDCRoxpd4jJwq9/vzk
cF9ga1u0P6AOyBUczI3/eujG/6209y/rwQ+YnLCu25dF85GdEQjobFzIzhbRLI2+
J0LqrXNF2WkD217CcUFLfqdAyLKoD4ZPKoP1ZIPOrakF2Wq2T8UDAgsQf8bo455x
1NuTsy5jUc+1omRBMyKlTkmqg/V6NOmaxpnL9up+JDczjaW92SPy8uKtthTefMYn
QN7DvaQMafCkOjW/8qaNlK9Wr3zHAi4b3kWDEYn85YPGmE7bESMRfYZpFxFUuIhV
6n1burcSeH8AG+yAz2sN9KKH28bV0FeJuJvzbY52aBFA2afjHuAfG82DUqAK2Mmp
h/irp/LHh0eDCfhwdgOyRSc84LbfOI23nfhoFgVJtmJbw2DbrpJyHbNJ4NZc4Iaf
ONUci4xohh5ZfYiWRLiuF1lVLf63iRPwDyMWlxM4XwX4HDeynnIIu5rUVG4GbTY/
JbmLCwlY8nAAcfnf95jzCUPkfWDrkYaCdNlaw+w9ISRt70GqJK6nsjDDKDccApnm
bQNz2spvmU5gx4/HCPIk5/eYtOMweRdmAekeW2uq6fjxJy0WmOK9+skRFnKRvDzN
rl0jW1b94XOcMz1lOfmZrqF1CllGWACShGdIG325zT41IFVa8qQdllQWxI4Hf+x3
ytWzosW5G+JK+TsoFz+UX9rE4l4lgX6kH7u6f528rj8jg7cUr8h3C5oPCG+HK6Wh
chBT5GCfaxNIypj20G3VsX6bdUSG4QivOByzHztjsqGEoRrH5bVIsBRbUo1aQ3B0
U7W8+GPWwbssd8D/6FRN9r2zngb3culdZC2q+is1UhKvPNvaUM7uhuD++z3txJ3u
vqbrDaDBtTywTdVyQ2icK6QAQC6AXtU0TN4ZM+Ci8HKHDAmxrJB6YmFABPB+1Pbv
DqMtuOVe557tTKmvKUN86ymwEwGZFEKw3KRj2X4sIbk1TcCLThXeAD35cwsQ7m51
700pIopfu1pQCBgII1HWlPmR971684/PzqX7LsfHvQ0OoOe9He+SSzB3bkTbWbbI
f7tfZn6f5oUPoo7FDQ/GfFF4afggSqyOv8oT4HuE7wJK30xnqzBBDoDWB3U5dnSc
IIRpQS8eL/QaH+U6bnFwUpoTaHod06w0+wqja2l/QhcK1/dIzETS88DwdnZBeSXY
BB1zvh2RI2dy9trluKe4gewpWboELG38lKIbzvHkeUdAUJFWOGFj32fPEoVBCNf+
gXEVvA7BHkuji4O1hEd+rSKdthxxJioo0KiUDbkXvPFiCSj8UYG1L6oN141eqO7z
1+3NIWTYbrIbQdLpx9Y7iAAZdEpbT8SCUkWgf7XeOyOZkXVkmR03RgSBGiiG0Jv8
5P2Nt2wlkk1wHboz5FTn5RIPQYTw0t7WUfYJijf6d4lGtRrgXB4jVglK5pNvxyXZ
BIcM8WNB26154R3QAzpiIeTUeIUnu8yX4hd20HekCDZhiREhl2qRTFIy/H71aS1M
reFnsFC2wvt60U6Vfg/+nvIIm2NjXfkmK15HIO37LNtsuJjNg9tA0qShmcJ2d+Er
+Pdbk+BrljlkHhS//l90mICN20/rpEI2Dg0Mq1KaDxNMp1HtXd5oJCxm2NPFYslg
6+nVTh3kuaI0nuwt5oNOc5DZu/3rqRiLmJI4Tg3n23Cf8JdBacHt7UPtggc1ZLUq
qM8ASp8iNFuXCubaK1p+uthUz82mMCZnKXik0NcNj17wBIieH8WIiSAhDrHR7tLp
MMAhR+T9eohj+7c7tkJJ6mMk7fwYJOVk2mf/os71zu3jZP/carp3fTjcPlSbKw7Z
My8BPM/xRLu6idtWBMgIC4KWlT2r9kuz6OSGAJVpQ2aPxC1aCoOid102JdKzKhv0
6xbYs/QWiityGByT6F22d7d8HSw02z3NVghWc0lquONNwinAKhcO4ydp5L3aDvsF
fnRxUz4CzKEpJM9ZT8N4qRSaSrF8byWfRCWRGk1hYnYP/jYJ5/gqtBru7mTLfkJJ
JsK9rWU6kCbOmn/aVMqmmRLSBeA3nieI2f5uMfw2Knv3HAgVTN5DcR6dwPEB3OCw
N7WGcVAsRaXfK/ERkaQgsHSKm77HKhi+BSkLtEQM+Rnz81OJqhXJpyLOv9moWTHR
eoxGNcoes4wGoh+XpGiwlX+EkrANw20pq/RC+BXbrJMk6lwjXnIzQryXw0M5J7Nq
Q45ENwh7PMwLDXgDJJcL1gjOoia8NxC9F1p2f6r4k/c94DkGQqWdCHtKhsWNHp3X
YNP3GBOFh27fbEuwVt2z3+VMWsoh5IKBgij4YfGa9g12nkRyyL/RR5T5N4xqqpZn
Os/Hf294mul04u28ftkp8HO3NFPS+wb1wC9MznB1hu8Ok5qWYAz5P3pTtST34Ljh
A5dXmGJ3/PooUCc6Wob127fQdFG5AHbJGhi51Okrm9kBYwRU07o6Ll4aI58V/Grr
UIQAv4w8DeM9LaM6UjlLiJ41KBqwHyplCluW+I0ptbzQuxYfGO8uxsgIlJ/jA9CK
x31sixWG4RUAWAiNVxVxIq8Jxdn57Qkkzq+BK/eOAD2KEu2Yo8Z6/7XxWTGc2tGX
hvWADdPdhc4Bv5Z+o3qvBU3QAMVAMRwVO8HsLrZrpNuAZlZ9WsPAqopRtIByCJx0
fvMLcSYHSBgBi2bMdEjPzSZMgcT9TBVt5bLRXvB5CDo09vNg4MCJLTooJkMlkV0t
ThwcfdqiR7jVUamaQ0Whic1u4wg5GocNH6oq6VD4zQGo8BzEbJ36lEpoUNKEH9J6
hgP2vkDxwv0iRAHciCC4F48NCy/JlbLUlgxeW7Mk/+Oern8jM2kgIKd9c//bQlnj
LbnRsOted8Dmjlhh+pF/YvmYbCBzIZeHwMt2huwIQ0Jt3Wws0jwEY7k0NltEmhKh
Wx5KQ6hlfHksX1iGMKRWI/WNvuijXI/R+QfjsmOQjAnvuCILcflTX/o9VK8L7klx
DiIAdofVp+rCm+iToaCkXq+fL6rjaD1R/vVCNdu7jCXqkvooLkI+5u8tLPAvw/3W
z2Na4kkzC3kCcHBfTtb96Zo+GW4Ey2o73QQK6/OBWMAumxE/K5VUKPhRV7dJG7r7
HrrHaX+VkiE3U10ZKXnFUHeJqAwugPBQOV3XM1saGyrvYLtxd1mr4kCTiSrhIhCR
pAnvWvHQgFNb5uau9G/H7w1zUmuI1XfiEzPkLGcxyKeoP+HCV3Dzy+KGiapL4D1T
nEbxN9IVwOUS4IrM26Cd3ZOukWrMcS9YWqxWgjDuW/qXeSAd704DAiqj27Hm/ZiY
pDNIvSHvKWiwfmuKBxaO5eyuVw4CMok8cSiENYm44bca6l+g3OER43/e3ZBVjz7Z
hCek5xNHslJRDU8oNN6i1o1RuQFRwotQHeYzH5CqhNSDBifn7ispJkZgKcWuXrlS
KW5juT+pg7WimPDHOAUdW9xHpt23VT6ZptH86iuc8m4oXNSM+LwDQM9ra+MwGt7w
Um9vBJ2hODPN/LMfm4w9UHNEbzhxw5I0rRHdq7uE9WjjUHCYsEU4h6ydBsCSTBiv
534kSP5mX7lS3nAeyrDcpN8g0y+MzvcjnzyU5VTsNR4h7D9+nElHtbLtm69qM+Ot
Kdfp0xXWLX390WS/x8o2nR92XEgWPHoyFaE+wFv0bqDF+7M7nlB9V/98UBgcU0+v
v6BZyXEjvtZzmyW9lW75n2k89xTqAkZ/npUs1fsnqBghgAXbDPS76u0N/MfunZis
QgdNJWZGQuYQWeUBa05Dcqqtj29nSZFieWPT+sPB+UXimuxt6Qx9AfTonVQl0xno
RJyCTx/NrHIG3eeYkXjAWBJdS3L/xJb4CKXlWAXzOXE3OLFqssJNzMn4JOdgo2eR
tM5PQQLAFnqHjxMyrrCFzI05/pUi10NUAeFao8IWKVUWLaOMfx9pavTcveaS78B1
2hAOFiOHtXlJcAgtaLEUroXHEmDil7eDBlgfurW0Jbv7l6rQX2xpxzlelP4b4RZX
MRqXFuDGjMIz8ANIKylEG/D+rSnODXzUjrJUz1sh2qmADPZIfAYs/OKoSandvfRR
8jdfP6p6y2HVWtPTWZhnX8HSWmF4z/ipQuchnGpRLX+F+y2p/BwZr7IzVF/SEPlK
XHvd9Kvla7DxfhGdsOljUkTrFnevmwqZH3XyVRsJkBgF+kgNxu/ePszT14wEFVmb
PrhG5E8wDzNM2BLS4MgykHvwx4DCic7Jc+owtj80w7AMUNlD6CgnlvY8Bj/jZW+J
hKQeTguVaE2C7dWS/A+PE0HEdSijE/p6Kpg16vEiPDBuCE4drmVaaRbsrIT4XvLl
uLyT0wEkBo4RDj3Tz/YTP5IGKKB/f4H7b5XSkzAoyCF2A9T4t9who11/LInX+a7J
VUmw2ymli7PLWZz6c0tjNeD+jXg/+c6IleDnOQrTsiggP50/LsNJQVAJuA2u6PLx
EBpPBBh7/R/WwZotVTOneLIvvNG41a9NwoWIPb9y/RlE1bwAI2D1LLdeoD5diFEg
PD6RGzdzhPY8JDNF0aupK25RjqjVE1INQanj2HI948BUsFRR1TZfVDu5MjCECeLH
cmpSTUf7cJ5Sbmh9SlmMSb3SA43pe/c8Tgqhkpg9LWxrSb5YOf8Esx/W7S0hnzmQ
ZoquyFg1EivMwBkDbJZD9iLtPcXw8M5eh1rwAv39mWB3rPHU0W2Vu4XVotNwupk/
+6prXuLN6sXkK9hOfUHBCTVDTifxRtuF4kY5IqNLY0JxqT27o6Tfm0bAYt30aw3L
reuVL/cdgKI2+LNQs8hNNq6YFAAePyAHitARoCxFs0rKbBNeHhjs3qMlXmWCVfNx
nhD83ebSv+4eFwOL/MN8n5BLGz4YlH54T6bxh1EKiWY88grohr0aK2dZ3Pchot29
OftlgddHcd6rlkxlIylJg5mtW675umjxG7PKjdGwrT55VTQp3WObIbeMWU758GxS
ju2HrDnzqiD/+Z5ZxSG5JmUVqBuBvqPSZKuKUiWyWCm5UvvaSyFQ6GMBYX650fBZ
m4PAL99aFFDl1O0h1Qt1GsKknYVTKFxKDg5z1X9fak0T0bFB4aSEZHFBjEvv9Inm
fF+ORo1/pt0F/CvW4qR2uc4RorVxnIRcpHJ27WEbrRAXxyzqKz0pOUVPCnclhWeQ
qjJudamYb7ECKzsGkhp6BvcKXJUyBdNZAMVYmOXrj14Pz6iU45THxO00zuyXPaE2
Fa4Fun4cXAt71Rr5Sy4g6ugAoB/Ap7nAExXkf+IeOP5EGnVlnGD226JXoJjAeopS
WLflvMuFIgMiZQFq2zlfkh2P3HkGCJ98/0M3S5X25flNpZUXWgxnvx9oT+v4jPLQ
bGPW3NdBVb5eVrge+AmaRg4eWuuJ6gPxAv//nwuWZf7BAonL4F0YOTicxJMkth9q
RpIiN7KIouCN4cLHUKHxWhN3c2NTMmWGznDseEjDPMh3k1nW44npUlhCmItgFXFR
ie5RG4+eSp1aavTGx64KxlWDWa4MgFYM9fTC8b6IuItJgsc9agigY+cDup97IDTA
KiLq2L1VXPvuv8p8kms/BLg02NF28Vmr2UKFUFsf7VUmNS2EKN2P3mWc475tw/+5
JcDqyrgfClCOU5OOAiyq7BblK/5QPnun0KR9nSxY9Gw/D4jsZeXqjAP5ygEDrqJz
YAcl2xM2S2v6pRUYeuxdb6FOp11Zr4YCkFYOQON9OrNlm3isSCCIV7xDU3OhzVHF
09Aiuo9k0G6Hrl08orX4lHS2Yt7cKVQbvXjiYohrL0Y2JdbVYhvznfTdFvHY8unE
Dmh8i6mC1CjBE1AdYtQZLlEEfSA00fK+SZfDI7oVIOYrTDckKMgfNixbFuD9Rp/J
ko+5NG8tn82x4qgIXwruJpSFLhV1Rvz+WgRK5PJrg7JVwMCrA7PaKKQurYY1ISlb
ybxpt3fuCvqT4vp60yOy1aenTN2pkBb4XGTIZT3rEoTT8XYwkCiS+9AThtNjMfXA
YBJtjHySm7zF6bR1XXyFRVtYjHmXQ1KgPE4xW8ZF3oy9spOg5XNDtgMymbzmJejW
WnE99imWhCPxxEU9+PvbGJpHel4Av82xv7GIcqhkK60nwZpL1/j/op2MTvEk6/gj
3TNJZUxaWTiZ4faD9mDM7/LSUPUX4NBKzooPxYMPDT7e4LMABbQYMjoBc5p7d+wJ
mlgRb69OErksPTNrl987Zo9rvTQGWr4UyZIBYU1qj79O2F+iWz9oluFyVbpbIPoT
XdNPpkcxBC9rdVMZQCNRanuVrDQPHX2rPvx+UmTqdQjAKVH1z+zg2fy8Ant842X0
ge1xHlBOtSP7TR21bMHVxHsK1RVeK/NSJg3mEGBGvc7uVKyo4+bVDR22Xn136sN+
9KRu6n1i7tbwD72qPONNKfxFdoVev3wzhFJMomXv2+YyvM847WKZYPQ6MJfR65lF
0N5eBSdJCOQsuKv867fYSRJ4MPJTtZlLxlMCUX5M9puhv9fgivHldW6tKJ/xBj1z
hCPpdgrwp/OMMIhTC8UIDssP1p5WVj4W5DD14IU1CUrfxQbH+G01JfvPjv5h8lvy
sY1cZgIW5g0f1XUG5bJjqkn5n+b5l+KzDDS//O0T5N/TkdoJ0ID13JnHBNQm5XWT
I3EN3mz77o3F8l71acS2f19mfvucPqg2Q488JB0Kf5+5MXpGa0x04dqev740fs3/
D1QhqXmJcE5XI4KbpL5Wjrrm3M+ICh6Fx5cr3RCyxREuXGLf+ze1367QjSwko6U9
JGKnWCNq0pRG/sRLGW9flBjfxBb3Xzj7etO5ZJ4wvEu92d5+vwVbcMnBEM1CJXHE
LCifuGQQrO7KlKlFMqIN68RbvrQ9j+7rBApuypOM0ZDiUryiBr8AoahtqS5pPsXw
ZxN0KMT/eSBOxpzufMzJGtXKhJefEbQbLomYMpBYVeQ=
--pragma protect end_data_block
--pragma protect digest_block
+v5n+UUPQk5WBb0DN5bQRxuT2n8=
--pragma protect end_digest_block
--pragma protect end_protected
