-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
a7j1YEgqqv3ALDNkE4ZlyhDC/SQW7sjehnEv8RUGvq76hMk0tlHxgUr3bdNg/CaD
I3nuurzIIWuHgOsK3lRYWoyjkMvsOyeFHU9CwvX25+xN57/RI/lDKYpoLGMXg+QE
kqhF/ng42/ChEcCh2uiidiAYR82gzf8ZW5opxyGOyrRmCQ6/qx9Sgg==
--pragma protect end_key_block
--pragma protect digest_block
AURWAgvDVdHQ7IOywgrzmR4d30M=
--pragma protect end_digest_block
--pragma protect data_block
7wu77jYQOCoFRRUVEI+zS3bjKMO6A5ytIMaJOYwKOq5sTFKP8yilPGusj0Wr3nk/
N/l8CfCwKoLlACEMz2G8pXhs9rO0INzvsjsG8Kvv9i9ImWt85C1UTZJzMS33T5G6
pzBZry9NkZ2rOQHe31Ra3Z3uPeNB08xYzaEDcC/1TPTaJGGj1ZjSgbMvv+bJ3D8v
pOcCZSCEXS+14RffxEH2eR5mKDtSS3h7gktm1/hFSZsKzHL6Ux8P/uXMU3qjaO18
uhzzNG1aULuVCcCU2VlDo3bNFXFBYPqwtaHZtfjT38j6yh9LyhTWWsAjv+B+WrDw
1W0DZUsq05hnJFVAnm6S2BHjYmSf2qVR3Ld+XBP47t72cw57PiM6vSTjLwURHLNy
5PL0qt4Bpfet3pDStUbWUdDLR3qBRGW768yjA7vGOKwcynCNK9/HKqaulJBC5YvX
4GBPnEpOeODz27e3U+lKbi7WVUfPSO7uvwQf/xqnKsSiE3dIowzOGmPlpiM8Ifkp
6WkPk6c6eN4eKLfB8J0yNvy93hSx1FadbJGScYAa6Zwg7Jp++qhWhOQ15dyjJwCy
L+ulwptAgnp23S+WSOlw+jro9GpvGRJT/tY4sAdv9PoeSBYvgB6xYk7QFE9ato5d
EEGooed8hAW0j/CDM/vFyHhZeEYH/MOXCazjHhxBsKc79WoxuFpeIWlXv6fmKo3b
J/mCcOmG0HeJktUJM5dyz7hSQHK36Rd2jyVBAJzo3rZ/SIxEJthitiDN0ex/UdQ7
bePHIn/VMx63y5xrAzExVZTi3+mCmwS98SCr15tDY83Qdo9kXc2QXWTp6Kr2CcqW
I5XJXheF3Jqirq1SxIJ0sOyaxuXHq+Ijf/6YECfBrlYa68R8mWrNGi6yKyGBeWvD
aSVoq06cn7uj603Gknke3cgj5P1rVB8kj2Zb7Vp74YzEZQBu+i3S7Q36YoaQzhoY
M2Zp8NDQq8V6wvQ3zh4lc/J3h4J0Rfkb/ZHOcnzHLTmFbNRjs80DqqB0GNlaTbVw
negCTXsvSkj1ziwSgxtl4TmWdS63SA2IxKLtaCodrMu9s+XT+8tcIBYlDXMIGu7u
CdGzajVBaBEzovyH/+K6qv8kM1i2paS5CjEOwe4vpnDehEduoMO62qphEXPT4Hb+
+5FeoULHfXNuMgjLAWM7r4F2B29U3wZZMpFBbbIPKXbKET0dhCU6h72mBRjnxje1
vMG4qJ3CgwNgWHps+D3dNvYAKQ+JjYbQM1NNFgrozGI0qmR/u0Yb9GUM+wW52S2g
6bEq0iRt4vjl6AKU7DPt03AJFvN482u7+fDhmQBqyxvzNcCUTjmrrPF+zYm00SWL
1k9trY7aniWjj+YEED/llW8nmHJMouJ+1iPOb1/Fts/S9MTK5M4Ra4uf81SMY25e
9sfKlmOSHM1FdynKYLFMc8F6+W3MRwEmnZ0g9Vud9+CIPCaS2bAMbh5riuI2MlNh
+NMROGXjRg8LKLB+tC4220QCe8FY1Nf7nHd1QUC3YscAcygGk7fFHYqpUbj37mM6
Eq27kXF9Tm+jGwNBBnBSwwrOHXgvA2DguAQt0E0eu/usZCwuTUu4B0sIZX10SBXO
URrOPvBgkUQvVj+8MFsEHTr4FflDry7ZOGDr5A3o8hYYvmrt7IzMroO7+SXeVxKK
mCliBPApBa52IcCTY6p++7mwBb0i8kRdTHOWBzUHmAVDiAwE6A+v+99grY8UuouM
jvPIcydILHYoWqV/DXoxUDT9VR5QmQRWaChpIfqZosTeFQe4vqe8oB2qhKPL9b2n
YMTfo6jbbfSUsNiV6Pv3WsNM0Zc4cwuSzxWBsdAxIuD1B1S6wqLYvXE09x+dRGTJ
wpcg590XZLbUkJqN1Xxe+nyW6/9jvKxIMa62WFrFtkgP+GrU2I5eYhFUKRqbfbMO
8tjD78p//kMttmBpIcX9PuHRHkmc2lLi1CFG8tgOJyJF5rIdTjm+mqW7T1d9oXij
L9JraB+kl1jFLLNVTt2W/KwYocnea4h+TE3bxAopxnUQ0bdcgnlBdMRWomnXiKLY
zGz/UkJ0tYDl4w6h9/eh13eYBPcq8OUMRsyzDLUjf4liYAoAUf4KbGFZjCNLPL/d
aQ4ckB/qVpmhzN4VLdvHzSK8wYRTTftGgJsYI3mDc5IeBOeZLzd9ktCkfGEsNSfO
I0Up8FE/EHyVMPWedgbhO0u/NjY2wMiRaalb36Q7EhpgwxBUS0/f8t/PsmEP7Hy9
C7hxgTG2HbILi3iLoN2sS0D7Mfmd2QeBChSo9/Js8f6eVc4wZ5Ag5ZOIrqgd+exK
08pHeairuzGQjwkq5sWwLIqCLqIEZDJmf0eGKV+2+0OYJj3oGr5K6TqLIg2D0AxD
BJSe8Sm3Vc7Kj/xhp4hNAH+tErtKNXcofmYeVQH84ua8g0xRs9kkNJ+oJOJmvM5w
3UAW7sz1OUiUOjUowyzW4DjLYdVUx9kfVzB+v/KjNkhIuvQecD4nUQcCG4AqPDqP
HATUaWnrfcN/7ETWt7swsSxtqMqPWn9PQsjXuzo9xyHR6rlopQJL+UNdG6xhWLQG
7zIIzaK6C7PPv/EJWiWgoBYilckeA4nYIyZSjyVRaU057FXjWJ9bR2+xkLZd2JGA
5RryXvr/SBlAy2E0+xC/K4IYPYbN7ZVLcw45FY/jIavgUFw/jIxJ0LHbkZ8XNhA/
AvNrXGW33SWh9AK5lM/NobPffpTpadhhASQuitsWFImINObzA04+8PfN1Ajf6gGJ
WiO+k6QDqdhJHYcHBTMEHO58Rnmkr0k8r+hmVxOqOwIuShlY2Ti4sxkYoZ2rQJRr
DyRfh4xBIt5ModYvErLxDXwHh6B6E0XwBbIFhkm+7LUaUQmMm0JDSTF1WzlfzRW3
X6n5CXIICx7aA0TG2O7q9+RTcalNvVtgX9tQ/hvo/qTqfdh/bGCk5gzTVYj40Nm7
I/GoUWSGC9+s28g3jLwqIABxhaeiHl3gY42CsxW84QUCLRyBovYkkVtnTmE8FvRM
PbKoaQZXMuD4gwtZwFsK1lEiWeyf351/TMYukb0BW/4K5M7pVJq/eeG17Kp14VBH
GRrDOtkJ15q0AIRLHv9+Q11X2gK3hBz1YxGDJSTVygWLJJm5pC/kqOs3kGu7TPzT
mksnv77fO2EL2dJczwCJb1J+vKvOA8/DqnA5DDxhIzjj4sbrFjQm0KCadRsS46ma
VEqwlRTvpTfSFx4rUW3RtI6l7c15MFur99SBko/4E+AInU1UtRYHmVBXUqXX01Aj
eetyTHVzd1ZVAEV9x4nOnP6Yb8O37oj+34R4qi2QIJcDdIf/g/GgmsTqT8E2sWPN
VWiLBUTV7/OouFgujpZLWXL0zh9Gf1vFcukKXlBwjOTW5bG91SJF1RzRBSk5duOk
oaIpZzKx/7Frt/TvXtS74krqVoO7jJedc4M/ROdgiQtXmECZJt+l2UC+CscP/9D7
lBDGnOsf3UiCxY9Hae6np8Pc9q1Y1AUg3APaiNLccFii6daUAT/8VooUkLJZqxM2
rnmcnRE1pENoZZ01AhUKfI8W3kO2J4TyqhEog9UXJ8bLWddXsXjEqAr4BrfpkLyb
71bFABxixy17yT93nH/Mn3GR6D17SRqUefZCYzngo0vPTPLSkFvOkFtP4skYt/SN
OrEOb9CVSQzJacq4CSXKctB9OymErLavyqECmLIbpmEHUxlI0SofbcOdVm0uFmYI
GO3dRUSzg/WPlPd321bvgaTFT1Kmxzrz8zxosiE95xQdKDR8L8DyyNr0hlFCb/KP
slYPkfVhrmtnmlOWGfST6WOsc9iXTp8ZpSs7h3v4JeODjjZ8So4gVZIxqhmsiLrW
pVenVp9rMvzspXcnstxwRgEH6TVQTgr16xOmd/CU2bKve91U+iLN2ASrvyMw4FOw
p3fWseFAz0WRLYwXpuZP0RSVfcEKHLL9sojrqfb1MNGyuR1LJc/Hl4ce890psDtH
Q02bEfINPo4+irXKWT9paErVPtxeoQ7/4BNHIAHtltF+vEBtF8N/4pe2ExIfq7K2
0nTwpTmIfMFo0jUCyUYBrgus3PGrPEbrIiJqnUk52gh0SHpGhWHvwZLxbhM/rzWM
GRPtcSh+pYRtmosvPe0O2C1qnwaPEiHsnmkdQ/wG97KvnBqykT/U7mJppy5naBgB
Vzi6Cxpk8X3Ct7Nwoo2UQSVhdx70h6JQJFpEZEiimOR0Zy/h46CguRn5Uu0BFLNs
XYcLgaRxVz4046kzwuEuG7wGRhSAorsn/k1rhtACk0lH8Z5m/11xHv1NzmBUzXkt
4ckuZ4l4eSMJcmwdWv06aUrKchEC66aObBVj68xzI0G26ebC61A0fL4SjW7e8KGp
LWZeIqE6VW2llXrh9sjuXqL2urNUMBkRiAJqDQkTXczpDi2kcSNERNaOTjaQu6mH
BPoffMVBtVRAbLpKhoTtoW+LtesjhwKUIi7p4D2rygHfG9FKDInil2bVnkgxycNg
ATB0KP5M5UgVrSVxaZ6p1XhJIxNC1ZS6M8akwgcyQaiprbE1lHpbycicQuHXAC96
csPF8gN9kUJnnhzUmGoj78xHTFsT1FHy4sPFdV7HJ922epB+fjlqO+qRAjKKCFdm
SRHsx2WE5DZn5XBQLtjSu4SGDk9HH6aYnZZNxQFkRrHxUc+fBxcPVCwzAvz0f46Y
ICBZnlUuw3ZdPmqjFdGrzd/DbtHb2Knw+ZyNzYb8twNjc+vv3YwOm4Jb5Zhhu6yI
hflCaPUPM2u1+7X/0ioDsQiCYC33e8XVAgQ/qPPaLIZRX+MQpqWtxZMbw1Pb1Mun
170zqWUBtf5vkrFMPxWgYt1pWENC0aSOwz6T78sCvdN4M1/DzWPAvIFk3v6s9t7q
lR70yogn0N1qp6nACovb/QWUS5e/vDoVNbGUeVEcup6lIGHeOc1K3zcLKqnWuEhH
5kbICgq+IJpo54uKKDyMF6PCvPcNoBkb8AnZN2m0VvejF3Vg00BLYKzdOeCo03Gr
XBWsTOQiF8dHcpPFTKP8l2d8vNoPpjefFOsATBETKLV1OxZY5BiiJvSNmTS+1+BZ
fwrHdzmxo/ayKcBy/x1xOjkx4rCokjS0M1Chlzr7905tOGEWfIGWU3iH/2OEY48l
Y8dX12aJJekMwtZFZskKtU+HJeQvFbBaADswEuJnnlym7TO027IrPN5p2Tx0EB0/
YYXnufkRIDt6lu/TIYR4TzSAd6+x61JDOp2O0o17Db7JYqyt4iJ0yKOEaun+wjeB
40u/fbSNqd3Iai8KiJxqz2aJTYWNx6BLjnbid6zVdSZAdmjSuYDdryUr3o3Iwt7o
ehh/5PxDIKeYDjO2hdEU0rax/qKykiiwVnLk5kdksRjYqZxgAyCRjvFN/mMSXEL/
XA/vGrqaqOXkwT84G+dxopX/437cDUmAyzqKQxJ8jpwBj5Kgnn8G3yn1O9RUjr6/
3kL1XbGA5oTeYehWirWx2It+L18077USJcjqieISxAbaJ0JbonEnn66gnTaI3hwd
t24wayRSMj+No8bUK0S4pu/nMfNMjG415iomrYBxXFSLfS8O3nwIfsw0Xmc7LDrA
rz41K9aFbppxboroJmzIZi5Y9yRDLh6nsmsBNmqanyZjSeogIg4lAFPqGZiwLQ0m
REkmcuIT2Tc9eYVmOntHiA2FmrwPBE9zLWADkpwXdtmLt7dYpAFtoSa+hFNNMO3B
vx6fQGUstGYlqQannuTA2f5f+OUNRNDcUoMOISODDgZuYTd/j6Hs+xMW9FbDDf7e
DapM+4D0ufnwBw1EkMV8nka3SuXAEl+tjxuFmQiw6Rj4DCLbtleUm/48IGvI7TsY
B4enZVrU5ppOswmVZZ4iJia08KYEPb2N7tizhqLkb5TCQ5ZjXMdMdLer6p1WybRu
Q1wWGunhfJckrT4T/EDcHopmKMsPikTluUvtgHP7twE4Qd8T76r4DpaM9mh7i9LU
cIwSHNYtqXCrD5qXAx8CxRl+UPb4AjMCxgoxOE8RUMk3nVIFAfD1qCF+mR7Su8lE
iFIY3aVemFIjk6YIDQRAJO8XszrGF0jWWWZ5A4RfV/fJT1xk1pORW+AGzLsk0yi1
tpBur6txMqf7axdFtCCh0u8CHaPxKI5ae9CGiqx4PuWYiBSfLxGD+ge8da3ED5+h
CiRMmIc6ZsofKCnPSkevgQISp6QqpbZ7rtgqZP1P4lP/KFDaQpugR6VTvsYIa/Qr
YzZmHCZyq2W23jRchZ/IFqRzFOxyIeX6I1VBmaQ/OMyENAvDNZb6ph2hA6KYk+zU
XniOpwL/uJVEb3YgG+NS6zzHas2NTzniuDrJp2d5mjSpaZeqiEDCXJyLG9EMHDfC
Tvxqarf1yg+xX2NJqpd9TVDkZ1GelWHmW1nHSK95FKL1TIZJIL3GKloJ6Qq849c7
FkQvuMUD1yZh5Nquvdw8TBFpOlfy2l7p44JpN13leX/kfCVqb237PvkEzNd9Wet8
pgx1dQTjEFoVpZo54cewyLX+VzE3ZvNYaDmwJoRjYI7ov9hnMfXC+ltV8hn2BV8h
J7wQg/pYihpmka1TqXyFCFk7rVEM+AdT2SuSAfcrY5ZCAxQETRYIiYWC1AlkBlkZ
NzHhnTjSP+bzWvd0H6BodajGx5ooeJJNPihyy2AcRbnCPNYLLg+AQNvmAqsT0oQk
5HCdZTzfh/9qKEmORRjlALHFTBXiy+6qZk1j2kLXIF+MS9/Jw041TcOQN8sUMHli
VUXohrb3Zn78B15e61qUtW6QbyIss+QlPuTtllN8edBhL4lrn0ke/LgewIqUi1SI
CXHEk5fJqcWm9dercvlKytdVbFQxf76MNsW2Ja6Tcoe7Daw2ySlxD5/sLzs2fvj+
GHWHbc+Y1qFDZnxjQVAYMamT2czsU0wPxmcMLrveQYY0BB7E8nNzAXQP+YsuML6P
OIBTeke6WOAQPTkMFR9sUDMUaIOgoME8nltyBwMibzTWfCcmBF3dFy2y7fGiV2Qo
Ij9djhRSXYRB60ByYhG9ZcBwULiqaE5uldM3Sx5Qtv3YkUZN+m7uMOKQ7KhTfAYQ
DQ0XGY6Rx1Wjb2leWaBAMTcqTS1hqnYH+FuRBc/J3VqzQhcZOXieF39az0d5YyWx
DhvJvSx/Nx/ktyiJF89jA95cSi7s3RyXSIJIie9MXBZ9w/jGBjF+KInlWG28bbtH
WYLvxMqbx0YXzPYmOzlZn9Yheq8Ruw9CD8PPCESdlB/qH8XL/imExX751TMLvHjA
uVYomh8+Dh4ceotSwX28cWKDR9OHjqFEviZwKv/jYBRZPKGmdK69RU/22chb+PTH
cIdhpQ3zuJ5aD2gblX1QdRsmeSTHJYpMfG7SQD258K4PvJsK6L9KwNIVNdqLMZzp
Sa6zEyH6/OmINfuZ51QzWMddXFEkLS5Z4SicYUYTK16ECHYhxqY0o+HDos9xZdGn
BCM6ceBOxhrWHA8MnGO1ZVTSCwJt35rhoe3gNc7SU7C55FFtA1xGYJvEFjgzAbO7
ML8Hg/+9fH1XtsT6MyxHUnU94rol/2d5cOkG0Xv05vzxih9ZHa5AN30UCXHXQ7Ba
cblyuNMTBgWPnRabaQw749nHAuV9tLVSjfKSW9YXye9xKGiQO5Z73SS9shqE+0if
HzyoF7jZHYXPXqY2iPdDGUZybPxq8e7Up3kBGXwX5wiWuycGETckIgfogXqUPHUz
17+8t1KFuT3IXqYd4PyugeYzqbDBnlmh67Qm4Rob2HjWQoh8OcxjfkaM+S/6ipOB
msIt0yb3svZhLqBVDa8BXqNk50njVss6sslHgbMpFJnXnXoWgo2p6iiE4h/j7YHh
L8uTysGFzncsGd+VjXaM55OhVnHNbamhPeva4x4jE1iBT1JwL3fv4gdfn9+PxCB3
fDBlih1Ih/gfB+zSr3wLP5/M1TxlsTwoNMxIe3ZEfvIzcqjTHr4JbI2Y4uYKuP5X
jsGg2q7McCpDe0vz+uIbXpJmmTlWbKol5Fg0qHw8iRRW4uMEeyJ5yWuKcuYgzOzO
1NKhBkEtx1HLFNlMBUKrpowUWZtpmQmI4ig2ReJWpgzqIjcvpZJ8XMShjfaSEMgQ
zBiEXo2va5s0HUNwlCmOinRoZ7XFYRe0/IXMtyTrT/FypyGXw5qIRdZwLFW3rMiW
HgHGZS7BukvrvzjrHfI+/4lO0H7ekv5dcTnVcLiJcw0QCGzOkeNSNYCtbTuijbHH
S1pehqtr29q30Or9zRcGSwBVIUP+uQc10BaFAwtczqg2wPSzkyqW7yF6+AJNVJZp
DOtP6dnhXEVXoqlhLkbO3NUybPwn3gBHgI1sX4lDlT+pU6USoA/8N+6Wn6GvpLpn
AbcY/vG5rTkOT8SHcnwuOHQlpUsjXFhOB5zmZDvxb2u1taLZHICMH8ZT35OBMKMR
8ceY9H++c01e/d2/vA6GQz+iExjDnjkOKeGADNKn00knTixXD7LXJv4O5y8lh8OP
HIE8Pe62wpD4GBBWuLWEnOuqRwk40QJJa0sO25klPAmsGtBsjyzaNWHZXBj/yno0
P396+pZxLfXpz9S0mfTmPRsrc7UTRoj01whIOP5aFLB/YYjzH8lBnxwHPhQKpAN+
cqGsT0v159B+oHsC+Kkdx3luyz55Vh7wNLaFD3uXLoEbun9WWHE8Eitxjhm7CQBB
x3Fh5RnRWfXGIVezK0DekoMPIhxUuGNLfObnW4e5Y8A+rIFiOLLEn/VShvXx2xUr
0OVb3frlrMZXFCGSpxaHsUU44MfA46rcYyv5hiUXtBjJi94F3Qy4WAKmRigr45VM
xtdnKXK+TBPLLyFyX1PzxPz1qvlXeOiHAMg9REeQElqVD79tYXkUNXjA+EbBTiqO
otn6SybV2xAQNR/jf9uuyWWFp8QwDKmL0i4sPiYkvPqQGyTkOH+D0BVkIU7fdzbj
Krz9QggtArByrucFPe73kuXQ+VJNxIEXQj62EIQnaO+LbDmo0xXFtBlsUfuyGXSx
6LbX/nbZJ3G7cN8c/iwp89TN4QhL1UnrUvlLYyR76RSuulHlK7cnCegx5h54LtYN
pmTtg2v7++l5R2m1bMWd7rOqbUS/wNc5H78MGnNh/KWjD3D7qaUmz3FwMDXfcm8G
dA3Z8H9xMTeoMw7MFT3weDHZy0rgvZiY1fTmZr/Bw12+NJPVX/7sKB/cyHGKPwVW
yx1/80WKXZswXqFRFDAfQJLZ8RQxzG3rFf4sCGvyDbeeJEqp9kUbrjGHedrfhNty
5DHzjgyPzVjBOYoJt8hnOOkuNZrUJrvlJnn2jjYWGV5fGt5ABpvO/k/M130VL5jJ
LzdVQZE6rMiXHAF+1jlYpndyL9dHXcwdkNM8VjFPed+VBl2qo4BtdBKd+Q4+rLka
6j4RwKRe8tAYSSr3NGn/dUTqDyg87cnXlHdsqRXf3y0wQW/8OczPtesR0JidBxoD
o0/IS4Q4FdZyZT2t+vhtFyzT7bDAAkegR/BOwJl+3mp0wzdIvuJN0WpTODG/tc/+
Ik3tmL+/P+23NqYLEXCocgM9QuImks9zDw9ostFCDVazBk2OFnJSazOiYXR4pTVd
WES0ddMs65r6h2IPz93DvK+pNeyhw+bgeEGv5SxvDZUFN+V+6WpzB0Oa4xDXjXeW
CkducuAASjCtsWpRC3vnFmSgLAVGkbpA1HehZWNe3gNgyuynWwIIe9kTs2JAM/bN
KQ1CmCZGWqFk+2orw7lIvAedWwtoNoBu7Ms7mWp1X19SVkmsSWEfd/xiwhuUAQqN
Bo1MyTsjf6RF8Aur+7WMGuL3yeuV3xOSa0uXJyNAVzg2Dou0xePxpwZydA/UYQzQ
wKO/qkx44vIj3Ppt5SD8nc750oX6yqtw22dw6ZMr4aSRYR9Ol1qA1UM8Ha4FGqyG
RY6xxkrYgh9q+mmSILvIx+7zAh8vr0sHgttJDv+mNMbMXwjfG2PeVpO/p3cGqnDU
G44Qv4X2moFzr7N3oXuE5qVHOMqUqLkVekQkrqxoQlwbug7ntk1Psvrlt1IJLsb9
4LBWcEXs8vAqI7fF4sJLIaUC1le1GginE1Ch5NS3OoyQsXqJ8os/Y0XZHPdbju4k
xHAJNt+W7umjOTzVkMbLXxTg6hbGt9yzOBEtd4/eaP7EC/UFwH8QadkGNJciYQfk
J+yQS3x/jukbHQrDOpccWkbgHk+rXDvf6UydoCGAFIIGZTXjiyS+7IkIkV29xsLg
LUstgS4edJ5S9tSX7tVSIMESKiWoCk+Obf0S/lyiWrhFsAL7I4bQ6WV9SOS3bfsO
waj5fSrS9/fZNmGrIfDDoUxc2FV4hiFpMVlcNNuU/fPtIfM/nQNeYZYv3qZXOuUL
VG0JE+T8ulNqns0LZMr9rrJtAQZqdNCCVTemG1S3RzTGJZITyea39K6iyexCdNxC
z0Jg2Nprkr6WLeL82Q/0ZijJEvr+s0XrcRjgY9Ense/mj9p9V0lecyQxv1ZIeZJb
0G2QsKrkop+6vPi9TiiDBSofcn1FI4n1JQJaZ+aBIFWWT0YqEwQR79atl8UK4yfA
XwajB9Zb+nUn7U+5fI0wijQCPH4MMhEYeik2A59p4hv5EGzbiMl0cEQE8EnPvLVl
rbr2x8tW5uXAEhnks5vfbxzXi1PuPCBPdMKllKbuQ5FrtvX8B5Oh70uSENAjXChy
VEoWsW5Vg5qQ5gzut2pA/aGTqCckZzrDeyZP5oY81dqUkTFBAFXQeEzzosrZd4a9
jZZ35pzBMjeRPmRAutCHTI94/r3UU1a+hSD9jPuygFa1UeMkC9gnjQjFEWJy7tgV
Z9KpxuEs2IPEOkKaFgFLHq6asnc2eFsG+ocsW+N2Ozf+ShgPu1Syfm2bw0hyE/Tw
sF+1fRtwMQxV6GKeD+XZf4qZeNNmtTFGwkRRjudT0LdvSYWVyn8d9ToG9ceJadaS
5byv948X/vx+sv3/hYlyhKixw9u8fDi4bBXCXtG80i6d+IR9bpUGJYmVS35hF+oN
aYbKwUPlP95hgGLqPxn2JRm3kaDXeGhmyc+ztILHkOGSXIrzNn3zglCLCKGVY//p
t+mfHzlWbwdDbmfD8PUJAr4w3gcS2gQB2Lyzrqc6gd53hkidiB5FbSnIDoxntU34
T+icMfvoiEdX7Rzj5X3t6D+bYYcBJeiot+n/A5tYJjbjg0jBPO9c7N7xoSwy2l/2
Ya+MIgJmTJrmzcYs4IE4IZukI+RdXfeZ3SD/2Vbn8wvx2kHQG/2tAapKicnUO+iA
xOxhiVxgxmsNZv1ZMxnA7Dx5IuX4Ly/PvUumA5Y1xnQuS03PCFcpQRfK5cHGdhnX
7SR1ZFRvuUa4kge91C4ViuLqp4GNRTcqHrd1+9HjtGUzT6xCE4FSZrTAeKzjvMPQ
n6LQgAxQo5qwdE4yOIB29xXy0a9/J6WHZD5spxFwvVtH8oFn9u0PDohmwkNyFtWr
jWPXCq7os/nTCypypkOKw/CahH1GQ1JxHeM8l1Jrdz2vBbUBm1jbBF3HP91wUM0R
gogcvDh0J6bgTG5TGELLLJO9EK+iJvu0xGNLYPJG4pibAR2+ylCPFDL1qR5HIxI6
Tcz5AcbAMbqQ1xrqys/wO3WVGA+bGDWFYXvMfyNO8YB9dxyVMviEQagssORFxorP
Lc+IrVYL+EqKsZdr9MmL5urjgwUfMxOhnZOxCpsLIlCy/m8Uux5aSI+UaGXsf6A1
CwAyDNi4OCx0fRy0UZDY9dvFl9Sm4UI9F65poPzKrFDtVT0LXwBix6l7ZzX8DSsN
ChgJCLPl3SG9koo9dQapWpkjhdLrkB99Cv5L56soFfd/iZMNUBlNFLLztiH4zTwA
uATiC8YYGkvtL201RhSnDcigxRxhMl2eIo6GJGcsn3qH2nwixJIMBkB2Ji2T87uN
Nx/BvdAh9MBPZ0JYETD+tUVvfDEqGgBjwvagKbuFWW+Gh6nxi9xaQP8qwowgHDVs
o2xmywlVh+UIWIF2w319ilJOs2vVHTjhBgPl+bOyJmQUVAUmLhzBQRE+M1lNDnOE
Qlf4NHdpPm2PTLhqE1HB+7frkwN5y/nMDpTOU8Rp5vZoKqKI/IKSfDllN1yoGi16
ngPcfDYrCb8SO+OeTPa6p6TMKO6Jmk1HUPPRbMdq09TiymeqxFfGLG2aLiuI28XT
BGRY6dUSyRKq9zL6OUQ4o4QF0DtmvAQpnbjRzoNyqIm4VANCZ+Gxuz0eCxQU0j2H
BvSiWgmUY+rS0ee1FxkmiyFs40e3+odRV2cFICaYZFNqu8CepdLYkgbwMzjWWNP/
14Y0ipp6fy9SRjHLYhZYpKsUyoKFTx6QL9fk2cpOqkJojtfUZXfPWWzowm3Zdgqx
t5QM0GXKze3tHk/JRXbMDrx3dUNyz9djZUZ8puadN91/BUJTz2BaJB9M5Qb0TwNm
I7WgP+NfJpqsmmPw+e3lmE8wy8u3z2PDzMJZ9H4h9y2pxJC+D5OBaVNtDaSWSQeN
PLMzUHUtD5KqcH+bB98dH0k1tETb8LIzuXsoiMkeo7UbOv5BCvabTVQCc6wD+x7G
KFD5tD6k4pwi+viAcUIYhkl1wtRjLa4dh0vD1x4hHwsWBpmFNBqo/8esAuhzNcPR
huah82vHR/MZVyTKA7AOjpCCpsGCkujs08iB+w8762E+3lSuMg2t7nFq3cZy05S1
aCD+S8XxVpLu11WXOgx8ku+rkSVQlg94ez7mh0wxKax144SuC5tbRwskripXRiAl
jTOALdSoAkgb3jjdj8TusETgLZ5wAMjsscg3gMPF7fMdzFN/hodAHVAsQw+lsOoQ
RFRAFNxeC+V1ictRa4qrFp9AIjwkOfMLf0hrk5l79y4Q91I/GercTxmTNMFQqgGT
KBUm2qMJXDUSAZd4KkYU37R60RvfaOQhWkqX1X8any6+nqFIaaj7kvzucR9bugrJ
cQ2S4i8EVp15GOaU/r0DP2xfzKhpf5wkRgbZiNSo7Mvdyyq5fi2AUYOJ3DK+4yHD
U55ZbSQ0xSNNazQUt1aGufiXZjIYfZ7GtdJzrJDSrIhN0q/WMxae2cYX5vu6vpG7
s5befvPAfm8DUp4skWek5+pZAX+dPyhyMhtOiBLzUO+qi2MDzQ14Tle83ozb3lJa
I82HKi7VnwWrB70hTFm3LIli9e/ZAhpz3JhuOOXTvJxHa7dPAmASAeRD7RlerH3c
OCs/RjOmGgqK7vN3Y07PWmf25BWzWAYwpGJM1skLVScHrmDnbsG36/lGv9DLJu10
2mBUWq0pjHnbkyVbJj/Ny7jcUmF4Bnpvuufm1BSV08WjE2lFgyP0Z68Bje7g5+dx
vRR0c8iJO4CahITMGM1VQAOZWjlL38Vfu50JreyOVcHmhFk9zFV1UnUIBYZ3afpx
z+MWiuW25hIRri2ZCkW/eSgGpNfoLwTYlmlgzhT7otM93AlHQrnoOdwi6+qumQoy
EPmi+WTojIegis30dI8gF65/1WDCVwlAY6MRz5tN0olGD2zLT9di7QFlwwoQo2VT
/m5WiR95aOEPKwGMuduKGlzzYg04ord/VYnF7oueQ9nJa6sR9vsebajCIkHRbVjy
kSEvAr2rYEcDCXYVceDJbWvJzZeDZdtVNfWmbmsrNr2m2FuLRkAj68cmfHk41Bwl
DvtRJzep5Vp7AhQmc5yH7jT7KtCJoB6iZKsISXTVgFN32E/gYHc1Ln0L+O931sdX
PtTfB8UKrmm+KMJqd4cu/1Xj0viWNiF5mqjcKAGYKLolL5cDD3EQRERNKUYsdnxe
BgwiBcIER//mg/Jh6mCoiVdW/VK11w9ZhZPom8O4apOil8ZxulaiK/bNy2N4k6PT
lLkSKvaHk0q/W1ouHIqg8WBjEuwKc08JFc2dD10Wv5nruwK4dXTcvbeXjhBlviV9
KWG/2YX/Pq51Ov0ZplHsbCOiH4tptaUXY1yo0rbagooXGYaW+nYJ8G/WxaRYi9oL
OgK6rjUZ63pjzQNs+KNMu2SHkKyb2sh995WkrvCBzpUxjARiFITgfS+TJ4kQ48Ru
3jvXB6jmysTEeHSOKbYT1hLXARhW2Oh/DRujzEETtFPHbUTZ3WjiaZoxMwfQX2nh
lQHp3CRWBieyySwV8AvpcE/bir+hlm537MMNs3Yf4ydqJuY0cb7rX3TpVetSCX/Z
BnmG88RplRRVO8x9Xwu7ZFyJZHxUZcOrQ1W3mF5cv31YigwqiZ2UTABAj+Hpmv/3
65CyfWG9xdufVIjiQhKhoXt+ZKSKTH7KGHIPLNHLob+jLp0YpHtzECOL6jvtq9Tt
isNIJN6U3scRBI4AwFcQYqr47aYJAesZg2qqjcoeyRr1iiJPCzQ093uQyNNB/bnD
XcM2BCsNSyZG62LbxSFqiVhbj01YiaEz2TKobtAu1PMSSIK1EozwrIzF339b7MoV
JSmKTEbh3qD/LGh5OwxVs6mogYSQOJjd68If0OK7nupeleqXWAv2j+4sX32XVaO3
SUR6Up/BqBEZ6YnCZ+Gdhij+0ErnATKSLi8PeRJ92QLhxWU9QZW4XBo2KHAoQ1s6
g4+jrjAq7m3VQMLS9pbhY9JmNFo6rD4Aomb9sGiD+t26pKREnh0SLStPLQKQnrTf
5ZImKgYc2pFGgWh0+oT9/8bhp/VQQpDjr/wASg0pH1/jEvVgQ1yauuAJ+HHEkpAV
UUeXlhKtPcySIFawYOZyRz/QTyJZ5ssOPgt8qmN/kuVbizUhCWMzIVjiDowYPrhQ
5RO9PmtyXzo5R0YHFdK3mk8AmQpXjRPENDug0NHIuwVYNXo0RyKHzAQvJthTth1V
liy6BicXrJVc1v8CBmLqDTEO7Rn0JFSpvv62QdYLBwn65oU1556qOY78h+d1vvdD
VQHbmMK2OgyYemqfmNqEFpTUsMKg2IjSWNuG/rdhvATLPeEEkmLipe+gIOe6rkEw
TQqX5Gp8jsepuizQvxIHUGlNLlXP6NUGi9YZykWBBX09humcH23kTjggvxKqTH5e
E2tQtf1+MQq8ViNZc5wuevsF5GgKUm0VTIy9bzrzepDAWDKcPOvnVBCalZ2qMo2m
3ZuoqCXJ9TGIkK5ngpOt/Y8F9+iGVefTlSiLncRT0xh8MvYvzj090/0Dcf8JlZQx
r7W0uc3LS6VyVyY8OeIN/h7DGyoHhXuoTu0bjKdwBUvfvAfXcCuWYX9AefMlyimV
WH1flaqj1hvJakQ28qFlU6Q2okd6X2AbAhqNHOdvJJWPT3xqThFBoSr4U709mlVR
ob8UQsaVT7GuMT7g+DGt7MS6XoV6weq12Y4Wnt8sUtoNK8cdxeNITjaclws37Hqp
vN19+FhetiM+QI1f/VMBksgMju/Rwk3RViB9mg22J1m1pgqFvgTYMy2oOdaz5AZ/
AzZJi82zFC/YDSjzvkluzYHOn7wKprZie47Jd7l1pe4A7g5blv1H+LW9GxK3LklC
xVvRTsneXXmQZ+CHP+xQMfhWLikhu4x+nCkATgDl56ISF4gGXVH4ZtT3SDd/zX8i
pCkAk8K0bfP/7HAnDUE1K6HT2dxAEzSxitY1pwSifrZ8nIEPfL3N1NoiUarbwur1
rtvsb00HZ+d5NnqtP9FUkMteAsCV4YL6VUAn1rGS4scG+XDTnzOaSZXJjaqMQ9cV
WOQ3Z3r/NK+9bzzEsr/NdIvFm08RWdEvEzIq7gfvxXZRMww9yNdtx6z43a/svd0H
4iIRLJpYxFqZ/+s6rNIMRlWSTBMTa+R42c5YkM+Ns086AteU7d2JiliVzi0BepKM
MjgkRgM8gxeMhcysg98EvAuzXMiySPZC8M9fmbN8iDzawhDiwifUyRn+50RqwJh+
IEhCE5q4Z3p9tyRZIDJQDa2yYJ9U9ZhVTFdiVeunqHuwk7FNdhaMh/N/a7EbUneA
ykDYdWg1Jtrd+bYCKeENaONYbFU0sE1KFToWU78KEFZEZGa8wM6kGvkKHs85O1u3
/ETvXQi6zuUFsMyKyzYKt2AqKNAg7qFc2Hz9dfUAiJ2F15DA9bN+j0a7+OnGa98C
B1C8onuKQ01c5keGVuflNED/A2lF3Nh7wJc0MEtO5Z/uVB6agpVVx/XItD1Ibl0r
AlT6D/LLY8RCkUN65sZmVzZLEZyouAZL3F2K/hX1pAoFMYN7cw29i801ZHdmg84c
Of4P4tqUHQC1c4SynqN0fnkOf7zNLrGWBZS4PXc25UwSLo3ow1geiLpQetcoD9wY
8MEpaZmwsa42kqcW6/b/gQHNcaX/T+1Z2Dn5ETett8cCLJ8kpSSflzPIjf4DsBRY
WMFhcMNVCuVseWyIabLImNGWPeB4y/LYJyDtul5hvwyB3QRgubXl55G9tnS5QzRQ
tByrB+gfJUPporRvnTq6XJDaadf0AI9zRpZ7KFpe55wLhlknFzMTD/p+piWfNzJd
Q5z+bY6XLPxfFJYrKxMdycB19+nUZ33iToqcbno9ryzDC++TMuDwK9PliWqS9vU5
OnPYb32w8g7RYplunf0UdXUBQOY0JjhXF8DwrqzMyqIaVZtodRy7NZxQ1+lZHv86
sLR4SGnwbUCd22ffdQHw+begB0GAmv9UNNXB9O74IIBw85MNtVDAhsXaN86v6WSY
ZwukFx22RzZ5C1vUqDvRfZ2iLpgDATa+z7NXcvrkkLU4XpKnxsWj8XaBK31bT252
6VXXtdOd5aqlKjCXuwb/JrT+qAEjo+LvyzkvTrDUC8BWNZjGK9OtqBvUMIVqQtag
AyeXwAFS3MW+gTBOFXV7wJondpc2rSN9rMnuIMpU7PAo1jClomIJKv+0zR4ww2PY
P1OenwCdBMDSHPXtVOGknTbBTN5kHJJO1gjd2JRp/ij9zYrFJuvkEieKAYj8g1MA
DutckecZcQBPN80R4yvo31P+JYpe4H6KFcSC0NNN1OrZcf5pPw1os9rzkK41y7n9
DWYz7UuzyXCVtsISRxrDUMPeuOeBXGPJwIFd96pxqsih7SqjWTJMgDkQgQkh5lct
Wv6qot7N71DiwqsWMflWdY8TP9zqBZhh/9WK9Y5JsHgz4m6K0aHQuBhU09vbhvTd
fHDe2kqbxIzBKW4psLaw0c6eLhKDY3N6OnaaMLTYdlBjaI2AJqNtNz43svQndadS
Djq94e0Glh3wzWyMNgwep51ZBHU6kFxk5BjJUAtBHch4Kops7lsojGXaJaekASW8
NRFpfqbTG1a01IVAEjYSnUfNPyZINtJC8Jms2O/INx+mbOOaWN4yJs7A3pPn2vHY
adOwa1k+pC7b2nCPLWTXKmJYV+Ar9EEWNEwmwYIKSMK8vW+aw11q/dOEGmbLlRk8
nT+W4XD5PC+pXkF/FznKxYBZgSCIzjZxlvvbz3Im21/M84279BxQi6bSClTnnQBw
eSR1SUhvcEZo+M63jFS02QsYlI/+SfRykM+naF7tkboGnFmdX7/f7ZwP5vtDd2MM
ucUsr4cTRZnpe4/jLU364yULHPGrjvsfcTPz+4rQlrxjowt1AemKu8PTyX8s3Fma
13ejGYZnnvd40axR2UBEnLF1oElu7GVpGldwIHoF3whsSwvCe8pCD9kixbjTreu4
ogTj3+4dOS+OhkaT8akEccmg6MUX6xnf0Zz0072xXwcIwzbOxvwyXt5Xsk4vX99s
bbbnvl4mlXHpn0IhCHmSRkTbaNNMCJu4S8DmjEOtJPiGPVbf/bNcGhPz6t4leGBe
OB+wTqvrdxi5y9+7qRQrAWqboHcbbXnaFnAn6bralIvEun8exx5o3WhwxXYgE2Or
WdsCOuUsaCX2tZ2KspLM0uTPr2lYHPhpLZNAJUpXlnUAsLhB5PUl895A1txSE0mB
+IHeqbCrQr8nk17WNs9fnLCpZu088FJP29YtgpaUTiKohbs+7ZuWkeIHRKuUR1k/
hvUgAloko/+F4azFAk0/cZsjtO6J6yVaGJyg3TyKa0Ag29owpKfVTgjQ01QJXzUF
S/SiCL8RScLr4ZbL+LnQtyeCetmiGJeaNNs1/3n9751id5GNH2V5NITUzxnw7FGu
G9O1w1kQmTgrUeAHWvmMaIPoJOzNiVzg2fZa4EGp1uDHgFpFoaIUuQoEjP7bC2b8
ZdYYVvw5JlsYO3oOwrd51xWva91cCcZl8PHD40iKvpuSfQoVymCwriXyrkHhBv6a
quN/pQuottua0qm5PyHB07NwHMUWrSpr2gRwarLD3aXEEXRHSR/MdLK0f0qJIXHr
6nBz05GBTYZ1JQLTIPV0I4ePs2HaODCUbPbhRDefLrkuWaogyzx38xIV6mIKiQY2
SpuYyY4uhyI2FoVPbOqvVahSC/nvV8AzyVtpjLUKyPa8Iz+uo70MG9/oE1mL6c5d
heI8rzOMBZTub/5vf7K+SU0QN8nd82fFCL8lNUBEX/n7CqSluQHsUUHgJhlT0FWR
wdWBLmz4f4xW+jSXNPtA4h8FFFeSKnK7lsYjW+OYNIODwx7Unp6n07iuuZskkOMd
9E6Nv9JyXXn685YIMMcUyiXlRzmUlvaEBuShW3s9lrHPXr2lmL53OGb5t/GrUrNP

--pragma protect end_data_block
--pragma protect digest_block
/ceHlX6pp4CAK2VFixg3MKLnJ0o=
--pragma protect end_digest_block
--pragma protect end_protected
