-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
0AVSq0CIKoYK4MsESHXEt6Htj9s6ulVZgckziuzOSZrjF+l3vjRnIPCrvP+5MPqF
E+ws1Ptdpd37mZp0gJjaka/pKih4NYOOHhHPbnugI6CmQYhi7O+4hFlk7sms7p6g
UYNF7c/Sg7G3Y9kGedkdcYh/irW/KsT7m56VZzK45W4AhFB+zdTBmA==
--pragma protect end_key_block
--pragma protect digest_block
+nxhmskvjyagNF2rrO6Tbhftn3Q=
--pragma protect end_digest_block
--pragma protect data_block
OxNGukBQCaoHjxpFgpMJ3MPsIe+Xp4stYFxMopLq4200fhWJ+Wh0Oh1bVU4uq1n/
c4vRmv9K6qwPTmk79rKW1JOkKYJPtvTUztxUY5+EB/MhRqJR5vT7sz8z8+GmrKfm
7s9xdPYvMJI2KLJLcVEc13b3i2Zr76KHENA6jVECFu28aLCo98amyfhLH/qH8GDi
tFnWcSBMYHHuaOpcU8LxIHA2l8GoYEFi47VIQFJfJ19CrqeJywzeeexnywBIuwRa
RfgWJG0QpJtkjom+rwiUBEkqEI+VnzCeFVoQdYVibBepoAv29OTX/z4Q3kyR9B6Y
SJymzATxbqyjwCkpo7BwQH/V3g2WXkPGv+xjeY3TEiehIcDnmA/iLpzJDsmqomVS
jj/q0YagIikeUj8SdZK2/cp+lvQ5yZXfqYjLQtnaD09DLV8WD7GXRnbiayMKw/ZZ
JNyfMu88Y1JhOJ8CEmHqo06HWSbxF3WTDbfUtsK7BOzdC0uPM32GQrT8uISrGxho
xjvPHylbGAj2G4s7ngc1bqubjYmJt1Hep1gZeX71dmpzv6Rivlxj5oQ7Y9jW94to
Od8rZEwR1PeoMPVWXrpOiCuMpiA87m09RGSY2KDQYeBX3WBQxeWXgjQjkLRiT/LY
PJNClhvQBr3/feWgvMNfHi05F/hcoX+qk8FlFL61lO1/Jesbr2aKzjIx97tJp0bB
X2yNU9aahpn8ojmodvkyDCVbB7rzX7A0orIkoE8DaX0jWG1qFzNSRZRk3mGroa2R
bnlrDgIPcVJ65DPc/03IKN0ymK3xZt/DEh7nVLmUOFapl4JC5R1a3B4i8Mklk/28
v2TB3pyHMUOYk6ceOhZ74lP65y5cv+WQnzKbNdeIYK4s+nbJhPW2xVwpwPURrLtD
H/71KKEOT+/nQo+MmJMYqTdzB+UIOc9z1wNoqEiaguH0X/CJHQn8N3f9W4xH/+Zs
svg1kZpOvhzx+8OpFYIeVnAxhmh3jk+KsLe8DN6hw8gWFQHkbBCUm9EgvptCYSmn
mSeutaFrKSVWE+uGzg1Lj4eLYplvvTd2QizzcMZLLfH3DcLEBjG6p76WUAAMmP5c
IxFVWHfRr1720T8aazMJt/+AxVW/85brOeE1t5sBTuzW8qnAwBV64Bxi1etEZU36
zM+oGp3xBJr/r1gFY205TLXBXNhwIiI0TIU4Qyfo3j5gZ9PhYkr1a4ZgTmSLUgQ0
GiZoa6sl5H/YMBeLp3vJEPxa/kjVU5xNf+5Tk37vU1oC0tI3f/pxU22up6NlBjUn
U9TyrIYc8zG96NIjlJQQjVG8zQe3krd/HEvXaLTZXAboszPv9D6J1/ZR5puNLSOx
keMhkT4lUt5/+LE1SgdCx4MhqqvFOWxs/WepJ+OZOciow0iBBFb24hYgAUnj4s3d
tQYhJg92qkUEX/CFlBojIatlGhrIq6nCJ8zJ1XjE5rzoG5VUE5C1EbTEYdUxJgVp
BoZqTIVUjtsGl1GTQlibsKO2yNb8Euuqxbs0aENJwtcPtXrElzRkSUFLXYwUXQvf
cv7RduWnCNSYJ0+fnzD50k/aYi+wOaGwO3e+5+MXgBu/NZrThyUC4ZsJ4aOLSjIj
jqO1SrVDRrg+8bk0oIhvb8kGy5fNG/G5YyeztLBAbYUBSmpQNhAq1/aWxfs9xhwQ
nW1emwaOPbKfK4NxOpcCIIRR1NgZhH2QzO7CrEUnd+cj3kg+wrTzXEuUwGoXGGim
xhoUboXxzBJwXcgFXup8Gnre2ynue4tqg+IIh3hGBgMzc+/kmDWIw3q7OHL7PCwk
wX13D0O7qLZgR0Ag0nlYKFPhALZM++qeW1fr1yZpiAtFprXEGR3JatIZ973xonMv
/uxf2GbZz39M/sI6RUyU5fgEcDnwcnpW+vgR5jdAHCYqq9LIlDydvK03jo4NLr5R
Mhw86MNJ42NYXo2frdl4mHJ5Fd4+fADd7hGEeN9vjhwDGUKu4s2sPi80mjfx/mPI
SSfdVMqwhKSCO+DfDi1KzvTXw2NL5+3jqV3GW2/lYBkqTuEUEyOXpXjN2qeEN8gv
7c3L9CabTYoI9Ri5J25KNXR4EiaIlZIV9oT6cumELBNDyCixCwRG7GV9QMHfRz8q
kWPkyzfBGxr+GFOmFDXRXS/JC4VQAX/ZcQNVqZvdjF/V7kbsNC9NXilwLz1K5vnK
jq78eM5EIeENoxJYNrpnPnzbyuz6dKqTkykBNU9cVXRXLqcroexI3LP6Je0hJFZM
r/XkhwhA+0ncdzJGQs4uBVKbjrFF2ZZzPtfpGJYQtjYwXTZMSnBD+6ztr6Vn31oV
oNL75XC5VOo/tocbHDkR+fsWxZPoBG52guD7wrTWRqmCIkrvleUzwpmleUjCd9nc
FvweQU/feUOegEIDY1oWMLmSV6xYJsAVX6q5g5XvgxzxAaEjcDwdB7+4olWZs9nj
9tHXUzLoAqd0ZlqXq3vLaF/7gm/4IgIHGf1hbIyEMWRjU/62fMjvTKYaZxetUmEx
pnaQpvw/x/nw5Ae51mrhh2YrI8zYH+mnIF3O/3ufhtpHWDjUOZCaeSXWiorwqjqx
0qtk+e5Z1ikR275oAPFIKZNi6m8vVyoYQ2Jg8ttwYgHT+eLQ9rNA/n6XPPVSYLJT
Zw5xsgVYccli4+QBh+dK4FnTTPdxH1QV5NRLQyZGsoOlqemssHgtEiUSLfjuJ50t
SBR8Q8HfYI/EA2yXLmo+52PfiXAG3d/jvOeP7aQwCtc6XVAy484fvcMGfUbx4k7j
hpIBtwB4AS/7uZqTqtvsOZlVEz3ZLbhOgOHcJAZ7oYSASL5ntvRQ1aQ1Q6I23Jy5
6NtiwmFtoiJk9oALmWgmY8QnAbC59BWtgvFg7d0W0IU5KfefHNOEvj6n4FiKFtLq
sij0A+yjE9tMJHrzloKxlrTMlaYNmLkNXTYwf9oHnmXlFB9uSUfaTM2oR2Uc95tu
ESanvpDGSr79IdTVlm2Il+5OTL3WsWni22C8HXh40bh9ZDHXiQ//tko8y4MqEGfu
dBmWY/FqdR3JMIGEXxX1xiM2wtvsfllOkfWZrAaD+jV8ECXWs//cJij1DexurHD4
vfjcOeRPkrSMO9ckAE0xTvZM5Sm3SyeX1P6UKzBMWtmKeffnT7mnRwprE4lVvGUn
eRxj798lrpPOM/eiRTlKtytGSlNO/IrJJzpk5FM6UBP7gqAcz8CYYnZ9ctoowlxx
J5ThVsgYJRvy0rwGqp0EdR6mpGSge0070ar+NHRlE/DyAe3MIUSINaudRi0JaHM8
DZuRpaCr9L0wOUQETU2BO2MQPMcjkyCVmZ10q/thOr5y1KOzpsyAMLDZwozB+C5r
NbZ6xEfr5g6GgAeTd/14zE8NhYtdfPRAwAukkTJQgE07ygZhuVxMsPamFVjyYfMg
frCx2cbsirjK9z6Pl1lARL3GgMbBgxF2xUHWpYP5gHXDjcXHIULZzQG9MSY/8puF
2dzTFhYCT7nqRqpkPw133FvMJPnwBJLMFRWI8cdbdKqVeL9yHdTR2Z/dDw62dPdI
HWTSiGSPH1O64+tAEwusTTyJ9NP4JHOqb+YkP9t2aBdN9o0INsQChf+uYbdgkps3
gu9NzSeYknVFGPRmjSt0VaP27dAD4LtBi0Gis5rCMyhRk4jyQBybMsCDOgP0L2x+
KAWdb5T2NGuxGTltdNecJp1Ac2gPKl1nMgPmhNcjVohjP2NCp1pNX5Kt9zKzELVw
vrwFOUoi4tYGaiBXZPX1ClMmaXMOKObcKEJhftdOreatiETerhqa2KmtjP7lAlz4
RxHMRA2y2PftCs2wsBKoxOH8F52MGtGYt645JqZQf5ZxwZWue+EAOok7ca2BweMt
rI/Wdus711Ie8EOGRLH8fGqLcFjSYCQ5cI+rjLgpgmCV4JBNHGTKcWBYaDDTI/2f
XwhcNYlzqzpDM2XM45HVsiaw2ePTZVfn2dgAUGqjSUgSBIpE/VH/Y/Ra51os1oxX
7L4iGtWZSYm1yX7KzDJfoslSZ6voNMhMMcHJkiqV4y5X1LXuRiSzjlJruGsU/OJc
bhzMoaWH88Hti6lXOomUYe2LIXRzItUFIzR6X+hH+RIchGbWFg+eJ1aq09WyDcpT
8JE+w9+ZjlaZeR6GIOy3sywrOzdku8hN0wwrTXdg8/athN+c0d3jQmJkkJIWTQSK
ARXUyiBzeHUtQf4c014KMejbuaVnVJBzP+7vKUZGCfGRgc0/ftH7w2A9bYjaKyEE
+IDMzHmeIYmr59ar6ii/CpkupCTyEgYv0OZ3AmMPUpeUYYc8cKsX5L8xZdw17NGR
nEazqRPSjarRpZOLY+9hJJtkArfyeBylck+ZFn2RqqPyQcJNnjML8sGjYPzkj6gk
o6nadtcayZWGp/68nCf3hKBSaHCkfy15q1aAV4xPygXSqm/481oQ0DO5LtALupKb
dvf4nksAVcsq19kVce2ghAWTErpXUAM+sZbdFTNIdd529Hry28A9PU2n9YRFosaM
aL/COXrSo8AbHcBGGf3ajeQ3gbMvRtWOtHFbg7kmA2usXbXTrQKWGJlNZGy4nLVz
esRHaOJ3ZExb3iDonOlvd0P990wXBbez8Sn2zRxKR4LNBsHIb3KozyxOvIWukv58
2ZCHy4tlM/HfV1Elk+V+H87vAmPBJIjl+aGKc1s9CQz9uc1qFTo2jlNqMFuDGYqr
7dgHAMrFYwZUJqJVyy9ALmt2rlJudnrDtaKZhgI8P6mItvXnDU1z9NYz00ctt/53
oOBq+rlb67oaSruTs8i3DkZpB7iSa8esLtRD/rColXczNykGZqC2wjRACAQrfzbg
BaJvUIVSki1FH6j0vk/DtETHAqt29Al5J6x1J5uldkrU3sLY/TyekpHGH469dg1C
BGthSgEnVH/dYinL2tykmXPxlwsrILV3pGGjv06zhkfSbu2zGU8XPNdKhELbuVKJ
thcMPmhD5GjqNG+QsX60Gd5Zl703mEE//zjinMnkQc+TaUEW7GuQadipD0ELr8N9
OI220VtPSHDPf1eX1yBI5WuuwKnmUv5RnRPAakKw5BSc342EfAC+XLFTUFmDi2id
99xMF3tIW0yTCaE3bb4/l9dwzsu+w4VTxMAXuuAsg1/hzCYMeOoV7n1pVbKEw/zn
GgesGAEEaTInKgZU/dh5KXk5QdKxCB1ivf5g2tYbJPWd+OKH4I5iiQ719sz6n2U5
/7a+Ht/8SNNs4Wde8ElzRxIVsG+WFCcuzyGPmlfzjJ+lQuQ4AhWnGE1xbjDZ2lW2
9GoMPPIlqMzbcwZQkDFmkEao/ZEPESeDH+NxRjB2ZNtNFsMeTgtp7IkcI542uJOm
jplBKaGzPp7Xj1FCjCYc/ZEki7sR7OsDg///ZmDbZQMURyXjhOaVO1E4wkA1J8ea
LezCDIGRMgz0m1H9lMriEjen1yE24w7NYsbH1dAy0ltcwG0Aleo4R7HHvmZ8aYTT
S9OJPz3FQeB6dm06xIFEnBo0lRfGtEfFQ2gjih+ZP/KG1kGlTa8JWCECryqsbb+B
6fX4PeTPSxeVHs4bTsDE1393I+fgWp5vUc14xFFqIw357QiExCpOR506AdraP4k5
yHJ5ptY8SXelb6qlN3dDVTdEKBJZhEMx2S6JqsleYqG9qcfZyj+hWK5+gnqppOLv
Z3AtxKPVbSnarmMLvgoza3qgLcaiyYxpfuW2r2pGiwepLgU06pkI3esi5/iOeOUX
7RnPTQdBJjzpRo+kUhoyH0XX/k5/jdN/isM086Qf1LZB8yOf9ZDRpP7SsWcbErwm
XRDCnNL8RV6RVcem7MqOtsMeCHmoKWEhDI7TWNd4cQJR9UVGBQD3B1TNBExxL3xM
6xfyJzcL7MQ5edb0PhH7GbyUniiHmDjtpA/fDd523Wet9K5txcalu25Vs/aZ6pmx
M3P5jPbv5vt+CR1siEWM8pMF9LgIaK3Z0W4V1Lt9mVg5PMNUuAaMgCl/Xwb8E5/W
RbKQsgbvlAF4fJgAAx6cqLzP+z3S/vegX57E2B/xLVodnJuW4TuusEZxI49A7JLZ
0kq1sDPPFfxVfu63noxFKEIIUECjrx9VFOUHvj89p+V+h9mXq1ToKcvJfJllQ/TG
kMZn9PUc33FeB2o5hvxjeCFOvYDRLR0TmwJFEdAAKm/2BTwvDcsfk9wo7yUoZ3+u
XafW9QErrTQhT/lLYs2O/HkovcQxGbtFGxpvsCbSzLn/MWaP6REqfmBmSYacoXzJ
xm5YJpSefBIBTrsqJVHg60Tg9s0L+dnOs0NrEF3fE5GKXQEkWmfaF1t0uuPEsrxa
0JCBzXM84At3Ouulp3Cqq5Fd908pBiEtipIYqRcXpaD9qJBqeZv+A+E+U6scki1N
YKx0muO+PdBq4vXvkZK2cuB+BBtmZd6iAJ+tthDCp/BATM0e/bO3gZYWuDZqY6ZR
5Ly4Ltb4lKPpjw7tOPdwh0cBW1hmlpHWpRp1XLQhhcLQ78t/kz1QAAOBnJwNJHsk
l2Anx5QjY9PNpYtnAasHZNzoQJ5AZXx45goOT3sGe60tUp3iBXDQEsIUbifcjZ1v
+zFkCHW109gQcdQmJRrCLmP488xmqp4yVfSH744Uv4UM0jNTx8m0o38oLR/IjbZB
fy+R4d7vlarqQkJ3bS9yqyKeX/h0my1B4DIz6OqNTZ/5W8kjMAUbO6pS+0AOKitq
rR7eitE7VJNHRE2ikwQznWDs9y1bOd9NTZ3PJA+jg/vyHTPP5CBThDa51g2Rwr1j
beSJuXAnZwbcaXWiflhIuTa/wdF9d0ctoWwpkxNxYAXvzCTANUDqzMlOWfFEM3pA
3q2BMz0ReBR5P+2iaqtHAAa8+Y0a0MCE7bgkeyxxUXrzmMqcny6ttLrcuD0T7bfv
stmEyvjuH6RrU9o1L9mHs+nIspnGZB/JBie0ina5oZL/Ovz3dzSDM09jr/XVdGk/
+2Ta9ltWlmDkGlMmZwI6V2nglFQQWyNSfThUV8povuJny/JIxlhO+AXAn140Z5Ae
/z67xzDvtjtT+ROoJzGkdJYyO6YKY35hqTgxzU/SzZ+inwKTASCOBWSieTHrXU2p
g3IYeaL8GH4l63B6Ro4EZ+6CCfp7TfDu+usfyUG1KXS0Sz+Zxki1bI3gl714iZy6
3bO8+wgn1QTNMvTOlK+3V69JVv/bd34xIjLv9FqM9SuYiwMgSSBm+x3osEyia5AY
Mhxn6kTRzlLaEzf+zFL9H3hqtxhoV0oCWr06Ltk6ojJUlk2Iw30wraLqAybJ5pGp
1OngsTpu36yB9pfFNWO4/VaM8SpnLqlbe/2zd/nT/M6d0jOVLrcs+ugHC85GSAPj
VX2Er6W1/M2pWGY6/5GVopWy5sth6fOVZdoBxpaDZITAK4Wqn/FVidxhLHeW23OB
gcNGWagM44TQS5gCOkfxDwO6akZyUIJiV4ywmIOqLA4pjW6vlbZNrJC2fV+vaMbc
AC3G2BHP4Ug/SqC/T0maFHgY0d5l3RIcuBKvkvUFaMJU3g2lWMKlLf4NN5IgUo7z
0ywJKzD30o9vqRvP7Amm8tPqWT2ld3xNSDFp/mfTCpWeo93Da6teioDjZQpYIKfr
wGiDN+eAu6yv5HxICFvSQl5uFU2Zch/ZmYl2vqNIgC66nLwlJigRCjVx2vdQ2GOa
pi0R09nI4QfBpxAPpGv4+gJfRAgEpU83mnVzlm3ROIdPEapAktjoaRaLxbVaLNr4
7z9IJMmr0RPK74CXMp43/awa0p0IbdiHEthYXeZqOFmVHUcFQZIM4ou+Sx3qjgeF
Cx2fgAevMgd2t18FqQS3KQeXD2ln2ygjFdLSz9oi18tT72tQxMwt8INLa2qvsRLi
NPZWSL9p73BtO3vqkOE+CrUFfh/g3PAMv6xPLdDmFBO2R48uTn8jUvIIRMBBicsA
JDVLawzfRVF/lAZ+zvcZGsJO3JiKZN2Y9ca8TYZOlgnm+2hB4Z0oLkwhnAMymfiW
uspbnpCAh1nulTMY28Whn0iZZm2AKr9oWBjUjWzpSsj6SPlOUlMg4CWZIh8AyEPw
oqzAcW2dySFW8Epqxte/Tq7ZEqRP8Vaer6/tm4Dr3+N34T4gZdYl3vZ5aWvDo7DK
n4RgduZTbI7atMkt+kzpougPJERPzxe3neJwQijExU9eCxUfbMaTbDQ/rjSXVOE3
F6rcD5z5/u1bg8ZZJ6MvvXdjfjC4t0rQVFEiZA/+dGniwfRQ+f7bpXqG2WuFDZvH
0dL0vKsvatwYLbnQM5rgTmlBu0Ejw/rjArNvmi4hTCECfhNQ82ALnkfl4RqRFRCW
WHzah8HQhT5I+zNrKLO2+oqh1DDQkGUzPhfImshgGFbfK7odnjpSGvCRiAujwj1H
2p/PxDn4z7/AlhAeahZQF7RoNtap149zKi3ZM/nCd5ktT3xc+PpijG11Vzwsidxn
QgB3GpwCvSDIgcZZ+jj3pJbbiu+QTg/x5id7ZGLAhJLuyfTTquH0Xd23rZbfmr1U
GN8c24p8ojY/sT7ucZp0BrO7dyajbF1Fgwf9jzcy6W9VSWg9St+N2+CTZBVPsLvW
ZAPwDYCM90ltQRP/p+INHWn5CsTJ8rxN1Y2FHoMq250XU/+0rswwMou8jA1uhxYf
lOoGqOcMR/vmCVd6sZR0MwW+j0LtPewYUP6AfoRJsMin7VA69iZ7y21f3QucRors
rcnr3KTjCcW/CE/M+4MHAF05Y10CEwbrB0OknQeRM+n19oDWFgNHsVj1TuEmQw21
7bxG+z0H1suojoddKZ3FpBLKJUN7LJqDkjZBxZt6kRsHUKMPhsdK7QpxmTm3D17P
6iLm1rj8lpLY5EqYtvSy/4Kero8gILXMHA9zLxCZDqgyEIOmbCjZAnOL2PH26Ses
7cOrcQ0TxBwaOhWnIYiQu1NBl2G++zey4q6NQ/k5YZzp1vvI4NNdZia+t0tkQNZB
1B3bos2ZFebHhhZduTQIv84zgWlING3qX7nRDO+GhpJ1N7jD9wmas92HaUQEl26S
JlwjCS9HSqDc+WGeauI1Fdqe6ylkuFw+zcqrE42xwvHJux35MweQiAQZ40Rq+aOu
SfSP1TCOhHazv+Fkfgjr71xdBx2MYNCmN167TSNlQHsq875cq48w8bQ5fdDPfAAb
zlJUpvtLP9r8I05dGEGLHfRUsPc9lK69v+g7oqjobLjMV5MGeK2AOpyRwFaOjE4/
Ir4KBc3dmcZrEUgDC6/5qOYyClfMAvzoB78ufimpGysFDxxEXdZp1mScIgnc7vdy
1pxxfarTQdvhenGfdUl4KNH2Goe0oH8kVTpOWTg+rUisvaQHR/tKGYu3OPkTiJkG
SZ5OsMTkVFY96iLru/+4Ax6MfTZBFTNazRDhCPMruWER9gX80F7xPni21B7xJ1y9
UqL8iIbxjwQQPlbngaMawTTXzaMJfDa+ZWisHihL2mMIwWzY59M9xk4wW2sOxwOM
cGpGdMPJm8cO6O0ryDmG78kclhWHxB0RcpUM1b70NcfuEyilI4ZysJzL0Z0MZcEg
O/HoRu2jCt34DLhVcu+cL+BqnilAmk22QuutIY4Sr5KhsV7FytquO7vK20WZrNGC
qaEIBQ09twKwmXiRnh/otPL7BZtXO6nBaLAMmDjcXoskka/58bMJ3rTA8TULP2UQ
lUz70IWrw9m9BMHR//QbPfGfIHjBZE7bf62yypkO4QVlSdGbpc3JBGgVY4YdbzB3
KDCmElpRFYzaZQvWNGtoVLjv9zb2WihCtwY+p0TCk3LDoJGeTCFj/wH8daKwPzqw
wfwfqvmE7aDVtab/g9rVxVwPOetkiJHZRJ2dHcbo515zljURD00+Z0wa1kE8KaN8
pFt+LZ83WMCtrAxiunhLSABJULUM0fNzqnS9j0zlAE3RKh+NNaS9YTneBZsySMI2
A7FAPDsgr9Spg/Q2ZlnvHlphF1H2A4OVfiHR4DHP1Q8Gcm0FPT4nwIgjheczeg6h
6DOIRe8m3/I49mCtpSi12xs7DgGkrv8747WKKGrMuHKhMya5wjwMyTNGp0UF/Zev
5KTXDfZrbXotC7a1xIuIpH0g+W736yCjGVpRhIW6GYXlhNmH9H61hcvBlDnHyXJq
2EJ0NWZ9SPVZwSaF/dj6cyEqzAIhTUE8BSMoQbbJngDQGLPd1tYo5ojFt3rfjdg+
V0uAcyidD1Hcjrrh3LoPLujYqUUxTbN+rdMahgAel9rITYE7nTQCeVYjHU6rh6JD
yQkLLe0mMCqA7hTr3CVFpsveITk03VXcuygc2P1kCqsy4H33pgTjp9caxKWj+mQn
rSJ+mW9A862xSPVmzRyHSunA4FH8D7qWOCsvIvdw/xML8o+ZbnKsy+jvxkLjI9YV
3KK/7hitQDy1rKx393HfnK8XBoALGv7U6lFoqEOlc3f10uSIindzQUuQj38imRup
TylISezFrM4sWPLubdSIL3BKNfsWFnGUr1aCB02gKIF30i1kZ7Hn32U63ZuY0x3f
cMzABMuvMSxP8P2qsjFyatZDxFTA3fOKUPk9/PDi411rJhjjrfOA0S/tmwpRcG7F
IhSm4PPEZrki0XodSrla5QIYBvij5/i3uTqMu8mmK7Z/u5tsg4+vif5i5M8Jey63
Zu1Z0ozNXfRixh1WnwNPIyWQX3C5omrbnV03lTdzm+DL8EwUsA+XpG2hmEVrnF+t
JuTkwQ3T3p927wTH3n2H5XkkKROp1s6u952nNv4tLYZcVbuATzxplSAM3nnFpxky
P0/+8XhFqnkUvoeKsojnFZJIFUGKuBo5KP+48R++ECuHZCY6hVOUX20sskpIX1jN
R2oIL5meZTrVp2b0HHugp98DaU9NnJL0WKOzWyI+MNi7DwpUw7gz7xz70SQXv5bf
J3XQTZ5z74pZMT1Yo9tHYs22PEF8Fr+o19toykD+ssUp0rWM5l55NlUKb+yPHR24
w4aDzB1JpYJOOd45EOU/S2EfNCd/KF49vgTE4bi7wHCtzupuxYcKsByjCUlArt0j
kc/F5YwwlkgFYEiwn1NMlcdEq5Y4mRJnwC4YdJIFvKY2zxdXWNSfN5ehHPb7s8nP
sZ/TwhoEYs7LqCneq01o9PRhSksveBeCFB+uqXu6QmpQ4DHYTxr+2QnPpswXOSqa
uE+pge0FlLYyy+emaVWXWdMKmFg8mOshx9/Co59KY2TG8l1Qdy/1gFSzjKvB7G+s
TDJZGtkUEmMjLOZUkdiJmSQ4PxHI6SqPhGXI3UsyxAvqKZd/UvP6jyU4vCGOErZT
gea4GwJ8lK9Ypylduihx4dEja/0dPpwwSJgdjxLv6RzL8maZBEA3vWVm/Zj5QYo0
Ysv5i7NeY1XYOd56CDSF/wFTW7T5t1lhfxOgCHVasTEtaRzilWuIu1XemiAgHpVN
lMAJY6AOEvubC8fxP9f6J2x3g5hNF0qeculMI2JlSMRPJtV4P/EVwkj4rYiltcur
J44HCSGbsFzxe0e2mW0HtNHQJuJDh29ArRrDQ+zy8vA5cEtOtWcih2duvDbwIWDm
Z7PV8Ss1uhv3UYtuGNVzV5IbvpF//AmV1+777jlgSaTiX9qBn5SCuzuvasXt5m7N
IT3/DEPIrAR4B5BmOJDeOu5b4pdSx1YYrpwtaeYWY6PejTl1qCcOvUot/Tp6j2e2
AVdbFuzlmiDBFEforE3+vT5UzWwD+PCZvPP0n/JVQ6FAnxx+htLnQ0hLqsh9kHCl
86PjKx7TyNanrjPxIONHlpbL/ik8W5gZPMws7jvANH8QRfxjR8MYaflqXuxKexfc
zFcUHQZN17a9RWupLLaTisi4t03bKDUzGDgim6sMp/1yY6hc1wCNpZj3STV1wA8u
yLK8HRkCu4DtVIF7IaT4s0BuNp80EiAZKRSWwX3ikjdxnQS8fydyEWOnmKPm8wJI
6I+NJYhbb600Lp2mXGxDzLjhNtj4R9iCYNDJbbYFeeyEYa0/dRSqjwpVuprluy9t
KKeYhnhTCjsmT5hqOYIu1zSM3Kydy0TAJ3XFY3ZJcg1G9Z1crySCbpfJyeci2Mtv
ZnvKiIAnWg1xg/vLSyMeMwslnhC6hbH9eE+2Sl0Q2rtjtNQ4XyuNYY0MLizoX4c/
g7vQAunLDefOnZYiMRIcMZchONz7+jGL6Bn7DcGxUO99LezaZma/AgAaKNPB9wUj
A9DvBZk+ODRH7/ID2BiJ9Zy7vcnzH2wIc1vnefF51EwP+oSXa/V/cAPuveVD9jlv
RziQ/9dThDUBdHUSGM/8mqmHHatMpVCGIYEykZ4pvLc53HoSGYsWfzHg5BhxUt8K
cI+YW1lKQknUJXkaLED0o5dFxQcmaau4R/HGvlJjy2e6MgkdaIyhgcd9eksCLFWe
P27HhmBz6XTiCE1JmlcNgObTQEbyxIqJf76UQU1QYC0QR70Ed7ZWrcQrSSVjBpVj
XJldCK1hG/whewKdnKtv2En3UaVLKAj7nbPVPvfVv4m6LJsLnGYtes95PaqsSWY1
SR81dTqck6k/yzvpsV7T0RuHTvYZypoFmsyQ488jpNNlwJoe10kbO+ghpWqhfCre
jnxS9gAXS/+tOeAtGyHffGzustQwKUjDvhFsOHlMQ/j9WZpAcJ8IvszC9F4GyOVd
SpMtpWxMLTxe0jk92n5g9Cy8mXaPEGbAjfsUXL97zUGMiNu5DIB9fruDhZHDGeLA
cIb/JeSunM/KLz63u7oOtWO0IRhaiAlEXvnXVQXNMLq/NSTv90Fu3MBiV8pCTFni
JCx8ijTYwK9BjuLv8Ftd534vkNrUgzccAcv6xyJhmiZAf9En7/1HReJsKYwqZeDW
8Iovmv6SXP/QZyH3OciQFCpIVUYioYq0/lGOZwqePyMBLFrWCfVOQAZOZ5kIwBHk
giK7V20L6ciUgGwcqskH4/K0d//a+VOWnLYRNZ+86PeZbq29f4fNvP+ibdJyzpj5
cSPIg4DMRR99V8E0V1iMX/G/rb/Ce/jsPBOuB1o6N5/XuZp6RDHQjgFhrdH7n/FE
gC2/2tZsojy695bb6fehBeFXwTUr+CV96ZN6v+HC/u0XajvGJPK2HWEkwLquFHuW
7Jb7UgYk5TT1eA/YTWyzztRceobNMdOCbP7grygnFfdpCiK3+hgHzhSexDrQkv2t
VjGmeqRH4u8zqh0K4yR8afe3LrMHAvtAVVD20ZYU9zyUoqfiGK7gZ0oS8LAZ4hfX
ExsV7nDLRDxDtsxESgH0XWCJKeCI4k7Vi5PItNN5UKN4d3TEhDhYbu1bxyimryB5
SQKGlCDTXXCtz4oADLs7m9QnCEkA7Eh9kH6t/EfBbg8M8KLGLOSrIW3WcET96kqU
arFRRb3GlPQ0iX8QKvB2qpu4pAxI5As/kS6GaEOKRV5HiFXgscnAK9TLKV7UJnRV
0MBWNFWb2nAmFEvu9wOMT98tXAX7S/vU8JNGg4WN6jf4exqk3jhPhkInUCNCyP+x
eaN7i/90WEv9ht9+wl49Ign8waOckiESZXwA/xG8qBQvA0kSfhdXO51g0YjA9CSI
AdAxspGbYmk1BmLf0qekFYmacPjnkOrr1DjlK9mPpjnpMRziOt51xtYjZtFp9Msb
HHjN116gfGeub6BKNo001s4TflPIqRiyGHb46gsJbKWpv5qwOGNI0iqWF8XWBhlq
s3ldS4sCd4gfKoKahC51a9JqUCj7XgZ60nBQJ70rz8UT/SZnPtjjduJon4w3Hnfq
q0+rUfdg2ss142+lF6/XhcD9ONmEtXFrgik4/7G4Laqr++Brw4HkdIycsC9oXjBO
Qb8LokFAd3WBpYSiYneB+M+HPnd7lATuVj56W0BNzyccMbvmbtVr2aLhMpUsBEkz
WJNVw5a5TZbUi0ABlrPzo1zaEJfeXI8B9LvGs3kM+xSqVM0VYSNVHQPKwu8PO4TP
JPOyJJ/7mNu2yLnYdfFmcY5wNHVPsCrxOBBLVkKNVHJWH0nunPAo56ZGvpLfODUV
eZpZLWwZbm03VncwEL9jhPabRf1sOiDFZKfxryNostWeEzCPNppE40Y+OkY/rOZQ
6Iwxow75H4IZ5j1bT8zeyWctZ+cP/LvBro4el2pPsZXAmLMxME9GxpWaZSbvjwPu
ipiMEY8nSQZlfmHv4LgEYa2SwZbONsPsE25+a8FfKmvpLm8ybwiamwHpeOigBVou
CnNbTjK+bWfiZNJKAN/skBugxl5etr1LTjHjtqCOV6BdnFG/ukhpELB8Qzv7mgpW
M/0AH/Pl11+SuvtQyd/LNXn8EbWvwYLl99DTT0miRLAsuCcwuPe7SwGc7IhYCmcj
g9f589SRsTtPXaVfJZzp1LqErS7dLBw6iIXHdMI1Jd58dtrkid/8/4j1jCemo6ln
vMlp1ALbDT7KKvm1wvVNbIVz0+jJZtPVX0PgVsh0UERLJFg+npCRO5Kjxs4BhOKy
GKuU1L3o/1hLmBBN3X1mdSLiEpWCX92WjOgKe6kYysW15g7JaKD5cU2h+pr5mSTj
wvRgyCmWQBezZaP1N7tHTFsq91JH+ywryIFU0vdVeAook62CoZVvMcoYXlHEFFES
EO5U47wYkTSO8oMzIOrCF30/ZIZvdH+et7ZHN35L+nI5jrFy3z4MVgOUjwdHulx0
uFV4JBHBBrtIrxX/75m8JBV6JUCl/CQadhNvdWGzjVcOWEJAbot/XkEARRSB6GKH
U6udqnod8qVRt6qi6XpTshfW+6vTHwo88SfkL1JiQlD6GDYKTZ/w4GRvvO0HempJ
DrR7lVGV7FVhrJ1A4dy2O89RxcEpHZiENsX5l2+ZFARun1T42AOG+J/gr9r99c08
oReUz0K/QPCgaxaiYkpUBdoxX0tJnf1Fln3NQ7lLktjW+Jic+fxa2vYPasufePHb
ZERMQKc1gHhA2GqbE3oUDTImyi7Ia9CAh3L1qJs1Lzgnkpqm2Lkj15sTIPXzhMQK
6fruUmqg9iPZL3bWEn1JAi4avu8eIURWbFU7dTaPtn9yRHER/RFQUAmsHxZg43Kf
q3jwIughno0kXQ9TaUrlRbMxqHUVgVHHpUybU8UXk1qq8l07cf2ytgcdyX3rk+Xm
Zn16TezyZzA/8DQVHuc1rLnJ0kM0IllqMvR/R73Z9pwnkb2ZQSkRE8whG7glFoPn
DbmZWiHpff/cDz4v43Jg5Tn0cI+4s48Bz84pccOv4XMOFsvHl4LUIrWoe66I1n5R
b2x2AFbs4xvNys4qK7mBjyDGZqMltNQrImI59ApLBGcjQboVpyBlEVY/Fp0YEKPL
Gkdp8GVOiR6A+3QmC8QmqNoyPM5ehTb8l/FZvChha2mgemhe58tEAjSKZj7BsW7C
cqFR2DsjGOH2Q1uCz5wtj6g7bIHUtedg00iGqi36uy4wc+oZDvFX9Ez4VXhW4Wil
EQa/+kPsEmuMVeBVwrcWHwEWQ5yJHo9sH/pyUMm72gvF/MqmDNczqYlImWhpoazJ
VK0HO41bj24eZuC6S6nU4AWlLE8DdYn7Jh5cYb2wlPPaLlZ3wkRBnrkYe79OiToC
rVFV4N97XC1lgVC2zxK8+4ziHiia1PmlHKbdxDOt+SKPMLknP8qLLY4a/zJQg2/T
sliNyRvpU5ewY/+7uNLgvHuEDjnuEjCiOvINghmVdCXLpJW4MtsJE9H/G192mzkx
4mRUNDq5bQhcq+XXa0MUxoFXYSlM2keH1dsgJfCjv4TYznQWvugQ2BwW04c9vpHU
6w2xR54H1mwCfergj8X55Wg+NTiHqTunFpoqv2/DDsq7Wb/ozgyzfk1de57FWjit
5SDjh59T/tkHoulfBTc1unuDubqGIMsOfbIjZA4IKsY=
--pragma protect end_data_block
--pragma protect digest_block
FntmqZEbFco+C4n6eyMQZGYylJI=
--pragma protect end_digest_block
--pragma protect end_protected
