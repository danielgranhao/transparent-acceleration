-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sfQ8EJBJVJ4mfkNStYGJDOAO7keCQ6AWxKi0EwmHWYHAOhUPrNkWOuNlHpk29d5N
eSRIsvOjsTGWio3hZ/nSGBUlwkzqHhRN5fE2ECvBbPb5V30avg//DYxMF5saqvQx
/j5znhFyqeEuKcEFbDUkXQ5Y6MbzwudPu7wcN89AhAA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7616)
`protect data_block
HFaQfZSFwOcbSNtfun7HvOinqvHwyAIv2wciNLzMVrlln/1jYtARQII38zrbEzVk
uiwOvNn6GamJvUYC4Udy3pbZNC2X5R0jAgH4dSsqz7j7rZ0Accek/2wutwqb7bh5
ljh0XU3Xibc++eXC/1xJMA3BfzlW+xbS86sFPrRzo2f+9mJ/MoKZ6Tn+HSOlnosp
aj792aiHIrO05WN2JrVB4a92hKCqOV048JAYFnAcvl7lNSD/BF26jcuzRHEvrrYD
DlKbyrfoCIPrk1OdMWHhbD05uHlTKuMJg0Vr2GhZJKbKiNOGw3LRtUhQjfPPf264
Dzu67pEHKGuyCWPfeRhocT8GBFi+H1E+1lF2/RSqd9zvehyo5wkJjuPSi0y3UOMC
F5UMxqpX8vX+tLDjFXya0utCUgxHrmtyp5Lbt5KE1hqvOKUEZCRKEO9b2fNtVy+W
/hOqUU6z1KrqIC3ci4YpUSgzvR0LCTHSUFtej7znQaXLH0dK6GXd4ckNuMxHuO87
dH+pSpdysCzjAlLa3i6evBG+V9XTsqNkq9sHfY0fl53ej6SCp2l3Xl15yi4PbRYN
SYPJt7MDRf+LE98+0FXBvwVU847xlRfkbXGE1Q4e3xH9LVZM6SZ5oNQ4Ab/HQNRx
dG0QuBXxR5chPpNZWBJwZhcYEzj16kuzSH7SjruA4OuVnyX+xinxUX2uclFLVquv
hzJusZV708BR7HDMdWYogxwIrXkthq/H3zt+LOG7BRC1sR8gxNVTB4d0w1YzLar3
WbNzHTwFw2iwR/JeHGfYrJcJrd6Eovfxaks9B20Ui99vV06NKj4yy/AtBaP+I2p5
gJ/0YbTQKRsCY/lClunCLQ7OnjdG7c2QFNb9oYp/scnK30o4C1bI9RtCKBeXDUzN
lyEEaexA9SWcKtzdvCQa8Iul9sWhCPI3eXK+SZbPiP/Q5vracm9b+Ji34dDKDPXq
B656z7lgDxqA4p4Iaq0AO9wTEPBIoln3/oNTiaUJtmMYuZQpsDzLrlbDbjOxwl/w
npScuFAV+Pf++aPmheQogsZGAm29rE2mWrZXwOsQYBCscRzIjS04+29ZJ2ntyWgL
rVeEt0ZZ8h1T9Ghw2l6LX41b9IfirP63CSmVvBxIG7x821/3Kfx5jHPBwcoeMbsT
7AvrQkR/y+k/0maq8xYPGWTWmFtnEQZEbtsVRMumg775BzkVetmDK9YCoBSgTSpF
9SkKT3YCugvap25yQxKjlvM4N0PvYFsuzTmdiGpFI0jSLDEnU+5BjbXX5PewOFsR
3czkZSIvxAFo8GGYIeiVZV4fEoMUaBGwLmpPHFqiYLGBeqJtLLM1JICom38B1KVt
B3agJPiXO2udzkyYJUTNYe1QaXW3FY0TQI3aPd5HmatIAVayHteDLMpD0pf45cRU
cCuIRypJ2rQiUdLXPaLU6Tx4b/he6a+f1hdA89+JJHA7JjROJnGopgT2JaIf0dBw
rt/J6yOPoT223BDUs9897lTKG4zQJbecv69wMwLK11hN8df/WJb3CGJLdI/E8MR4
7uSLHVKBijQv42usaSY42zbcJNSGCpDcD4jnTPou4SQMVUWl5QgypE+zlKEtXfg8
jzEoXCm9vN9lb+mi4jmpcKfs1c0mR7HMWEEcDRkNl4ktyJAoPMWMVDBVWXnxcTR3
+kFA4Oet+jDmSEZhxlA4o0kvbOhVWwO+Ie+LwZc0IeVFZTKPeePySFidoUmKc6hY
1u1UuhM6YgqD5vgC50jes4Sop3OMena/1qAzl1V4tHincYRW1P2fhsM6GcCe+vaL
1tB5RZGtw66gsU3/PdKowXgt+qRLH1v77b8AcDp68RUEIRoK4Cjq2zQRavfMBkoF
7QSnUdHmQtIN9vD2EQ+BMedd0WytjiFnlJlzNiEHwVvcr2MQFspPix9PLk2ngJxb
TJuDLeInjZ8HGKQExc4hHZQQ7W6gN80QzycKZvsZTHTSvEmln3ETmgy81f/gRvXU
PrkTgQqxVlDNiWp2QI7stxjp+JQF1NN7ETqfXx1eqMWFZfEcQHFIedOxvOc0Vy3X
2kUJWDdwvt3MyHvgSxWTNpZT/todoXTw0Dn5ihF2lmJ+eA37v9Lr8itWknDR8C7B
WPU5GxPQqTnhWRCT/qRnT90Ut+3AnsujXOedfQ37N/3/jlQ6Xxn2KXsYhdIlVJlc
BpCtvV5A6/rMiJnRoVPX/hWxzvNAliA4KphHPmhhWrsenmeQ1t/W6JDWjFml5qVC
V7X8vmkTxCg2LmmpT+KaYKO8HlZh7aaqvFKD0dR+Ee/3/nD0keKOGY0u078knm2X
pTDwXyz2xxFFwCKv0dXH6ihjb/6qkyF6hyY0qkCV1jfG1h5218M7Ug44Rztq7AFx
Ov8q0+ytvXkUsTkmWjUYRluO5ovsY4WFvtcWsPuu1418VFutD6qddnRKE4wQLgum
4+q0fHwqGnFbJGZeNF6NurJGo3PU0/Bb/szh+I5vr23iIpBGzsxZTu6q8A1Vc5/Y
Jr+sbRkJ6kIn1N989+oXWg7/sAfuD0WmCDwEakEKKrvpbEK9YOPvvny7U4Mi2Vt0
9ZAXB5z40BQh8l6r9mm2m558yQ7zUprwQmQvTEzyDWqFshMop3fuVhvHw2x31IWQ
KkUzWQ9qLh6iSh1RHZit6mwtZ2JBQnSlY7KOcgbSOHkrVVuS71MO9yjZkAJWQYDy
YqhcrPOAiK6RCCOAZhn5mYTM/hTHKP/BoABrqOFdF7x/8MDPOZuFox1auDkVMJLM
01kOwD7ae0xN8oL9CerlKvQuHuVx9xgxNuPAGjldIaXjSXOKQRxw/MVsmgfHJD/b
Qr4CvrG9/yDN0yt1cTGjXi5EDydMKeZA9YsXdJ0hPaHXlFhup2271yMOUu9DbkPh
WwLMQyyGxT1+kNtrAJzW/XzYPtUx23+nhrAPPKdPsCMLEJPvI6gxNpTvc/R7QWyu
vnWiqDluTCzFfrUbqKuAos+32NAMIr+Qoypyar/nLztZMo0taCRAq9pluwejKuuZ
fcOm4xGpHeIXsavcDOsXtClD+psVIyxmqX+5++7LE8lHoq3G2AZvSk2V8KTHvYAs
ZlgdQVHtIwKC9zryIswminiA8MBH74ar3i4h8p2wiRuBgoWSivReg9AuOH2mPHa6
qtHwSIFIvY9CWiii7YTmMPYRoWBY5ofPE9aW5VN3fgENBEEkWqZQtjXWvD9WWjwH
tstHf2vXxXWmz0Wr5QPtTdbI3wg8zFLCggaKUtdckUAXrsoCU3OdYJnYfV1KyffN
EP8Rinw2HcTlGuVN4m+D6G8gMhdRTiX6SjErbw+aM0m22zebu/KZseC5pjrcU5Pl
qKvL1Elwq3a9brYZ9WUBbNBKPGOrhIGbH5hnYxufk+4drOGb5SlEMnHou12KTv1F
8bkBOAKyl7VzNjjI15kcoc0VEWXx84RGKld6kHRwNheeOCrD+wCahOjo+BQOft4C
ounNThgqoIDy5XKiFIs99ZyJtcCi0BSyV4p4APPdnykjcM9bm6WU5EuIQOMdeUww
cO3Oh2d2wjkaO7Cr6KMFls6Wkl8P7tab/i3T0e9P7rjsoripds5njDF7FR11PkJC
lNMRFtiF8dO7nTiDJjYF4H/8OddGQ+9T4IH68+mzzZEnQWWQteArsh3tXx7z7ByM
BHjQVusAvejUZq8ScKQBJlbhIZodE641vMoXxq+SL7FV3cxP5MU1+S1ddmnt6McF
7mHyHSeEox1XaGSWIb9wywqSedXGxRGiDG7Q6Vnj8lYN+G/RtKR9ODuIJ5bZWXUe
So78ueUL5bmtsJdgxiw9EnLCyRkAluU72lFhWTLUX3wsXr5ajABElT7CMprNS/+l
oa7Z+Uy63d3IgTQoC5x2FvI6qlF07n33EZWRYZYDyRexuG2hIh9YG2SXLQgKGUfF
5HNd79MVnG/k6Jz0mKY/3h46NATfg0xJYY/xyGu5ffKyiLgyGnjHflp8WiwLw2gx
jyN+gQJHt/dR6eFGS5mBSK22JhbxSAoevW8R/tiM7YvtblE78Z1YHCaDC4ezgQ/b
zDveFmUiQ6Yx7FBlAjLjyMcP23INdS+q8g7tWFBOswdizoxh56+SjbmncDPC7m4I
y4ubzK7RLnM2tYpxJ+yJjyuXAuJ7hk8x/elncqRu/kV916zluYSAMLU6mKNQU388
RE1tIa+xZ17JOMJ5sb10P+xYjMv2hLPhDIHnCsFOwzJiq0cKfx/qjn/8MSl33uX8
oUg083r2bIPOJUSBRXTghO5mAqJO7qYpLI7w7lgdtAADb7wWY21yOxTywsO5ZNmf
ikWyA6ShN21iRPmQBHhd2xYiRrZ/08/nBpmN2OsP/puJDSKRl5x8GnWpkwMINpFJ
TEAz52hAdRjFekqN9cHXChWNX/jYKUvGbJbcfiqiU/EbYCYgntUPD1WyuKaLYbCu
yxeeVP2m6jDwC/VZZqqYPWwt9xLzaMlnfQIypbicTl9CeKg0kKm5kilJIZZWtxPj
BrGenuEaxbalkn9hY8O+BE0lpXlkE97AEysa4o/lCpOjHnYjTK3WlTuc76e2Zj14
68IKqMhEy8CkIrMumq2PNIOrXkRWqEb8Ebw48rB3sjd08AbXSr8fCKo9dmWsWgVw
jSw37XIpXZKqO1TiKWUj+0MxwkS4YkHEBTjhJyl4QY1AtZT4PvE8AxS492r++PW1
Vro+9q4G0782XJLgNFhOhc3g223SquWZ0C9RuvPxdQsRARXaV2MUjMpkib7AEvNu
WXqL34E/WeuRWKMrp0JdUEO8WkhrCr0oNT6zPTmToC/wzmbe5IG31rQEJNXz8Cpj
RHsNdROJSV7ZFSQeIoGEvkKTc0Qml+UXBYvMQneLGLl5UHet0EZJ2GW2kLVBr06Y
dytXGllgnO8uTOpsGGzuZXCoOVy7nR/0qr0g3lSd9LQSLM7NaQBFVQGJx3AgLVGx
wL5VsxOrtnhtVP1/uXJQ56q9OuHMtcnTeYB7RyotRStvDgS6NxHXwC5UySTBRVN8
Xf5Hz9ydumanc/K4ITvW/XuWi3jM9zXedCKi5wx9tq48zxIQV+4sbueTpULObqIs
CnY9iOzzADTeiHg0Jp2FIr9zeUqRAGj4UG65X1n0Dp3zkXoUBUr1wwLtldYBHy2n
6HSDGwaa3iR/b8xF5v300JLKkFN6DM6r/xfPrjG2TwOC8Pv9xjox7Vlq9XbU3xJ0
GeZJU7AXxMt9sRKAT5P68OIm9pbsx3qLZ7se38YxxlRPFz5nTPE+jn+v+AUuYRYM
oYBQqOHaFxqq+2kHaS21d2xgpIfjqSvNMDWCMgHSpDiSyChwxaNt49RgaFkqmLRX
XgWwV91nY5DjXIVG1r2xEAcAvWHSQGHCtOHyN0oIN/iyvYpS34KxPtyfteMEJcaf
hhk8IK2ngLw5z11SQDKuwGAsQCMCDy1qWQv208uWyku3RijTcH2Su5ujjhEOtY+J
2S17PylY7F3va++YzbIxFNqPY9fVXZoskfUG0FxuGA10nd4aU/3EZ3TDfVT0qiKF
EeGPki2bDCjNGgjdykQKuSiACrcyoBbskOqsq6GXjlY84Q4UH0M3Nh06632kwewe
cZJqf4Gs8mk8M1FwhjDdlG0djwSBA2ChjrsDSadEw5vl7fPwxG/9SRYZk7KdU6xl
S6WuV0XYMcmzWRF5C3/0Rg9el+EL6/Kmy911BWhqAov1d8GHx1CkyDgWbYVaA8+Q
oiUKKoNl9KyCHZrpBz5PPQgV58NGwrWAPNeDTZskn8yF1NhsGTG4LT1u3TKk3X6w
a92W5sMN03tk/vPeqC8Avgar6YB8vG2ZlNtFVfzgZ0PkBZT+DHLxVdPfOYccXcqt
yxTVbgJFm3uWzmiEGpU4s1hzJfEul74LcqDm48VWy3o0Mc9rYO3BLoAoF/5Mu38o
5Ps44ldISAxqM3mnEL9Cgtz/XJoNL0P4PRn407tMqsl3/8LnzJL91NAb8Wjp+kVK
XNHNRJ+gQvliCFs3QqWkeSZHj5yJIqF554ShTRuNE5ON3Q4jd+Wg3CCp/wOeICrH
HBrRVxMV8UsRzzydFn1J6df6rcmJDTiLmWgVxI+dsygRiqmj8jkbY97nZ75X/dAs
LDbktDsDG653K/UJUqu9B7JD5gtukrmeApCrBAVdOXWVW35KA+vwq2ExJZYtwoSZ
dn3zyKwWvhu/Bl0y7hkaP8xw608djqGuG1WM4TQXSzWIZBqCCw9RvxzVqgFxZLmv
AyHEmJvzWRxxXW7qPjRlXoD8Rk0IdPZ9r8MVJr+qEEmsEBLJ4639IEvW5eyL/UAY
u7bJT74eal8/W/wYiQ3uEHrb0wzYQl1t/BNp9NOq59b3v5ZN8uiM7M4HZ+m0MYxO
DLQTzICRpUffBSnUJYEkDYBLDqyXNTnxl90r/G3wwpnKhHwMAoiDwIdhTRJrDYa+
B+YDNmXdPwDBpPvKWw5E1A6+K34nxuVuAuFf6s1jiarlvdsdpGyrojLdxd7i9Hml
gTUjdAu7Xb4Vep9+nS6q6CsZYIkCJ480+mui7jeXpo5iAFrHjTOZWHLiL0irLfUX
4q6Zlmo+fqtdIyK1N1Ic0ViThr1ebTlr/l25revseFT2ksAksdojfUZGskunqKOW
+ALv7TCs+L3AWNjEmN8/cPSrn/t029AQ0nsJssG1YcGQZ8A92SOvFzDO0XYuYZXc
DkqfUc+lw6wpzA2ICFMKsSmWjrfvkP8ce4f+lcxp1D/GdvxMBik0ncc+a0xH7eFH
SywugjoOV1Ra3V3Z53wMihb5OZiDHkYVgUSyr/WlNSj3q1bzSLkDEt21gOQypaG+
Z3pgMoJt+/+uIKy3E5U3ugN9ihhiV0bNuu9iGCbL/jYYpLzuvPLY1OPUrneq0Rmg
8AocOj2OGnv/3a8CTNQ5Go051gZCByCGY/pEOrDWb7CTIrS3P+VTR59IQ/6ZezG4
IWLoQHqXo2+8KnBPvCH4YWVjMCfjokz4RMHvK81HUGGQDbXz8prZeUa84qURVtgb
xQ2p3y2ffe/YyuocFdPAv+dWIE31Aii/peuIFPosjzujqSvIs83SiLAa24DUoVSq
Bkfh+Xj6VfjLMVRMEaLDs6RKOMJTnuL6P46jc6sBJkrIQVSwYjcU7g/RNaTzspoG
24e9tDqN+UrHdY1/Wj25vNWx0LsfVXfofLo2OlFfPSrNaFJACV0aQqjZwa4qtS77
B6fVzZJBDMm02naxugoH89ByLfvtZ/KkhMhLxFra6NQUHiGi10lJ36AWawQj94cU
s/9nUwocW2X/9aulgJ1QxWcza++OlWJXRKaztwVPAK7cilt9ygp2RhjBJ5cIlSWV
fdhlPKSTi1OZ7ao+OdUQqlHbf6T9BZgmIu994b2bmkCQLrxjLOS6rFdDDjN+jM/5
6CUuf/meLqZ4WNY0QBGXbfQoGbzdWHsiGMQlC9Kf6stOIOOGTT/2VzVJeenLQdf5
/0xIYQjMt7q59TCUkCBqe659gUlJ87LCsjG44s0Tas3t4jVD0kFvegWNjVB+tTAM
sTBabMFweENyxw1qNmSen7kiRYaHw61zxCOgva9VjhLG7lB6VC3axSy4bhep3sUU
bWf20/0Kg1b+6Ped9Ho8JM48IAGzwb1U3gXJ68z2BmTO9mX3X2gI+k5KhvlHBGIw
ELm/TsXWynO5USgQyT6DSpDwmOyQm44MeNAsl4XspPOHdUDYBlE/FpR07iqDyoMp
QmBEj9fGL82u3e1a+LX+WVDFCfZQy3zj3+CTQJwFmOkpMqR6ZGbFifD2YJvUmxvf
FNa1U60XHpjJClIUsiFjfIMvh8YPuA09aYzx+PvmBuSnprt10P8q4jeoENGnA5rd
87qlBc7Zb2MXZQJKqLIS+rJF7jtqh2zt4k4XcQgQNAK0/W7kPL1V1Wbozo1FI9P8
XYOkyjlE96RywgWJq9NNlFq4Y9OL/bJi46oPcdC/bNG/Ew5TabXDMM4OOLadLN9X
dW12/KocOcC+6hmOLVMrMRWAZ9+5DmC9K324uBpWE4SGhSDeB4aITH24oeZRhHkI
JWAtGw0J/Dhjrbz+iljq4k5piENXGzV2gXEXoXTTfhZ+T/pf547sv+EY94W336AK
Ju2pdT5pQ5zxaXZoO+2pQDXJLBpk/+McOZ2A8tmDEh5RCoeAeAJP7tnOi2+HhAft
EOnT0fX8vuKabFnirtZTfFDalGzz7E0X8uJpdRFMtX4+Jhkp05cHBUxQHmH9nRqi
MS6M0lHqdArBftF1g91nAsLfQi7Bsl+heVUEQUxdUc9Bfp6B3olLV0IXSyHyYQE8
EnRlJEk552kllZLCydz92btm79jWqFWSpB5hOyi5khO6UHi8dUDB6GnKB1z4UYrV
auY1RxTJ5rugz5oHmoNRyafs5Tt5G/h3Zi9XFkpHNfII/1UWMXe4TOoH9NE68V2j
uYnTt16LPI46QwuE8dbNAlKxj1OvZa3cROLknPMiXkOXnXhpjvTYoK2O/BlcZHit
QEunU1FyXrW5rOik1w1w9XvjNxh3hl9e2G8afuDTOIxfYjG7Hoo0oJ72h9XQ9nLN
ACIvJDXu50MDhleN9N2neJhW8Aq0tfx0vxfS9Yg2Qysl/IL7doHSeHjC6xM6dmZz
ll6IAcV74oLgHQD6UAdm8eEo5ptBK5fAwTIKvMiy4Q8neVvmwd2y224qmNj6Xt1k
XXuVCfypolnjNrsLb5X83NXsiqx7ZBIu7V8BXhVLxijMNgAUHcXDjt9SL2f1A94Z
RkWBWx92a7hu3U8GNTpSfmFp+2+JA7dBXAcQOpdSU2NqBagXYYZqLM2vI78oyWP8
i6v5TsYrZc9okxeTv8P8ysg6jolP2hs2PsEsiwfU6LPnDRrdhNRH8LuiyBIH7hdO
AHAtXjNrqt79ZlISqipOqXNpTjY/4Mmm7ZWkk1G1lt1wuxDmA16EqmQJO/2552IP
iyk1Av95Qj3GQ01RyLkA553BXb0zsEbVZ+BmBWZyjR+MtrH8Hq6s9kTeoZaOqQs2
oFDMTBKbb8LVL62AuuM2NjUPH4aGj4Ot5Nta4Pyx4S+IGIjxsa7n6eqh633uEj2L
uqDQNddbiy3Y5zZ9D+S3n8Ltx25TaFaKotPzytN0mKElpcZfsgYa126fi5Br9JkA
dPxJT4b7L2HbMIymTfD5wEaTw7sYx63Pcvd/g6l1XAwJE6kijItK0T/jx+MFGXww
tOcxk968uKAibku1f6iJt+sbxsw7Yp3rp4a8wBvKyPILKTGG1xtJ4E3A7VFC3znc
94nh/Vjs+ermEYXc4m9kJV+k0YfdDUvgn2K04ebLscFoVfvMT1vYec8bQlXY1bP3
qakM/q4DdfMLs8cYrBxVC8mfSH84jtg1Kz1fDu31S9mRz5sXYduoGbu+N48wz9/E
7LngB2Tnohhi0O89HrVh2iLwBKtVk/CVhH0CaMoOFBJoil+WPYXsH5mEGT9Z8o6w
RQdCkECqTydhxj/9PAVDmPRJL5Un88W0605wA07wNYASm+D3NttbOao3BWQg7I++
HBUYSGQWw6RTayWZmrrU53l6xfZvOQjSSgcGVILYilRubDjFnobccs66c+AlLHY6
pQRWwSS+OJulO+4W6ok+aQsS6CV6GlEfwP26bp4TkD6/43qghmVRCT766MtKxez2
OdK1C0M+BMDyLNNsjPwTBp69SZzaNXyjhb44y53XNN5OYzL11anlUVykZFZlRAPV
3ND7h9p3pwQgHJfiklY4we6FP8AoKlvdlcQv1BNwhY9X5zDp2+IWIApPgjuQTv5m
MM684ki06xS5Wj4shWEn+5vWApV4QHUQ9xAuzzM+z/69qOUPxAE4iTFpUKOAS1zF
tbNWLZ1CPaWRpvfHWPEG01QIX7/CGNXpLVWusjPZXw0YJtaYpCc9C4VarnmCP0pj
puVK7YGWNIedHHcoGH5tyMmPIqtdrsasL23bQ77/vq9JBxNliJdXgqIKJ/+VAdmt
23dYtwciWNJ7dGD5WXJdF/YrtZsAcS9EFplCwSEfcPYwr5XHToY+whDTzBDa42AG
nytFi8hkKfL45W7sE6FNKfpX78jI6fr3+7qiK3k0f+Kw2v5kgVkAVQE0ysUY2XzS
mItdFJn1aNRffrEsh3C7gbpn562/PhuPSWsJua8LgmuTeO6ZITBtIl4cqzxsqR7j
0M3ndfh1mQGTAzHfMUWCnguvUeaF5RrrZF04A8KwUgE=
`protect end_protected
