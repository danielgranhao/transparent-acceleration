-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
U3cvnJSjtxI5i4Afx6ingRush+CfcNTCAgRODXkv5u1mbV72AY/Lag/YhbeLBJu9
vyEJ2vq4eg4vxZVnh/o5TmRAg7WIlGVPtkzPAJIwoD5D6TJAgHdv7fRpTVGeIcc+
Gf+0dcTyKukBJ8XTkXmVOvIiyKszH/XiFKGkzJfeA+k=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5640)

`protect DATA_BLOCK
zghiSO2E1cY/RbxOnfJd8iHlQITdgl4MJOwc0proupomyLTTKsINtYEatfqP0pSf
REEdojrBzz4GdnDu6cqPjObYwacFpAXRgPj7HUpJcOeOO/nvRFzIEgBg8x/2eOY7
wZqdfoc2yySWWJfs6j1MIR2gF+IE+MJDbhwpHGcUrG230FDqsyz/7r2eGPPj8xwh
80yliszxosa4mP9H/+mj1R0V/K10eE6eNs47iiN/BgH5XvYwog/dr5YUXimrujdj
fdjtdw9mkgddQCMBCpg8LoiYMjZzrXP5LpTEmgzzJfVoBWZGxXsdWqNAo6h6271c
82uZEaAxr/tvokdMeF2XBc2m6TbHwUBUlT3+h38ScA0L0KL20u0Ty8O/VyQbtAmp
6AET6nxxo/+T6AJu8dIWfquMg6Z7txOmkcJqn9wizEb29CjNz7JfVsx/dCmmKZpl
iCnwnZWG693xwbXK9W6TWErhC0j1k6a1iq3i1XOtNulnDfd5h452whvbwJNOtNyQ
RELtYtvd4U6n2yFZJ6TfElZayJ/YaaZ55Rv78VbvcowsFh3S8geT1og0ak53Vv4x
3CyOjWLwZgr8K0kzAXYkPBsmPt6i7+QAYlZWr5ne+Suw87sC+d04D1xOGmsi3ImU
7APELKu9hgcXw4bbTK2CshkLp3htmeAiazDWxMfUi+dWDSYz5mWNPXytOpLLoWMV
f09shH3A2FN/42elQk5oD/cKW59wsFZcZia+Hn1O6vKnNlFNpDQoreqNo1YvhN7S
ACRyZZmdPatsN385ajhIWcs7x0dxkmB29fU7Q3NjeMMB4ss9Pk9pPA7C/FTHAgZ0
vNPQuI1+dq6camwbFFqsrJlGwqaePcE8BXAAFJlSB5yPfqYryj7ETZ44QpD/pdlg
t8Rs60L3KGPhlAwyKCwsqfPEFeZxmC6EDyQfvZDw9yF5fAjZzrp1MqXF/DxImEmG
DUNmYr42U4mIt7cSJ7GJrcwjR9V5FDZHN2h0ZxkzlHpCmeh+bnn9M9keX/1XIY+G
AYtJ6S2I7Qz9jXAk5dV7ZbBLLbdPi9Z2pIbMfmQ+5BjEDgc/j4ySY0rA4UpWBx9c
AKbFqFljJcfD3jM052Ed2Bw9nNOM+IPKOkQZjFVJMEtrKYEXyGXfkT1Wxq4VXRwm
UBtWiZGWkTE/GtecbDDDvr/PmG33o2Jb23uFLhm8oFj2P3A94hTk2y7kaJFOnXXl
av69Kwo4DPaE/988Wt056K4GVCtjvQID3EWumsLsTLMUdTevmI/5ABhdftA52psB
ylQDGZ/Ch4klXa2Eu3XNOGE63divUodrL2053KDrFqmXbK8x0dr+ucKOP7w2+pzf
2rutECFDoGUDSvmUc45hdq8kpNAacZhpVXpp4rdJD1mJKlEmYozZ0wCe1BS5HV1o
pNz+4A/qxsh462QYm2lAlJEzk6sg6kwUxuV87o59rAjKcbZHrG8XCifdHzbbWd7g
Ahqn1UuqQFpiyMVxyKJ+Y9xc2T7sRfiqXrKYaav0YXJZKLAa5JS6jqHv3N+ovUDw
YsDrEGGrXbLpipBNGNViiVGGJsNfuze/HzcA1uRdUiJgA1gXpu9PpW3Byu3+QTDR
93fkfhLpGNv+Jv6v9Q9wrFMS75xcKIxkhbWrHXSgKawF+BX8xSQkfah9asGnQwiw
7Ix4K8g1Z1lkndBYiRrhkRFCETM63p4TKv7tKRLlxuCy+TiH4gukLKUpwx171JMQ
plD6AviImgpDzITMNEQv2E1Ni0WahjW+kTWi+kKgTNLjTD2Cxv+EaFO6WYLxDR8U
exMeot+ayO6Ks05JjQ5VWc+JE7w2GfIRpmHzWcicbyV5onUY0/3a+8YtK403uYqC
LvyU85pOS7rgEEJ1FWM/scQxVeQRtjDk46byWazrXWjDjWkIQ1hsQ5wxYenSmU2s
TYSU/XmIq5ZR6UxSVByzL2L66Ol+sfRonuj7VuZKVxtyf6pfZGzZOSvljNQgCCc6
U9RmLX0pQoMKQ1kJ5opaJJe8gr2nT4CgYr3JEuEOdTpqTm5WlBC0jMiqZU7I/+Hn
IWIOip3RAREvkcQEp3sfCkvnpnJ9wm9ka9R2cFbe/RR6ksBIuWVJI/fHNRsHTODb
lxH/aOh+PoTbksedNLxnTslw+NNJCYPLKCf7HagqSfdqIlRiRZFJU3/YI699+zIM
/HvTZFIXdyQQMgfsJDFAByOBug6KEhFOW/VlaztgrCqb++OeWPHGpfUzryoliamT
WtEO72/CrHTX8vTh0XuEMXLgVx0o8Mw6hSvIqmm6c0j7IXMFJ2FskKjTEZcJYqvJ
xQYzMqPXRO7jBEMUSQ29NLVY/1QS1q/s4IraH7X6gFeCNPlPUQiTVxi1U9Mz/Frb
EuY+5lJbhGZOXWqT4wr10PzNxQ8KKzbHLjDMKC0u98MqIt9tJyaXSjWgKzn272tD
LUB28KUpdwJpa8ogopkAo26URjN55bOXpkSPl7MvZynzWAPqr5SrT2RjXP3d/EVs
Eu9xAVzZITShmy8aIxvHW4/rgKDTm7UO8hzVzoRBvtK62e+Z61xki4k4xnu5ETQL
UleqjvP1oYVr3J7KLJzKSc+AunRKLG652rnFJT8Qi5VlIGWEHOqkf5IzOTVe/IBE
a3pYCwva5Dn8EphfSHFu9hzV0Qk+cefvSMuZzqHAprD0aSJsqDXnDAetb2nBgYZ/
In7nDCD0KZXj+q7OsSTXz8oB4Mm3GQgPif2lrzr/GNcfcb0sGwheFa/qsRb5mBOq
UMtM+PGltUBPLmgnnPwbwz9FrA/ZZFsCIBxIYEWdjM8TpJ/4iskHotOy4pZUCxMc
8Yfn81YmPF4mhg+JX3OAZIe+LM752L29jy2ACHCHiogONBNi6XLFYdF5a4Hu5Uzn
gzHJz3UdP3qRfq1XqCrNEtZ9q4hvYp6YtDFPvPSauT5mJYQ8q28OjC+xXC7b7eME
Cjxo28rG+9EQ/8QxlAaYXbvE/cEiySp8TbebUcdXo76Je3dNlCmfC3yPpCdl3hpg
N2kVvbr+MIGiScuNRj1BLIntlwnKbsGSX/F0T3gzy5GCpdc/PkP4VvukgBvA5Zr9
D3dL3gzdONTyKoG2pArnCQnQqyMr8muTpfTh8ypV+EkKWNQeZX0Pixn4MZ04mtGY
zVkgVJMv5Gg8b+SiP+lv4BxyyCBzNjfVZeUyysuzua363UW2nN8luHIkI8IwXOWD
N+U39S3D4MbkuKy1kbprAe2iYEoN4El3Eypwl/8oEO4PSqKCd8OrHZeTQ9bxgHs7
OR2j1U7uBBbXWCbc++MY0/t8zH2GhoLo32FrX0jqzhe8x8ZDTWsNkbV+s/TP4if3
beue439X1mrUygtRCusu07MbNKKnN7iPL7yf7WQ/21hm1DHsnps0sa5ym9Et5OAG
8kDDcoOjfxQeGFpSAAfuFvfyYPOyGmykNs6PuKUMPkRC9AhZOGCCVsKokcpZOBiU
TWMcw074XFfjs3Fe9NhLafbQGysDtQ7HC+8OBdushmOOT9EtSfH+Npo9tGZ6+oQd
p6AergHEE/N+anep39zPuvycal6CEl+wUGrz6XDixUm+Po/cHxOXqZMu9XVN2bcp
ydBs00D+94zlhxY0Jx7ut64lNKjPbznWnUmuz32Js7oBhDtbtYYYebfuAJ7mTHiz
FznVFjCMCUaCO5AmapRenB1x1P4mQErM17HFwI0BBNivDPgqCG/osVHVxIADQf94
RGXw2XW6nVf8T4pq+R4dzZYCiKPfTuBRSKHOeA2ByWGhBXNmxkBEmiEcsl/ppWy/
SsX7rbTxfrGWWxf7uujNFUxZBNUty8G37AIIvVVS07Ns4gAlT2XakMzmcCuhCozP
TxL7iAPoK//F4Dx+CugESHMPLDGSozmU1zNUc6k6B8UmOCYfZgBLxXjiGtuRFGDf
9Uf7I8kJBLysY8X/bXlAldsM4xz+C52HQC1aaY2ZE8CmHSahUW8EbHyKW43y+M+O
c/vMRbYUV43rReggoIziCsDyYfXprIFDdHni9Zh5c5yoEEFveq/939Bw0qOnFr70
vJlChBLlOKS94neG1w6xK9itIyLcLuX2fnq0Hh3609kHnuYv3MQDCJHxVzBdP5gp
GCF0HPI1++t6OsR/cUBK8whagNU40vFXAx5YFmr6J7X+ZeCZEMVZIOE4s1lIo9Aa
iYLrAoxsx6AHqbHZuDuLkIjICfWuMBrpBH3XydOfkMb1ILwiX1LpOU0MMN45HvDK
BLMvYYSfkC5TvPCJQaGKhjmG4h5ULcBF/laph1V/yjH90SzBHofhx4qfPTnvXkQV
9bALenHmRGZEjlGgN6yS3Ofp5notImUOvtz5ypKqiurlcDUWp51wLGu1TQl99gNL
VirMsB8ZtUL6Unrm+F1jrMn29R8E+uywCYfoQnZl8mnepDB593m21hM37SDwj4rl
vgpdKTitw0733Rj1XRUB1bCskS8iVmIyXqVTmVL9UW2xon9qT+bMHKu6rhQouxdp
13iE4WVy0Rpq+RjTZ1ecOACH0MPz/uEyFtvQLQnKmUzrPnmxumYPQbKq4weuTWp6
k0Ri/P/J2Xmok34wq58GEtRpUqgeqauwvP/16CmD41eZsWIF+YgU1Hcqm2j9Sx4r
yQ3/s83PEjTqr0mlkB3P5SNjuueaSC8fld/O/MH6Rcs0uv9RjYx+ce2QQR0CV68Q
LZ6eUcPW5WSfhFoYcs6qVA6/YNvPrqMF/cptRSpm9w1RTHwehHUawbC1jsF8AOLK
v7wSPJHS9jmakIIriEo0BNELrv1DOCGKBobIZe3BJvS3mbxdYIICG014Wl3f3gEF
frgmdzrC1ULVXKbHjSAOUn5xen75pt5uyy/O29RxNyyg6VA51SJIHSMCfKbEKxLM
lsOo34JvImojwCcWe8ADXXjKUL5RcH5mis9mMZ+1j/0oDNqa2y6h54LQHGSH8N0M
pnYUr4BSrAqJl3+Jcz5Lyh5rgzN/Tlk2AbJ1kX5paIOHn/7A7cUV8jaD9VN//as2
1q3rfES54xnkBiNFbf+2r3agDDrv3Cwhe6F5ZoEYokTINV5t0I6nBA8rQedsB4G4
pqGagX3YJvY6cq1jursFUU0YtJhg5/61jSarIoANIGUcdc0Izn2FYLSR8ipR8UAP
vkCSr5+AR2bpobBosCm2WSDQCFMVLS7WC6SHQwZYe2P1amZExgTCvvhWa9i2T+es
zIVjmRYsFY6HfOtglX1fbbfHZ3KbplcuAt//CG4TSHEOz912J7yKHe8VTwXFZkIK
UFkrgsue/AP9wShq228T0ofeBn50bwJR1b1nZExtwwZKXKOLqb3RPILZLxanh0TP
PvkiROiGQnH91jyvmSihTwSlctHWw1L+ZWQr6zSiATXWb3TjnmL+8vs9rfhEu6a6
A4UGLrHHyaycpvWF6h7BJSN9FPAH1n44OIS6AIQyrY5DH7CwlC/jW6f0EYDkE12T
uXmiYOCoC9cePq75RuXk2NxyhCuq9L169uC5wIyQkmewwpcM7O8dOqwqS1Mu0E57
PzRqITvmkiTnAud+i21Zp5BXhEI+COuX9ArkMbFjTpXQZOI3acwHxv5Oab9M930/
d8YUqpUHDGHieUDKqk5+aXamJPUyTMe+eHr3as0j0obT7H0a2OQ5AqM+Tm5S5l6H
xVg6JyDSqi21tVms5Jz4+BGPWXzKlOxI6Gq2PrhzMFN0LUQNN8DXXdewW5Nkv6XA
ZqeLXkIliTAuEkOiLF1sBnWZ6DOLFbVNweXrRZq/vlZuHJgE13VN99Y0NscPnkBH
v9UjssoqP+VB+W5D738Yh0Gw+bN89wdllmwcJdadZxLKIoO/urSWsSmFpWksjQI9
d/XkTBgcLmVcGq5HEys0yX/AL92TRsmyTZRte+sqVQo1KPqTTJ3u2CiOf9hxT7J7
jCQgMSAoO0AFmDRb4L6N5iY+kEOgxqA2YZQ2J7VnrxzQfzYbh79JEUSDrGrogjeN
E9cntCUNrW4aITDxNJr6UUcZ3NT4MANAbpK5TXOrT//XCrqIpO0TRMquB/tVVa84
bcESlVAGbRKzcaECGoS9wh19sbZk1N7h5sORknYA1PudaJEhKqpOVNavMPa4wwuA
bNYWTGztIhbppux+kTUz/9VNWmrwpIndtFg9oklOtwT4q+NJ35XOD/U8RV+khCPh
0j0X3KBK+P2RsUHsTaYDy5a+uGWgbUHEkbG+Ll3kVp/UDalm/iNIu/eW2Kl5gLZ2
hSfv7Hbw1Qvf26NsZnBOSV8HqbZfcjfK9M/wanIyMrxDi/UVhMls/kEnPbrPEPry
KOLckTI/dkfHgMzhSoMTfD7G16nr40CNedrvCW/Xrf09JBY0adQEg7ngHD3Q6bQI
+WQ0D0B9CquNoT+J8mskeu1E9EAt+eVXOYuTF+ZAyGU///4mXLMf+h9pqgdf634X
PqFc8+pMKlyrUluCqhm2Gu4UdFCoxTsG44UYK/IeM76j/Mz7Ua00tn1VFdkq9Duc
Qduqjb3waoBxDM1o+WAuC8sGKoCCjZlQBuyHmnTwspxNUDUu1UPCSYxGV2HXsid5
55JX1zOSHnb/F34EodF/7L/uG0S3ILDZ5DcVLXaRYunBumoSz1n6LeYjHf3lewrI
Gz7zODtqUqVtUGIcTctdn1Gynpxya4WsrG5p6EYsFhpk1sIYOg91OZ6WoM3h4hBJ
ZYb4dZQ7nDkP+hRAZSuU5WqJSbCLmZsjN8ThRZc8vCrKe5Y3Z67mHmWGQUAOPYa4
cPKTDyX1ZyFDzX1PowI0z8qoq+II4ikuIYxTTPgL50GPJN2oOJM3o1lgzlY4HBvK
JpWDyDRG8FmFQzdOlyCdL9Mo5tPThnPQh/kc1TGfz4p0XRbRdGOyZqkGEmohVWg2
/Fe5m7G2A6tghyNfnXizeQiscCMBnA0ZHqwEnxxSSlbyqUZsawr/NqzE+Ualksxc
pLFGDdN2LFQsJeotzmaE5+tV0Ziks6fjJC+a7hCkcJNOEH/yYPr0qX+u20vC2fRv
MnsyvKWl6Ai+txZBFoNm1v9q90aQf4LOK3N4L1bL8EPtTifH9oojahibY+e3X0O5
roYbbYeXrqvh3AGy4TVIsw8zY1PuaT5ZJiC0T22qAbfI/5F2Ya1yBg6rEvbwgD/L
ndl9g8D2kI/3RAdrlrKz4W6p5VYdf3qGSiVfpSKLrXensd5MHh4qDMnRixZ4Umxm
VxAkeEcyxwlMurWDLYcCHzXD8YliCZrJKuHMxa3dpdJExW2SrI1ePVpGxyuNwB5L
DL5/8sSgwEOQB6VYSb9Ec756UMJcRXBsDPS+LUh8iKB2UoNa5Ty4UrqisGGG3/nx
FEDUrNtSWMCnQTxrOMakWYRJi/yGTbLXO2CKJarQrQyShkM4Tz6/IUKq4zzKein3
wUlN7ykXKm0xQyrz1li3YmactagkWB1YvqXzBb+NZhv4HD9vqhEKywGxHtuybFO1
uVVizIllz+kH7iCdBrypifKhRD4FoXZlJEuWteoJcePx8qpDbVsQw/CrW2YmQXil
hlQDqtv3L1a2LjaWyZ/jyiHjXDbbj4zzwf5ynh79mgn3FaJBVyUv3sPmxbf9Aj8O
`protect END_PROTECTED