-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
L92sCUR3i2T81xtPxZLItFQhgJS1PPmrykB1Jae+2hamBm89x71pTqxKB4x1TifO
jx7h8CQGg/UQ0VBF1yVQnj/CtyTe40RDYYpKo4e16OeTp0RlRRJxttRzTvhZDAV9
9C2aJknHXiiYwbyc90MiIQRZqZiBDzKlCvoHBTZq7k0=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 21392)

`protect DATA_BLOCK
5fXdMIDPu7dWNLZEK1AigsAfYIYPNGHQ5VO/SlXDIMbvy/UidLTYiyjrS+A7ieJJ
KAXMoB9h3S3peUSNJ7mdyFzoauXeU/kPYlyo7sxVzkzwFqbfQ5oxwaDoUvefKbfw
PMbQXa+OX4QnD4buQ0oaYuuVKfUX7DZTDy1j2DdqVBGXs9Gu73A2xY5i6C5KA7hi
5mClUj2I1b2m+e60KKdA2LQ0hOZOLf+0OmAxLeKFI3h+JyPwo3soZ0PLopAUQqRg
9iHsrTEKS6LUf6EVYnQDonfFmuljC94E6+fQoa5N29/tpsM+XV3YOll0PHf4wmki
zkft92rSDPomGR5ZpqR88/UnDsp52/HZ8IVmVxRB/HaSLXmtNLC3fbs5rILpODL8
zyaPJdN1npfsD/P7VpxqwOPukWpX5QEfmzU3TtuR66K4jcxeocRxCqO0ABXC1Bv7
LcNtEhivRz+zBmdX3F49eKgfHAczY66GeJmBFGmEOubqTXH/XT498wtOxSJ9iBkr
+RUD4mzfAJ+AoV2F2Wr9mUH/JgtGi5fkEQwX8Yl1TZszyw0VOzO9Gu2aF3dBkKxd
Tg+7F5jtMaujw7crLVsJxYfDrszmK4ZvoJh0CFhu9LiEFD04otod9nytO0j+DQcP
Ny/yXfwxRJ0oWAXh/esgNSWRylvnthEF8qA5rmIJlpjWozwNjdbQKUTruRoXVWzO
NNkheJGJIYBcKZLmhz2XetiMLtqW6JpOLuFrkxm3lqhb7VbIDVqATJF5KqgG70z9
y2OvJ+BMSNgoXJMBLhVt8Sn3cOTO2gU2dPuOJ9PqJCC8FDcFoFHJhTy6JGOUN/xO
pMRrhZnThHtQQxdLfqb8TffDFNeXZGQEdg1/Dk2+OlNFymgRywhKgGiRxdb6Y1bg
ag5L84DKhfhSleFx8kY9x1omghGpdPwN17dEtJJDFybx/ebtNnSvPlTOrms2SU8d
dPCUNVaAr5Jel99hI+JG4gAugKv80CDugUxMSM4p5LS/8wlfw8bU2xAVoC463ezL
YzGLMF1SDVEb2Gnf12OBssaT3warVWHtYzjxrQVmbJmZ5+l5lAbU43/+C7FjvUFW
TkP6gSQy/ehS9Gp86XXL1U1OR8HdhLykyCafmZJD5dsZMqigFNuDgfYIGDuIyZwz
tAMSNIrindijeqURmU3n8RrU+Vwn5XljRkaQj0VrUgxtuvMEJE/yiz5SmjGDpGdD
K41C66Tfmy3SePYf2GHlVXHwPjfZDakqKUFylqSsDFff7aMANngUhyHEAj1D/NBY
MIkonacKXGlEs4qDMe2564+kqzG4vIjtTH2cjgDXnYAhPiR3m7emwICRI50yA2Jq
Idi23Rcdg/WGrWbH+WvbNTNuAfPTgjMLmSgPVni8UxusAu4KyZjQeQqjuV64ZF+f
4oXdBvocHfOxnGueZ9H7pqVM5dSJ4ES45fxz9xQSBYEZEdbDR1/23NR7gRpnr3EJ
GIz1cn+GWK4nAUeBuIzbvA4GURQPUeI2b/ovzRzUTG1P5ZLTEvddUMpM0m7Ho76t
FyY7AdIbH0hRuEaCit3zIvgG5XzUZZREFPcVFiFzLv7IBFNOrqgVfOJr8UaJ+W5N
i1fH7S4sojFSMJ9h/DzNdzgbOZs65t4e4y450kNeWkRHwyKjGDHa0iqgiG3DteUx
NwZOGElE7sox43uA/gnYbLnFyA2BS/Rhr4vrfd4ItvDOxXeM1uc2abwcZLXE/0A/
4f7XOzBQJLZ6vmzVsTCxhsohI+YFC0LfpNj+/F29GfkTxiPNT0eU7q8NCZcdi4O9
6eywVXXKQT7fCijFWfv9ToJFj7glClEA9BoZOy8ihhExudyNTXiC+Ey+J85fmLBV
4KaS9/SDozovMQ+DT9LwCGpBgiFilkO/bSGzDB3QKWOYmGHppBQc66I2zrarhwqL
Pqdu5tvGzFNVnSNCi3N5N4hwxhFa0NrlG3LhSK+l1ZaQcaIGUZ2YfcEnU1NtIiY/
UYE1fzrVgwfEFepIlH9/L5pHMimoU1ai0t1OrkF4uAjnRr8W3aHRhNwGc9Ut7gLL
DDeF075njUHvYVNSMaPwAWzFzGZ0u5ACuYwbcGssygSUTEP/Gt1pYclffdXg9Ff5
UEBv7FGV0QtpwQdC3nI1vkCHrcZxkQQTbXLTySY2NjjShYaj06SK+210VdCHCQZE
VPm9eb5kzDt7aKFHG730pArp1hT2p9VLD+PbRkR84WrtzfoO8+iH33QuGNzNOOeA
whJrzmtSL798EjW0TP/WbdaSmZ6y8atvBvUWwGn3SjHpW97o4o7ZIfe8+q+6XOY1
xZh/C6uFxeDQp1+lyIDKr2E8CNLGQP+ShAy+lCtUQ3XyJBEx4/wnf1EU8CXJSYDt
oyOJtV9DYL3pfUlJ4lrrW33k6Pcd+ItJlwx9E+secHII/uqCINzXuzrS391bLXsa
SDow3OsZucMwNXDdKHNlToWVNNvOKHvAIhnGMSSsaonrzHhjJ5hw8Ir2ao5SuTvJ
F70cIgFrTAvTZPuSUqXd9kXaJvqlfmVZCoUYS2VtROOHWQsLSVQF4olofYSZ2HXb
9SHsx6HXZEsAf9yZLNMQpCiu5hUBSLJ5DrDiHQLxe/km30kx+eqVO2nHCmMjCPwn
SqJHdDYGqntap9ufgw52b6eYIFvEO/1T6JibrInGFXSrUbRdEt2MIGJrqhFYVI9B
F7mNZreXhYYxbjKjcNgSfGj0sOyqSul9PTrKnJOH9i7pxBhlQvrNtXge4tbipRlH
fOF86lEzAUeJj4r2n6+hi7AqbI/juZCoZXe7Nqjr3YjVe48Uw5G0dusX5USCYAlu
9eeTCly8SivZo1M7lAmOzEH6wA5L8ojL21CXLMdN6IOXpUmGL1eBZB96cNhRwS5C
+1w9beqEm6KTjkpPJVZ/jt5w0TTmbjrNBVSLfOpqOjNi5jWM0tlaanNyr21ZmoGh
+1RDV/UhieekTFIMnVEBPV3wFvp1wCW9hEYL/eONDXZ3d5e6DSpcR/mz8CsF9cAb
AnEb30ji2O/5GMO0augoFtNtqWsr6ntXQmT2nl/9dgWbqPuDE32gHkY+EuqC2vin
6WqHtsgyMr4DS1y5rciBX1+Ki6zcqxZnuIkN/1RJio/u0q3M1LE8kJK2mvDcVzVw
Y1dQcAfdyhUOuEo04/0cHuYKLQqISO2T8jjHoyNVs0PBCjvy0sD5AflYmnaaUM5Z
KqF4l0IKovxCz40sv0KJeg/u2nuBGSPnp6J8OWnLe1gDTQ2VoLsAimsN83wOJTWO
D3ICpl5VhsnOTVtejsU5heiTRtPl2M58U/vIlSDUSg8jmtPJqwUl/+MSGHuocjqX
h9G60oyAHaMUJ60C+5bqZM1vje1Z/yzF2fnh6FCd5dl15pPhEC1J1hUctVArpnKP
1hAV9pi3kpuQVyTy0xWTaAEkpACwRchvIJAfcHB00FElLR/IZkUUv0Juycnayt1z
gxAecLpGzIppm9MOgyr8mHvJQebpA5HLZ5TSazQMNZUg9ZI8mx5UVhE6tzd5jhRM
cEwhsc/rNwdG5PkfprkbhxW7eo1hHNZpcAo0dLdCCyFuAD8LdJvXy1aR1KKM8Eis
q2tsTDF5yrDdk8thgvYlTkJfLpHbmHt102MrWAGBCh5GW2jKVnv5CN6+wEZxdasQ
hjbLIbSiqJ9fAy1EHc302+j5t3Ja+02mL5Kq7bNMR1mJfc97jCKTJfIosTMU9Ufx
YdChs7CTPXTZ6K2gxUI7WYqIiASBsbKQ2Q+A2X5loBPNUtneNtXoEOfeZY8AbXE5
2dqpSxm8LcVCMoabDg/vDoK5WKAL+XezVVgiayZ6HdUBKstcnNetE/V8jb8PaLBL
e590QVTJ/WhBMFH3MeSszRKcABIrhTsbwxd5vxlLbkWPXv+feshCrL/ILDcjNefC
VMdnkZrdFLqUotWbx7T3ZJ+P9hhXmS8C2+6LmG8cIxdecNAGvv+SjVd5xO8mBizT
tXsDv8rImeA5caP59vPEhATc6kaHNQ/2sCF3ynOGHUpQOaVsWxKjalK3NQrv+Loh
S08eZvXqVOzAn5BIkwPq6YKfuenT1b24p+2fn+3FT2wv1VlukT+zeIrmTKaVPG1Y
05c/T5cESKFz7js2f6WJBtrtOYwpY/qb6oAoiRpPgdtzf/LW6ZW8r+nzVFkpKCa/
wy2BDDPikBhgEYMWeqlZ2HRmxZ0UyQQgwrt/rKtt/B4QEhtRJOMm66IhadIZ7cUl
HuifkXXCNKQCnB9o+vjTFDfnfFLLU/l7kZIPY4lKY/V6jed8KNgFSCUTIhWPw8nA
BhA/t8bl7FSjsYmkVGmm2j4RrzH4SeF1QsNu7ZfDHNDGBQ3qi1awrgQVDeerQXXP
Ee8eULajk6van9z7i2IHKlYXh8Vy13ryNmrNk3o5uXj815FHx1Oo+kwYOGJ9XZvX
Wvt2ROf+wuxSlL8t815QbTIQO6Lx/Bv8U+T9oAaQpJjTjodMwxg1x4/zXenQmEDD
rrvqCkq95Zsmg+ljzVlYNhgFbl+nPUAR3OIsKMWwUIvGpeXvrDbyOB0ezzqgx2At
tokW+5CSfvQVQBEbvvkSmo/Onzg2ZJ0nJvb85CotznPrVWKSAtfwq/kI43z3xUQ9
//uQuWqax9POOWvjwP/oH1e5o2oDDtdo7JVLXj3QLc5Gj28EvU5eDoYXAtsYR7PP
jLJ5DZ2ysviobXduCRfw3jRo5WiJBTFB12W0Nz7q5qqCN5N9TcZR/6Qw/rTK4fZK
Q7P9mEKXgxyN9xs6b+h9huZH3mIZ/Z5IE4cUuhyG5fjirmMkiUZF7bRo5Z6D7GmI
Ngw7F/CBs4gaprPxqA+qQD6C0OcYZNbPehAt63CwdzTOPTKQjEWw7ZBKX6QW9LkO
T0DPBagj7xLPx2qCC59fBHM9oUnme4IL/eKyvHgm9yYn28SpkRyi3QbEKiyg/4bq
h9/QqwCkWy9wUBlWC++wTwF+k80/rTW39sPhe/sY1fXgI3e4BgojEq2cnbCB3cSj
a0YX85BO2tT+teDGazdfz6FK+tZKl5Lb8wDz/gNCcC/bc5vz1VCcrVCGqLYVVV44
W5W7Vt8y5JlTTo0DasLzzXx3xSEXxEVBMzpNOz3+OASgiNPMOJZGbn5BPevRrzq+
cA4FvvIHxmXlBNSITM6sv+XTgqc3DefU0et06Yk/eQtHOVq4wAuKSXgvyGuYv0U0
L2Os5Hhm5d8hI7GBWQIOnJHVBJIK8FhHB+pR2sUbh1yLeP4TXt4rJIstYYtCnFCS
MDHN3apLM/DRmpOja/DYInUuie2BANLpXZixscVXlacPqo/QMeD5BxN5BZMHFJxi
qIrE3/NMExYkYtycif5F/lQGDQghULA8Qn0IQBQoTQrht4wYLG6KQb+byvdZXyog
5mSOSsBJbVsdGQsiBAMfQb1Qs0PumJCX9+cRZK1GetT4oTHQ8JlaIJ5+9lNjrQUn
gXTzYRd5iLyS0JR/KOAg/25JLeF/mTfWV8BTvQ9YFIDC+sU1ogUJ2y+7tczNZnRi
4qumC8ti5nR9Y32c7ZaqDHO55GfmFf9CLItUq4BOJ0nNyH3xW9BTR6zVks3E5jJG
aOp5zW6jyu8kXFLsalrdsvJRTkr7k/rPrYtvMM5qNZ7VXbKs14o1IQhmi/VYAJoF
cg746roJUuHATzmHNgs1X90UdrDUyxNafl22lUby4tz3Xxl+VmEVs3bDsEfT8NZX
ahiq1NDkXkURNOJ5OpJNgoEkLy2/z+m81q7UGj0JRqYEMfXg1tt5P4uWzFZ7aQ6l
dVevN4RvEyuQejezMOnG2YUJpJveI5t4lrD6JUNkizJhnWgnT4b2jOdG+3PtrDA+
MZKqGE3mUX36H8JGNaSubv0wt8gDkIkdby/xErWXiy/qYpfOFBmh3PwSOdnRiRCV
pqlWjW+xrNUeCBX1xJGLLTQ3dYz8hbImwKUxrd73DxTCWwhCAd3uJBfRkJTWyPvb
cP/dN1phskc72/aSQHUtb1GgUJq983PvW9Ucjp5oc5r4cQINczSjGgmZSYVm+Ns4
cVjY+gjTjfmLdVNk1c40cCrqtB29qumEMw+Iw8DSnOwDouycn6OKFWt96aP3e/wK
zYrhBTE2StqW0ovT3pQ7yxaNDsmJ9KCt+ojWb+LwbdVcgpo8ogzVEbxL3L1EBca4
pVqpFYqr8bIbREvI3sXIyAB8rbqkR4E3KnTo0MrjYkOT45tRCQ4BAvGNvtYyJHZV
YZnJ+ryfMhThSiwEjQFhN+0kAcPGHQ8pEpc6xTu9LvvlK2/CpUqIh1JT81lldB84
G8EIYb3fYWi4wzoHhXD2OqLdypl2xdxX63Iau1H1zjo2sOAPQXH0e8DFH8myBPZq
xVl7Ma2gBJBCtkdSp5WU+eUl2iMhcITsaNoNE/kX5y+TD09L0CYbz8kEv7tqgRff
JpP4bnNR+4p6/q0FvYEDrcUYmVpsRLSxqa1ARBFtRyKuO05AzZkREq8R6SJgSiSo
CWTlfCys1+nqZFLtfL7S8QULCoXy7YDj+MO5JXmRWv7KCpb7qbnYdbkGd8dFAUxt
KxnngEZuBb6CQhkeKelcPkTFZoPmuDy1bGfYj/DJ9X/ooe84cNYD5KFKXx5N/Qcx
kaKOccvrVEFTJUC0O9ybhLeJWuOKvdIbKDQqsf/X+j1yMYi134WuJ+k8f96RRcjd
LOS9I2NRgp+vZGdrq1mGz9vCs9LApHxqcWEqdj2KmtdYIO1TbRqCEuJw7zLss6rc
TX5cjw7Eh3iatNMsKEgINJPkwEOa/mip5jFkeu4mAd+CgSsCLZo9EkbFv+9HprJq
gzs539s0XQVnISCW6ISmJj7OtzkPo8cgk72AL7QbnsNUVHYy0Dp+LhfDCXydoxrL
A5qdkdZn/45PB+13/XRRLv19F68JQHjixp5Cra/JwK51zE48G1AifSay6BCBN5Yk
IfaSOIEAfsLSKDfKqyCcBvzeR2zvIEdEvKyszI+DAVxwkaTZq8mUwDkKoRC1/tCQ
CBStrqHBRHMummQjNjGWB1wCVOC097GHHHINJNHvT8cP6FhCoe8V8ZXtP0WyT9fQ
KJiIFKOEA8Q7O1lvpJH2TuG4JZWA17M2Hw9XxBct7JYJ9UnbXBeEVwpSxtq8AZV3
fwku+dlexyg9bGVqQzF7jyouiY80k7MQ6RTkX6dCzJz7D/tf0lJBcj9yHMjeAFoP
18/pyj/9oCVmSSv/yZ4APKa2RzUfmHCfeXQNUMyz7Ro7uiy8Sa4LMhaVP4N6Sois
vm5WTAiI9syMKyUTIPHnMhRiLftW4R0H+5Mh0Ti4XhHGG088BUzV7R7hNGYHUEwS
yqm8cRFhZzvRpc1Z7SE9xlvYd9oeDCJvVgXVfNK61A9Vph7MasouloJSCy3H+JMe
PS5ZYxkw4Wa+qAnSTR+sls7NBtbnBNf0ZR1gItUPwIrqgKh5dfN4s+6uQciStdWo
2PRiyu49sAnCzZCNA1e9oMQIk57WNoHedFMF/HJJZtHpcVzWsw93SoBjy3hNwxGM
w7/1qi6HJ2m/jR2QaxKjrdPBi4j6C+WRAU8cKlqmb5vIA87e1Cfz35NbrLosfmy6
MbsJrSmpLg54gR3wEf8qJzQddpk+UGma6TaXVOEfyFuVA6Xcn3Ek+ZnlwBxEphdi
TO0ffvI+VgDeK5nszYPYUfPpsaCfpTh3GrkuQETwUFjx/twQQIEPIwichi3DazIm
HSBX5U8+SI3x4uVqGj6WVg2ukZRKeAMqxKVo04XBeGB2kfV9aegam4Jii775GArJ
ZknXbeeoKutOGVITTepjiN3bQTsE11J+/3SP4udDnJok4yGhQ4jsiyrNSGln9mLx
e7SCc/EyjWWk0azTrFEN7DHmwJbCRTZM5RZ/tNF7QaNq56Pmq5fCZs8bmqEiFc5P
rEQ6/mr3s0mF6AfiQ7fKqJgujUfjPQcSi4IIKIPFMr1tGoaWOGjl7MUvW9c6kJ9v
dF8Y4tJa+/pIBeEuI6ynVdVL3/ejj4E34HoY8IzFE74/HZ+SBBVjl5Xgo1DN/Moj
F26MExvIiGISymGWvT9QMfFzqrzfkbF3ExE1e1SLfYQO/GEAZ40ZIeNIqhxqepnd
wZH1B3fpd5lfL/MrSCJmlBf8PxTwYFq4D6ihzIYUJD0G9A25CcFzqVeGF4WlUZtC
tpXbINiXLkbQ5nlUFk2LrrOxuCIgJGtKwTgOvMxMEUYlNwLNltY5NspJ57Ekg4mO
Eau+Rd+fMJU3QZ2/0bJ4IbpaxHbT+rrfGB3+3c5o22F6NXorpOrNc0Z6bqt0C6WS
JriCDXQnGsavy2WI26jV9mQhSlFRTpvtkOQHB9dZg0/JzQBcezVz04pRlN4ktP6G
hv09nr3JsuFqZCbpLCip3Nl7IsuzHGbkAgBqE8NfmT1aZytzFX8a8Dr0oJeqjQH+
Jslcqxf+Aj5QgDJLEDX7Z+gPC7vBc2+LQqXuR2m28WjKLamNRp7lvGoxa3EYftB3
OmApkS5qyl450xiz7VQcLYFARRqlE/6gYdCgNKlYUgDaQcN3sDIJoerf0DtZXHhV
ogzrZicoEclX419W7mTlosq+klmF1Z87N/xFZAAPZQs0dqCIRQnr88uSlNcKnGzd
jKTP65WMBQBgF3UwKsGPhnb940gGAf+wNDuQii3oV/uYNkhFX4+USwah/mVNosA8
Kt5pAGYEoa1rFG43ein655rBpQwT+MlPK0zLKGijfNosxjKjtHMhRnQzr1zNoHrF
pdPepEPmFTxx8tHqDv7SQtq3BW+ZQBniUPGP9YN27Z4t6VzceYO/rbD3H7xzAUO+
qovSOJWfo8xTaCP4SZgZlt4TrddPi5UWvoosKymsZ9dBIgKMq57s649Vn4ppRHE8
csNdIAzlnnjq+0BBMP969OEcVnfaHbotcAUmBlUwPG1a6e047oyKl7uw/0bC6rkD
J9dcvd+HnT9IseydwGIfrKl+6JD6675hluDhHTxUHc2M0S/sRHQ3DXW/w5XkOa86
V9CjW/wruM9aTt2e4RKsvTSw5Gr/acE7pYtavT7x1zrI4fuiks4ny2pftfqujzoH
EsxByGby6lMwatsVM2KiZwSgJEaVEeV4md8FzKpXWNmAsXR210NTvo4LIbHe9to0
bxevrOwCPuIE8NW80ENuyH0UOBeS8Pi9hnjinPglSGixoS1b5h+zV6gFfVaowyoy
n4UBhsDU12442t3hYMaykDrBEurRCxOo2Lv/cA5rMNqv5uVLGQWFAfLGJqlFW+aF
WBoMrRISK7xavG4MTLFdV2vh+7TY0H4QbqtlBDR49ICl0nymLzRkHN9gTc1KQnPO
4YfThMwX6pedSg9kb9/ru8coaBCal3z+mv60O6cBLgjI0G2qcZKYQkq1ZMLetWC1
UMV6fXAq2DtnIOIFZXbte4Lh88e84M7Z8z5XrdFy/l5SzpZKf48FG+9yNB4TrgJO
P1Ie8LRNVvoKBZBCchRtKRkVwUhEm3QGjTiWmJnXHEtiPYGoWubMf7/JC8F8T/Bl
kutZS/rshPaHrQEn1vV7YOFGxo/yYUOEC4KFOGv1vJcsOIAn2Fzp4flKdfpF6Lw8
Z+/lCoD5K6ZJMLBN9j+O5bVddnZjTRmgK+25/o8wrXhH1YWMJ5fwhhdChv4x5ud+
tAI8iZNiDg91bQeX4w93YMc/Snqt4b4qrv1iTd7FYR4sqA58MPqMDUTjDIJxh0vR
UWzPJoVFnOr3fQS3imxbBrmGyWws1NhZdko+4lswQ9iM9QT7+4IOovCpiI7FwQOQ
iBRb+kehDhrP7a92As6W3om45bAe7I2krSIVMIFbSYov0X7vMODa+l14AyjF/WKl
KN0Yi9sM8ANxIvO602UbJw6ZaqzP7JCfq2MpqgMqj2eK7C6n658Ead/pXNM5xalC
RtK817JeEEAxF8kTFtGU9tGiJ0O+ptu2ihw/jwzzFh0JVYvTDIdhXhbRCw6TV1dm
Kv5SpbqxHx7FH0UN7xpYl3iMrW8VVpAbk0AFb5HhCcoywv+NZJ+9wCIxPLkWCjJO
sb97BMie35LbYD0XZGo8EtmU/BpDGWcipupmtBez4XyoioX9B4ohwnImMlsUtEQR
sBHKUZtpfmrSVCqxUV1af+c9BacU+7qxuQm6vKSRNUNtkdPfdyulTsBrWg5qBJe9
QNAG34+vy9UTTCgC04ugH8lC4+iM7qZYixsOsQjnrBejWmLAkSOazVpl9Qn3tKUM
03nMRPeKFVq5H9X7GZqCAKu8Bea2oUPL6IrrUB9MQs8s6dO933+QUT2OphFof0Ok
sbf3zAqQdnJnrWrmjn2Rbdw0hS/4rWLk/30dHgb/o/LWUSrZ2uY/Micf5wPwHj/5
4KHfR4B0cq0hgxSy0tGs6c6qH6LW4iY/FZfBHl6EhAOb9l+zDdFhHzrGuEwBRzW6
9ObtIOJcALRGqCJwTkXhEHO0djSgfrp5oagelAi4ERC5p2FI2ppu6hsdeebbaPa2
gkWGTCTObRyRTm2vwl6a6xeIk3EkHA3/6VOOh+zIhx0Z4npBJy96AWfJ8ohOjcNw
3ttZHTad4r7eE3Ah8JRLC+/g46YOt8iKojzIb9aUNRSo0c4WALcZzD0RoWkPG1GD
V5LsRzvKOyqObFWzrRU2zUT3CC14Pj/FGjD9ZI1IPQ26x3UWKWGPp3hFG71PhVUZ
Qm0Utq0KLKRp94neYnG2J0qnFZVnWXBh7vCbSVJUq5dB5YX86Bu1A8947YXNHqII
X+VvRLd3ll+7NqtSot7uSm13PfB6vuQO6z95dX8TnUMTkYLL0mBNwsifCNutNBeO
O61GvabQ9I21/sGk7+sHm8I4uJSnsu9f7qkN+rikCO95UexQXdsDHAfFzVjzTXYB
ICGOWIL8aqg1NEEZZwm3jzNc7LtIppc52dF8FammbmbvPCUz7ATupr87x/MfpwSB
BjboEFiDLJc7/RnaoHMDAaoxlbNL5/xAAQwsrL9NV9Xf7GtMqVN0kDxKfnierjT6
kHTsKpRSMukzCKLTBSi6MBEEF0MX1dXQHC9zp2GMxDqPq4x15BpUCY7N8/SKRSkP
zHlW+L3xqyKq8xbwkl0FP2OeoFXa40MA79ONUx2r3RTus7CY0F7hlsJuNGDlzkuM
0zBmOJ50pAkBH1q7ZFHG1a77klAbyEVogXeo3fX4oIKgSZImxKW9ehM1V9qT0PIP
DUp5QQFcSrxqJ02Vj0yUo+ZUUf6Wfm/Mr2NiiC6dPxb20kjbmOls45B5DXwf1RlB
m2bJJmuh5sCKuYDICltCfQF9WSvcvdF/gGHGtKmOqU/y5AMOzDmw13MxybvfXDoV
O+E2ADzyhVuc0EDTWtmUAllfTkZWaSQfviVNAc7MpOcwmFTKJ5LaLAaf0/Xd2wKp
1sMHKSIm7S+0tCpJeUvUJbOH/Px77+KhLYg0Thudap5Mags4OALaSvyMPtWgxWS6
pO599IKG+qUGCJmsNnann4YceDQDvSc8dtzkY9QKHZqI0Vy3ON2uK3hzjGMPzk3b
OOu707QfddredqnPXx8opZl/hE270f9BjYk253Ts6QT9sSE2Kb+RDx3O6k9pvmUt
OBBIXVnT1MtR/uKcdM72TNJrY3qKRfRJKXJFeOwwaSh6EmmB3UMyhtqDzSKe5Otz
nkJTPbIdx/WMX4Zkkxm7INyDx4OpVKOAEbsa/N8LLkFt89/Ohp3VsQbPbdIHawMP
5yPynmz02A7MZwC7nWbTYeJsa3rlTCibXdHrUTXR/wPX/VdsttVotaq4DehpvJ0G
YHlHi2vRoTEBsOxtI/g39uHANSiKeCoaSKMeS7UMj6y2+BTurYL8p62+RP+PyTBM
sv59YQ/2tGl10jNgAk9Rom+PhlgvzRKmCWlmOp/ph/qKBk1zx3VlnfcRPBx04L46
Kqyt6J2UCqFhTR7w2aLi0gXuT+5/k3ovY4gtVhvtgz0rsF8jDezbX9s1QFmKfq95
uruF/uFbkl6NmmWO9aze/EOZdeyCnlHt5ar3seux8W9U+2kvKP6+PFwrLArZf+sb
74DfMPGiVt61DIOgqZoPT5ETCiACzjNYzG9H0McSDZmivN0UwNvoM86dqvMNHm6c
vb25yODwdDjgh3qdOTKtxqu243IlBX4r3xqNxR/i9wLW1fcVZbjuSRfQIHXFmMBQ
XwXd14xIhaYOQ9idoMaHIlQavMrsZDCkFpC6C28g7Zfmsq2O/IEjcdBOrygEwFhK
bvCzN+fyAEu98h4EZ8OOTkjdXYB3MXYLZOUZ0J6Wf8vcXSPN8PBp4F50tvUUb0cr
iOOYCTr1aLQcaUDedNTgvdD7QI4piXlttllp/cALwKETC4uOfGLuZoSdLGxSZQuL
e0aG9iH7dwzQnN2Bh1CE+Dy+2OKMQnHEODoaUUJIZdQ3ymZvdpB997A2yNnyYORk
sZXGPk9K1tcHMAKB8OtDnOLKZRiAGgGeZ8WOQHKAH/82nMuv55KkZ5+cPgF9E5CD
Nsv4VF7rsJ5KY6e0pRRomoRCiX7su8+feBfycQ4OI5AZF137hjn/EN6cPwKELuDf
h9y2gnW0KdQufhtDlH3K943tYtbUESXjcECYErjRG3s6rmZ7K/tT1lnaMtflLXDQ
45w+9jqEBHfPx9KuMTfJsPH7Yu9RCNsxrYArxOZ/8Gtf+bpeAiAIWDrkcNzcXyMs
89vHm0VR0ShxTTxdFyKmnziKx0FjwJXpRKMRRel5VJ4Zw4W7Z/hCMUsri//hnhm5
UGDQ86co6oHfub4Wf2sEPEeGM/qurGfdE8Aq8JW6HZ2VEiIFJod1um18L9ZENr5m
7YyD94l7PQPb8ip96f7srP5awiV0kmpm59s5PuXvw6A3JxgHOB/usNICqb//+tS6
Wtcu35NAF9JthMmUZ4alhcZnYhnjSAL7T1YbLL43sRsL9K5fUL24ReLPH80ZSmz4
uTPh4o3RmVKqiOlq8eXb6l/7eejkEsZqWq1J3yVvPgyeWkv5GNfixrMiYlYluTad
ikQbglF1VY/osKgLLhqIk01e/KA1ecl2hOhzi3rCCn0Xp7s/b8UEf6jCGRtpiww/
jk01t+bwPKk2Eeo/UONMMk8lvCL9Z0tjZBE2OTk9lypDINdBj2PzL8T+gLUN7N81
HvKHRNhBoTSyqHm0m/gG70wSmKd1HYEKJ3yJDfPU0WKBnOr30uQ25ccabJXs5QD4
gX0LXy/PW+m8HyrBklQDogSuTOPzRKGQMcD7dXNBGFJoYuxsGYID6kJLAcb03ntJ
gpRv3+X/uHHQZP8uXg6vt5729TQ+34EEuoVBmaGXrq2uOXRbj869OFyVy0y/G8Lc
nWWTdm0pGbS0r2jI38ahF1P9nkyqvpGuP15PHEbpSjSRfoMelHVuof7upnYB24sT
6FySOB7wQIEVDwhMy36DEwvEmRBUqNoolMbWbGzezOvNjjkCQhvUlgo8Z5ornVIO
FgWESBGmLZsK9V8S6fIHAXuGmU9iH0aZUZxdsA6Z0qa5xTl69y9OzJ7Ph1o2eFnV
8nLX9aqVer9bz5290A5Lay8gdx+QJTk5iFF5JDHJwoLV3SS3xDAYBdIJ/x1Lm2t2
3B5M6ZmuL8aapYLLRdBtyMXyiZajlvB5eedGIQ6xHjaaYGOJx8jhCoaCZncMSc+X
Ln38hX72k+lLacb9RzJKZzQfrELsSfetiylaUmmu/zFSwtbrE5Hmn1RZGMBqr84F
BaDsfdcRlGkdRTqEN+kZyn8hZWGedTJiBA3XxfbvtdYOx/53WR9tE1sIyFlELgVI
gBCDUVHv6kLVV44wWyqRbByK92Rec2xraHqxH44yn43jXam7NafeBCoBHiu3kK0g
V3qP+M0uTUQlkmXtFTkLTOc5SycPsTklx3p/zS44ny6O+sfRMUqICy2fwQB7xkCG
cRjK76Y0DgubE2DkPZp5XR7fU7V9/8c/bU3FxGBuKOcRzb/xNXfjBX7MrshEgTd/
g5pFtJue8K+KKAJMN9BgqwKmn9jagdmorpmkDsMIGVV8YqAteUuiRJ9jEBlw1Gpy
JqwDaC3QRAT4+uAcq67dsEuwrvFZJcDNrQ4102Z8VVWCle79vs/weASkBWNjc3qM
Bb4swz2T/X/gxOrKZKxRkE1mtRjR09+Aqzn1OoAXoOMwjme+25977Vl4mF14gybO
xNvG55lLB2zGpXuSXPQ7f40OkjYCkkBwVu5gpVK4D4Cc6KGtrLmx0Fg3+Jv4CS3Q
ZtVA/xwFJ5tLU+l32NU7fkOTb/wWyTfABOXNqWvdeQ0Lxr3n8R7iOLQ4UQT9L4sV
ShsIlrUdsNVKYGkf0SAx+XQaVYNFCElUZNPysGNQUzs5T/FukE9VbjZ1b1stK4k6
vLMkMuUAKgssMqHjd7sfL5ApUBYphj5rAA9pI135JDW79EqfKFKQQhAMHylLMJmY
tQvOp9c1htGvyOJJ8Ao+0aLhss1c3Mu1+RGufbHpA+F9T+OLdXN3tWrB66iYSF7D
S/DjXcuvk1md5lEfXCmCdhECW4v/XHaIqGfkiLOt4OBMu4SE+ID1Eo/AJuAHQLZp
272GUBf6A/IGaNqiQ/oT0MVeX6tkkUlaa9HTMGCe43cqMKfFiLtKUewVaf6UOYSH
Qf1DI74uNbGDActeJ0EePF5XltOu+/B0Y0EmMnBOQaJuKBELT6bakxfx3k1UjvmA
YFv0efeJ2kbaG/juSrFTJIzweX/rJ4hufNo95ynX+AY/cZhYTpFwW07h4UW5kQl9
t+5dvI+00tvtZboZs8EgjAnvUJ8zzUCyuw9UmQL1iDMuA6TvYKFaJRtpFVEWqB0L
LZFOss5Tubi0uATvUbItEUaS1zImLYeomMlR7SxuIVg9kOnTCQ0qk9ck9iGb3a6k
JRhdPL8Q9ixgddWJFu3pPDUrkzLuPZdvlCi0NF8mFjyHnuUKijPRN7zew0baC3s3
EfORiZpZiUTbAr81WblbuJbxWdKSqzjqxYsqPLp3TGHeppyQKmvFV0ms6CevG9Ws
pzrGu/Wcy05as/4T4hkU59OpTBIkEKDkrdl7/YV2jmp1EX7yW3xbIfhKuptbqkwG
UkecAxBtwfYLpHN08wweSR6tjWvr2jDr9Hf+HM93EAzT2AcrqEgF1FRXq9/HMBdr
dRsvJTKxHtB8LDkd6NWAU2lEufuNVyZHkZPw6+QaBs98/Z71mvRrY8KdLX0idXYH
/ZbzaDO66QcS5d8sl9oEaltLSBCrIyPAXT6LkYSHIH+6cfuld8I8NZn2lj5syFsM
LHNdmsJdWxoEu0u5vXJnxV3GuFP475M4xQPPwGcerSOm4GOEF2d57Cj+pMB0rhzB
ypnLomKQYOTEaiHvyrAEvWRGY7FxtBv8Zun+GYaQFXdnduIRGoGzBWCHqOlftJFy
58pmQavvS8TBR70iyr8pMKCFFa+sfSHJ+ZgKWPwO9VY/r0aNzayykZTGb3mX3w7E
wiHo/0VDA5Zc+vBDCo0NYznTWS0AAModyeNQr7YzboBLUCBJnHp3b4gMeTZTpNzV
KstTXCLnRqlnJecU9FiLKGNdvTdlG9I+ROESIqI3u7DHS43874hva3c7fInGXmfD
Bc8IGmvAjASpF6Qreeb9QuvDQECUZ52f4dIJ9EsDQ9iN7lSGskgHLgKbamCGmQ9b
aXgII+iBeM2FSeb9rGNcpiEz0TEb2Rv4xKzJEuMUZFB6v3xZbOmq6/JjkCriYR9g
wfGcPiL6BfVnvysvQ6+qWJYsmk+8rnZeM5H0TGWaltDkQjHhnB37aVTwbadu+HFj
jIWQBA9qy65LWdndeTCuS5BQLCtwQyHdMA7e2iR0PpM9j40gJ7+UZO9nD+M1McYh
jzVUnLUcW5KshPi9t7+OGGd8FgxVaoG3YwxcLvv38ddywXxXPHdppRHWx5fyR/cp
jM5muPH2yaFArmjpGphZGCYHeESodUHR76WSdvxKcgFB6w/nSf9A9DFwFEkT6EhU
od/+IfZFz0ufEB5LUVO2qhldjJSWAvk/hvuopqPuvELpB8d3v8Ve5ZP9w1biFXe3
BPU+oShcxlvots1hmN4T8e8MsOh8L+h4iCuykpK85JddzG/BKGtzS1CV0elYgzSb
DHucIzqxb4uS8kfiFhRoCe9DVPvKEQyz7Dq+JpVOyTrM8GWms8zKJoixlzN2RFPk
gEe/vGl7QA1ZxmfItNMyKpgh3a6TI/65lr0MfIDVHaJMqurLqqojZxtoGkUBvIai
aRQJpoynK4/RfFfb2gzsPnk3P07JSjpaGYHX+c4mNSnzXiktl9cpfd3G1P6p0F5h
wgFeKSCyyYMHu4SXdhYN7EtFX7fiIDoiW32eUwO6NA0q//gsXZnP6Mh8KVmAiZ9x
cwJq0O4gxIaOZ+t3HqnjAamXrke+AHGymuhjQJENNDnQitHD2zZpXIvZsuRbQE6l
grzl2TNiJ80cA1D4xn7V0aYzDQnnkSeQAIrrRhV4ZE+RKSxZ+aHJcZZAgUPT7JUB
ElBAKkBMvvceANi1S9uYL0VyIkQu/eRLBTB6x9/lVL1dgbghJdr0uwyTKSLXO7Ee
0nkiRycrHo1FO1lYJRH6x28/6mZCDGZcZh/NjFbI7j5VxoPBOH6u4xT4J0MfhMyh
Gr6emUVDN1OUMc0lG8uU8KVICGNsAXT1Itp3gsCdfvIKC/DtCfrYzEsdBuUNAeUQ
B1pJmhGR10wu0vEWbg2OikKbyNqu26MLKR9ilEsRuGl/Pp9sOxMEHhTwPMxHTRk8
G9BbbmfD4dN5DaKsvTxLxZRkxMPfDWJ4A/fCs9+PRm3ev+DsFWRYudJFvjPgtiHL
Q1xYBu8pbNPJUbW5VeQYH75inlQ1AnrV+pTkyJK7y8cXBnxErBR3oN4BRbkjrrQi
hth5DNOtrZKciWcyjUfPptyo6+EHU4QIL5EtJBmdEYPi3RvUCW8jMPXo+AIug8G0
6e6bzGW6Bqt8PwiwZ4u4tkfaYeWXBEQAHeiXh/KR0KtMg53Of2S3OazJDwpVsCxq
LF8cv/CmlRq1x1ldMG0vPIqw23wyyrP8ohv5JKtcsma2ILH433GjilMO3u26t7r5
ZaqHDMNlaXaBGCybVKwEtMHOxfpbXctTIs5n/e6ixdiDeGad1CBj7XWmoJOYH9/j
6tZ/F07HxfGxM6R7elcTrnvv6FV7eCLvHSJOujufrqx+E0Ymn2k38k01U5Ajgzhv
C4nuAGbpqoik/Xnxd8Y8+7m9SEziBwZbnkqBoF+wD5g6gJCOiJoGOPwsWv6VRulr
ptj2VVbUkB2bZ1c6Ge5/dy2YEW2w7FNkxFXdveP6yHpBLDJzVwsbMbRLROkwxMFS
LF2PwLZKJWmF+GPX+PUM9ZVcH2JM6QHqwaxrkkH8SfHnIEz+X/8df4HAqBUT4Rd2
sqTg+u+UPtX5ErKmhs9Q0BskCYD2JtwJyFRENc6rixEFCxTQld+Tpjp4dW+qMrc+
QGZBEN334IPg3ZB6696gd0o80I5PcDE8VaRFa6H77e95QSd+wZQYNOF2wOlqUCN/
d8QLTvTYlSsdgc09P9Lk6/nXKPMQcfoXv3ZSi849yIN/8kZrNkXkS9xYuRmAGZKg
v39ke7yqSH8/4Bbhibvlafi4lB/l8Ms4LN4IVPO3pqUDh54gcLRwM6i05QDIf1IJ
kqD/heLxfpmOXESFFzteIqx0T4zPHEDI+S4O5OeljXdt3PsNYqjq1wTVxL707bSN
q7NBAxHhMe8njwByFR4mLQr7i6dzvdnGUC+dY4FZPLVkP86TthPUNItTgyt21QEQ
BD1E5vtgzm8gZO1Ho9oPB4v9cx2chC2hF2p4md3hrFmfLw6rf/lPjrZf1+xynNRh
KLRBEUR5MOiQtz38SuOu3/w1ifX9NoypRF4quFFfu5ONpkn2EFe0qrA1tI3z6HoC
1jZngLI13Zz9lHMxljLmPi1wtB6bv19eVCIbxHUe53ig3BQpL22RyEhJ638yQ624
VLnNEeCsVfq6cKC77e/kqPHh/rRGe65w+SvSsyVZ82tQTUhBswXMSsbRaRx0fzzv
m6wvQorwHaVFgIK4SKYvMzXunpyPK5w+fsC8mW+zSEwV+yBwx7rAnrXz1OdXs81I
NFiWrWf86/vjf1cCbboSDS8b8E2NZroN05tezLGbAd5oFuGCVM88Ha0kCNZdhXLJ
jYciw0Bd06Qa4h/YMG/1nnRgRQo0m7C1Yje4V+UCaiw8oh5gDnE3pFWolCnMK9VH
0ORHCWgaifTo9S2deKLK14K9mz1lmqyM/tT5vLR0gwc+dsde99oGKVHqp7lK9yjg
5/EIozvLs1JQdOq6c8tqdoKQ3D4JhYI6QeCEtK2D+poWoEW5GDAULFzf7XRRUscf
3OaEZ2KMLBrjS2XrwQ2eV79b0q0sHKYdQW8hQ8ZhHi+UHZmbQuw88PudfW++Ws3n
eMKWSHV28X1BUD5Dv4Cs2jd7eG7hntVrkSZn73rK1ll+zmlUexZFUJM/P6Ais+j6
NVSmQvrNIhg+LMiFE2TYCISCnPyByKykhvO43CYbNniiKXd0x6mX3RJq3ouagxjQ
XS7xU8nIktKkcQgSomBRNQKGl1rQA9A6MS8FjkedvYme2ajAAqoB3lwiqK3ysrJe
TSi6IvLS6gLl1fOaetYxlsaI4MC5q1Er2OX1rc8VbZlhvQts+pf71+pTVRATGfEP
QUmQp3sT9rumMJ4WVSNpg992Sx3u2DpxhUWDQ/0YEUh9tUURTNFFBh58FOozEL5R
0bnllKkEdxaqhIu1QOYJd0XsZeCeTbOXDJis6CEbJyX9ZqL525JIkuBG+KFEDIKR
S8tZiI1Zcl2SsGVo3PqUgrTlX/kvJYOpLDa86VTQYHngG5ctdNXJOigQgE3aHUsg
cxIp6NUWlQ72is+al+B4yTnfds4hjq2BPv0yJYYPill+k2O3KqDNSehJQFHnEZZ7
JuN/Cz8P9IKObqS9St50q4GuiGYxzG3pYuXGkXlqqfCvWF+8DbEBIXROZJfdFPnw
vX+JSif9ZT5th+7OJOAVY5nT+GL55iVcpVTjMMzHARTpd1W5EcKC/ad/q6kjtZ1M
gky2zo9fRsMERgSnZPk1xyWrKnVm5ZDKzYOc1lnzmU+CFwMBSW0P4T1RKTQjD0v2
b3Ngfq5zJDkd3IrODpbq/JoMfMkjCrxwJsy7Ld+lMM12jMfQ7bo0wF9AoHz4hpsF
XL89ZKXwOUxTjsWr/rKFtScFwWCD825TMxGnn/Y71R+hTGQSzrQOlnEYMEuppWPP
lAjJYx9s/F28xKmVqMbBgg3fTb68m129q69wMpW8FvyKQX1v190rrdRpmA/ldgmu
Nhe4oG2OfCJfIZJ2bTYRViXmLYjJRh1hCPiccP1zgUGtuK1vLKYIWqN70tOpn7vG
jNQbblqkzcxvpUQUbworBMDpedutirmqksnMM7iI1VA+TlBA73U10ciT4Q+pbQxo
GVY8z8LcmWpV2E4wc4xFDmmMmfqzMKs2PYdg6F2FIeGAh8I5Q88DX3/QX8Z7i4tU
y6ynBbArMUBP4SiwBjfunMIzq71hlh3/URQkGRmIfjxkAqdS2FssaJNTr1YF1Pvc
QW/8NUE7wWQqvayerU1AYglnjNNt/UXzXYro6p4m0nfwEZh0jWNYnE4H/QThed0y
zQ6M9z1hN3PlrCh3qUWlcb1wpvToMPfedSS/OMkeBf7fgHhm/Ju+n8iT/K4tktK6
vIUpvxhZd2kcTvVIZR9DkBDsmGupsIdfxInqn53cz9B8lDW28edsr9NkWgxqWtQH
hZrJmDiUPPr4IQvve3Ge+tj3aL7X3eHK3Yv1PyRPllq19D3czYHdGQkdtp+uzpYK
wtShyK93fQcKW99X8lIgtwtccIeD4Ga7DGR/XRXfCwAW5cQkqkkGKvY92cyis4Bs
GgTKj9VlMiug/layGSCUK7fmaGqWUgE4IkVrbUhE4986bb6NEoyyeysYn4D618sW
9+G/BgeZNRAX+KkgB3L8RNL22FaYAyKWPAs+JUAlGqIi31rGQikkNMjkN3R6dHbl
8NrMYRxRgP0yxTuqfQqqbHRwRnOb42kvwFMOG7nLhcW9E5kQcLNYXeCqpH6gBMgs
uEFl0Ut7JyPiW77wsdAd09uj4ZPXStl1/hVUlkaBchuE3Nf/j43rQjIs7AmwW1Em
MC4bO9VJhUC8QAMMuYQ67r4p+RDSaK0f4LfWllKrEQdW2eBETJMKBHOhWOOSM+vd
ZXboexcE/YsaYY0xV6Q25an/H6jOIa8OE75MB6Lj1Sk0lVM2lup0MJ0NtBFc5mN3
cQTrz2b882MTt+meL7peys8iNGwPf1OUr1GbKMq428+I4Qku3ww/Bb/U5iI83qFV
VZIK5siCPox3UozJKQFPHeJ4QBiDgC0hzPGq14JoPDkruyuAZiEVtEl8l5K0BJVS
kcDEl/cUVybe5QmkvMBdTdEOiB2b6IGIodstU1QMT/NXySm97EoFMVyDrNJqARRq
7aYs0ayS/Wvgo5XNMA3Dbe9CrQa1yV8tXvURtRFz1l02qE85TOcPaTDzEcDYv7lj
7nfDWyvCl+wc9kHwIGuSKbXeyZ2q4Xp5Roseb2Glg1GnNS8qYtBIih+7tHNkLMkJ
HtUB2iNz4zF1O9KhGKJg1fKTsUhqL5MkzJEPfXLEfeJeh/r6Xc+9p6DEobMT0b4h
g6ks+u10lKAJ3MYGzfblroOxrDS23ulTNPjKkq/KlLyETAxh9Drd2SEJM+GBjLai
m1dw0s1ZXcWFghM7T05DAm2zEPcf2bJeI5YYHgiDQjlrqmkLPH4VQvxIO3cs9PbR
1c6SKqUQz3p8VpKzW0tmJhi1CQfiXQGztxT6nXG9wcHTfnqIppLt8EJg2duRNWqn
dHjchbJUnC6OiljghpmVrfJCn5Cgj0R+xVfIFwu9jBfAfZF7hLSMgbkQ4qf7PYv1
ao+PqsA092z7W39mSSKLYfaof8f6ZchpHLtrXDBuN/MB8k73GywK434jmwgg6Q9K
BrJ6Y5Jb3HZhWpGRltcSs+OeLCcSWfWGwFZSsiin5hFULMO9g7wXh1JXjMKVlWJr
AWwy2X8d8VNAmGcGaEd3WuCqicHn9Gpe7VTD2XufSDrjWlQk0rX++MYgA09Kk82p
+BGEXdrPm9wI17621WJhTi+eM4ET0/raBxVXjsj9+RJcvTud6kka1ufclzh93Qyy
+1W2FBu8iMczUY11jbK/aTt01wX/NO023RdUh3/R+MQT55fwWwoLgfpIDmrNIYON
BOmodJFIYbddBdUpJjK1YDabBNwva9IruLv/p07bLmENcFngBbWA+h6kgP+STzJk
An5V7vvfh30CxmCeVQaq8LcSKKEUfvYVDrpt35TF7Z7lTFIXcYEK2LHCA88SRGFR
uLQxCvBUIydf2Wkkn8vuUYHd8Boq/2Z6KiBguqOPShqKJ7QTYbHzk4aIwJmiaZGW
fQRF8V+fIDxeiy9cN+UaMpr6DMguDjwxF2X87GH1C/rk6D7F9oB2XF6PySVbn+4J
vWzXPPTFgD8WEIShRqn466h1PknvCHgFKoOuV5DWymrPmG3KE7vbY5Gbc+Qv+AJb
bLEUHmbp4ZZcBpRzJ6Vhe6Tx3ktSU9+hXt3ToTIItFbe3NEgqXMHJbuQ/KACpkt0
Pp2ezmULh2xz6eaAeIFTuhu0tOKY36qLhVwtCRaF65uNnF7oteoRCUnouYeVqB9U
tgyOYMlQc3I98hDFZx1znvBPaocKYP5uddDza7htPXli0Tj2a4IcM7FBdXddVHd3
uBSMmgcPq6/snoN8Axb9AGrfp0vFZ/gpIftJ+bBrsCWhL7+r1bVRxpXbT0gA4/7D
/B6WKYu25MRU1Q3tnSluQXr7vdlumj+agXYqUmNTfV3p4k3+4+kBTb/PR+y/1ZCu
5yXLGpkdG+hZWseY6bODJb/bFf9rUoQ5JxJNWDX2TheBuZGDeiktybKeQD/SeEZw
YjZ5ZaxwNt9HvgjX0V9msySuRNS3+v6d/SXfr7i8/re7iuncTZuI0ovUDky3uCY0
TEowXxRsCLgwXSlNGGavhPnsztRh5YcvmZKwLPHaKk2nOrxtQ07KtLryKZPsMcYL
813XY8syIlr5TUeE8g2gUR0/IY/KARKDLUcDPpa2NhqxQVgjPJ24F7dgLrzspoBK
YaD6qqxn/PFFz2zVEHys5fIfEEYRClNUM0bv9H8pWRcwJG7RROh3bJiMR+FOf4Hr
FunysS5R/GPLYzGuj59x9uovM9b59plwDqH1c8GNcxNuYTPy+3uacnUWGkGHA7mk
iVxOZ77alLig2BE8Q3HnR/OQFfYZr+J51DaVE/U+2siL1pPbba1IQDFuKxPOxlyf
0xx/MYYtiqJxE7HaW6SUgPA5ckhxTPG0ArD1A3v+/J75lp+Vr5YmGR5Ec1BRKsX3
AvXSaCCk5QdUHLXqKULIQB0Sqcu+YrUcwJEdpiRo8YdQGpvdEJWfqx8t/vTHydQB
rAVrMKrcElKJ0o1UgLCZN9goCW1SkbWPH+Op/vwOZQsalpVeiKomBFGxd8HyU6Xb
EyQRn2t2Y8QEa7irJ96bHM4URhGEGRJyvlkVq2kr/R884FruiTiS1EJ5faGeHE9C
FRaZJBB9Gm0ucj59tn4JS0uiRgwt0cf1mGadq/tnLQEmhnihFWcn1Zl1dnQjzsCr
dn16cOP2Wy3Aagwt6tHS3XTOOPJ37Wa5wo6SnR2GV5PHAbStDz29S44qASiJ1gqn
KfKQCD1bfm4lwdjaPxUl0m7iySiEfSPZBZzVe+io/bpxfSP117nR3uTP51cPPJ6b
xbZ8c52/OLKZKuQsj5720bv9+z+JrN30W1ZXs5LZuy1OsQKUSaRP+mZQOQoySylx
OP3OAZyQHyN/sAJvxH5KPuNJaWksDRsFky1z1ceC1hXFWB8o5XVza6THfBYhfYqB
wPukwwPsNOri6OTFsXfUlMGQPxqaUPF6Uj7L2eMFCVj9TtY1oH5EkyCd0guGNMTs
UC1f4BOqk/OQGmQhhyTX9vOBpa58XC3xga+rd0M5Y+VXuj1mu/Qpy76qgcpgpfeo
rKGJXqZYDO0RIaqeH/jmGTZ4ZPINL39aJ+rxGb2/moQMDa/C8eOpK3KX/WtX5rEV
Uhp9hOsjEfnb1E8ScLVg03j83AJGLUbByO3TzjH11IGI+QcZ1ZauTYsAUyKOgd9X
bdSRULugRT1YUiVB/z28pkC5Jm6R8kdSHnFIe2xmMccaKZedWoOSl6dR6spudBmz
pSrhEnY4UzGcrISVxw3oyrzwHO7aqukY46WE6sbdCuiAObp6LsEprR+Un+96h197
W+DIbjZNqtw3HauO03fIAbEXI3uXI/TZORzpDuc072Ah4BVR5EIQxPC3hT3x271t
24RqtZtdbRah2nDVgdpIUdtM7i4v/hz7o/GE9eZPoOuoImSRHimd3e7FHTDQII8K
+AXRoA8KbY/iXe6WaUxTv0GKWRTd/wSjhrJ/ulanFcSos+5G/yvz1+knm7jHfDo3
1Smf9NNTniKtS2NBDhkRCeJThYqHg3p5uCPKgkvxbrbAXlS87uE9iwwASiBtl4+n
T99pjv+tyspr6+yPi0NEXJ1svbr7y4SmRanA0D13hpnkh/H6csOU4m+z1yBVo11Y
FOMwDMOScsYRIt3tueYOcES/Rhnm4prG/xUp3VM0FGYe5VwhQcivAsopmNj9/v7j
t7FWEv4ms0C4PLtL2nmEv/VLWDsQje0ZHW9kvnWaRqH9AbXVJcI1RZy9XhA8MS71
ZKJ8Yq022j4QjVvfMS8VlXNEDThOhJfHnBOfKSwyEcf4JczbaK2TCgvRru62OfM/
pk97rzripj3cRwodZT4F/pVTxRlcknXXp1QEpEt7RS3qcOADG9lQCbzMMzYSato5
lhsLaudbHXcXGxbw7M5qGdGD8F5RV2rUhE45ka7Ma53tx6+W8Z+av545fnH4tv1N
WUJLnD/TGCDiZ6iyi1DCIV+zNZ8RadwoyfJwWIPfx/j9/Rk8Rj9Jtt/GqMMXuf7D
ZKhatCNjdYDQrOEhEbkvjpeY5YLG1E9ADRBbfEMWwUGag/053vlI7UAia/Dvo3z1
GDWA2IM7Z5sGp0QGJVaXnytmQsFna5WSmfIaBAskcgjEAKNmfw8NBosY8uMoMoGN
/NZK4sJI864vRA7iGsqS18+W+VfbpvoPLrVF2pqNuuSfnqs+JDpLqCmYGq9J/Lsm
V9cLqEnCCZXJ4PZ/kopomRbX2oSYoWEgtCjHA5lemIflO8lraZaXN4tnMJYwNFcd
ZbMR2/+rSHtNf48Koq3skHnI4JCo9H7TyGeMOp+WTQWM3fqH3nEk0ZU4yI8ewq5V
GxkFVAZxivvp/N4rUbpqIrb8F1x7lEDpFttv34QBaNt3mJnb6lfOzsTnSDiN3CqG
IjjDZsGRGFUS1Y9Io6xyp+yXtELmdSA7sh9eEgq2ZAKe63fYHhUHRBiMTYX8r0EE
tj4lWFbIewAutuR2PcvcE8PFI4TsaWnV9/9RIpTum7s+MW7i7in0SVnDNX/kSO5U
Sq1Hk9QfvZEtK0kEMD1eATu4L9E6jILTe1nYWb2qQxCmztDLL4PihSbQoqdmsFrd
DSITH4EX6pfQeXzSB0XPDgCPItHOWjZ62/bOBvHROLKaLOIbXRLw+uOnzxbIy3M7
i1DjdGPD57sPS1zgCNWSgqKwshsloBFoTbk2hcvZb8Vv6HSN5RoMF2cFX16R3oAv
5aGAGym3seDn+RqAJZ3TPAjFxisDT/I8AtSEt7fPxtxDsQ6whgCSa/xFFNDBxzqz
ob8bjPdl5ihERQRcXVjKp8YwFXpzq9MGnA2b7iQ1d/IViD/LH/J2FY7WV9ddccmQ
26OC9349CVAKBY5LRGOqUoGDcxsoom8hAEnEn7bhlpTaLPZpSiZjVJA8EUty8hkq
AuURiEKmutaw9AtEmBW1DtF2AZqSXiM/lu4VF8TY/8uaqnceazB6DA6DJ+yX6YCo
uQqDFbkqyYOQrjXDE7TJJ4MP2Ll070kmLg0KRmJiVfmnCnL6qFeFATC+N+SaO3x2
rN08l0MhWWX/6Vl53PVD5M9Fq/tHjtPo+7h3w/0e+2I2DZqC0YT9CNwU55fdx7GU
8VV3f/RdqrDpOXD4i7p+H5qTO+c63o3Y9u0k4mXot16LtfK+eKAeMG6MIM1PvXrW
+cwmTF77bRhIC4NsqZszq2jL0EEjvEDBQflCjhOuwM8xQ/IxYK9SBrZFLRRd1Wi8
3nBEHR4N/R5oK26ej3+ikxHjz/3ChpQvwWzmy+jfWy6ztzlxtJSubl3JLlKPYxTB
hnzGza7GXwMoFv+bZnGXC324VCIEjLeii7Pl8bK/1W6AA0vCzFFW9o1eISpTpBKq
8gavpInsUy/eNPI5ZebgXeDJR4Zl5iL/my1pcBL+p3ljwufkF9iIGcIEZ4BVsvhw
0t9RmvcI8LQ7Iv0tE34yvqMjqyoAOzjRuBtPrBQB0MQr7nrK9halLW/OAt5fCCXf
dRfspxydcRMOJvw1EM0pxN2rHFgMt7BsaZPIlvnMjpd5kUjxKBYgJpFtBq6GEA8D
VpumDDUEECt9pfE26xQHsmBal8KMtda6GYlYFmyHAljPt0GC6z8LHaUYLfaTnSSr
YSY1rAhxqJsGsH+6nZHpDcf7IrlEAKOwZgVoO0ahsr8l/2v1ihvyznumO6vGvj43
V9N789WiXjK5MQ6JM3eRE4v8OJSTDZ1GA4gXoSZWsgo2dlV0kO9S7F0Oi4mr9x2a
Uqv3g1YlGapLvsMsMkDQ/nCAd+w4Kdlny+0IqgTyeS0USzK4ICSZIVa8uklAmLFv
LZdzs+f8TTRGHkzs7zjljxuC5uc/puH+wuX4mTlj1MgfYa2Tj+y/rOJo5T1nlUlg
LQ4z/q6KtDjTrddn6uIYQ2CKueYR/a8n44znu0yZZY6+XLyaWQvWdiD0pPGTcRjl
vFjmE/nRkuCnjwJJ47CpjOsX3h85ubZHXX6E89jTD+op4l7fo7EL7FREX4+orJxO
ARfhM0rvPdfKzVQfZwlNkFXbKHBHOpBCXfXTClVKD//DrBOlO2IAKiiYtenrhpgO
sHb7StGrpwH19SVesxsdoPYHeSi3Y+kJ1bCgcIxCsoyyGnCJe8DTAuaPIu0+Uj8E
0uHWE2wCO2zJR/+in8+HvG/RczpHwUWpPWLuVHC+6nfcQKqzEWmtbt8vVKjrj5R6
ka/ZAtIv803+QenT2p6X/Jg+49jcEWqVtZ21jcArIz3dw3fbfisUdVTY1ELnbNvL
OHbox9+espyQFPnLKKpBWllGc/JtdQuG2FkvoDHpu9huoDdNgvoURindOP3+J9sI
QCTIfWF2XPhnusIBotdJP4Jqn0gLVsz1R8CWvWx1GaCtb9Hjg2YYoio05b7KmOkJ
qlXsN4cmjqzPTRiuH2lKoQ2tX0TMhiaeoLYTfDfx+VjAwf2J952LP2/1+hE7b908
Xfdzn53IpBGHW2t+9pb7BKFFp+F/bO83deG+7MLT/ez3bKsSiUdRKhBCLjbZxPuy
LcZdCbqov4/2moOVenpzZVAraIxkBhnxRj+nydzndR2F64Odapu7Qx/Z6kwWxOI9
09o0WFoBfBTFwy5hs7OfEzeiX90Sqs2z3pz1d2xdqRBL5DIUSIweaa2YWDVgfM9U
a78fl5BgjJ5193Arx1+doGCi/fhxW3ATiPe6QLOPFhkBV6LxsNX+rxba+rpXgkDk
nJILuLL0PPL7EraZ3gE2g7d24irIs97aYLHgdH1n6hHZfYF/YC1auTKkVoTC0kSG
qBpP7IneCwdsPJ3uCsW/LnK0BngLhTfRlJLKMc99guqG5jv+4RLVwLr6a6vTsnuX
+1tuKlg4D5nSt824hgR0R7AWU4CPUaI0cWHsZgvfoj8UecoWfK3zKEygvIwmnG5s
zmpnbAPzANOhaf4qkEnt4GQbaXvK4HWQnFu9EMYSgE8BZUAZkTB4LxDBBKyeJqkO
y6Mwx/wJxB0EJaWFT8MSxB3hK8T71Zq0b4rEJzpjNw1f8o3sOJU2s6vt7nJZ1psz
f9wgvx2BVnySaBFZXBadEMpsFJr6mfUOEK3lFmH0iMGAqposZWqgzVaBf6LeRzpB
GxdQSL+ITWfMdLAU4MbZMuLb9Se3Sji9xA07vYfeKERZCXwHe5iFKwd3kOCMveBF
Ire+BwQq9m+N9G4f5vzRc9q6u+R5uD9NG/KbGuX+XRky/kzLdKR2BshWoa0Vrcoq
WVuXibSmR8SkkwzDlr8Rk2jqdEaHqePSknYxAJvKG1s8sO/IAutnWsAuorQNbNs2
17MEDrypGYRJxlLv/lUL3y488TVViHpl83l5OU1KC1zmgog8SmENRZEVlmVyELVE
8VcuPBsnjKeuUOPL6MwkndTDLipFdt+jCgzL9WQOVKYcjH61GX9ziok7IX+vTUEU
Mfgxuq3z3m5l0SyqK1Bf2ZsMjZU0+8CtM5ZM6VWg5oxHVjf/KAgojnDyjRHPb5PU
/tdfc2ig5mgNzv1bBtarznnrq6QWoA7MinokdJfRNRSFbAPP0kPjKU5VefIsw5Fh
zkzP52VV1U7PIET+McnyIc3hsc3yNWpAfFdTBB/M/J5t5RbmtRqF2/TVIXU/VKWV
7TnUjENZqISh/nXyvyk6lVcON4eDrCxvBS7cH93bpTYZQnB1BeXmpFuuQ7iZVFm1
FXJewg27sx6v5JgJT4sbK+O3bclGORDU2dZwEmP+70/mmpgQsAE7X5l1D2nQvBqx
242a/RLPSd8erqUn9eYTodmnR132JMyMVAHkZXrp22v7pZxwXQdRsl5qdg1Ho3z9
t59nR8WZ2awsuyMJZ4CW8UsPrul8z/PX7h6AnefGXOHnOD8ueQgTCapNDJy9i4Mt
vN3H8zFg264piZZ+anwBlYXCa87ccrHX6qcZjHwC+elBlvdqjqifRyzH+0oS5OSU
pOIhc4mZaYOfEyAZlbQC+xglOaruiUr1sKOwsBtkjIox/1fYtDfKYHHvCXIUkU5O
vCpppcy5ONPpw+ujLB9YgiGAZtH+Ls9ml19mPyXnH3Gz14DUP3fkf1o5qNGU0tQ9
fMCDOOdFz6FyqUG24/YrBDGf+fC7kn0pazqdlYhhNw90YT7Gx9jUQYKD/gN9YtgZ
Un5QuEtl1pwSztqWXEeT1qnecx5eH433Eypcm4T1r3W+aqI2YVeN6w1N59oLkP7g
58RF6vOp9ZlXZslWVC6Ukm9dyMKLtkuvZ9xYg2E/1ghyp40+nWH5XcUrQegDtkaJ
XMgzcO3GEcoGvJ6jCeVf4MF/u0xxXTtGizHzGhAvbTvPijc8jPmayB9/xo6qm5hD
ut22swpR0VXBr7xUefEDNgX721cLAXzJHQNnmO0tFJhY6w6fz8OA94qTktwn2juG
/Yi8W80s2rjLYZ8vK2hZNYW9jBap3dQgqyubQ5aWkkm4NF3QMd150wrkOpe5kl+Q
H5qNBHvMgmB4FneLaEve4rVXI2nw9/ZK+goGZu89+UY7uKjZIHB5fpArehvzzHPL
kZHyXAKOrfCAM4ay2vIrn3M9Ex6RwYbDB9DiEvMcfe+dyJsbJXkMqqG9vxeRis4V
k1G715vA6OaQ5uwv6UhYcujV6eSVJFcxJuIl3ic7bQRH8PKZ+NE11GaKR6YbZ7Fh
3gJAPd0VUUJedI2Jniym/1G4QkdNWQEmbHw2XkRQ+0xsskA2jNLL11vGVy1Qu1/b
UICOtXkiUE6dUo7rC2O7ww==
`protect END_PROTECTED