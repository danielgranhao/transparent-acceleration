-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TywCOYfSDCUnyKB8B3UtN3ycuFXnEyGe2y/gJh/LuOF0u9P62SIC8C4WY4Tyhcptchtr9k2Iqikc
0k8C+YGNzHp3VJLXVujeFUSuenkaBfr37gQaCSG94n0FgAWuhnSil0JNHAerhi6tW3hRVY6fZtJB
tkc24v4GVo/RbfEnVhYRNzyfy1ExFSzBhbdV5YljQdc+h1IyMn84/hhxpYuAYh2xLwwOvGWhskmq
O39z0SkYU9lkGZsfkhLBV3pFLmoQxui2Oidb4r6nFPr+YygCyyzbOi5rhpvgTPwETLGNpNz+qY60
i7u70VfJdceRNLUJztq7Rr3Hm9O+D08hdOjbeg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 19728)
`protect data_block
qdZkopsn3rIKN8i8mBHJSrA6+TOHDlY4lIBFxXrd2A8XmdWn5sqHt/wP3v8tgOu64bX4eqPvyY7x
Z9gwa2p7sRZkx2Ov7Zo+x5jxe+3wY9S1gw7mHVTORsGstSdFzxgOmNCe5brDHXU4ywCeBrK+9fTy
6fyvtxOOwqNMIe+WEDXc0j9tbUJDvhZvybKSMh+aFTo50jJuIWAUBdV1/XDOD/UyWHbICw0Rn+Tu
hwCOd8ViU7djTdgQtdI8tWHpcHghHj9TghO1NFRc18plfoHt1ov8SJDAoop4ZsLoe+BjXbGbZUkK
19GZPvR8AcAineETZke3slH701T3WWjLsowh/e7xVESIIWrl3imOs1v6HqfvQtNUkQ2wFYxeOqIZ
skt+qrfQYRaMwgmdx/GONobDW+fXd7EBQ2YbC3bDaHU4LAt0hjlxwscYbMMqogHX64scAc+CDsXb
xRerpww2EvOkcyo5GycIcCFuWnQa2N1Pg+QOhxMkLC8RDd77F8rcTECTv5LfRycwWX6+twdFt11b
lhZBFDmiPjyOHtTACD0dDIjIgX7rYNPKbHh7egBy1YwbJPaZv8n7i7KhYykxzu9AzxYT1oU5urOH
JKMGhMwPGv6V8UF0F+RZPb/Z2hKdkygv1F99cOnTXId346K3eBt2815y1qmhSeyJ6P4Un1YPiG2m
UdZAaKDD/JQjKGY8MmIT5wM/9LH1EZhJFHNV8EG432thleUFv8Ca6tbOE43bWFuEPKQmwmFqIf1Z
2yFdrZYTrTeNaN7SLvyfO2s+RGj4cfmmkmU0sntvDDtkciNiYT35E2qYVL624/dBihHS8NrLf2lM
hM4vJt6MBVRBap2bARYHRun0pzJrcXVxMTlsOgJJxFr7gzZDF5tWHTokW0jJ19xn8Div8O5ZCrsq
fP6OV2uOfLDBmds0wJsPjhFcF9PFPxc/ThahKBNam3OPEAh2nUElPGvkuvq5Ods+1qavwFNQRXk2
1LHfu/i/uXSkAXkdrMOUtNWZg0JVxgAHJPtBKu0XfaCw5Y2z90dFjw+UxQ4Yhlz5O21Uq+eXS7kJ
hgW6G+5BVqG6mKd3YJ8nxpjjX68KASUgUIn+81d7CPFVkdBiTK6+X7qxw6IXhi+RAIec8evc0eX7
q60pKohADyqY1HdbqSvh7MzDY9U69RywgTD03DWD7LEblsPN2l/xgiPPuJJa19YSrg9yMCUo/eTb
B6BRXkiYeRH7/gTkotQx5nQ5llWjVEq4KvinM46MxEW4oZ0dTyc7ikU8glMG3KghaYqi807IsewB
KY7WX88QAmNwmRBeFKbG8pnsI7rZ/PgzIQySvrUy1lVI1X/+wDH8lB3As0uJdoDYojy66ohG3jEY
hfy4fXxr47scWkePIQLtEkJVR/Ff03OQLBYxdqnJpqeHS2MqSAH5qp/KihmRGcMWbGvN2LeIagbt
4euVLrkTkci329DWpw9IBvmD9+ifmK6GTOiAKXmKi4+aY0kTmv+2y5eOG7RbpcXGs8bMtL4SbNqL
xv731cI4K2sw2no+4Ze+7f+708uqQjI0V2iLplrGy4RXoyKxhOJQ3zNrSGoEidxAqzr9mf/DLO2D
DYo5M3GrrU1i04V/NnIx/dvWtd5s3jAFW/1rmqCmP2aqLxBuh0xSk9mi8AlJv8ABF6UX6gr/RyuT
fOFZCL+x47lqpfVnW9i7vWCgsx414IT2LaFdA0EE/44rr0S9povQE/qMDz4+wamzSGus23OKCvLc
C2Dj28rp1V+N8l1+HF6QF3m9aeJK/hkhTRxXAbrq2Wd+Oy0HngnvAAsBvAGvNEAM9zOn5/iHYk0V
s0WMqCeiZJs53+lEMB9WpT3EcrgKZYWCskL4dWxHYsxZHUrE/zSM7ydXmWXvUDMSx8R2SsX09Piv
JTYcKyh7uIrpAK6/0x8BAjSe1XxtZP+PlE0fVAhd6EkxfzPUF6Q8Y/llTWxiJlAfZxiMzC2wCuzq
NI8gh2EuO0BHwNigPYnVQppIMFNzI3nJ0AvCSqrb9fZUlmL9MDZv5Raps2qxj+jDQfaekYqguz7j
H6L2hzZidGxYQKHtaTldX3npWKI5qpXJACl19rnmjQNH2FfoM1DWdRO7hm0dq7X2eF5o7mzPlWwn
gkNr9yXF9iJ/5bo/2/e6FKbxvsKUJDC63qRE28MSgFmQlDYWuUWcWuCtKuQ2sKhmf4lyr8d+3D7u
NrdU4J2UK4cj7stuALtfn6mVOYFewq5TKjlEgVzgD++R/6jhLJQAUvTJFBtYdWcEAI8wkGIzZYdN
tgqDwILgIlcksRIofrAeVtXUjEcJAOh9OqsabwH0dmVv11VorxvAGNCyIWn9ThzF0QhJ+KFv5rNX
sC5B9UGM0AAKpn6Y74BQCKg7cntKY/Im2oe1s18lqRxLJW7yuZ7cX9By+hJxQJHPspJss1pWNxNI
YVPeaXLSUpTS/c6deihmyv7VaZWPO6iacihCQzLE592uRIyE0M8T4Vzxxsxq2RZxuEsPJqdR60N3
IMHyvqP1RyM1bhAbVQNaH5cSWrCG/kU9r+DDi0VpFbil5Z6krflqGkThhuEpbnZiNq/Jopif4ESj
5SthHEHaRn1lc1tioW/dzRa9FEI8bgy543OT0+RBR4WDyOskNdw/tQMavuJ+RCGZnr3hYYDlTM2f
ySlElBnjalSwYAiL5RKaLjLsMiILSgJikMRDEZxouID8v906++cWnaXxLAFSc1Kru+hynr24soNn
SBgJDTOsjyh+gjBmQr/OSwLq5qJM32P26xsX5z5xlZIqulad3fXzhvyysOyIhVDpRPyYztjuLb8B
+hZo+J4SdAoWTaXEwzioK7Wgb2FM3Nw0wQPWx0ZVNtn47nN3v2L2n1ZdgmQxay+LYZCxE/Nn0viP
e6Yv2ykzepIYn+fP6HvElAOD9CdT4YQ/Cj3DjkD8wedM5AwIiLMN2htuYj1BtiYRN/OpYB4clXtQ
mCMrnudYN95/Ix8hPKZx4JAyGgNA+7X8Y+xNpED4wLZDJD3YU7N4GQaaELXru6v59Mvtuspnetba
onaB5zbJX54AIDDu6LePdpfkZg8e9TRzrgz7cSgxohow2GoZpRXDLoJSrWpFDIf/ea7PPcUPjufa
TvXYjO8ZI6rX07/WnOAPJsmJdDknUJk/0QKJASuR2k8tyAQeroSXxKmoKZj2xROxkZuo1+ijq2WV
HnPhoXsScD/BIjGNQ8dv7CuXvkY6kN/waisAYNsVyIGNZxvh3WjRDAfPgegfwdMQMSROjGh4FZAc
iPbcJmEhvjogXdRnaIUV9BfPFW8WqcWMMzdWQxu/MXecFoNPqO4EZWCmyZte3nEQxdJteYosqtz6
5hp5jVQbVj70RMnH8tHaQuvPdLkExjxCj0PTiqZSWm1fOoOe4/M9NNw28VgpuzWKdqPyEcnDGOhB
KwdNTszfKXDzdLuXLbZcOeae6IuXeMWnEtZoV4wtCmAq4s667H1pdPPo8S6Vo1qTATF0RHwFuDdn
GwzVNFuU1a9ImC0MJUcbhQM757GMMRp6odhUY0jOIUV6P6+S21OQqUpqf57r1RHCYCIuByhV6SNq
Pr/nkpUEBD9+lc0mt2kORJqDvMGsCRg2z3pmypBFVpe2d0Gc9w0cSNsAs5Kcnq8ko8Shrvnrw8st
JsgKo4T4nf4D/1YEtKNslPwTTEm/lWBPa10yohnDeRDNEcN383HrqstVZVN6+74oP8Q2GKNEuZth
BzR+m9gF5VRvFICV+CJY41Ui/YekpE8Fq+E+LnGEaqZBmNmdyKdWi86nEnq+aqz4jC50byDgmjhd
QVHgZMExZjBWKxox5+kgkCXEDZDf3M634iuJgVDosp20Ie2FHp7V0zvlJPrivupwJFoCASb6yDo8
yCnGE5+u+ssWaVGAd3aHA/5u31XIc4QLWU4fiz2uav+/Ca9ORo+jhS2fih6eblJ1YbAsSs99Gznb
RJDnz4BB2mMtBQ5cwj3AMrdg62Eim9ewpP70YWT14aiRk4SY/GAGhAQwyuUew9mc/vsiNokK1vaK
IlZ4NCtfpwt7ULA+qr8GKIZwvpxSVB4qS7bc/9Vm7bMeONZpcMzyfhAalbpqir6qzPlH586M2uzr
d36MSC+Z4zavTlt/p16kWe19mSSW/1Mg4Rlw+QzLZwaADaBktzNC+Zsi9SfLplm1wX/XDA4h346f
kiALP8beJ3UKs5HWBvEfUg2BM3sGpQCvVo8pb2U+hy6RYZ5sl08o1xveoigmwL2w/YanC4oOIPPY
rkudCWcJwYai0foR0GcVKH+4YxQXrsl36Yu+26AuECmKZ6+2H2Fo34OqYWdRX2g6rRkMuVmx8GUZ
3iK4wJZzvdY8ZYYtjjDio4BuUWXDf0PcCIKBO2RgOXRxtk1SwowQaILADsrC6vpqBkyfDt5V0ygc
NqSRnDWkmlKkVre11t3wjP9NGqqCtIIHxO5apKVQ6f8JbblcfNfQe+KkM2gaUU6AXEUkCGDK/kyp
r+OlZTECGy6oboyft9rbinHX1DrrhLSaNRkXLuTLTUUi/0IHHJPMT5qfCh1o6s3MDBG78NpZnr72
3ntHjeXnN1FUhOPx6ahoqmGTyADi2d5VAQyRYFDPel0MSmimy3qGFQcHUIvTWAt88Z5VYPSbNpWR
WnOD0hJoa+tHrqaTQ3ETKa/+xQPo8n2BolR2RAM9VjpqEXk8ldDOPBXwFA9v3rs1XGHss/hueL51
OlpDcmqvBSuTa1+++vUz8VH79KTZHQ9enhWirOIMFoLDOgpb1gpbPCKw8tZ0CaB7bV2sPjVkwW6W
IgUNWZ1+HwHEoy/1yOQxtP5cfUKK7juNiWwHWWXeNJg0F8YJOzrji76aFzUoEYfyZWBwDBTQR3tb
O9IO9dr8x6zBrF/1zYjBZf89vxKEeXheeneBy8JIWarTHYAet8d4aPheAmnSCaaF6vKyoYCjyU9z
nBEgAc+lM2F4eOdaHKfB2laHPG4GYMtfpqG5y6bH/mpjvomw1BWd1//GXUOOo6YJ1KZ/GQQK0PLG
sDjPCm3GLGxPHJ7FWy1ueNl60YTCLp9vkgqJGue9typ5Gy+2rwM4+LP75ueiGFiAfSWewdE2MwoY
GYXmbISthOrajeddhSnj1pQ+AAyneB5S+d1Suj2eLhJdjnfD092ZB7RBEl6/g2BOMI3VgZi4HyS4
Zzm0R6tn3AxdQT2V442RjKYMY3cO2gg3msjRWsNNO3Kb5y+/jig5Cp278v7Xbw14iA5k4zhhDg+q
QXdel5uSkQOfWGdkLa/93oEW9BswUx8h8+o6VC82E7BQRnXCDSbghoFrv5dgJwegKNyDLIPfKLNI
msb+B9SLFmZE0uQG/NmeIQ0JlVJJ4lU+KGqaV+vydlvLBU08Kn6YF9c8pxQVw/kkNe4gMl4Cq5Mv
8yaDB+4jBUNK4YDHApGisONkS0Z8DRzikIS1cYXNfgQQVAUHcvS7cNBaofPAoQ9ct1fjBhV+KltV
0Qk0INOJEWS/bAfihUrAV6gbut7NwcvJg7U7d4QYZBYblozqBIyAMhV176LZbGMmEAFZFXL+1iTM
8uhQpJsn0y2LzMVEJB7qQPv7r7JEfyRCfGc1aYh96rdWrLJMvxi+d87IPY4rMl7sZ7KCtCGIx3/D
tO3BxgzwAMOecudWGJXrBhoGxTj8hwSAPzGCD8SKF9rVk71ESyJ+zQJmpBT7adTHFtFaQLZFtcCX
lacaVoyaFXpdaR3Lo0PGD4MJB12EZ5wb8TnJUB3v+82ft3FxF4fIu9uNYhLXOXCMyMfHrp3QPxJm
O6DAbRzTPPADFWqo1fAYvQr7h8V4oISg6cjeM3qDYpQ+jcJLvgX5Kv7rbAbAwGVwXPycpwJUxI3s
PWzgplMqZvdh65FuvnE39EvwmjqwgOk17EcAnyJUDVOmhbZ/BGYY9/pGv4WlJU/sUQnVU9p9tY3o
X+N1a3Fws9BEE2RAJ0IRDia0jqhox7LCzLB4BNe3eG7HV/0SH49ZzYuN3gpNoAAyFJStiLEXdRy7
ZEQqZgnGkG5Ao0QzqJK3l+s3j7LqQqQwfdbQd9rfw+nF9NNHbFnBUm2drDSVhLozqHnuibqx06c4
rZnVZK792W51Uox+GEKTvRRYPpXQswZLsJnJJTwsCjVedi3iDmls1W6SHCIHBTpYGREjWSgSY436
Ka/JM24ueo0Dc4TfV7zgDt6FjTiFXUkAu7UXMtLKwc0m8WdgyDCmr0ur/3TNVCizsBs0SzfGn+RZ
VXwm+hy7JKzUiVu9oqBvY04dgXeQXzUx2mhE1kqYnCnbToLxvTN/qsCXLV4+MgI5Pa1z5MmyzYBw
uNuxADiHeVk6qoEnfPm8UtsnbPsQxdyD8xdei19FLv8OXarAu4+IRLtyRIsm/NmJaeB+hDkpqxQf
lN7YjeijsRR4bIFPmfH52mc+r5jI5vZ5QVZxf8dbM/eosfCEuV3audo06f9e3ok9089No0b4ZO3x
yJX+Vg+RmRSBLkfflAkkcgDFr2nNfWhW25lc2cEsoA63OFqPyudbqMFPn6HLRKLSY0BWiVFP4rbq
MaeBZECQ0+YbxLAok2s27llKHCDX9s2v/Oc08ISAxhstd+POKUCqyBMgrlSjUzwC/DyXkcAXUqje
ZI/aDrmmh4WqPEw1WXmRTRekwOJNJpv1P5pVITJZQMMYWfbbF84DJmvRpJ7CtmVnXEHuP4fbU6sU
JBC8mFjmaSHf7H+KhQqi7pyfp98j5ahfIVLPUiz41T93HDpsqeLWYvkr4bJq567urbrtL8b5egb9
ZMxh4UNcFWU9r7oNDEhWk1cyGEW5Z0iawkDzQsGdDj1ithT+R2untptGiWOl5Qatbk4f6PxvjkY7
XXnxo6u2oJA9A6+B7v1KDnwF4KHbVEno4K4ky1wdgYcDbyYVQfGM+vANkiTbfRoaC0xVJM/HyXOo
3kQv1FOGtd59t/CCMQhHKAzFV8k5yxkgycMptTDoaMkNhVp24awhdy1CVgiQyMwlHh+fAfv+Sq/L
gpZ1vF/0+qmV+XhW++Di7/cjiLbBLJJ1BVn5f2YS4ZvcVjGeo/mkiAgxOkyx5L9qsP53u9iBmVmK
d5++jvCNsUWpVG0d4GjVuereZKqmlyZMijW8qeSk7Nsm4T7MljYcN8SmrsnKLOMXlSx2sVudJY7R
u7IrttcFzaNvjwqOvlA6vA8s/bzAAdq4qiOpheOw85cTC2KpO6UDyO9iH1iTUfMaWFNjl5xOIkUy
5HR/VuQunOwXLnpa1b7Kg0ZNLaV3/IYOcM5PCKPPa+AZMy7PElxGMkqeffn3zMvd1EicqFvar+Oh
PRLQNAlsHCecTTgiy4jr/W8T6QpS6IGbs1/j2ieJDfqN1cQR8W3NFZMAoTEdFIdvRn/TejomwRHX
Dvbbvf9aEQXFWS/yfikqQnfe4qdkR1H+KjHhP0RnrZBpimuyz5Qp0nVgQumAsIHqt/k6JVTLuly1
PiUzGtw/D9pGJ7UlhiFpOedUEgzyw0Oxo/9TsjcKbg2OiHyPxrt2KkR/GYzOwrF/oSj2+NMitA79
xhcnZ4gmUa+AWJ+8dezPj0q1il1nxibS4kVkHgv9jUGJaaLLRIMh4FciEyyb0fpH72tF3NMsIjGd
3E+ktWoCMefp/w0Zv/Wh1aHrya7SJBCk9yH+s34WaEfDpNSB4F/dtasqx+1Le82KaAQjD0p0TeQE
76wpGvn8X1hj3Uv8VlvAGywPSEugguM+LJNFe4gohpBpmhHfIK11YqzOufz4Rs/sXFJIsT4pPk3R
mX5jxhwLMDxj7heIWAdDBMBr3c6tkP/dFDetZWHwLy/Iq8X/TvQr1jMkbptSfCkE3B8FWaUr3wKl
Xk6aEK90H7vg/Ctc/ejzE6HEyckxXOjr5LQQpMJrVXlPvJxI8zH4BHclY+g7sX15j0zQt24drmJi
xhWawwpv20LQR2Vou7mgvAi/ngXcUKVG0/iJ8sAC9xwDpsEjK6AK2ib0WNSC1kdOJxhJa+QYNqsq
3sW1N0aDHU91JX+oXrkgH6dc20tG9svDifQo8Ar07th2qpkybO/aeUuRa04hWWV14SeTSQgIJ9zO
m3IPlM7fzOnrFsW1rHMarrTbxKRhBQ+4h7jR0pdOdYhfR+2RQp2T6FrwHPdK+dihAhmzdb40Z6Bv
O8y13eptjSLZ9Gm5I8CDo0lhfjLzwCuib+NaLVcWmHoVu8B0mDupaqnPQf79+I12WDUo4T4qSG/V
z5MBqHFvy0iYwSFGmebiezD81uDP9dPBWxClZ7DTimgXXcth23B3iqRqOx3dOTTCTZX02q4dYBRB
oRB1uV8dxX4Si+06YYIqkdcFkGh74+1va4hxa/dh5ozp5VRgZ2C2j0BaSRmgbmYHPBeC5Gu7olKr
vaPZqIurS2aKGIfUGQT/QoozNy2pR3O0pZRLaknyJLznGb+8w8RCbzSNvBEAtvq9G/yNMvDJ54O9
pX2gW8q6AzcwdiNBKgI1rC3pOxzZDCHu5BeaJi43sN2fxszpv2fqK2hAr8GhF7lpJtVwS4w/v0u5
7DXCIhrua5xBLaebWdYJ2jGYyrLQWw9Rnw+0PV4RG3IObFqGBT6VYMfEiaWHK+b5znT0YieKDevV
Y0WatSwOpjo+k27i8XSIW/rvPGfkL+u148NEQXZ5uDkwjhpGLQGa1RlA4eR1BpIadRuxIKscghD+
ygctJGZYoDuOuY8dATrE+azAhyvYGyAT4O52v170nVXy/RWYJFzsR2KgFWkBITVXwJlJ4VBWdNmD
InmFroIn/mH4Z9okWiZpK47YZNJJYOjN3fJJkPFNoGipkEqDT0V4fBfMlvOYHxViTh9UK0NX0hDn
skg+YQzKLMC8fb2+M03eue76gN0cty6OtiJ0gFIJo5d+VlwAouKEpn8Qw5ig7rtkzitI5RZRp0TJ
isag4be+d9wcAMNDp/rFWIHAg9NFjaqxpx67CpRsRmcarDAz/p7JC4Mh69k+nvbNzVrJ+WdvrGwY
UKTBCIDR31CfSK0keYU/LW0UmdIOdlJ3ObCwM4Ox4y3CwdcNbeCQN3QR1nHdmeL2QdHpKOfFI9nn
xw8oCCI6MmXm32nFubgLqW5M4XECgBEi9VvPFGCXwh3lJeRg888drresvOvTDobthcIsiT3ETdEM
GMtOwnoNG7LWNArOVfAYIl/DLunaUR6U1NzRQ1hlwJ806mCF0ZVcMVtXE+EbwvnXoy4Nn3e380BB
L3RLOjrXmKaWoYrVPYdQjUwmwA2q704R7yUDLq1KOLtzcHTYBLfuObJuWwFEMdH5PQF/XP9xmE3+
/pSi3IyG6ytxhVLdPTnPzZrVeg8uwGN6H4HrfqqCJr4o2s+KxhBkw7W/m0QC/S4AVL3Jk3Bv+2ok
vKqrqldXY7Oe0q6oM/iHOhlXXtm6SRGLtUoafyqRUbnmY8sGqQonF+tx6W/PvBL6CE+4RInE9EVe
YwVe5cew6p8m6e4VtInVUvtiUjcOc0hjxqTJk5Z3zVetxuuknDh4CXQM1tx5dX6aTONz61h53Ovh
h1MNFY5XS8bMRGeLtisZx2NjbFWmhi53mbsc0XAua3HyWuE++MnvGN5Dg6JEOHxTSbTy/hFQh70/
OfhML+wSYsPP/gk34Osnn4n92BBuqxf9hUTSAU9pFq3NX2u+yeD2wUQsJXm0qZHENLymWrS/fEfg
1e61BdLg+z2WOdOACu7ORctBsOrxeNrEk4xA9nYJDUpheDE+o/aklyjnQX1YbIG2oahDxAScrAZ2
QhZuwRc1JYEeOsVGN5zVGhlXAqV79AEYNEMkpG0w0BRBVOeZY6mp8PQI9sgfszrfC4FxtK6C/kA6
i9xLrwBYiLBRj0EK9Mj7FwMx5+TrfJB0m9sgfMIHsHOLICJ5Zydw3TZFzpKK/wLD43smv1gtUKM5
9nfbbTI5YcwvH2231+HUI/L9F2FjvWM3oUHhKGsFWWr9aLYQG2WmI/XGw60zZIMgEIzOaRHTXFD+
mfrCIQqBhOWl+aTcg3KAv5ShGMtFxVdiM+qDQfoddn3N53i3YHOB1nSG7mixETFE4DmcsevtZfzF
VOWz8epmYO5slR4ffV8ajbauDIVrxtyW5AJquHK6skaBSAdIDiCVU5ZRs/3II87Zw34UHkRuQn5M
oHAgdAbwIBhjJw5KwHzt+wJJhSYVEpb/Z6ZD2fZAErW8Mt1q/eflLch9krDX9HQaOwky59nKfFc7
1S1+lOYk+2eF0lrBFrVo8XIgsmToV17wJFB8ZYuwgYWFkCXGFogVkZgJjnvpT9hEbLJY4WUdT9Rm
6w5Vam86D0Wp/hMOuxhuKrLXjn6sSMYY/uLs+VIQGLzaNniSsF6n7O3fFlF/kgkMQBffAX4wAGFE
OltjWy3vdiLJdlBe3qoYW4PJfifIxhxaLnyX6sHy/XtYzPvYpxmyLDxVRalnreGqvzJmPH3Eq1oa
V4f8i25xFYmxiLOBvTJzMeaFo7AVd7V9KgLKUk3KnctadrGI9HtXMZamroFr5Jg3ODxDL8AOICjD
wlhnhDtH1Pz7GsvrQBj+ZpHdM64qcubvgQRy5azt1yxeBBEzg180q7srmphCicx1Ch0kyG2sQK6M
gFNT0iR7hP2u3MeY4IiptkdEJnk8Tc5shZQPFCwRLYN4O/zCM6u1j3xqgth0Vpe87yPdlywqzEjX
w1kfre/ehJJYDlZ+0KI3PXNZ5vjNeRPA83cYZaV7AnWS+eX0nBoKDyP9ic4woHVXCc1bniGCskx4
rpwuaWPDc1v0VNTARWTuHHAd0jxjcYKjCt7TSRDTnxPTJnWIPtnEJ44BvIrbxcrItmbrrNKeFMo1
3XBbABExdUz/NKxgCN5J17G+bSx6Z8b3dp8ma+PXxRIDb22GCuDRYzliRgYgxZ34NRMGURwbIp4x
ds5FWFJqmwuSmTFFhf8TJMaBZ8mBZC5yaXFvHkYd0cj9R8ET63OYLRyXaodvjmSivp5Vk4HSY2RL
EUZBOrGLWHPnrePFwh92YkFe6+Jk8vRvEjlRRI5MSOSxR28BnTWSS0rHg8t5cHjsii5ctiQckoCk
wccost50ced12ZNkfkgpU375kj31YPLUhlyNt+yeFCzlaf4OughWt+lqZ8trIkVity3EmKvg6WB6
RPkMSLAVsagP3JDfXgRej2JsEVr40nJQv1dpCEORB6itV2XXdPIcyEX7oMpWo1XfHQpKBf5raLQP
nvFGgpzxPfKprGBFGcPi67W4zqWFebhL/9HQ63aJRMXyIrJD8CqIQn8nb7Pt8FL80LrgzSWowMD0
hXIM0shj0j+sbv6+eAAfJPYQCrmWf9lFq2I90HDmGqUK2V01G/T7YnscxifhpRFX+wIdgCvQoW5Q
kRyK6eAbH8CMITMm62v2fn80CNznKwBAAENwHe/eAMTBTXlQ8NXBO/Ql8uEx+9kTFXpW9tuo5SGR
hznzlc6CzsmFkQDeLgglYpJO/NoTGk2aHwPqGSuA7cE5J9X0qZx3OGHhxHZ1HRmbI7JRz+lRDPa3
99BaK9Ruu1xmZR8zizmQEXANK5fbVHy/rg247bm3iWH9mehyoyXLKcz/f288fAXIipDYYA9G01Gh
hrFXozIyCsnzpMqZi1JayeQSMCfb/zm63jj5a1y1t4O320+FvoiUQNhuxwp+m0IFVK/siDV2pcPy
Xbo5YAxRsZ0o5bZJKMbJSrVGVcXfjYA8llJDQC+8BiT/ylzXmmbILQj4DJlCFE0NbKGwezFKiC0L
o19xU8g7qxZ93kRjw1+szXAg/Dpveb7A4hA5RDW1UUy9Ts1iqYsX3kz2LHQFFPjmmUZuealg2XEu
vKud0cyWetPXVIBR36vPjUna2ZE8dRnDvR21dILM9reTv1PLJpn5JMZGK0dk/P+ZavKOULVTz9eO
ioeXAWUnUS9W4z15NhX6KvAeLAX03AmXlGK6ZQT0h4TQjaLNouEAnNDdgIK5+wIGQ16E0nSfAT2d
NL9xI8ErHFXY9gm4aZZRjTNnRKH4ncVNJW/7uWmbCjcwwV95lf36vTIG4693VN26rh3hzbT9e9qe
dfnE8EKMGZh2AVS0sAJYsGu58P/KJ9gJkkxVBhKeRGiZeHRLwWRgPRdxXojuVFoXMS5O1XDbjnfD
u834SpG6QtGMg9vJatcx604X9KT1XNf9P33mxrMCpSJN1NRi7ueWZqLAe9dIQrvZvOg5G4L4Cife
F+LLxM+t1tcPcx9hGKyFCujSo7CXX9+poAKC/IYkaKd3ggaqqzjvNmznQ/b8E+l2MBFoHpw7Cvty
vwhjARgXD0uf1f8f9DdQRfh5pd3B9cRJrB/eImR4nigkyH8G/cnNKiR8Gy9VhSlQlcqlQ8X/iKH3
2+8nJ2tzLDECvbfxPWisazl7iHnjBGpN50C49COwxskYlPk9AFMv7TAwF+LqRNV763+d9KubOkEx
f9dduG19yaPmdzOPPHmQ2NPvMZ6+Caf0TE9GqNlSlzB1Mvn/CT+Yqq23wDOeMxfnsrD7r4PW3JDf
Wx7DTcIRm3uhPmLkqzYSIfvHWosqR0GwXuFrN1sMtsPFNEP5yt5JfpcaptxNpBVhiKPKdfo6dhrp
H6XSlnnMjqHg5PUoIDt4jTW3DfPrFlOzjoN3l8HcU259QTgVC7SBjnT/qIv1V4LItq92AiSfXXzG
rZBnVPpvVBBQ4M4yGgp4hvMyF7DuAM18clctJhER1+SMHHbJTnuAaBUhIuhTsaBzY7hIPKniisIv
3fk+EW6C35tkEL/Tv0vw5cNZQ4qxOrwb65RC/SWviucRgV68fgmajSz+QOtLgyumf8nGDW4HVm21
TIR+0wLJE5njSzDU2kATu0xqYoviTsCSDb4syNFojixPIW9GMmUMYrQTt+ubD+wUsSx0VTFuIdQh
XfG6YSOAyTzt2kYffpEGc8OPrH0/v9GQ1KRA2zSalUcLscMlFVpuE3pOG17mC/VM7iArdvgkABbu
Zc1nMT00IpzgzV0cAVSsZXFUJZGX33cpMxpCeoLwWQNQKkkM7jFEvPBrKgnBzrJ/oLu/SnEyQ9tC
nIW0Mjw9cyE2bt2teIGyLyzZ8CknEaNCZhPyQ4cWmfncx3pV7JhGHTYDA2o8QGx1akogENhxqrcT
f3UQ3jR6M6Sf1ZeSf4HX3Gr9FbzsMFGdaQV4LdBa415KyjWrD+mrlmonaJ7/kF8OzChxI2eXqhUy
+/++x4LofNNwWt+SylXyXaRnFqGKZ+htzFSwv3t9ZjJiNfF3jw7i7AbQMLYJCwNytnJ9fe4aMCNO
4Gg/iHc954riF01wd/FyPeKTi9mO6YJvraBEXvV1FzRKO0bkjfkL+gftjJDj9RQ+WwD1uwivqURU
XHEefPL1b3L9QoncKcYpnJRoczsK2hYIwI/L+OLNvqu40yigbgW3mkvYTXvuDQl9glUNLXns/R6J
njMS8Agqk4/nfJByt9Srvu/8uyWoOubD0RMrjrhswHtVJEs9Nt/Bzy2mlTKAEpXvGTP5CKxaqkya
m15mL4E/fNs2IoRSjupQiicubQ9uNi9D2LFCQFrkftW/0x5Azf75Hmt4OlzBX4830wJ/Uyrcay8G
QFwNExTSzCp4cSqPFO7c8WKw2WSmDrLdc2ovLzr6HiKaPBoVzcW76xLpJiaZVaL+3Wzk9JLRPNL3
lvKI8wLDbKABGwgPi5zNaF+p+4eX1EqBvTk1FSxt/3UhRnDHEQgmgIkvvc1MKcN/J2CzSRH/u4C+
ivoOcRyMzYJOHSRY+5Q7WFGPVVqO/PzYDShb/L/gzX2sKpFnWQBBDheNA1dmtVgyYf3KSr/B9E4l
0roSxPAiIi4/C5qG3MFsRxKgmNdcZsZ6eAaeZEBGMgrCGPuZCuUY0QdiUv/7QQJQ3+seU8BgYyAg
mduSl7jAgzQojtz7sl9RK50oEbBZivmMiuTWdt7dyeMRZKBm5Mr8QvaZMjA4hOHf8lpJy1t1X+sf
ZdghrmV6Bh7xlsnhW/NDptyxww27vGucOHaEMseP3NDKpJsyW7TmWCweaO0AJRRyoKTnRcA8331r
wksuBoOyhwK2iDpx1dCfGS+u4GQBU97SE+F5rhgoh5omnIlRTbrh08OyDaSX+HURPcmRlDrqCr0f
fNZO9hv3C7U6vRmFm1pVFDGvQP5sA+5EfNwkZ/glw1PO5AxbuXTlsHypixkLDYaewt4tgxz96mwg
WlgFksJ5Gc8Vtzsqu9nMWBhpmKebx7XWciyCWqXkm4NZ1aP3lxtq629FxxhI7U+zhsk6maDQCkLc
u8INEqeGw2CE5Qm8gzBGAoSzbtOps4T3QV9Wi1jjDgjlMYyS4+/TNhWDfEAgQdhVqr1kpcA0WM26
dtDDOAI2TCkX0CyRTGwrqVPIzXBtSJv5xSVeVFn4oYS2c1mXykckjQm+qGLxUfWfQMtEdr2t1cLs
DQSy1vWJlvfGlPWeIZQ3M+gqRSWPpSXK3XfMktkFUaY/d0LdihEdOw52oPlgClPwRuvgvMs3odES
x2atvXym+K672bWoxuXMF4DXgBYT977txi1GhD5jDjovH8prx41hFmnLLMkxyeimxK3qLzc2Xej5
TNCRIwHE/UCVezOzDZOYOYOUEqTrDrv9DwgP2/9/dBOPIEiqGLGQG1TFtx5BNoZGqHFqeC15YUOA
TL0HMmCRirIB9etExUFiAtNA7puTpR6z5fXfM6CSPyrPKEuhg3B7xF82lnB86KLg3FdfXlb4eRvX
XJlRmoDLsxpxMzjQSsFiAajpg/xPknLUU/mJjYlajsk8fJFRL5sr8immNPSp+QywVbOVzWqIcEQQ
Tva7/R7QO2n0U2HRZZgbbyPHjbKpLzXKKziY/d41nN5X2Zi8Q3aFIX5elOH4Fd+rixIgDNDTiN0F
YjNVvR4lZsk0LRX/LFvfeTw2DI/HY2F0JoTCq8MStrXodeWDfRj4DD+loEeB1f9Ryycwphq6vqAZ
5oQrCWw4EgvqzRXFSbVFO/C839A6yfkT/cDd3ZY6M2cMq6LZ+MLfFzWYSnKgHpADGCb1PbUS7R7V
xEO63cV3rBzKUPEytlQBnsEwfRj51yQvvTgLcdA9uF5wrNcjvGnqLoKqe6xwcogE+ig60lVDEl5L
sO9WwtqlHzSE8c25XfG6wRsfVt7+5qW9qnLQPMgAvHbF6esxEeavpJxF9VFCbsj7rd0AQaAFdfXz
YcqyPqQLxWPvtFblc3RqOTBTkHss//4S7XR3ZXrtYdG/OFUAQQwJJUhzvDuTDCbpee8mrgagAcRQ
tUzIvZHcaA6lLUewnVbO0M635BmlHbwoXxTDRlB5uPCwfzWzIz5dD88c15NgmVJSzQthUQms2mEJ
toUVsurJRv7OL7xnXlEZEwWkcA6SlblbG8gnyW608X7QB5H9FKum3f5bSGiUSc0pUnZ+GFJjom1Y
Oha/xNP/eYueswvh1ppaEEqINi0BnBTcqRolZDt9oC1tT97weXA++zTfBPUlWYmmzS3oe5FNh+ip
Ay/fkRBqWvuUCCLgbuXQ0Ovw/vSA+a1F34nUpaK9PnRMsBBvAR4iSQrJR+Fr6wcbcjLg1Vja/guY
2eMDW3OefCf6r0GurCbjRyoxGLYIQiXQJ8Rzy3qtfJ0S4iIFJdjCkSjJolsDa/Q1wXHDr01cdMIj
0JTA+6lAZhS2glx7oCViq/T84CrwfcwBAAEUYDJcNe/Do5WhZB4d0ZNe/rUOzkJz7bNVtJvPrYYK
bXtH8VBagB+k1nQsYYmaWjHjqLhqXEZoyrlUOBw2qb/voxRc0ZW59vBUKdXRJqzuoZ3pV48gqlQ7
vmb+YCawiUoENOhnr1+Rhk0QsdLGMI2rB4df7SP8QIWe/sOcz7RV3dBwrVf+qP3iz9V9vEk+SY4+
w85tx0y23e9UedJsiCvoQzSqJHUnlwHamabCjTLMgL8/QZYhRhEGLZKMq2VElzmZX171BxazNzd9
tsxETCtCYlhzkwk/QtNEQ7UqDnR9wyUGs6m+GzvWdS+bIUEJgHwWSY3+L+gO5jJG6p8gSF61+3jm
FVxZzr/I1H0wI9p6W8zBfHzjA3TmjPwwyCR2n2Jrcs/2xJmuPK/WOpKn73dUQVXJXJfSGrmMqqkN
gf47H2Xo21CwdgliWrf/TdojIRwWgTG6ohuQww3Q+XNm/oRdgp3EMqWPSTmkk92eTMzGg2F4xsNP
lM/ve5t+NyfodV8VwCKixzFqEEAcuPZlp0JNobCDs9ZieQKVMoSqcVLnzE0H1eJbFtaWm5D7LWgw
me7ee56YtwLQmYPb4hOsEaZzEhelc1RWSRm2XeK8fLrL3ZdTFfxTeeY464olGuBb6kQGlTvco64o
CQHiOgVCw1Lyz7u+nPo04zEhgAHhEdC8kZvf/vU7ZZWPQRrqfv0X3WTJrtFC8xpP+MqESw3Zexn8
fu0W9quBY5X15U/SXptVusjf2ETWISKNrk9vqxaRG8j9rI+i8NrLYLr8cbKIFOPk7dog+r8INCWK
eXppDxKmgbTBUtfKc7Xf4ncrrri9kG39GmuPEiwzsTBBp0CVpM6ad7vxaZkQ85eoREiz1MmsoT0j
+h0W+ovXCnuadhUZDoYf4mVb38PXetPzm07xZvHQjhOQ/OvI2jqGSWk/ZpxlB5OMkvl80hm938xL
NmmVJht4ROMKcYGv141DQdYsDe8tAqwS9trg0SfZeTKmx7KPR85rnkEzFSmNnGwvCbVxy0wU2iBQ
SWE1a3MNrJHdwmYdwZKHl+hImeHtWijQaC65gyAkX3/+E9J5DrU79evMN6covkkKshdBjj0mLdgN
pJ2z7LomdZ0KC6WBFWG6gnmrqEd4586vfZxQGHobQxMvwUcRVqvvizbQKfb929N3AR/JsGfXEWU+
hIM81hjbLNk3151OX9MQavKQILVQ2irKnSgStqApkng4+NBqltZlTMeNop5/v+rSeO8YXCo6NdbI
KWU5z2gDRI3QMKNeAXDu4ZEcB2yOC8GieUnWcPzcTMxn9+BPxx2iPvIw1fGPdNHH9i5KUtPfnl/3
PYL3dqUzK81XZq6C/eQyIcXswpO0o/UE98O4zFSG7gN5HgzL9LAT2UNjilXz5rjznr9ahjca+BrH
F+rTUxHCF0TiUateE1MeVCJtdcXmQLFUVFKKQB8Njao8yt0zSUF6toP/eqdA+5jQvn+NcT4SzYTN
IYuQJfU1rWh16Flb8O6G3u6mijsrfMoecoLaINrm+k4RT69dxsy+hLP/iIyDtNrFARgQGt9Iadnt
9bRk9mhRK5mFelCHFW17ahnY3Cx1u9FC8vq6AUsG3cOMUloMNOFrO/kiPuTsCZ4GqiWg2rKgADYp
J/CnywdmTxVHt8SH0M28noAfaEVLZ7QRBFY9J9pV52Ibb40WKgWtf6Vu++dDQAYQZGzNYXKMPegK
cH+tFCJYHj5W1J8zoLUlXF/wC0N42MXwU6UMvjXCK6jj5ihdQ4bt03Q3p5HRXTVAEPTXBFrObLo0
q1V2AX/6Iuq5rEtscSRViZwTBHLR9ZTzFXTtgG1Z1LHeLZo+2Hw0q+YK3Uh+FDnb0Y6PXM7ww8Md
byQHPfZfg1rb4QsIYW0M1QuWCAw/Use3BGP/2xCC9bYlEciSF9y427qJ0sQIRuw7NxR7+7yGearn
T63uEL/360nE9z3EkD3Bk0/E+9CjOoEjOhpSj2L7Rr9Swm0vFoD8wwv5SClmq3zBawD2Y+bFxj60
VK8QIM/Wma7p0BJyZ2iXhdsc1m9oJOfaldD78kRaiPZLXRYM7lSrT3LNRNJGC26Aw+jRTDmoWYtx
0alh2qJc/2cbrrZQJloxJfV9hKf8Vb62ik9PGbA8EsJ0vCtdmLnOWcRlS1Pmbw9cjoQQgwfRLieN
qTT2HUOElcsIcE005VsiCHHT++m5GOCxq/b9zl6/dDzjIDW4o5/GHIYPkqciuI1vzIFsE+KuQdHh
RkVSGuhWNzY5YojdcmQ40yXe5dJXPstfL0VjGY3raiCFGSr3qcuW3/cFtBOc5SKNhSVGBa92bySX
mWj4MAgkryYo0Xgspn4mUuFjQn4AGi4mF48S/oHk+N/B/hI7J5wPSPdS0qslAkavPDU5F3Nzl0c5
YZGcTzlZE41ImJ4f1vjiSA9aG3bQ7Y/oRlx+zd1732+xCx5J2mSBRaTuZsz/Ef+JcrSKkroYQeSK
oJ3S5xrOIUTUwcW0nW5sukV/gUNe2qMcd1j9pICf7SwzZ2Z1ugWj3j6hFlHPsFpESQ4hnn0zgXpo
MhGd2sO+qKU1wYsWrzoCtDeC4zl3p0oZyOKGkHs5NIvvK/UIAdXwS8S2uipYabUaPL4ZFxbuwtBC
wus/NJaFR56pqm21I3FbTfXMGfvaOU4Um55FZahuZXdCuwZf2ecPEQ5Y6t/+P2An91W5dsuENPCA
MQmcQFXRoxFTUeRwVLryDWi8z30lKHUQC/R/bFrpsOXaTYRALM7tC4ZmPjrFAV8+KiE/MqAr+Z3l
5Twz1I4kFuwjSTl92zzCMGL8Qrr8tJ3m+vGQpPY0QH1Tlp73YhVy79ZZrZOOhI6oj3W+UXKOuqs7
7xlgdyvO08pxEmqXlCVwc6v45+Hp77xhDS0LZo24UzGFBugJw5hJBKAohYLVNHDcpooejTTszNfK
39OFNZxPhMSM8wjFoj8BfBxojQrg7uFecM4P5xjxxjvu4+E49C7uJByqHo7Q92xmUwfzo429WWJ7
IE2TNmJkCAn2ViBVCZFw3hCA3PKYYnAAVkO/ERML9h7hcmuUkD0KwDb75l46sjX3zyrAmpfN4mvP
PLpGBA8jyAdri0Eblp25qh7RvtFTPSZHCoroD+JIenVG/wWFFLUcRcDzcNfSr5D6yP+XEiWDulTk
zRR60UGK3CeWBXDSTeHCYaryCz77pCbCqGIOpCwVcYNrBJpjhd2Twk8jBCZOo1lheyQaeNkzCeA4
gMzIUpgSDZSc81v44o6llJGvBHohoQtti03ubI3amrll91FI85m+EG79+dn4LvLePZrkRgmSMcla
Z3jLqxblazVyR6BmcoQ5MLe2IF5QzTLia9Y2gOl/KbWZB4Y9xxSEVkdvq6mpUflSTqnOxRWlkt5U
aFveXM3zKxwCfqcH+9kHkUlq1D7ynAxVYNGvP6f5Delp9B40ecVshFrp5yHQLvhlVOWGMjeiBh+/
A6WX1R8Ivqb/Qa3m2PdHzUrRiLHePmdu+Vh3MzMHEZTMEKnMJ6DhwDwfLOW3ISaVd43cud2zm2Kz
CmluuneB/XxD7LAPHxFb/bu/7aAUMj/ZNEJM1vq8g40IonzOdbXTxpz/H/1eRdZiI1GgPFNx5ubf
B18YgE2Kak5iXQLbhk60/I/nVrOvV1/d414LOOf7I6N1jeW2LhaZ+5MOzk8rr7wfflsRGDi1nCth
YhKHaLN8haf9mLHhfWyGerjUhe7bRVo1cQbP/bclfTl2TFtfoiECA++Gjy8YjQErM85VVlFRjzC3
Q0J7Qfl05rdOXjYZTYU3Z+9bDIlSfRh3cytHIDL3nxyf5k+/hYl1FOftjazKp+juv8EIoQZaVY/0
XB5zfAg0VnAZdTDMW/lCMIxEiwjQlSCKkmIFk6EeJrQAD2CKflVuYaYsj88p80H9m/WNHvcHUISk
LAonWKha7VJEBzpHFlayIjRw9EV/f+6KNDnOfY3Sn5Bt2MspjBrQUNvtGuN3jbsL5PrvgAZNG6zA
n5RpkhtDS/API8/MPkMQtgHEBW4NcKOGOwztpvo8B7ExPR/UEFgTE1xVMV+tAH5OFcoq3dz9eanC
lfn4N9K3NAmC7pDthf0MZFMZVg0MaaCluKmUz4MC4jQIwtJHcgm0rVnQUIqZ1BLJYV02bZtMkZZT
X2cezpyqzcU7NsJ7LeLR0+jneUwHgy4/uxZ4CUh06VAzL98h3+wF8t7r6jtyzkVVlxaefF7V1mFI
LUqxPWhyrOOnS3Wff1G964uXu95tHmKzNrH9avqrgWTCyZTOlKRYvmLS/K1+HS4dm2ceAR2pYEI4
OasPsb3lgWvjlEaj4MsV91eePPphjQRzJqLeLhcCbmMmM9SSh5+7h4DthhkulXVIAzahqPov7ua/
Oh6EVfV+pY2Eim6ODZhsV6E7mvhs6gB8+X/6SUG2yEfjwzSTAQ1533XvWzA91YLC2zHrX4X3pRhe
torJ/Rx03uWs7IwABTlWerPzVxb3qUQTiW6gMGIK12x9QK8dhlIR4wS8GFH/AZWEeuiMjdHA2PeY
Ire1Tm4PhzBGt/kUTX/2dbdYwjbH6myV1lEzuXNonjuhRydqmYgaeQi1jOhFBIEASh2uq/9CoGAP
o8w4FweT0ZhicJZhWFLMwAqcjU/mN5EtIfKX+jucsJmOZewNQX3CSwxnbrjfvCFIGD0qB2e5lkXQ
IqcrW/9d7/Myit17QER+f+PjbHJ6qUTYBgfqziCrS2jX5yb2d2nul73lxgVMg5wBA/wurjyP86hp
06QVkt5klrYiRj2xIX0beZ9Y/323P5q17IJwtUjhI9nSzR0JedZKt+eJwc7JXvRPwjsyKjPPZEaV
OJ5KXVTK5os6OJBd2N9W+/VHukrGoMurhioyM4/jiYWTM04xEtH4ljkTQWsPDf4LIjk4Hbyr4L8E
f5f8qX93ee+CJ59ra7R0Ag3JcLmmi7+IG1+OpNbS80tJ0hS1wtNsw2EXfuA4GSkS2FQ7MhzlwYSh
r4QQhh9fFDfZ2wX22E5CyVL2ZvSwy3XBk1mg62jJBsraX1G19+hcueZ/nAanpMkqtCOnsdqeV2Ue
3kf40ODCRBmTBHMS8YeuEO5LlfubZO/NPH/VSM53LdbRbz6wlvyk4NysUYXlnY45MtEKGRqU3vlH
Bler2WP5tC7qvfmeeZxSPhYagwxn+/seX5itFMY6jM/Wj/XGIQRiAVUqzSaQAPOJ6/bHkzlfUq5V
twNaGeMqNn07YgQ1SU2VywCoX5EocT8WVRCYgeF5w3zJW9yd9hTyHdsR9zLoSHp281R9vwW1k3W0
ZaEns/o39Ygd/xAMAgzOZFm+yREDDC3CTK4NF1LzZkF3Nc5ZB/yKUfJEExbbisWEQc1/0KAF2iAl
kWalLULZNSuqQ6Ee81FouHQJ0YnwUWfZySHLsFtKJ6gXuxvwoWov7oJw7wxZxeqbBM/c/AaRBpiT
B6eozPd6bHjDCR1ws8HJHf5FnjiIoWn63EBYuqqRVPEFLQe3UaLb94UoTiCjyWsT1nO/8NelKBzo
2DZiMu5+xFvpaboUUJho97bElnbCnQqZZB5iRw2XO1Jccvy4gqRvdA2lbLPjWM6Ze1tgdrpf6Jo8
GETLwKQcWWGOKdN1nevuxWTQ135ihAgtqZDz+S8q6U/svBAUT4yiiNn/JU1S1PCeKLQmZ1RSiI+1
s1w3Qnk/1YIeleJScCSx69VbGUIjt0ZLdPBy44iyhLwo1+DYNHJ04WEtilIJTIsGCtqzJkUUrjV/
PUTsMmRM/lvUlum/dX0OE6rOGdnUH7A0+utt36W/6k67z/56XP7/CEfJ78AsYlkjcG5Ti8rMd0ol
PfNMLbWWEuiBeXNM4Qirh/ssIHkzzznMwGnDwXPq0SstOFItTBkZX5+GcJmm45pRZykeics92A4f
060KY/xDkihdl+ljxGeSYEpiyxf2lKRu22B2MbRJld6uKsu0JNv2S+lWjVKfGjh6O3WdMRY7Y1gU
YNfZCulIIdWrK6gABaCinoo7FkHZMBZQDPNBN/QYU1cokOqzVyWaVsh8mH4LcJoAZkgRi8WK2LXP
m75dMwirfxM77lcdTud6FPwb8M6yUtUOQjTkPd+gztPts6RHIx2GYpQKcLsxmS1YKxdfALmLH1Zf
g52z8sLz8n4Ty17x9VoSmCdTsDE4TXAtU1NsY06Vj2ENeKi5LggPTH5E0moSbpKFfEeIXdAxwXUi
fYqMiHd7MT1SxmWX2GtC+M3VT8WIWAZiBaOqnUPY+U590mobzIP4vfCdVEZfMFeAYKHJSYWuxEAn
xIWMRMg4zn6rmWgPMUyAvELm6Sx0ZpBOCXHjkvS7Ly5GEHvNKmx8pq/2C19Rg2OVSmvPRkC02JBI
tqmjhMGxxmChFP6e1Gc9rVlHy19v/ejg2FbqybvHAblO18fQKY35vsSf8XZ2nikJs1Vzy234PBfo
KSkWeQmRvyGaBgb/0x+CTvsZOZ1b3jvMRcvjcfzx431pKPZQQI2XWE7fgHnX/lsB2EscK3c1v6wM
JRM7+Wu79J+d8YKSIcy+nbzofxlgkey36VAYGRadJppb7ML35KKbfcoobMan2yquycYI1Cui9EUs
TkcKorB3JLohdqTRrshSU9c6W/3Ppqpqgqql5+XQ1XLzoH0S9qh8PP0jQaOFiGllQPm9L1EdD9Ie
p+a+DaZ+W47QFKF8CrV27t9HkYuz52fBE7ilp+I9X2oANIXDBvPTi6nGpg6//INevKHHLP/0k2eA
mFJZ1ARJAdv4O9m749Hf823DK16ZuuqK9LmEz5pj2SO9Ig0dhq/YXuTaBNqSyFVu9ZnMvr4vCV4U
svSbV7j58gdTuio79qHBQWpr5k4tGRiQzNQHQ8x74KAqGQs8HtBdxY6SIWDaKL2CgUWkLeJHQMPN
H03btnxCMbhjqaYqvJi1bMSyNMMBVR3wVghv6f1b2DxVH9xrci4yWNxTQnmGeIUCmy9HrxiC1/FR
njaw1N0DGGB6ySA6clJIvHe8RIKZHu4e4b/0yGJZG7ODT58+sGuW0D88+Ovz0DOBWUJyGqCIMoXk
cg/GW0ZDer8XtygBzbp7779tzDRctiGSOgvZzyDHhYbd9cgNOib1bbHzOMUjL4TL/9noMU30HDQs
Gi2p2UblRUHP6JvYimOchB3jmdPbDKfGaZF+BkNxlVIcilsA9KUSanFHES1qKoDynTgWSKQQVjsr
halEEFBqEmvL7vSSGDhmGmNhCpx9Vmp9cuFOxSE1Q2RoFin4tzLwNFL/+1M9LCCTYpOBq7vWok1S
fs4qfBp4vZHTL6bN8vk6wXT9MVqFCUGrafPhRzlE5CjbAwS+GbOPBOrnvSwSEXAnW+bqyOB4nZAx
oV/+Y45CroBMla0sObxWH7AnjBo26iD258P3DLs6HEAO9BlUoGTvwmVhVcJ6o+aplng1rMd+HyGU
PGj7+IYMPtVCGoGIv5O5UDd1oFQnTQP4/k5+yj/9ycJS8gg385kYD6jhztveJS1YWdpmeTlzVlJq
2IqMX8YmvJSiMEixDUZrVQMId1Kpn3kmyxq3cENci8UIrrvSoPjbQ7Mi8YoyO6U+OZuklm/mwqg4
1SjJ90EVbsn7zm0sBKPGGW8ytftAVv6S5fVoxrn59X56JuNxFQIqIzMV3DcGggc5U6RcS4EjucVK
tHutI1kGBPJ1zaqfINMFO7ENGdew7rkuHFCoM/YfoNJXSyGPyUQeMXtDJ/PpJah1ZCwfAvQB5xJM
76EkI+v7w+3dQVnFcrrGVHe3XByXNkdMLGUO52B3l6/pG1NS26KCkw2niscfH/HpG88Ir79yXyRV
ygxoGzPslJqgrTebzOfb+RMgB6KYshcZJJOVxtC/N0d1HxSJpo57y0Nmore2p0aMa7hicSHlQ3XQ
HseTIWxiFAGtdNsVQuRqeMvNDYy/OnIRCCgAczAieMrgV6OZpGbcxOyBs2zshPuO5ey+9uPIG2mH
m/uWa3gZzoT1FvUtH2drbFtEVTC6VqIHOQpAL3tsWUjdzPwFLbDSo8jSQqIhsczmSkuRP2rGjoif
85OnumM+EucStMriG/l0yNujwNB3zcFsb0ogqRQvRgsvV5EBCzLUimOb0KVICn1XplhfRQizokC6
9ydqleIDsWPdyXdx+RjgcWRvl1W6XjCjeNLn8Ujcu8BInzMnC6DIZasHPgO+gR0QAb0AQeLsbXBW
qqPLmOGmPlyb9h3OJzwzqBKSSZX6rxC3EFAuY6VKKGX1tRONCvbkpDhq7V78yrqmdPl4di4okWWA
OQ81AUHgI9v0Z99/E+/L4aFv53rhEo13V6xW8X315bPYnAfGl7VlVsoaX38rhr1smviUAtxmYzvn
pTmQ9GqUsWvQzbbbCN/oZN3DaY3mP04f6NtvfbmhwP5DpjDECmBaNXzBJ+6QKnTwprUfsZOqOVg2
3Eiy2m2HiQvicDAjn/V+9bbilyXE0/OerFsL2rTM9+tSJYPL1rfwmmbxTpM7qGk6rtpRrNzT+V7A
lCt+JtNyCY4kF3UtACDLb4nvI6DU6WO3orvs23VtzcWgc8UEcS3yZBIA8LwOv2cdZCn3pNOLCvtb
suQk6WK3naj7xtGtpfzgq3bk1tC6CCuNA/PF4Hsl1IUXTPA/+2y3roiy3famKVXdB2pTxfZK6cCS
KKWu29A6+4A8ikFTxSrT0mj8V6UOhE9LFyWyItWT1FsWuordJzW7wpu3mYBIW/BmLbZb6+GfA0NO
W9RJlS2iNB6+mHZgyxvX9KG8Sef0/6XNR6af021UXP2dapVT/C1e4XJO85YrXQgBShuzMy4DkIN9
jcZFD1FhX4jHjSpQaC5n5Ga3tgcQUl3okMJxGByRUthd7LBAjbttPm//AjJIOqw8garT73tcYjni
Fx4hGXIvJ0OlwoceYAIrvfFpsU33PdqJ1nQyyiMQ0O9zWb0zClAmKgmZeZJ5DS91ENcEnGEgJD/6
66y92fhvFtlJKBln5ywB4UR2gGeJ6Q9Wbanb9U8ePkX81OkMCeEtLT22oeRHYe+7jvukoPpqClhF
cPkufV3XU7ET65BEk1Z00ih+rTzk0xljfArzWCUyfBe5lPyEiKshuJ4zeyw+tkpkDW9HJgMye18F
4BQ23T9BbQ1RblH8yGzB8DvBcPlPYUX8KZaybIv9XzPof30HoIy69UB0awebJLo83whYMyJ0YGoZ
/Rw0Z3EV0637FERuQUY82rRoV3WE6MLBoh6952kWGbhRRt+nLs4ImKLM3P2wwpazGY0Ksn/bhi2O
xZhksQjUwq4a3YyEABWCKMKbU2GdLejNlb3S2yFFysCWAujFfDuTslISd0uZuT3qjoq0+olHne+j
WboiAzbUSsd0RtjIGQj/8ygnuAavKpk1+jo9MERbWsmAOFLwBUyLrXqRnyVMqFelUcbF7jQxya1y
M5G+g7W615TA9wJZk9+Hr9KjeIrXHT+JdQ+u5aOMoyA3SipS7AVq/5lrogKwROKiSXh8f90Z5zQp
RGbF3/0tMwQ8NlMKk+7zHcgmRd+q4clWCSGQZ0fZ9jw508hO7q9oShoi1/3HHzsAWj+k9bZV2HRD
BkSA18LPEJ7wP5lbc2xvHnulQxaGvoAeS/Y3mZGcBvhsByA3VzEW6e3icOBQGyUCLZawHSM0ihBD
ssN31Sq4/m0hTvUlg6lLTJkDaM++5zO4y4yCQUFALXX7jrG9IklTPmCGGaQc81GWlHKdTlPmjUl+
ZmauuJ4vZoqgTGQ7JqloyMDQlQWXqbT4N8rLs3HwxlOzmxF9hR5bo7fPkcjyav6t5dbeKJ5eHO+7
Q1GahuI4PMK+/BPkybz1SGeTlUyunHPDtiFeqcj50YfVh0nRHT5I3unRSS5D3Mr7ZxwaKG/XGbj9
pwBrXuWb7CvH3H4l9HfBlsYMoYxvG4vOXN2TkaeX5HzuCxyPj7QaEXZiwsD/EmOWmJ2FIGKWSPu6
NjdtgG0B0qCygUatPPyVJDrTGanCA+Xp5u/CzpcnmHJjChLdcut1qIx1mzFfTSy2QRoH0hSK5JSg
hlDAYfIHTda5/AFP1YiwLxd6mVtbs8lQr9M2Oi99HruPvMJVuk1HLE7t8r3mG5A1SlT/ik4R7ErD
88r0JEVF3dVT9KmUP3oN+ap6V4eURANulGLK48Bt4vyFWd2UN2/L0eR2y0NG0nHsW8j9WboWFTXi
3SDZHDaPczbqf56SoPNUaVeCV+y/8WBSA7VLRn4yQK0+3NJnaDOjB6CklXVbA4YMRZzlSaH1tTOS
aKXQv7Cg7SZ7WylGpRrJEO3yzL4IfKHXzW7VjUPlYqopDiD0RELsAJnP+Z6RBxGRvhiL9+QP1W5n
VaaMakXoWOnldy/u2uO2/+RCidiA6kGe8V4FeY5BdBUfyNhOdPF4G/zGbcx+fruZwhALy1EvIfbm
nnBeWyUm/h7lmshZs/sahvOVvLt0No+3yJMc/AfW0O6Wpyr8uksQDIgmlJ5P0YAtXeFkw+UaYrJK
/jb3DnlgsBXJFaEV/gwmFuIxGjQnQx+ss4dxg2mA9/aWsheohdqbWLLP/pvMvS0Ay3ceGPXodh6r
zPJhr2UtxyEdQTx/GMB8XaS5QGq7aFgEz9In716kOIpOB/3HiqYvV/wD/84ZyrW/IDd3yP087e9p
wFJ107voXKDmDO8ud3iuLKmBqrbFBwqa4CPqiRda7q0Yg2755iDYuqU+uu4XZD1cBYih0jkJYY33
d5lDrmze
`protect end_protected
