-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
w605iD8n5SP+mI+gv+67iPZ9vg2RGRP7ZQBydQ1KXtukq1kqAAfL2WDJiQ4BHrHR/QmFNZpCBtfW
bNfdSRQOpxggtSj4M82/Is5W2O77v61wic7hRSNCJa65YRba5YxkjUo+UYim4IQ+aKlCFaZSGyM2
PHIcP26Zdg6iz3/A5U4Frh2x9DzYbsHHEk1g8UXs77kJGPpIaKzxagdeTKOFWhi0FED+9SvLzYU6
R3tOO21zk3Y0hTk5QLUYDbX9evkOAjQLgv6GKuPLOnpwI7TCysQp+dFIEND+Df1Vp2/tKu2C6+tS
mYby2FSfoJpXImIVtI7Ic3M0zdAGqRrvBVf4iQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8848)
`protect data_block
8hYc1nDhGYdJ7I11a6c/vtC2TTNesIDkLnwlEbahmIOWzOEmH61wzt/BAzstHu6NthkFd2UfjrRI
UZaCa640FgE9DVbkeNUYhkbUw3K2FrFFXOc91pRS8KugNobS66PlLih/ceP91hEsGRv2HgGrbrFE
m8oJZYjWIezFm8sbzV9/3318l8dAMOBs64XtCqhJfSezEwPDkKd/cwFrz6Yo2M+tJkIKzsJSBq8M
zuLjvK5c5p1uQj/X8F5sX83aurm3pFdwEwWhiNkyzHfJCIvdmztJMSHyXbWPjf+tHcG5NO8xiv9P
33N253mu5yTiuE/LowXMp2yiQPxFQJQkUZIGbEbcHY5Z1OQLLEgeET/8ns03Qaxf7UK2RzZHcDC2
Rm3uI/ga46OP/u5rHyOJu5NeHpEN57b4/eTpeV/fJghn9zWUaOJE79dYIW6GrJKmqhXubmeGpFRF
PtlkLzoipnGFqeP7QTvrzdfYxkB5jCwoTDlFgbYyaXWMhXbeZ6yAUOU5eNhLteyepeM+e4mW3Lla
pSrq6drtLBS6WKw4azqtuoIku+d9B9mCZInXkh0XYrEvgaD3SURGgQKXDTbXlATeAst7Xha7L4f0
UZbO5w5BaOogCZ1gD92f7sZoJ9NH/3mm4KB+QVbZQrG/mTFJ4FSw2SdXOwRxXw/JePpigOtLCmLl
MQE1Y72hur0uk8wMYJ7PtcAiMBKGjOpnm8Te5VkkCJOB1M7VXo8j8hGu9Yf/AL0gAuKwj0b26Nea
s7rW3BnloVGpqvmlkISzC4eexHXNQ6ayopUXpmEMH8CCDmJy3Mq1Z0VtiCH32pZn+JExZQ0GdvRP
AA6ajsAGpbr1eJxGv3WOKWGmxKBtyaf62106vb8BbcF2aI+w3LMaoUkY+XBtYBR1mpRJJYBUbHQi
YkmVhcAa0NVAsCB93FyeIbS0HGVsaMmTyueeQqTY0n86njtkjSu98bhlr5O/0/gnOmFHRKlc2cXz
PT5Hq8sVTCdLwRnkwBjymdIzGw7HcvU7332zYqX90oXOK+T0GPxMjLMV/ida/sGzapCprkb5HcmS
4cmirNgG0ciQlKzFyRbiCPe26c7ZDCbnvS8GNlPItbaLCWXS5wtBaFTikYrxu+AG7U7S+aLr3IIy
GmYpYGYZ4K1XUQnD5T4BOGLI5Kv4HBq2olyicldUbOyySkvUKYGmjULu79A7i0XG/wh/jF70ZujW
jZFtso/pJMtFOtVtgOlnO0tyMjtq8GvcR+2pmDkqOTLv/lJG4+jrncF0Je7wQJnzW+dZ5WVGii3z
R4FGYxDAY5CkFsDvMjjO+/riPMAiFuDxGS/0yJ0TtpGEGAkgLGsuI024DFihYvkuJOYaBCVBo4iH
O0kwBgLf8RcEPu37qOthZ7SMSF3UBvx4UbRUlni/47OhxvtJos9cmv5fFlvHcEDxEE7pKeJRkL1f
6B4olx0pDKzgqW/mV7JcMbTnP1P1NfTlK4LeM0nSgRkfb6sZh6233a/yMo+uxEJlfu+h7E3x6PPT
e+rECP1f6KBlUvqesBH685EL7KPrPZ5vqQt8ZPfthdEJyQCKD0Kj8CYEy4ApEv02B5lWZxoSDFtq
qKBAP9SxBD184aRL2g4xmiMxb+Mg7QMXk4XH2fbmyT8Sprhww8E3mFZs5zUtGDaC2v4a1RR7ZjF3
Ez6xZfvLeSL/Of8/KrAmy9KbUW0uM/M8qyDqtOk/4pqnbkTa2av3aAYXw5dRCaP3PEh2V+MDKpH6
f0H/6yhrLddXPV6rpB+KQ1WtUK0fGqSiSxe20fkm+OosQDnr9eXnnk3tiSt/uMlp909cmB1+TQQR
szJq3LShxx8fZHW2HPNLkci0yX/CbVp5ZqdZ6nWiTUhAgDaCZazd49F+Fs1flJGHZVBqSr6VtE+W
+n/eG722AkdsCO24xapjSSOifdsDb+gcNlJ5S2qLIqAN11X/v9bER/I8Y+Ji7WI7eubcWsDHDwq/
1lP/LwvYJNLR2QIrovA8iGjYbDai85FQyfJIrMw5Z9kV1ot4JILhcB21tJRjRSbIdFelq9cH61EP
pOyw5zgJUyKWR4VLWoiP2Yg7ZWWAJ+YD0jgO8F7HU7pjgaZdUtXruDS9FgaHsKcDregp8z5ZWirN
mphJIJ+lNIQiFUOO/1dOgULIi3sxXChAQQDc3JCuI3N0ax6lcFoOEn6PXco/EyBsAyE9G64UJp+h
eFIDnFcCW4L3ZpuODUuWXjMdu3Q1fe2anKqoJvvRoOibKGxhn0QnTaNXIy4CNNLOENv1i0Fc97OV
vKJj3SRu+A7jn/nnKRkuiKMYpEKM383I7HVr5JwIYo2sZ2vlNf8rkcw3QQb1M1tRgfkFktwVPH3g
V3fTzu0RlZjpAbs2sAp+6nGFGtE9iVEBdLk/+NGBK7ck2P+YKWjaeE7XGV9x1V1r6H8xBSbQOqdL
1aF1JYiZA6zOUknJCCVIz3+t5xQgqvEvtpwJWa8pMag70OIuje82lYugfePm04jZGl0g1qAw1Vtg
fAaeM9VQYNzS+0vspKYJcdqGiUvQaprMzDN4qtSvEMiLyUrv7grLkhhX/VFXVj4TiDREB9802Aof
6Mwsa5Gb6wwseUD9Z2d3H+jm+a5OrnX3w3Dx57dy/PEbPkFGy4yPKlnKI/zqKlKu/qv2jNIaOC32
DqFQHeQM1ZGxbR1rNBpQZmOPRAm/q/EfSGFm8hYuiKCM+Kcodoh9rJfLp46kYKEIHgBzsKrhoDkX
mpJN8Y+y95BCtr/sk47nvc1jASJOa74eGtxJ9giUwEpPNsx5LAwE3w8jqP9TH5tnIhIA5N0i6rut
XaPM268HXOJmAT0c8v6CMGprnrqS4+O28HhyNH9c8pdaf6I7HAhP10in/VAbU0ZhjhGrVPZIyN++
59GpPCZfqbsDP0rzasMA38VpVlXyrjTR0dTRWJr03zCVwxFa82QqunnWquDoEmBgOxSln8rG8GQD
y/yuv8uu6MoRjCMs9GH7gI9n9Lw7MugaoVGUvyN9oYt6T0DGA+P/eMhEBVK7CxNXRYYXJE3jvFyM
nFbGNXBQP53uZYyRXkblcw9+jJ4e1vPYLugHjLyIh993TxZDZdcBtUpa5sdHmk76WGKM9Ucjk7kG
sXJjtLVg4p5xMmRQqItVO+8t/tNquDU3O2bwX1NUI787CG1EV9YzWRhOYxJCunJMAyI1RfL6gk9a
VpR1tB2DSYhEiPv3GlE2jzk2zXtIT+gETV3FDwOUYQjFLuekIVELZr2JIu/kw42X2VhrgEiupqmW
R/YtHMRN5DEEETlgwMRLF5nlD5qe23W3c4bsAmooB2M6Y7IzK2BvBfObbpHzobYybGJspEo5XuNl
t58KZYStsggpW5twKhzl0cVQydG5CTBtmd5L6HkeqEAu5KKd4vN26AUq6wCw65LFGed9NlkorqcI
7wki2zoDOhkWyvEBi+gShaZR0QH0yi+FmR9ioYl1gHUXiVB85jgo7HRvQN52H1ytG4/1CDS8xS66
4ET+g1YQgrsp3ebJbSH3URzfBBHdMKignUZH6l0J2dZWZErDMt/tXBd8USiKbBbCHZCXKArm74T+
iESMbhQx0L0ffB43SsvgsVfY0B5cg5TZb9jbUG8yCk3S66k8LB9+iLzXRNe1wLm5roqFS4Yk2HP5
GIJKtToE2sJVmr362yrJXZ6PoYDa3Ks5qUJht5OQAhoq8eXLgl8hASmOT8yzoazJ17aZe4f8VmI4
DKUZUTmhkykRiQ4keaZTIW84OKO85Spgn344L9XCwcrIJUaSzkkK+eyOtG4YEmbvbgBkC+RqqYM/
F16MZeG3KZJwI4qMxRAwg5ur/kvuj2f+MVItXx+iJRwZT8pih6fchm35kfVGNyJcwsk/fJ4g4uoe
G37sc3CWhdPRw1d5bCrpp4BKKiDhNJ2rjlXkWrNg4b65VH52OscnsGSxVBih2BEuUfdutCcpAD/m
pENLa3sFn2FVuk8Rqzw97zk7oQNy0D8IuPslYlE1/hHtr6Iz75/Y++cGpXv4Ixeq7cxgikZqqD38
T11cwRDTaXrxQ7SIWDrFeSenaWkaQEM9r4C2VMrySV+kW+tMVmnM9IBq5/uKVi4l0gOUA/ZzEb6J
qjuDlG3eZzGl/cI6gmG26+7D7WHU4l7+TWiV8LecAfOcp8f9wwtfuOeXC1pLGKQvuZpXxVmMk9Lx
MJaD2wBFbvLHz3l8UD85Zjdfj9cTxcxaJ9j3kNLsUmVELkIh7RIB9sMnQUxT9xpD8V0/m3mWDymB
pI1Kv6vq0U5+RY6DZ9CoCz16S2rz5lzt0mJvQogNefpCDB81ao0dMvNsrZgV6eFVnlEBO4Be6BoY
gKGdbxaaFgBM8QOpuo4glbtdKALYNLnt7H3WfnIiu0yG5LuvP1E3ZEEuK/Pe6Zc3Tugn3XibYUW0
Smr6q+9hTxhgGNF/xdlQuMAFX61G9DuizA4Js3+kLCzcnTS2hXX1KFeFiHOj0slKuVkzx2AYuwwQ
AuEGE/kFue82YUy46WPfHpP6vOWiS3v7qpgdTeAHEOC/qiKwgXApgsYtddUJ+AGzBC6MW5S/HELE
9YQNOCiXpiiqlyT3ERNhF0VwR79LrO+WnBkmBxbr0KLQPtRX5/ClbDszJ0oxnZjaVYQ4RTJuY4qQ
6SNlrawz3aYV93TGARV1EJJpdEELVwy6+o1/Rk2kAZGVtUl90+Bmu4QX6jDBKp/GacatKr9bZdjY
Ijfm99BlkjVqvFgbbEKRQCei+U/3wLjwQOUrDp6/PGvIxvMhyjpKh26Uw/Jc2+hYgVgiApwyNREP
szQPgF4LRyGkbLk8+AecycCJv56zqMAEWmBzOZ52mKCgMBYFNR4Rh4yvLjlwkPFKOxXEkTIw3esF
WHSWljEhzrvuDL4X76xtJJgfiVH7Uxf2RzdaPxh/4zSipZahJMXz3u20PaQmUjHO4dkMIrKb49fn
dw0fMKdkZrNabZ4nhcEzLFkVwxfSinDH6kjAZXZditIOrHhVdlMvPHcjWFRRo9N4D0d4K6o2Emga
yD8BV2XXe9lDbOOO0FJ6i58Rn4P3w4CXYQ6e/lAjQD+bcLrnqoVFsUhMScQbioLCboUzoe0htoYn
o/smA5IkR7YGycINLtYc134O7D+ClXRV6vU/RMnXsJsMNNWerOzBsykHtq2nUG9QHDV37XFr1/wd
M+sY79aWoek5p3ozYx3iPXQ93g01izo/ds7LlreuXSHAdVNxBpx9sUJsbEYmE0R1TaPWpjomlOUB
Fd0jmNZjf13CaXP4hwctz+QwYbxj+DTSRvrPv0ryuDps43bgMXldcyJDlko32473ZgdjjGhR+cs5
eXZU/rM5w+oksMz2RpIA1XEs/zIV35hlDkoKVZucte2GedvSWfK7IkLmq23RH95Yw87/n57czGrZ
Nt5QICAiYCdAN6V47AlWWjZ+SknC/DQtVvnupYAe/t+p++5Wy00gdcI8i7vNlIoDEb1s6D4JREMh
pqmrfmaO7Xw1+2DAeAjGzyKKAxOg5HUcBRRU86xXhRqL7EkXvn6M30gzDDLNedsDRsP2iihr9d/X
xMS7vHn1EBMyYWj/dWHTkKJss32VTHGV5kO1Svp/rJhjJm4Gu2NskPZaY4PYcL9ZlEy2JFJ0Saxc
gUOHxFU6125XdcJql8ayDRCzZPPQEYUiyAMEZys1rV4fGWrs1n4Vgmho/Up38cWPvb7V6TBKE3vd
G9LYNlxHfHqk14mnl7AxO+QZ5s6puzlrnY3N6PAzPxDp8UtpKBHNTrdL7GRqmr3XSYkerYGuP+lm
/Q1F5j8QsGQ4TlgAIDEEkmC5cYhtjpVDru0VUtN1jARsLvFJkI2SZt5kksto7Qp38tX8RHgzpbH1
aZjVm43ZxbIBONaUTP1OKNFQ+bCVeJUOLW5nwe0cuSN4HNLFEsUWzUDaF5/kivRtm1sRpRSSFbaK
FFy6yQFGUlLYF3UhVjq13DvDAUc7i6AS6wwTCQoLRojRmqeiMxm2HSjsZjHKh1TycEO4KXAhsnnD
09SoYAYqr+IgshuVE7a3+R/afaupLzK4qf5qcAH4rmds0zTZ6mRFDMZn+yTGLlW6jo1rV82QKz6p
9p/NKeozNrgsscGPOwrpKD4h7B4b30FIi9kOPTRSi401ZJkXuqn6/5g6c2jftzDNShjHsQ6ijTWV
3rSZRUGewb3zPNNEEPnjkagEapZ3+DKY1Y6COjOyRzzj63SbJvEhWaJsExBAXzRKw0a/LjdQPREE
VYqEr5mz1OCfOQrZl0DgfFJPE3TR6W/c4vWjCc8Duz5wcxUWDXqMaPdVZuHn6iCZn0aObQN+3v8O
Ud0z+zXt5h3Q9tvmmL3cdtV9e6j1mfo3n4GtlTMXbZUk3tLSnRIuyiyjJUhBNaxlvo9Zib1Bon7G
DZNGgdtvJcwOyoIQN3cBq0p/kUZ/hYywk4t/JYt4Nv9cLI6pb8nmEXCv6D5PSQeIFnPK6HUJ8fim
Dv1N0RNYZj4KaU4nr9ZNT1B+WhedxC03nemOJUFlx4CbAohUhQ+vPERVnWo63GNmtQW0WY6aU5p1
CeBML/cPgOEZF6hFAsWTN/srD7kIrsiF7983UMXMb8lASXFsH8afcSoeh7rrGDMOwCLX3OeymmOu
8JsL9Uu8BFUJ18esX41DPnsmTgKAE7bd/rPpUlkiT6XDDkCKBflOIs6asu7XzOhytNUmLkgzwjqz
Fjf1FcvHP373T7XbS19/q4xZFd2mU7v2PsHlw3UjnVizxLIxc1C54/aOKT14bbU59byqq9obVy5k
OkZwF5fCrGW9uzo2wqoIsr1a/BWh5e5gxFo17VCyBKyMoGFSP/l48BdChK5D09idxohhBUaJ5AZL
3X8Wi7lTW3ffjzYgQIK4v9HcWfzA/OiXzyKtmzGUokNAXSDkFQxbSfeGuY/3jci2ANXrrvwfVP0E
mxLnNBAT38wtimkgRAhjmAWilbzA9fzCWeBZUoVYyDTXGjj2Mob38VlY7KZfiG2DrHb9UuzkRuTu
LsRI9DO0EGbIg61FULVx0oSOBuNhv9ag2YCg4ezqI/5+ZurV5RHtcyDaVN/qKD4Ez82R3dNPwBAo
QCo6RqNeF6ZRzXqRe7YxRf7MYQjsT/QxsoeUox7i3LZfZ9xTc7mGd9Bv4yd6WKoJduf/gfi2QN3O
N0wmA0QxZIWhIox9Lvwa/JVUg6iSNwvszk6bhdT3TJ2KGHAT/+g8uLCGGoPi3+WtpE/bEmhLBkir
N7jqvzunwXNdJ46N8h8qS3Bl+b0kBSncZ/oMR/YizW4gluLOGDfBDapqERe25Ck1h7v83lvigBjs
AA4906lsKYFzIa6XY2p2o7b8sWoWU8wawSES6zGfdVb0swXBeji9qBVc+z23FB907meiqPTpahyq
KfPj3Z9a3wh7GZCuV2J3oqNtD+65BfUIKWcz7CgGkSTxB86IUgrqmhdCtf66eJUpnI6vcvyzMEks
i2W4MlC1Xq22P6Scxh9XFIFv0lDbIF2+wDc/kVQtcAXapaJ8B7l2pxjwpXdCkFh+7FUzBdYf5Wsf
OfSVWBUZLdvB58TXsvR+5diIe+W41hscghcN37ZXP50UI7ObgTXtalauI+RBymvgRU1XqXKTdnd3
JE6OgcAcAV/2fmw6FsfwVWbUor8Gwt/ii/b6whrVIUVQbCLa5zwT/oBLVqeZnIjhTTnMrjWbbwtT
UFq2M9zhPVQT6VZISn1JC4kMXViR9ixsehSdgUrDqFbFoTY3KZdgGyJTiya+9Pvu/OIvAoWZXs8b
93rtoB+mpa0xpozqZWP9jQzP6VKTD5VRqO4eDYA0rYDusyV7lARnfW3/EU0Ig5NUf4yJDo8+bkL3
0bEJFB1u7qb61MWmDy1175SrdsWhXz0oMnBgBDhpO4yAeHdTVackjDo+Uu1vO+S0LO76qlsF29bE
MomS6MB76Kq+Na2MMq8PUcWU1BbROhtN/uFzTIr+twqUX7NnjKp4Svq1NkOnvbvq8we5163T4yvP
u1AMwLWzK9X3zPFZmKyXTA07zcRhUPrUz7hK/Fj2iwLmWXQvyEROY5mEers4Hr2tb9yXDjUYWqiu
A/4vbEe7zhz5+1P10f6K4eUsUDdiS5MWvbZvvyVA1kZj3uGWC/aoIWkOjmp8rnOddWWAi8Xhk5DG
zZgxFLS65sqjoN0xMFum/7sywVvD1lKj4MoTrzOSrR7Q66dbN+6vD6nr3T99WNtkBY8l2bGuu2fN
y3nSFHOwskzpzPKGbeqJEofLdo1YKi06ck1M/E2eX+suxFWsOg0mOPHI4H9bx+8dGrol0E9T6JGy
Q2xgD93RGtPy9PKmI8JTL4Z5qYto71RmcnLtCZdu/3GjN/0mT5T2aZjPX6W0ErB20Zndbfovdv6C
NGCbPRIrCZo3mTZsHnMDoXDwYSV95qco5ZKdo28X+XBn+ci/9HMB53UCHMNeZ96yWigBQOBvGMj5
tJWZpDx90mSi7ewOONXigEIdRFLtCyEPhunZmJMZ3JRO+1dDAW2aLf5oaJzn5x7Z86ueZ+dLyBDm
Kf/URXnzZuQ1xdoMRiolr2LspZ0f9lzdQnDiG1w1l9cjOuLzuIb/AMQGkS/qUEg6Y9IXCyfUfzDl
yJRLruJh5IK2K7fhDOODNmxaF/I/rue95LEm778GqtpoEYQDwJH90py13SqEvx3XhnhAbPf6TcNU
vtMDD36wBb++MhCR61g7RMr1YYQxBAxEhMMU7pIAVPf8U7R+KuxNJJy2FTB1aDy0LpAxM633b09D
eHr2dbQSZu7D8tO01dhQqFmF1hGWcsCcPuB7Mct5mT3+vrML33kTd7ctrlIniWtVb7FT3tCWhz35
oZe4VC8+NYBXl0L47zlUeiU7bbbxUrIfPBEMwKDqVB0cA8nlxuTkZCu5hhykxtQ6PTyUj3fCPO6Q
hxdxqpFRLzSSiKXy4Xh1C+QpLZnKo4BXIdAam7YxQFZ0og5WiOGO/cn9uFp4q1IvWaHhS/IzrEWZ
zU3FiAy/pmI2ep9vSNpiagttYUU2S6DF3NnyEnoYjlCi7foUVapMLor4N7CXocI+tVVL9hPAHcJT
4gMgPc0m3jT8JKKOfofSMVtUyvtaQhTqwTSQdDkaz84IDQFccztTgKTQidLeX6ilA6raFVI4K+uN
g8y9CK4x1f1Qb0XUmGmnl6aEWlEtNDNFhRk00XIZMNhKTFNuJs2Mv0wJ9xcjAHl87fnNFlwI+Xde
ihpDWbglphdlCVodsJn/YxEXxcBYJd6z/mAGpKM50GRafkqREg1WJaLtSIeiivjmXktn/GfsA/h1
T8tRdofmq1YzzHaSgIfkiQVUQ4goPs5g+rQ2NnR0iiYcJhB88+dr2NtWYoCek2r3YdVJb6Ic14+p
eN6sQuyvvL4E1g9C1Fui6sBgvouhucsWEds7LuVClnWY1JVYIlwa4AykgFuEa+Zhg/VEe/CK/VtD
w9XURL2DRwMDSki2hi92BfY9g/cukwbQ6CiXtFHXtjwN0vcjrg4mvKG1Wescy4+U8SQSdEnKvxzo
SIMitmXlN0WrYAt2gXzHgp3JaRXIA+9toePu0Drix4d3fhYdUUzhMDQ1yCwelZygvb+mxQCwrBD+
K4zOwPn0DrLAG5r6dIPpy1QoYNjH3McQnfT1NRkZvZJ97mTWqTTTNRmIkDvuG7rSzHx2uv2TIho7
jtIqKj13rR2fd7aiWo5gNqojsHEY2A0/zQWCwi3nn//oAy5mF+W4rYd7v8rRrhW3iFmcFAGvSwUj
qq12PseziSvoLB7OntE3dumm5KmOcda0ZE94tZAZC3PVtUI4wiQEF7bcX7yK0QVqDGep3iXzivzm
25GIOgpMmThG0JMfVw+BG6O6y1yIE4aoT73SY74Zu52zfocbZKSogzDt8IHrkAEPqEqvv7KuAQr9
ebzS49IoaQAVJUGixWDz2BYwYcdWx1SESSwcwL385YAPRkjdtU8TsOGVl9vm76s4oco/LsPCybq/
BhQ4vruYQJ7oJiGZes7IALX0P5Nf2xJOO2oSmkHrdNShwhxrVA6ulh27kImzQ+Rvcp/MLc4QLpBW
aT+6NggRBy+HBmx7/I8fOYb1Q+YQ5Qyid31oNt2BMDh+1UcRroa5zLrb39g7lD6zQ9hxWbWcplEX
cNKsu7bQpcLcET9sLZwOyPKWYMiUQaKMYKLSBBu3HRj1Yp+TD++LGXgAPgY7tFpcKm7S5qxyccxp
4RW3BLsrpH4w+1Hu2CcTGyFr2sHHJdDe+U/WV0hux8a8lPAAGZTx6oQ0RoiYAeAZLt/pHVq/QuNz
8JCmOM4Jrtv3oSebd/rTy61AZVFHLHP4bZBPe4Zbfp1O8A9wFrJ8J3UKSy15m6qVY8mUs0NM2bJi
JLrb5fl2NBftCJgWczp9azYD5Z8GgyG0SmjTlVYuvIavApgp0cPWaGjIuqeHRK2V5wh02GFaW6sK
o9q4dFQMHfEqcG5ahwCFe/e1fA1bjawQDaAggvnjyGang2TFVgRdw6WtL21ozWc22bI1KxR7Mt8/
4sdKIkCEoBtg333ZFpnanIMPzvoZl3gIIYVIkzYN/oFt6DLkz8Yi67KkEDljfggmTnSauyCchZ5c
XTPDeQv9SVOeWkQ/lfqmwRVCtfAthzJbTVqNpczMGE0iAFh+pZIbmx4e1braFn7H5sJtVeV3jG6w
neZljpmXWcwuW7HskUOCsg02hVMD5atz2UUIIo5+gklRY4ds2mieY7/yWFMd9I29+yrkh+zE8LKj
Dg+ll/WwV1wA8K2ghzmVBTscugicLP1s8dmeCQTyop3VMgeWx9Vt1SMAPYnPUUaaE7vH6Tr1h08X
8lfbl60kEIfylVLGf+z2HjnIyqTntRpEKS5EBps6imMdUeAUZJ3x0J8qPVQJ+dbKK4EaJXxjg/BW
TLiI6HLTbys0FFkWMOhkqWD4cc8ugn3u9uCVgQZzkP9EqoG+euZBqJa6DUfhWsycG9AUx1tQw6Wx
R4oaN/mg4vNZzyDHRT74uSEhgRNJslf0GeIABAuZEqLqLWQdhZI6I3UVXQ+xG2aYQWhmijr8LbCS
vwG+IsBu6rZkBv7BWQBHKPBuHws2SCr7cMcuGre+pYLoocEQ4Micd/VQuUP33Fl6ARuiQlrtvC3i
HJrG+GYQIao09eL8COVH6tWelO3RmHDzww0jHUp2FJrdj0Z2Q3BiQmxcWT3RDEXTdydXTng7vTxN
rSyHia6T8YVHipm+so0yvcIXGQP3iuxC87xwPrKnmaVzxpbrC9rejE7e1DfWGM9I1KDAHOmHlLHZ
N258y3NG8iD6vynCSXODQbXescWcE2lSXuURUlsnOuCn8RdlhRiCCZuv+JSV2QPt2crLKbXZJpu+
v0RRdW5RpjN8Im1W8zF/8VR7GRZXmlsMaaP2he56KOpT6FaZXG3Qa/AfqsaUtzhf7PNroDjYre2s
waQENQs8PVFJmbnbjD1OqedL4cVOzghCYQhaZat/EG97zrFWWAG6hrTn/Y+mQE7Oq8j5uXQt6kfc
wB6BWZP2XFW/j2OsTnU5tZbkgcJGeY5W8x4C11Egb+d2iOSSxH35ziMmWMIRBqlHWCbu8KZskcGe
vJsnHrlMf/qxm/PC02RyG22menLZ2aF/NIdiPUpenXf6g8KR+qhVMQylJH63u5SgL8EICd4o8jOT
8i9wSQiTQNZr5dyGOW75fURKLlQFXNhy6dpyj7v2f2RKT/UaIXjl6JG11XBJ6q33uWrsXQcnj0P+
ofTCOIHXcTiYebyRwtFDFUVrogo6MJuSUOA+b0C1VIJYBjX4zmgdi3qIIHX/ivtPahNzDgdNYPz5
gj3dhOFc1BcV2uyPyA==
`protect end_protected
