-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
WnddPBQBElZ1X8nCQ898JzbpUjOPbJ6WbpoD6cHqsCqrNYrymhTcy31lbbmevuYm
RNcS1taZul7sP904W8RHQ7xCx/Rwxz1U2NfanefFYRjIAkQTuWIe/TQICr61qAFt
Eb/TIiiphOYxkzeWx0t4TtoMr62pdFOFJ0Jdm9D029zLIo7Ma5th6A==
--pragma protect end_key_block
--pragma protect digest_block
y1N9JWhcjq+zn4YY2zEm8pqZm/k=
--pragma protect end_digest_block
--pragma protect data_block
8E9vvZQXlsKNSMHAYWIBNkKUAIELRFnvE3ppQMO/6NiL9vX496o5NqAo8okumAg5
Niy9hozKQNP2rnmj+4jfkR0bOhYkdY7e9tEX11yMaujdEKf5rdolkFhqgT66FoQ/
gMf7lbwX6O74J02wrgyX0n4j0ZRTXOY8HD3AI3S9BlOuntEDT76vdIxc9u6g4Q6C
tRYlcJb/gClI+Wh63gm/wKVNmCKlJH9j9vIeGNxXa8caF8qmkizy1XtorITUqmyT
DXuYM1kWDfpAMSPijNKEGuSq4750a234HPXwXnqXVx8uwTzuV213IVrKMTT6E8Na
hhI5YczCtMxquAwl/XDCBjWOWP9+pqeZpStd4TkP98u/JoG1IUM0SktQVpVbf7as
E6PAYPOv777nQWoZbaX/VQf7+3H+rr9ekbQVrhJVDDcFcMnxkpPKeGu7pCSbqqDw
mH9Ul6rgSEwYIrJ95Cgo6AcLptU+IK3OTbI9jiyjjcfZk+L9g/Rg46NKzvhhJwbH
ed9XZo4g+fRHjbk5Kf1e+q9gCLHy3oJjl32V1sDuYfWISfSvMDJVByoibJQBW8uG
4vtuFof5Cm5g8YZdgafAxy4sGcPzxr2syxCaVR1KqEhNdvngzDP8sJvuTcSQ8lpM
kcJ3YyxhzdVLWHjcTDeF6MY7MGi7uqNyOGlG70XD6/DfCAHoNkIImbAReohqKFNZ
HCKcU61pAFmuS1mswBRyNZb4mGQgzSD8VTN+7C5+K3NpiRFh2sTttVxWwQV4iINk
wOJU735IbnOy5xlqBBmgjjJpyHDgXbPyv7aDEVHoyFHo3Nq8esyJIq1QXtha0IpZ
WyqTptSoyYKVVksuQIDDd25bRYtSqddJb/SnvXYCN7ERQGSoDd9FKYH+23NKGR0S
iN0TfVn8D5nrLN2Xtgw+ayZuiJhFCchyqqJKGOXAvlZONyyfKCvgQ9vbIxwxD3F6
KkE4oq0a42icDvBhUoStU1tR09va2Bj9pMp9QledibuUyXvj2/w1HEALe2Io6AqW
cn4cOUXErFI0erVVX6o1DhLSMgQcFYzPdKDkwlBH1IB1qSKva0+VCQxvXaQVlbB2
8wenBibpZNld7iw/p+gBVtbZtZwf4Jpue0OsWGHUBWx1msD6VXs7P8aEAmmHoxbx
/FFTRm6Agdew2pFM9KFVrtIUUdzbgtba3e8nFgeGSgQi0hPaSgBm2ZvLLNqfSKdP
rMY7G03hDY53B0IwkkNsmYGZfbce65D/4Lncc2OMRbOXnX7xvqbnHOh68jkiaNIb
KITNgDZgeWtrr6nQ7qMSHp5iyVUtDu2a9IXFRyoX/6tMqnYbhOx0l6E+0vHNi6SF
SAH2wAbNs0epVME1GTL6Lzt/YNt6k/V2pOK6p5a3YfAskxe7u6ZnXb6tcLWV/Dz9
BH4NQUlZ1POA1rn2wydge/E0Cqm/ooCpHJKRtNpLD9zTnaIcrHjIVyQH9k9Z9rdO
aI6Wssb0dBSUmOOQmk+vSG2S8qEdAUyCrnLuHbMlMZF95qYEt+5zWLYoHs9XZlu6
4IELgYVTxhrE8o6kdoPAlSfyidK8lOWBBsJuWSoLVCki1r4mdhXtdop/ru0Ej6Z2
G8ZQgWftEtzr+ton9RKd5Z26TW/ytUlnAz/pNaNBE8fsT1JdeoEALR2zixm7ZyG7
TnXk/ogXh6gcYU3SMHfcgi7iQNBRY2nYhhomXpfg1ZWTeHORrtqQ8O214QFexDga
Xs8IOYmnnhfsvcR2dCchD48mRsLxIwocfvfkuece5oWFOaQcskGFs3UAPQ/9Nl6H
XBNgs7J75kXjc/15VtatyRCsqAfvg2hPc7rIVEzHLL3LmlxM8U6aid8KfiMJlC51
Bsw+jyboSJEygNR1pibqnbQS7q0hX1h5zKtVdR54MxOYWQUGKd+w3t9vDDvKF/N1
7ZIrXQEMVNZf2Fu+5SkErVRpTfN3BOMVfQOHkCaMVCzdD2ZwtlzoHj0RdDjPHJ3S
93HHzF/85UNzdMh2IQTY8mByeE3K65q4huMgKvbK6nwj/AOsZGitgTdtOFPXz5S2
/urPblAn+9/tmMnMoQrWxy1nFsEblR+Y0Ez7llTnsXx92eeEw/1w/S/mm6XtjQZi
dLbLZpc9NHi789FYpXGTHOFChS6O5zo3VrF5k8o+ZtQeclW4acs7Z8hF9TYvJ0MN
YI0RCchGhBk3Z1aw1gFd4jWnF2b5vm6Job7DdLRnU4R3WGVWLWNZ00/+rPmXLUfQ
cvnBNw7Gxo+khMIR4/bsKNN4el8LcmE3xoZ4eUgpmHd0hb4qkznNV2wr2jjVYBtV
hNS/NH9Om8Lp6/q2q3jHmh3H9V1onl2/GcKALM+9xyrUzNdVT2WgCrExkdtlnLSQ
tqotspLS6VC+8IAh7KV2XShLEp+iOSKO2wD+isrKZZDHIe4QEdIQabCNW7ekNMgA
UqgbLDs5u/T+Dp2PBoArgDJLf6AOuTcBm0e0wrTruZ9FPcpiRUZFfZxtihf1goIK
hs2OCFhQhexK6p3Ro7pRgBqPgDTyJR1i0FAhvExE5v0JjBlRPqqq5OL/1lf9I2Gu
5sYSE4tqjdmejGvNH8J8TQ9LwtQQ77XWYWBs83zMoKxHr7UB2j2NlLr8UOkoDXP9
1i9gO6T8gwCT45UHzZslsvVwWjEEOBclqUUsmr5Oow8rWC/+miIT6lIlqubXm6Qz
jl2G1i8OSqNsA5vm2YzJbvzzgjVop2bULwZMVKSlMjPdnpx0WusLs3fx+BEvgLag
DFozhbVE5RTAA87zkUWQgqcC8Kx1Dx3h8q/jBbaNH9YuEJd3e0ZptyUAgWSBMeya
/mIZQ2gZAjbkgfb2haeDcM7WDLzrGNurvJNn745WCdeJ9BdGi2ru9i2kj8eJs/rl
+OLk4gg0MCUxKgAAARk7ixt/bNgLSugiNI9H7aXQ8neoo5pPvourbIIwjSJtP+oZ
P9ubAOIEjai9KXiUEiXfYxsxLUDkqoC2TWyidE0BlbgASySIHnCxkSlAM+GlGkp0
u/1htbRJKbzRV9FF4Hs5hBVb50T8UED9Mc6si6EDV7wG+/Lq7UrNfGpohU6cZ8lq
NhmjBvbXO1Rq04JIvqx6EA2NTq+HgPYDjd4VMiRRsZB+KjVeD7gYhCTHTGvEjc22
uF7IHq0KCKMtPPum6FHx77uNMUdkCUAgb3+QyJ3V24DQLRLJCHL7Gpspo2SxGYsp
r4iD8w1bbUSZz1CgfM19GRlLr/scVGpFDbDQ0qGEBg/xTGQsB9/SfTUQRFZjmN/V
hQ88SeoT3JZDvv1KZ7Fepu+vYDR4f+5A8/Y4KlyhPfbiVzg8/XW7t/69gzmcb10Z
vuueyFy8oSnRmhwH3pIOB3spZFj0v7LGJXL5nR3n87me9XCgkdISb5wqURK089+B
3SlgQBeJuUkX5f81YGRquvZK04ro0Orzr+pSeH7WbLEKaFeJv3q0LOBNLjViD1m7
8E62cSqSV8pww12Hxhsd1GIK4bjVt7USeu8a33At6J0FmxYrYyYrd92feBr78D7i
Q3RfnysleJPPWfgSyktlAq2QyqtwKXMWkPv0OVZgjDaCoUcDOg5ICiWi2BavZHiE
zq7/6VaYvfTVyrHtOkMUWK60zw3EOkI+4K9Sx1v/ihnkjRhyUdpAZ4e44GYoPa4p
9TIRmkRLQ5r3ujcT5G1JZOc0a5jERVtol+K/F1lVX/jkh+wSrj5MbrF3llYE3vII
BdgtpHul8iqLDCZVrEYBlfA/kElJkJO/KNMyXVnwyZ6GkOU1K8mRafvXCQ/X2KTw
XROWsXFq6uJV3rIYCIo1djdEEqXS/yRovGSE2MLsBQ3ZAipkEnxaMt5KSkptKyd6
E71Igy+oEg6iF36a46EqQ8tsge89smofubf8/BgkMXh0BePkx4vNZMDgb/9XeF0w
kFzqB9k73yaD5wFdr9iL5dy5DDB5QE0DqdO+7ZOm6Da8CenzZ1sqQBSz6zlC9XPK
eGSxiKLn4mrPNIkHCJ+SsFxCTWsZAzNOf8Rc7H3ZFsobVQ5O/ckNvZ6hKz0rNgM0
S2wGwEjvVo+pJCWiFWG+odHfKQCcf2L/zgS0Z5KVYq85YP1YAwF1ryLggK5kGd3g
Szyq0A4zc8s873ohNYE7fp27DNvfbykZbyYsHNRMpFpvweXp1SglOujWncu6HclH
1+nm8Iuwi1tZQsNZknACxVBL1nWytIWwuMdryRYvKuV+Ay2WNuzAGwQiVJ/A8E68
wMSjni47wiF58z/JNsrTT2wmHs1KhRSa9Xt6FaabCiWH6wFJyNurt3K6lBaqxbYv
hzfNx8zuy+D4NMsnytmxs0029/Pd0aBB1+Xil65ySPW8w9CHGT8TtC35vy/lDAD1
ops+chfXUwbjz2XDW7EXDyYeLtFkawhxyjap5Pwb9SjwrIuFdpIps1UfKzBM9kpz
rOEyQl5XveNrOf9fSq87TIt8Cc2aeixAlQuNRd4T2LJNzCx/A6KfY1LOWLXY2A0J
o7qV6Geo/rHrdGColIWuJMDRdHo4RDO41nug4g7GbjR1lhp7z9gfLXY0L814kcGh
Wsf6YdWKkTiMnSNQm4uBleEPhY8jEOp5zgUcM0Qvd15xb/AD15ArBxbKUJOho37d
K15FXAnDNKjVRgDFyB5U3Ji5+/uOixv/FVHievorr6HAADWL0Ee9a5HipNWG+BEI
ZT1jGIIQZaMEeGlmLUV1KuBDLfl+yjWBzg2JmDwHxWfkucyoAmW6T3KgvDTNxSgZ
d+VRzGGlFQEBPRNaWejLMSo/896W6SHI+aqAoa7swsWjsvoH1c9hS3yx/ubzjFt1
koQpysKGtpC+HWTPguGnO9RuED/PVRKUplTmUTohzza50/anJv42gFmENoBYIeZs
XQlWmS7XykOOk/s5UHuJPh/xE1XjwsqzEFLZ+/HYwZAQuwZMdXQwKUv6i8MG7dBY
9uW/1vBvwnBOb9Iu3jp18pj5cthnnZGF67+Gc3bj/tpK4G0Zu7ZRTgDZ7o6SjiW4
7Ih4xrdnAMwhnWJ3nl6TyonkUNHfvgwwLM6XKpFH1zy0QDo+TR63uI5LZz1yDdO7
UHTMzB1L0TNmHoO0cPGvu0LEwjLFthUkwQcDugYMO+K8l2d/Ge3+hijQzMmIaJY2
BltmYUYFvFCZQJppjwT0L4TmlJl2sN4N0ahXOh2fMYMv8npya+vlQD0ZfARUi8HZ
GrjP0+uAG4moswzugYvULTOGMcfXhvy29FTR6ChAHjYXfKs3VOcJwV3N/ZU5Qd96
/Yg9zNM2LL7BTxAa73soxgulohEmYqzy9r1gyQhvDYyWPjS3U4qlIf8xyyZvwZBv
UyE2gAQIhvZ1c9/0OR0ZzTOSgasu9HskFGTXjxZdE+MopUiPcZkwJy85hRWJ9qba
cs98BYrJAPbhwUR3DNkN6/HZjScgnBf6xK9fMVleM6dr+vYHnTj1On4JNBNiEwrY
MRE1TrQKPNVg+iv5Fin1srQ8t9tZkZ1scGV9UA1KHrKnI2N74GjsbP10gnm4LKu3
xpIrxdPffqvUCXqETe4V062YFNVoRo9wais6oXYAqCVqIAvgggqJMBif3nXJpkJT
BTgT8j3AqIOgt7lck2Lqd9QDOWGE87Laqz5BzZ2weF8BbQSjl0K7HyJ/txjIBjGs
HSydWILT8sh8kv02FWyml7knaR4oOu7Dqf/rYVbn03VhpQiQND0V0XuqGgg1gir4
s0yeYTmIeyV9aYt7/ObKbAYTQ/p6kU3wJYmSPOnaHhYmsp4+MHZ6FwEoAk+lY3ij
EGbup36aG7TVJMa4ne28i0pP6csube/SLVUxMdu323vSNEvhCJY+MW41s7ERm4kH
x0eUROFcoS+cS6Dna7x0vqz9l0xyBaNvhTSaNCXMhPZqxTflBru/zG+NlJDVXcTP
DZqWSh5GEKXSIKUj+EIxW3/MqqONWYoEf740MTU198a4kHQkIeh4MVC/qXzEtwBA
DBWz1qiEJQAOOUiQVOi1D5R4+8gev1Z94FAQEfPJfJaA9EhAqQBHXzoQFNhnEWKl
iuG5uWqsLXHN7XxuJ3xIPNmsIUBf226ohN4So0hEG3ZA70xSRbVjrqR/NsCF5dDw
ho4nhNTFkG+pLLLB7d8qN5aUD8LEUcI7uJW8V0Si92fQaPW8/5FKuIpvg6GUrZjp
xTAaN1nYBFQ1KkBsThVpeeTr0rJ1q5la6rLnWa9+kbLE8bPMLukloGQRR3RtZLS7
YrLyYkm1PdWyqRwMrxWuN8HaZgP/R8O9/mdjZibsbFKvBnFaBuxZJ8V8BQY7QnJG
NQWqJqqEn2p93VjPwdgJUe8gclWjHdLEjHSFCicR+OCVXt+9Dp2+YKm/uJAAFW+Y
5HzbwU9+OaWzAW0/cj6Xhk3YMTdiMlHYv1t0vHH5vxKLKmu4e9cFVaa1N49HB7zq
nILnQRuNTnUnk28V4t2dyAY79ex/6oqESHPt5a0l+9X7W64z8vfNTq+3Thk6k2uI
uTBXWMAtFVKG2WptwsTAP4hXoNlaIH5IpbZZz8fhQ2fr2XsKnMxbbR5drFfkfzv1
xT55JH+YdFawWEPrTIpxkJAqlZkPdVfpsPNVsQGixmB20uiDOiAdVmEzgqeNqwiO
ru8wKT1e837QbTruFXAA1eabk6EkUvBAiRyYv5dsMqn1Bxja7FjLUww0jEWy+q0C
G8fpCCw8RnPOYhMA/5374fetZZABx/lbqfo2sZeDXGZufRJkLzhsbmdqFigvsbXE
Smi6DY278cfz8tkKUZll8OljviyA6101bce/LmDJulAotvaICskQlHl1DeEEOWcP
M5AHhTDB5KNSNCX1d9lP/dQQWeGso57ktuXxJ0kmm2o6GvxZ7bI1uDot7J6o/0tQ
/k0xARcqzE0x522t5lygSDAV8cROQXqyAtFnr9WBRi4adCym+x23dhalXObTtG/l
XmjGINXqTixGYabBjmeRnMCHNg0+0SRbJLROAD9ffkCQrp9mp0VhdiQmpz3dwhNL
09bhf2jxlztsf5NhY0oQD1ciav+w17bies/AgMW8IHUe0Ct9y9rQlAobcPOaFiov
HgJ9V/VKzac0NfVPIh+e+ywutbWvjafsZovmtANnRUejMBnvWUvlamMsRkmf2SBP
ozZdu+X9XOV+VdPNLZ5ejASdaUkWNx52TdQtE3KuYkqABXmbk7USwViM7CmAbaSb
2RoE+irU/OX4U+ateOb91ZxND/6C/Wxtp2dOFW7Z2qqI0lhTdJZXCnibLqPRLcHG
aqQ6wn80Pj8jIfDY/iEXhWmMjkvRroeZsKvMPaLs7Xr5NidJOPRe+An1Q7osr3vz
mwOpPC62h6JCD5Uhuo+wqF8JbHgfdHDUco4e58t+KO1TcgDSxubfobANus7NQODE
1LfJ/eDxJKFE2sWG7JvlX4WlWqb/+Cg5GeZlFx8+o0N5hvrdMHJ8U2OhBqq+vWAq
h4EBol4RnBrINbgDy0f+MirmX4iebMVEMkgsyZP3uROmnCT/Sr6wD7tOO0Y3wbjx
6g7D1IzyXgkJ2f1/DFogsBHSYuvswKUy5VFLANn4SkFQiPBkfawbCUjoHXWwUFrD
acv5ixsBMVTgvBKhcG6Vc7T24pGxChkLiDztt3v20HsKIJ8SGgl0rFceCeSMjYzT
TgVsX9pLXhfX83ZRmCedl+KydHu4j1xkNzAUI6qVtdPVOMCFh9YmuFL443dNYhsP
7T73O917FVzkv23jlDU12y1QKOusDuiu/AZVAKZo34jIU1vbSohBIXKAbHLy1FPp
X6ocu6sOc46g2c6Npu4GMMJ2ipZKGBXpbPWAaW6FBGeModV5lnp9fG9OXz2l1tbR
LBCYfV1skeTKO7AvABDd5yWlC4UzQ5ydOBpdEJZbPkpbdEUUg+7DY8WOC2oPw7bu
2e+55D3r4uTYXTSnwsv79YkAkJ3CNBN8Y81ZdM64LBI+zW4jY7I0hxb9Xg77kFjl
k23LhcKM7JrYkIpqqcWb7FCMJ3jawXYnH2Iblx5msc2kRQJdtQuWD4gE3YDoN4XX
34b7epxhsplXaLiFbARC0x0GB1q1A3xLk5MhZHUTb0qgATdFkybaz+HbNmvB4WcV
xwn4FRdVEZ3zYYY7dUi8QW3lxRAFA/+3OL13+QTkYINrugGIhjG6FsCUKpnq0vuD
lrJMTca78tOkNUkNENYb8aVFEItf0xgQ0My+6yi6d7iOgYOZoZNnLAZGuPyfaQ8Q
KR4c7oLl7M7KA2JBsFiDqnT9htjeV40mDb2ZlLmadenlG+UXBMeYC0swmNEXVl40
HXJnL4NWW/91DDq1vI4lpMJlpUVaxA/ctfbGiOQTbkzoMER7gR7ov1SSl4/hNXIz
7Y7PGH56BcXNrYuQkizBL18Ti0ioBFd1dMwe7KKT2AsA0DADXwlJz9ays9GKYIY3
/iWQoH3RaEm1ETNdDecq77blbJCZq93j5eJm9tl9ocRZkSJqmeRTtOgh0T+2EhxS
yQPxb0nvbpl8ESTvryfzHv4S+BNdLvvU3ZEXzkJ1TB6TYuMaXiTvuR/im4SlEpmt
4X69usfVcm7aPfpe8bFUgd4fsErMc9LWY8pSX2E7s9xWP8IBwvymxPYQfXHOEhgu
O610sQQeB/AXz1zw82ZX3djKlplSjl2PieOWsL/Mpax6Ngd1GOEaX6jl8nmVaZb5
teWsF6Ej/lTIqPLRHi/XtjvfbR9B3i9sdaABswdCjBPteiUAlJQoWiS7xDEwco3n
REWA3JwLkDfF3dYAs4dTvTHMg2+mXPGyCdI7Kb+uO45d1gMoXIipQW62iOJrPhUs
DUbXygAmWtVqEIJPnbBf1V2rSCEQMvwJ1hk/6Hto7KUpPW/lTfgksfP28yw2PpDz
+/g/whC8tLafW2obveAD9/nqRTN6jr1neJuPU7ykarrS0eHNUwXuF5C5NhaxVHBt
y93vuskDEQ4gAtGvtOQ9+Zc3OrPS5ItUqcQQZOat62Sd9l363uA9wE9snbM+RW9B
XhGYIhwuGS+0IByFt2Qm1IRFle5swOi8O7/nz3VxboTmdegi5uydDqvpWlqw4vjC
VPqs+1p4k5O8FPWElNO8Sq52F6+4+8BdzjwifWsHk3YnMW4WG6tf4yUO9DbSokVv
frYNz+gjwliA8wzFGwfWWgBJVAyc1apJi0XFX5I5D9QGgDOVFvXdxCqxZ/RxTnkA
VKGI47WHRxELIqMpdafShcJk8ZEmUB7jLOK6x3hBUk1xTMEv2ZbItpPop81wnD4l
dRjxZ92FmDkoGd/NjZfLv29YHhPrSk8XYtPpVkdKORRqC2Tz7vHMN3r7EkY+K846
H+v/tflWdkIaxd5zLn96RvHq2eeK8WP/aUfT0+3odg4NToHB8ZHNXoCpbjDte8/5
mDUHZflremql+oD51CxdXjI3nne/DEKQ6baBkpT4GDE5ukseAwcEurU70u2PBm+J
78CxEU2Sy9hSx6G5JSNpI0Gey1Nov44CkrEvzgihHZwwdCJxXBGmls1f2Ld1jWMo
rESJru6bpSdCKQNsII04F3P1LD1bBQnhFWJDW/0XvhUF4V5a1Y7EfrNwAqwv90O4
z9M6FmH5jhv87FdmyozXSJ6GgI10lpt6RN8jbbvTpaIOj8C5TMdyPfHXxkpvENLQ
JyDV4Z4MiJ/gZ0qXyXo+OJDYMwM70S+DWdlEC62VVOiQr525ktqXsgbeNV32S5fZ
d4YjMlpHsn2xSPXpWp/fcmFu4stTl16zLs0sbJlPu/vcW9HirNinVzqW4NoFPNVv
nNRhyo0GEq8pRrok21pV5MK1irWYoAJWLrTr2tq9n5FjODmcFm/Xp+Gpn3aWlwrA
t2HQlS65Ftb8PLXRVP4LZnC0vrJY2E1kb0v5f1piXzNXGpgfa5Up8rzU0xLFF313
aI7LyLUQVM1XAqbG+i3lAxpttwDObE6zC2vZT3MtcAgskHPhP2ae5AGpB469nLAA
rdu9wVqzA5svaNegyE6tYF6QZi6GMBgao+pdw+OKxvnH4P9hO9zABq5OVwpmnLzj
mK6seeTLr02fLYrsvUMjfNO1xsgrBJUqorpo28JOLb4JrKA7726R2XTZ+mnjSzaY
URbxWfmXSaup7uMTYL3P4zH3gwX7xBGmeTDXupuJPLOFT8mm+I3GBR1RO4X0d1XA
4wcA+TNOi7Egv2GiYkGNEqAWVQgtSSwpFwtDRqE78YRtVYbyBVcl2+UG40JnQD42
K8c16p0TyoRq+4RnU7zbpsCUcpMoUvA7tic6Y54fLya1qS0DAzpGHEJNJ23/cyZE
WGi6C0g6WcV/SPb9SsJYlMj240iB1g8aG07YbWGwkMN3aFpqLTP6/aP7TcjqyrOF
PFpTC7DFMEuErNC8XnGwWXLJGMPEUdQrkQ0K1g2SZdKAvduRT9/dAt0ZTT8ZXp62
6UUbWg7HqhDY3XeUamg5OI95MFHad/jbMof10qhmyAU38ymDuAX0p9UFLnI00ffB
s/tEqpvA9NkbOLA8tamkZ4lfxn8MKRToW3m3S6ntDMs/X3F0p8myRE8jvAOMHYYz
6Qm92xqGNdCVLQm5/Mud7J9v3PF4uTQgdpl5Lar4QFloRuai2WRlV+B2CpjKfo1O
CquXAMvcgwkmKDiYdbh5Miy+ZwXq5dLObAgbUawRBNoXp+fG5POpo+y1guUN/2g8
grs5VP/Wrm+uPeaHaXgvRsNcXEXdl5ryoZZ0bUx0fYarcNSdyUFakTcO7tyayZLS
QSA98/OtIhoeNzBVPRt3yhZvDMnx2yN9RR9IXBUPLJGxVodpdvpDMiJziHXFls6Z
BnJUuRk0T6ahdFAeySvjq+Rf+AgD1gdDL3ZL+kYtvqXr/5Oqz5NJ507CrDaUHxQu
w7bEVGLyrLO8yTezsDA4lVXdBMJsVKePIS/VwO1bZpK1xpZXBhYr0yH21BA9WPJg
0Xccmn8CDtItdKf7Yn+lTRr5jiCro3nSBorpd+tzwqFSZO4G2Ji5AtN0ZiHh//KU
2IYuU8Zi2KrJLU0Wr+LudVVigFP+s6WlySwyMVO3ofqiBV3nSphU9UQ4+2hm1iu6
k/Twnn+LUqo4SjXp4aIm6ObX0krs4r3ujT7H//1/G4EI/uvJrRcG3SZYURf4Jkoe
e8Z3BwMa1tA18WyMmIg4ZVPoFHTXmV+xeAP8FTYeIYdar1VfZTsiCCjfZ41PFzwM
0tI3zXcB2TvkgfpMeQfAlbiw5/5eF8D/BoV7MPTw9NhFRE6sWW4XkIhLQ2ERym2L
RzJhe5Z5sPanWiPcNau8EcQFddHZ2BdRZiapJIUBpPw8TelsMYgLGq3t+8MjFu0I
nCGecsBSWezb/YShik2WgB1mCffmndxpOQB2vHkK2NH2FMQnrepxg5AiXfpdVwYA
kiqAYItojdKSoDqQW/boi8SBWfvNiu2lXld72JaKRHNgN29ABF5WwJHPAyhQ0N6n
qZv6Qd4tyeTcDjoTbzsJrFLc41rMl4q17Q5FESJM8m1qG8jtX4YaBCwSUg7GAvRr
eklP0dWKa0qFtHWtuRTcKSz7mK05EoKYS6ahudDw1SGEw20GPkJ7QDDuEzCu2jxJ
fZ+H/O9kzpFavRr/cAQT6qrqlJq1JWLjXjNEFLgVBzD5MY0B7BhxXrZGDaGqO3ER
qs8CKK907tMzy0VUTUAbiA/nHIG0/yNVd8RxYQooFWWihT6XO+Sem0OisIOCMTdz
B+EuwDFwHOprvBjKCkwT+u93pIczg06mLnTIC34gDX6Yt0ViWBmOOqA87C8Nlsn1
wxuXqy2/UOfLIjSs9zsgcpxIbgSpYTBfhoUDPiHczEOECLy0k5nrzXCWkdlM4sxz
dZHPZLb843AQ+XoFqPuj31+fXCFZLVkCz0MHZ5u/q8dgVT5LF+Vk2tRlb13Cu3Xu
d+5QLqC+5fsOMk3304de0oFjsz4bi/w2k1nqYgVZPVaUgX362EflPRLC8po4YsXA
xAPuBNhO2yJFR0MWCM3jU83JZA7X/1RV414nb4j54VALodShIYUtEbElSInwWPaf
klKj0IuQ/tTUQbbNrBoK7kRFnFe9n6mjBiLbFpzM377hSR2JcSo63+/L0N5pnc87
EQtZ9z5LMA1HU8SqMem2aca3+wt3by811y2yZKcsJ+a8zUO49myURFlf7eZOyub7
qetRhyc9TrT8NPxgrzbPS/0xY1IlywM1vYyTVx7Y1Bf4AYk5sDEx7V/5kkrN4rot
95k6yCv1oK8j2FZzNXkETrvf2CWvRHNrs5YDFINRGDmsiZXdp2scWpeGIwkf/GtF
S8s6WBhGOC3h5Wl64YDyNWaAhA4E6OyXYtlCyBoukym11m5CJrjUW5nFzkiky3zz
/W4NIWSHd9HsszktihoK7svW5DYky0TOAoVd84u0/VyIyPJqnV55Vl96d78ZvzIf
p0MI4+SQlBthzEYCpRzhaEFLFhl0CrI4JBuUL7hHDRygjwxHh6QDA6gWRKg1Zy/W
ujVbGdzPpZllH69BjpDgFynocePpABxH9u7OnD9dP7eEhzLsn2U9nlVfrliuq2vV
Y6LhKW7fkmMT4TzYO41c3cUvvJ5Xy1KeMIu/a3FGDAX0Wh+Mn60XQQ4wsKz5wxJB
aP1cFoHL+73trQbQa5HsZKH7nNgcbF47ercAt2dONrAsftUYKcvkpnYOMZ1GC8GX
VPvOlO2dssvVCxi7Gs7Llcle3GDTcdDr1tCkzNcH+cNjvy/5tNjYIHEG89RI9yBx
V0X7ZCq8NYtOBb6P4fN9k+PgksD2kU1gkHXPw2DWdkxGLpqHCiohMODPcx/GwXWD
rgcSWQwtrdGOUu7MRHOPSZVJVxUTO0mbrP7AYe4d73jdCyUCHm+g0/Q5mxC1NYnT
byHR2MPS2B9JvigUe0yLzAxmviKJCUCbEI75fqc/DGVbEN+DkS0KiPcVRj0HzJFE
SwRyC1SE5KRRC8r3cVY6pB+ZdNKvB95vZHwZYOVyHZ5KOEoPcF1kpKVF+VWVVntq
rc0fSVFjglYzRabVqKra5eS0oNuFUuKxubEg2LZGQh24H+zWM7An6g2+e3EfVQ4Y
YK/wp1JdOKdWSl4NyhZ9TQbxwAxhtEBpAHV341ab5SBv4xq4eND267sZtZp9uPiw
Xv/e+7Y5Cuf0FcLkgYZiB0TM/LA66yWHzYIOk21m/4CBggoqodZWa+dSnVsIv6hU
c0KtPLSEV2mNKaur8ZvaHYzqThwA5vPiWnwqURaCkU6n6Nt7nK1WnTTpwXXfPZhM
3KQKjsxbdXxLcUd76p98zCqaqkurxQmosEV18oE5ekrPwvY8h94qZoWfSBz63Njw
w4wECV0Ly7OoprwCb/af4Ogt0Bx0TXlVzw9xw3VqZoNlkN/A2aeHzeWHhFmsM+Mc
RzHJy2g5lrKt/vGnRn09dkCRRFmhfG3F2S9HC30Ji6A6F/FWp38Ow9jA09Y9eY9p
k98FwJJizRGSK4dkNn8YjYEIWPNbdyOP9gKCvuD0nBlPKtMyepqC23A4B45Mq8cv
j8IojWfoKI+RG6CpOIN9Aw==
--pragma protect end_data_block
--pragma protect digest_block
axOHD1D/Xycts3M9TleuBVj7tcw=
--pragma protect end_digest_block
--pragma protect end_protected
