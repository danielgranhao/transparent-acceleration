-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
cxJkXeTR7pQQtjO0OrtfhuVZsBkXvAX9WwNgm5V9BDSFcYa+RI6abaRnFd5Sl/Ki
+uUMBtBwurXQGNwPo1EhH8nvWmZL5jdWKeC/79emzGpCur89FVa1Hk+T6pHJw4ml
VrppnjzLwFA7WaXh0/A6xHWcO6LbYDYOeZTijigBkGM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8687)

`protect DATA_BLOCK
LZXmla+pg4nvYbSVQretXtLeCdCZNpwgoFk6RLiJhxuouJfksqO7zyVYCUYrUYZe
14CneQPVEa2p81ebPcDNSKDy21bwMW+BMBsN9pWSis03E0Y/DcAv+XIsfYifAKKK
brxBVMpd0aaIEOVdl3KxbHw6+Eae2AdSZX78tUBH8y+umOtiA8pdUzndGcHfczWh
AfuGLfvroTaDnv+aY8l6ZLQzkhLkd6deomRiQywK1L7HP50SgigcnBYtEPEeBqeB
9AYwD9qPS0Dga/KdOxJlQ0H+vV7YO3yQyqt9OD4rEIhaBmbUcnBy+55zBTNC8bYZ
zeiltdJ/2JHoOLa8u44HUPfT8do2RHJGGrr0oLeoxhRSiiVEfO1Hk2MZV8m0wdWs
NCW/WM33QMPIhTzs1rUj9zYJYCsL3oBLrAb/W2VGMMPx2vgXjC6JAiDZqhw8P4lt
xvvR054p8vQQkYmx0SCcOMGAboB0/1WFod0hOR1rSF+SAB1Vmwzfpk9nilmBFDqW
twSJwhiEnsKVu1jDrEM/KP6+bcye6raR2e5Gu2EK4sqUcr5BxIGWWMoLSjQe0O8j
f5ToAOSA5FPGhVBrq2s32Hv7CK4Rnod15Grf6kMWQkR67TJjXs9sOIl5Amq7YDur
XThDnT0qBnAqDkgAmScO9KsWXEGbPKu1ILM6nAg6Lo831okHNLALJJ7yHp0VlMSB
PSoruCW3eQeR6UB+5rbWocPhZEakLQz/04TSPvdDGMUcJmAOMtUmcX3INsJqshhn
7KSZF2ahK00syKxcSXIoJWVqlakl/O3/dOhX6rw3xUtnAiCPiD2rKfuwVRA6C4C4
2PRNEJ+oxgKjr/vggVx1cHpgOghXybSwK/wbWADN1UujpXmhyz0276xlFFcJYkbG
iax0tTR6Wy2DIeCdalQxTGPQeGPyRmAbEQJ/tVuMdGbptd+7wYQnTc7AiTeJ31Qx
WgQU5KnUoSq7V18P+RH5TUQXKh06Wc/1bYdwVdm5EC32+tWRddn7d/tS7LVTztwb
0I9GGjHseVHQP0q+y6RB59Un+Aj07QcWZQDTBVBlEFWe+F/J9BDANZVxISw4T146
Dm+E0pf6YUDsaXdV0hxcWXL7d6HmPnZAomWXI1gAwlYGIRAr+S7zeHzroDU4m5fa
J0KyGgpVjOezVEGwiKwKYp22FNiykdSfU8k4uLcyowAiEeTc1ryx5bxYyVw9mp+r
gJQ0R9Fb1Xo6ASDhkZ0456tX8mNKS8J9MxpArkcctTPEFL7pLPT3kTbm5em3tGMl
Dh6n3DvmnD4CqLWRVe/76Mw1auCcqFZVMPSmyJmpYbO4F15GyubjrBMuAdTy/i8O
lhbWhURU448Kup3/ZckgJVEnbmtKURs7epZtZkf6kNWdF+AMMXmZgR/XXkGzHskt
635tlEhRNM1RBUwiprT2WPKG04oTN4zvR4AtJ87Y5DHtIL3eG/3GzYqngqgDKGK7
GoK48WREVBjC88FYPAv1fDySAjPFMo8k7iYb5cEfoLICe8A6yQOJeUXjy/jcvcpD
r6OmQQabR69JKXptEwexclpZRXE/Ns/TD53xQoCs5IBFYyzPglwUxWmlXWG6nLKW
3oYLE8wkXtOhbh0wn9dty98LZKS12DBqdMhnY+PqCN0Tkc7EJyHWpSXMdO7lPDeA
+n/2R9hBw2hXWbQ9C4YMn0L8vQfr81v9Y4OzGJp7Vi57sDzQZ+wr1aVrCkx8DRRL
GhPY83qeLZxRPagjtOC1pM59CzPmbbt1Eg2vq8sONdrzXsMPAG4M/UXod3IspJQn
7TBzkw+6z2U3n9xKrVR/yO7XR96Z9icZ5GfuSg3X3zA//leZ395RWGgI2JIUnjh7
mOW412sy+UkmgM7hInpIzA92LyHz469c6GWhE0cUv5YQhZzkXTvTMPxLthnsiixb
zUhhmXAkPidkbbea7PO2Nis4h+eJzxZIgzFHefxI0TafKnXjg49Y0H2u0ypTl5jd
LlA6Xh/e5BIY1kVYwjrmljUuvx+GegxKuVN4eGBwFxekBTgCGIeLClEIVHgwPW40
c6rDUK4BlXEZnOEsQl9C+5TPIzAzh74RHBq7t20bWVXb6LviYlQnZfnYE9cap/rB
q6kwbQBvB0sALHUKHkEJ4RawjsT/QgtwPY+ucY6xkmPoCZ+pwq3zWArJLFlGnQ9y
YrZAVLAyeykCMjpZFc+LFvsxSkoTcvfA4jSoCnik9hZYE4OTv/xiJD8sTi2dS5G+
QIeaaEq6ANcyOf8fABaLXaTxZ2HsEZDiSrn/BcPTLQMGCu89FAaIehLC33nhv/Wk
XVs0oxralCe5mOIIp1hAmLJTS+18X63WtF8qjoWHySmlBMNj7hvMX2fTewXI6f9R
DWw/YHDhJXVRzY+9qcW8XDcizgmaVN03txF2qmpRohKB+B3TL4p3eBTgPAbyRSoK
AlNZrozadxK5X/kmWjGA1E/NW64Rm7J8p3DUZ8zMBZC0AYkSdZadOMQcTo31Jrft
uIy9HRHcF9BeAmn4Eo9UspvEgfFlhv8b5ZooqBh/iDsHHkGJ12UptAnfydYvzUN0
A2KssrQjOjiTFZbT6rqNH38vPQQ2XLw62sI9z07KOW/5i59qE5fgflV5E5GJPFvU
Tz2xXUTG7o5AEl2iyeXLgYvs+BATOfRtChLF2DUUGXTMXB8lXQtKIJ3tKn2P0zSW
n1ISmbS9A2BknL2eBy9UQ4zHknQ+Wj13begmc1gBjC2ofJS4jyAqIp6cccDsNf+f
SMAR+PXXPyeoaXENNApHYMSDJlzZkc1BUiraPfwufYXTG4QLczvJTdi0ZDIZ8zOl
OJJbM/jT/Mf5WXoINr8L3H4Wy6RB3WpxmK8Pov8lnNIJVf+AOn50bT5aWeqGz2lf
3zV7sk/o4No6b1vnmMcKpfb2PhkJ3OcU0r0YqxrXiBJUrZCq/OYYKm2LIrQlZnHV
ncnV95dgy89DaVkJpg7rwRo+8rW2kF8kdomuE9jYmfhK+rh2lPXW6QYdGRJx4Gbf
vMnSzQNT12CqAASc7/SeI3DzLyowHhKsN0gHlAvayfIqioyfouac6kr8NR3ApVRb
BXjqIZuEaedEtHN3jk6CAyU9MQq01rcZydpdrLdLfh3l1F9ZVKdWZa1z/B2D1d3U
2pPNNQwQDtH0MB/KKY5VCsl9Iq+yr2ipKSeIRA7Ff+vK1NVURXHxtPqhhNAdn4S9
voSNWM5Pgz5FSqD0YQoiJczlBviB0Ww9xsAtQBwYMhluALtmRvyZWoFrllO1G7np
P6uDXSEcRza1SyCIe9UkvlnK/7Bl+hOa007m5j/VduWtI+ncQKHtcJol/3lfo3en
wXKOd2vueU6XX0fyuF3fQlLDKdzEBDLNNQYJHrv5zsHBuDdl269JVqipkqhRuuFl
2HqRQYFJFLmZ+aSFl9/wNUljCklJT09hjorDXAk+JUDJsxURTHX5B6IE2tcXVtp6
wa2FQGpkGK5IGbwhJj3tOpGtW5RLNZIyrdVMThKYEbelXS7HOQRlT4gwMQ4vTscX
rlz6+hkJ7YZlmhOwDssv2iXmRsPjvyj5dIz7VaxxvdVpRD205oojy9QuUgGtuheW
Kn0jcHLhdm9Al5SnFNDZu1dAI/5B+Qp3R1Jgyr1rL6jhCYJ+WJFyF4iZ9ADe019q
x8PeIM/HnExYTEA7HB5O8allDa4uh1JE3sRqj/Xff9H22zT54wmpsBwTn0zEe888
usbjVOptEjT9Xx88omBZ+lD+gmpM+yXfACurAF3sKg9gap7LVH7FW5NGZCzayE/+
4jHtFK7hh/EoQ/fvAi54Un6DFn04EHQAIGsODtaA0xWrpjpH9/RrVm44m8hDoYND
19GT6atLKyO9XKSINrARPzu1A7NCg5F3wqUnUTXsmgjklZZZ12BIHs7KO7wxXeyz
c+4BKV/YskC+VoEi3GbPray4+JuvUvy/blS0EEvR1xmGO4eT2drSRMX76vwSXMA7
iqzmewTReVv2wZ7WwehrEkzoxl+CHmv4ImLWynHQ2Dri15jjsxUmXBO1TfsmB2GX
lu28BoG4KuVT8ccq1VggW8HX8MUDOXsaHZ0G6X68p58TSOeTLVtY13rmjSsQBDe4
/WzzT6tZTc7DaniRnpoi1kh7+XzhjYW0NClbHk/Oxt9s2Pd8x+3I4DtzNnQ6WCqp
2XXMz9ClBRH5oL0SDv46Mzu4YYJzdpm721/ZxeS1yoLIStqq8CyTAUwddm/Uf1b0
Ejea+SJCQxpcmDwDxIcVY80HSyIk1sOqwtiUNOpS9uRR5zwWW2yNVY/0VG9Hv90Z
r14iHfeT3jgxhLNAgcrLGSYEnLwNeel6g6jdllCVRZQyAfB1xH8aqhtdj9Vhvh4m
nvvFZpemzb1nyEN2tRFHPUOBkBuptj8vghbLgCtZ1a5qI7Kg/aI+ASbPW8MngrP9
7yru0OQHfWzzi614yD65xCI6EQwN3RJXeWlaPnMkBoNqtNSzzUL/otzlVGRQzxfU
lDTSmnwhUuF6VNNmWtmPa43LUXizP+nzsiWWHed9N/fW/uzkqj+tuYm3LVv4LgH2
6qV2OFEb7Tu2EGiyTvomOgg25h1ZCx0btSkaT5MVJyYg6k3uhvKFSwzOrtvRA7Lf
e74QxawQ3u9Oxuygl1cWoyajQTEF0A1pfipJgJa7dAiQEz4S8LqtVE6ouGFoC2E1
pXcUDSFW1Ig1jfIyAXtvlYAOIpRusP3mGsY1xc87gHZfjUe7YE/0+LLZQNtm79ZS
LGtIs+N5VR05oTfM3WfRneFSJ9zoUYlAVjcT15ledgde65XonQWVhkvXzGbMwyjA
PFzBgt+A3kMJslWnu2sPHlRKkyHEgruJSz2sLMplQhu3t3k4yBIkO9/rtV1iDwlz
XgOgPkNQvkMN7DWDdEVuFf5w5xW2Y0JN7cvlkexE3Sb+cHVaHP0b+bnZtIlb4o55
d5slP6Mh9rAhTlx+JeNnFmJd1qHyhz/qwgLVCyaXSy5Rv8tOmc1hYadTgDqUBp8Z
ApX/5UggFWTPMovLZfY+8xZY9neYGNIEQTM6reFNKZI1f16ESTWIY+5setFo1dO8
6tS9OC+khBIREAgus7ehRldYS/bOfCxWIFqeOBYeHrPo1Ap4jp2JnUZWmP6kah/X
KUqeenA1CjHTLhiFbClDDZ3moMeuiDeQU/z2eXVMsgJnzcyZZ0pyJGPgzOt7g1WJ
XDijwvBlcvv46SlPqBwJy/39oYMroXeb4Xj/AWQpixY43+yCAbm+BEwVoL3Fl8vI
kLRlFyxTHe0oa7hw5kpUxO4PCgya4IaAsMnpWESlTrViHdJCkRxpKMSRcxps3MNX
s1bAPpTXFNKBfhDfOkYlZL2850/dqgkjwItJfnVtZ3vBtusrel5bBnGjm6BKAbVy
Nk1/isqXcImbgeUxFxHTjm+sKmvFYK14XJwAkHu055gNZfLtp04+RW2t/0CSzP2E
rHbIQegkKI9g/Rry5QzrvbOM0V8ImBt0upl7+Xk4cW8pSBlk3Cf23EHSbNC6sNgr
bbXVRcjFhGkGp+3CTw7+es+3jr3XIG1/O8lnpm2uUh6YVXas0uRtMe0f0DalYotO
WneTHaML3gbuUudYhLwUEmO6eRmnGuxz99MuGrtbMycUMIK7AFrU4PfoA/bxQbN0
LgkOvstmJBtR+vccvU4Q217BbEKpSi4gInKbShBNdMXUKuQe1xMlf9paQA+Of+Qy
3uXByHpEw7jqyHOCxPdtSXlEhlnzpj+F/16SP26GCKLCpbkwNObQl2+2Wg5SKnhl
1rwluq4OQfowitcrcGOWoe/Rm1uvdLZ3wk8BN2RA620j61CRBtKvQd3xj5XQOP1r
IHwgSYqCTfEvwoq/lCixOfIaGiAsrLf84OqiMW5Cw9tRpnU449laIQCEZpNg4gPN
jqKK1xZjqXvft/zFf0kMjY6TlOnLj3d3BWHlCllD8NhK86PqinnV+lXdksUcd5eA
+9p/LKdtWtIvwqQoOWcvHmrGiUsGzRPqXOCbfHBom2y3mIUKBreOF7dXY6Cj3Yq3
9JPzPMOnGx71pxJhBSgJD93ddxYpNhKuwyVQ9Qx0yWmYAKUHVed0UthT2m91MApB
e4EyUJNVkUPHxnvkz1RMDtdpQgnZNam60zZCUQiiuUUwvEmKUNRrzA1Ai/hb3RV3
xNYFEmxib/Js84APc0ENwGH/OKed3NSaOA1B3xeO3INcrw790ftYj4DaOkeRxmuw
f++lruOHRpmPAGqB4uvbCMRHLeTV3vnyMnXLZ7Kcq/oMl4VginlwkwqOs4e9AMCh
x0W6E7radhqRY4R/lezNZukCKK9P65BrVMNBCvZyLVxHyb8tWoyxzClbrUO83c7B
3lREP2TY9yd/9d6RRVp1gtJYbRqGqUBR5z2azpc2UthDfgdVW20jeDsSF/MkSezl
aRts90MieErA6gpXm9K1DUauvnAPtzMzQBzkQaxRN0HIokF86/ZIOuWs5nTngFSI
JcKOchpFgezdkz4r5Vbbglzd1GiffQ4dOgAy13Fnk4EgkMg19oYsgDHWT48+8T+l
sC8o5/RofEMueMfPIAkxpIUxHKhQ7wcI776vdM17067i/TBuISt1nldGlZSgPi0k
Kj/edQgEk4DTxBUDQqcH2/z91uiMuFNiMawkASCKtQhxtHT8hIrJl8xbZmS+doi+
K4/tUrDx0A3Qwt/puJdrAHRPWtbYj1x7Mm3YKWVlQ2jRetQsUZXhv+wqria5jOJG
MPsdxO9BayGLWPs2Sd0DBSAkOLGJTYHNcsauKHkCWzbai84AOoJubFf2k5tp7hf3
xbV5YRLm45BqF7+yQqU6LKmZ62fTcDPOSeWjQhGFZYVYc7NRw3lw+sTBY6KmtMJw
2xzsEOW6tT0y1u/FEAsz9Fzp2AIZLYz628/1LaHsy0Pw43k8owLOru/anWjdHMrK
rn/FS7j4SBohsy8tQshBQ8eCuykF+RwzzDGY9az3xivQL1FSBzkujZOEv84Kw7CX
BgjkHTWhsDfFqmp8tj+hp610mf++5MHBBAFv9CEz36cXoPVmZZP5D4PkiPZrR87m
rWuO/U6tnd2mxYp7sEvi3SYRnGx4nlhtQWfzxaIETatao7fyz4oIvMuoPcUGjRHO
vweGNXWRGFQIc2QYnGIGGVadgBAH8nNjrfowhht/YdQOeT8gR3dDewLxdGkV2MuO
wlpl5K3KvNhlEyh4qrI2xLC/ZcM1YXqA3A4KMnF/9Tpk1LkBWEgd9dVF6G9V1Lhg
ObmFJG6qE0XaM+Ae4n2KNUGIiIfGVsVxDg8FAdTJFn6cKzxRYUrzZbYSm6OYWexb
Rj4HHzG/ii9Np043KIeYNcNoh3b5gAnc3uno7RJWy4dfuk+3nJfpEeiY7F14fw7c
odjKOe8YbAN8uLPuk+GY5Nmky29UHy4IJgLdWiRu8Yx/1/NV8OHKi1oTScFKGIGD
rwZIv6HRcVS/om6/15WI/cx5h5vNqSYwFqiXPgpa9ty+6BiaKndvuQPUOpeaSnUX
bEeWfUK3urbUmm2gRs+OnCKV5gXcmj6U39aX1ELWAIOMlMRLDy11LlHrcAT3XjmL
smSRolCC5V3Gb8Xnq7DK8TklDUPfC6NROUZpZKFyaH01TJ05g50AYt/I3owYD0Ot
RO3hV4wtB45j3R159H4a99qdTqS+07U4Br/dfqChPu3H6X5ZMlSSEaaZavGCWDP/
S5HNHcnddUdRDbPXTNqwTM9tecFDlaLxbsH9duGo5LHg+aikfcfRIk4U9awCIlID
0DeV4UdP8CxkGcxTvmWk+h7B3rZsYYXZRg1DK2I5LXhvlAU4kF1xMNW6qNEvwFWx
IwMoEd6GzOSS4k+tLrHkFeT2aBqelOFPfL2uESWqvKkKFfvcZwNeG6b3wHxLN6NL
OrLq0HEFmgtF5lLduXUYigbwP1wxKuJC6ppG/kjOVhIlMzqTJGgI0C97MXRwExBI
g5zFaN8TdWeaFqbBqvZBjOd9FQi0MdkMktmf/tRim3KQVV/fvqiCV2wyVvvsXb+k
lN/5I12dD7bYH35OKnO/TtS2XpBV9EwA0y7n3ePcyMdIuz2mFrza2ktnYl0O9sRg
gbmWLW3qtJJRfnuaaKLy2vVvWwI4taJkq3qg2/e3slGrJjrZpRmNmEEcnfAnSIXp
JocsUL9AkeEaqeGd77crNZBVJGEV2ajKWQy4Q9bRx3LDQp4UQs4poBOT0sg2Ar4a
JfA/DO8+Ym1NW1sleDfwXfJHCbdHGSpegtTyFC+I1nNKPj+7+rU4ch7tdy+5Uqqj
8eZCFzbOoX8akD7R1uZEBr7Q6EqSUvxu8UIHXhm5bURMJFFIpJBUkPCXoOYNnwAV
lb3/xKQtdwI2ddL9C+8uOZy38a5kKmQdEJqzSghEcm1qZ1hdD9XGnbd0COC3PqYl
S31Y0MIw5UKQ2knqOt7D+t0JL2Rmq1fz51TDAxibsKUK90fa6jVsOUeunGXfbfHX
565/vqXGQ4SC2bW3vdpN/JzotyauEE1dNK+JS9cxmsV1MJoMjuCMs4QqbWnLphRB
euzWseMAUFbazCLiZT7JkkVZ7DO3ZrfswrTvhklwnLXZtVEAHDUU584Z99T5MGWj
iAMuyn91lIz7sIyVZyNCH4SWXSVsdu+8P+Z9BCVokhplczTlsQasMhR9/jHkolpH
FoNJfo9hdy/XnEnDCHfKyivBCeR7/Eu7tnp4wDtL9q4E0QhlHl40FJ8KuXzHKCdK
ytDNodD7sbni+Isv9PmUotUD8MipUmlvQ1VGk4O2WDyFxBp3Dlw9Id+KK4oowxo4
jYE98CvMolxjHY2KLlVjX+3XUe22+9vBC6R5E1es6ctI5nHgGbW1Xe0fjcLQ0lU2
9Vx33RuosJgtdjYDP8yI3XHGZ8B9NY+TzLpeGPLuXfKFeOPt9+TmT3h/DPXhIOl6
yHcDuOicjuDGp9TlZLPagde5Ij3WLqrgT40wGxX6Ej3wBBJ03XbxhZDkF/IvMGqm
QnFaOz9TNBFEfaFZhpQsU4XvjqgVtgub6RE8kQjm/IQtDRSDJPq+b0yLWC1YDwkz
8aZcdhnkPWdQKoZL1YnI1zCnnaAhM6I/JLQ6F0lno7wKqlFPNDFi8PpLZpv/l77d
vXQGzrtHO5xTyfUC1vhQjeDFz5GosPVZ3uu7gFSHqWw3sdBXpwG8iLMSaN+PX+fZ
JPb8+6Fq27IZh+mnW9i1ZhoE7h49cbTN1u3jKsHiLH0XbcRoiC1icZcunvk65r8d
LP3Iri1mmQes8TPwx3L71ns654rtULmJHewm7JFvsNDpzTCdRy9u9FnNLiNcPeff
NbulTeJ+lVO0Zlr5VmDOQcFpJbIFbpUDYG0I8Y15u3LYqk4hdbMqVmEfM70Y4cnA
qvetxUaJ8TFx24gYHBHFlPfVhrnj24Vry/LScd/Dj3MGkgaNvO8d+A8zqo8A2zLe
D4rTSaPpRHwNOckP69KosnmG9rHHn89aXbzMul1unoL6GhfUc/fXb6/wlqq4abKz
7Mo77j5TKBsRmzjpDZFWDSRKTMMt5V9BLLyT4RbETKEtHyp9E4u5DL+uBI1jYf6a
3YusTQLYVJ+ezyNGE5Ebk1K+Nq5pZogwYHITBr+HHQEjD5pSSXi10C+iVlVFnfNB
pqzKC1MWpeRIZV5EAsu+6g7q+JdguujCcgOcG/Sb4TaabSXBKN/LPqXPPes7MWZv
YivIR/AJiJGJOG3H5aRKk0kQzEr7Dx19bAPsoEfBO3kfZM6YSISWT3yC6yGp46Ht
8tCIxIqqjoBSIzDATle7pPyKDZdsxgON0+IW9ur+nr4AbEAJ2fJU4JDurx0jhuAX
/C76dfxNz2/VkHLPFA/WshyK3Qud7tu7t36mAQQCUVKDAbciWrTeAP2qfwoz8OgA
WhSFPsgUihqSSITYWejr4Ga0FBK6bkZs4six2cZ3/Zv28RZWqAKJwfHGQntWU8PR
KJAz2+6JRLpu1cSOiKQCMixXGhwQ+YJ7dkVwd8DhIr+RfXQeK2cHY98DwDR8qeFy
ZedizKce5cK1ny28GkdGH0D4dFlcuCu3pkfwABDBSQLhJ1mJTII55Jjup5bTFnls
Mhn8zsknXY0mxsgo5ctTyx38CktdEcb5O6V0EnobSf/S8nqJOuN0ikB5M34oCQ7I
BPWchQaCko0Q+kNX0+0n/gD4tM0VO29MEsg/DjAE10qwpfeVz0bgUAW03NuRhG62
xdXnIdoipm38KvQEEcl2HLTVu2ZOS8kOXjEJKck0ojpCOLdimVikve+mJ2AxJUbD
qliIGq346YoZFt/vcNjUPDp/fN11xFb12ccqMaaaqALMXPkm+bb8zjdiSpN78TUx
w5hBwBmkoeh2LQjoas+rCNc2UUFIBH3+HemsCXuySozFIY3wznd2T6RHzE5mDgns
T4hKKulBicK1KD3cPEY2UQcr58caugMNgWpIeviiZVpXnxElfq9gVRRgbcK1hRsJ
KdbCsj+4FtLYodOHsjdUcGPGm/MsddnpTCnCcTKPWaKKqRPLBT7W0E+Fv6qFsXId
bh+Wlv2+q3j5Nr5Yeh0AypiBrKnY2NKLAc/wy4LLPxHksEXLwi+VjPK1bPVmem10
YftwXLcV3uiIxECFvGrfsvU8iveAPEWoS2Toq+Bk5YWWn2CeMmvBq95B+c+5+c6e
PY4lRKGEVWOkju7vkUpPtWjF74fEI0V38Ee/ysI9o0HLVZvo96n2WRU372gKb8VG
ySykNK4+p5VSAeHg3hRIiOPGrxoLrK9fcAezXt+ZmqfI8OXQDLyBCIt3CCvFm8Gm
rEjiVHNt2Ka8lqvHjR8wtGSAZBR6z2C/aZQcvmG/txAl73vfra5mbltdWtqYScJ0
aQZ/euSJPH/Y801qdPhtwVY7Itf9oKs499UekI85G8B4aKHkHbLwfHbTrT8aWoyP
QfSTFPfDlfnJxRJFoe7UFTGTMhOoyJ4FSZPMTywq0CDCEMgcM8Oqk9epPvYsIFrc
S61pevLhhKZdc2L5GipDS+HNJiC7qveEyWFOeFT/Nybd7B5aeLFCEgh3wraOGNLU
255mbkElmlwiBD2UaHprb1CoxiYMiA1zyW3Gbz8SZrLHzLtJdMtF+py3/UwlAj0o
sypcU5Npdwi/7Iw0oGHgu8PTEwojbXCPKGB0pEbqewfGEJkIE8S3z6jlkdqdA64p
UhUSN92rWNjUyK7jKxEXLwGfsmQvuh69yXbBWkKgZba7YHB/HCQKE+4a2hzq0+gA
T7rEmG7T06Dn+SibZxNzStYlwf0O1Cdi+hdgXKIsaWbBED7eBf9BEUjeIIxHEpqo
2mPqdU8jfXkt1gBLWV3A0QKxi25o4PNnPYhhiKS02G0bffQ++aEgbG08h0TaKoS/
5RziI62BJ1X2KiU0fvSX0aKYWI8X+oMLN45HJVJkGfL3HUuZ2DzhRZfFAHfggTlP
j+iTs7fdN0i5/TrJ9i7Iz2nDcQ4ker0IgwlHI27mABbR7jSi23znTh8++1Fn/n/O
iB/AvfCKJ91P8l4lmBDI4/iozD4fRQ/8nBfF5UQqLPW4zoPMVB4OXU0ivkQ7x8zp
v2om/G5I0wtJOTZLvYtjWQC/K2HX4GT4YMIEHUO46Z8LuvFdHrotSUcj3E+elTWX
I1S7dwr7U3q6uEpCVSSveQ==
`protect END_PROTECTED