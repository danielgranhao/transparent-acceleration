-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ATkX6waf7auznxpZx/S5nSxtCMzZi06P0ptxs3QqA7Zf1yBjcikKLBxcN3WmSuZH
bjiN146ZcK+A6u2NoL3Deo/sTagj59arDBZy8J8yfhXksjKWbxda3sIC6EhWMZqx
cIY3CyWF5fbuQhFGYfjRJB6XuJXB5oISuxDc/7lbuHTTFbpIj/lNIg==
--pragma protect end_key_block
--pragma protect digest_block
h/kw4fN4pBmWGFkEK0cEC7HMDtk=
--pragma protect end_digest_block
--pragma protect data_block
nr22/2ylsnUgkQMJxUIxvKv9bj73rN6nJnMTKsU3BNZXKYJYRF09/9Fkhmn/gTjN
k4PNROfaUYt3qz9HlB4j3whRJgV5zDXRjClcbj1gSJideSladjGo8QZo/vrg1r6M
0sLoJH1l+UryV2rkz/3FYX9hoKH1+8Vlvz8oSU2Qoc418ySLJzx86EPvkulO+8ew
JgHoHYkkhLWS0z9/BE08a0GqUAmlprKfZnaLhS2MXAqhZulOkj2u0DPXjSgQnWDs
4J+fUH7aiobainvoI3lU6uoJGq+QUTV4VL7hGlyPYJxHGPM2S+Gw6nnfdbpAyMg0
o1Hy62jZWzzrygfrF3Vnl1PjSass0aaohSSuoBVAIrDjY2AtZ4mgukUXAySyXny5
3UT0Llhxk1WVpSK+uNIkTtJZ7tLvykcvJHeqFNCyvkyvsk2EcNC689nHpQFck7TT
+9h2RGRxKynQoabuxT4bgIoSyjOyvSDR9hmnkpoy90Mtj71U7WiXbpZ5fMLcACNl
lbvQ1ksH1CD/eTMcPSUG544DoJEPiWLFwh1lkM08XulVo5LfkDs7y9JYl/XU3y4c
e845a/AxbY257LJGS4uy2Tg8g+k7ucQg1hugB3CslLrMXGJd9Vl6Gj4Wu7yatQig
kAajv4LqVFhomgZmA1pZ2F0+o/CC4QS4GHJAl3J/CIjFRQjoYihb1f4dJnZy3S6A
byNS+r+5PQb+H37OUGbyK+A2mNyWfUltbUCVvMYAK4WNPEIHKaj86aGotiYQB9UO
7MrjzIz8tCY+VYxgMOkpS5ej2qAlamwZLHJxTeTG3mYfypw+jlEe5vY8tUDPgxPr
KNN+bkzK7VqXnfBBgkcd3rg0PMPNwk7SP61H/0J/7TCbn5topKFpfg0Ytybp7li5
2M+AMyBspVirSDRnRZnfs+1DvpoEHBIAzWdSJ8Hn6aTDoJnyLxSi7TGR/pJY7pJw
3KZNkfNaBhiioCOoy6rYl9xVeAiFyrVvYfD1dk0uuN4ZhNb1y5QcRhCx/E/mRMWS
SqHzcWFhnshr0AaXcoAxBAlGxTFX99D7DyQEJUHut9DKhN2hsmr0+26/IjLZdCOL
EORcZ2eEuw2+IO7cJ8/YXKkbSO3aoLaRUWBCIXE1pAxSifuoo3bxbn96l9P55LRK
MWZmhQU7I6WzmZiE25kIg5U3z3mEhOxC87xhPT7ZPTR8HshYrOhZicTebFt+lsf0
u2Rs4rw057Zmn+heg/ImIlCnv6Y+oBh8ywEQvwCv26rJXvyeIjydJQ1cFWwPw39O
n2ums1k0e9clJK/x2la4JmU5Pbq9+I7IZQPFkm/EezwO8/Zdu1t2zBEajRCNVa47
6gGk3d9hHsr2iaDWqMlV15F9GKSp7mf90iZ8mjKCKFzs10Pk6mDacoXWekiGezBL
5R2ZAHGIK75uVC2mx5qzyM5VC1Dh27g5NTRtugnzg2s7suIHZ78TyE3dSPSlKUjy
5I/4aAJ1cWVH2mcDsg6Z/JF+VbSngv690vVjPWdQFqyWDOZ7hYTg4q5mUEyxz5py
/g9c9hpAGpRfx1e+JwOhjXOo9UrcLDWSODpRDfd3tRQV5SnzeJh7tZQZ3tjl8V2B
b9BbKbvYp0kkqyzjtc+jDMZAUF4d6SXNTEu21NIVYj4dcSvkBuFozJSz5S7PQkse
GCyDTaKgQL2mUHKpLzg3c68SXOsP0yOZpBf76PI0dDZD4Wo4S11oQ3wGLtYPBWSe
FeG2jDQtGH9wFbFwQX3No4RlHsX9G0zxfI3gYFgiKtd3C/qnYoJq6hK592X26zcz
NP9d5sFeGIV6fXdCTq60ewlF+YW9YqC0D0fpa05q+2MyQY+o6iN+UN61n5eeVP91
yyYmmCray+de/z8crgElbaWCkTeYVilv1QqvNL57PppJqPSpQPqJJBQFrYEXbJOm
JsgTbh6Q31eh/ErqMn5bipT+N59NlCPw55M5a0x+gmbC/fCVzmpsfq/Tr/lD3wIV
uiGXsc4FLeIKh3JNUlN+b6uX5YoYxLf3x9avax1DVnkKYgoA9AeXSk6uRpMfYT/1
TUzZyhapJBsnKCdl+h6kpSnaoHERA/Z97RKttH6v5dKSwf/z4ec4/KHFuYikw8tr
egWl5dQKELrZfRmVJcf6wSguUCChXd1jT24vxLeNtUjnUeQNTpQhgNfcj+Y1kK+0
b6F8H/athG4Onjm4BJdtUUJR8Ka+L34j9ou/ass8FtFgqiloD40Y8ETaprZD7bPa
Y06O6IwoKq3I7uNXrj+HzWRSlKSnSTH0zkOFmUsl4GCs7iPEPQN2BP0Qi6cQ7adP
DHcs9puJba6QYkozsKFCtD+cNXgZu1APf/GwqQOuvWA9dYlr75s3XM6wuduxf8IK
erJCSgKi00wcXRO2CjjW6yu3SiJ/s0A29g6EwH2VnpvOZkZeADdmaen8ZSEIC5p3
6RCIl2PMvb95YYYRoaqg01isO1eEYW7OEeX9Ha9G7HS2jm9P5tcmjKdBvtJyW7I/
Ad1pvNiGWR1mznmnbaQa4lQfU2CS1GlMPUuPfJjt8ii1vrgWTS31VceP3Mwx5cqN
8UeJcGFVcQ0aqJElAxSYnEjNlt0Z6hxLxYPjwIaceGbYfXse7m+DL0Y0B417VA4w
ha4Ilgez2G5NuWW/LTNajDfLD5o+axs+jTv7H7P81AnGsSWCI/Mc16/EBimGLpzI
I33qZn5fU8mk9enMeow4C4JyD+qqfPJ4mksoLFRQSzALiCWx4MYLOE5ZXKQRzcgS
7iq+V7LQmQ+qOEWP9iwWIg9hgD0zWQ3t1mvDfSMVKgVY4wFqfnFwzNPon7/r6yqi
uXSmeronazHrd6IskrXXukwSnSo8yZESr57Q4Q2uALd/lEYkzXgMyjLHqupKv6RV
lw/U7sXKW1b0jvE6E8JfkjocxKHz4XcHpj5CCu2q9B8kb8RjTdmZlYqRUC1wT2xS
Es2lRwaYWhhHcMQN9s/a4wv+vv1tDWbmyMO54U+aXuMUrCtNPEipofMWClXtegqL
1PLPv79Sf1v4M+/qwxT7SwyDtLfxgtWrNPFv+mXBC4vSYIi3Uc1t6yp388kWJRcU
J6czOoXyhrNQOzHmMzwhItBh5A+k3SA2LkzJhUl40J/6j5kDqADNIyFbwY3nCGJU
qPmfcdQYhmjINS4yLV0Akk5X/hoY5zZAXATfkRN1wIoWVIyeMLMzk+W6Zt8lmQCU
reQ1uOQIWQswlVtSuG2m0CFIHE6a2CprmFmVWF5qnHHKX/l4m+2Agyoni8GvIG9X
0x3eWE0/EVvbJzc/lDTVWm6RrnmUDLcF4nzdX/XMKaHf/KEvqw9GgH6K3j2zycSA
HatlKzlevQ1Ti1UYy/cxPA0aczbWdj5746IkzANNrem9c9A/Rn3x2K7Gl8kdWzjB
N7pqh0hXHQwenwjziK+GQxCWNm+KPQpqkmey1qfRxEmhkXp1a/HLu9H1i69aymSH
a7YTZzS77pNU319gfALV6LL/OeBKtRzawWvMvmAiHnuHe21CQc4tIVFt/7uRhqwu
TQAJaF9xs65BhWrzlwoUGJdek/MNJMJ8+/P7F348DCr3bmlnwnVtm7gamWsX4po+
MLWSuj745B7c9zTwoyane+Frx2wu6UExLzPrNWY34LZMWR+sv6vgbMBmiqWeJx2b
kZ7fBoCoDGy2mxP9VKwiIkCstKuajjc02U9cW3huMMZjgoUjyLXfLeuEL1hZL/ye
kiw83E0Fl5XcI/4YdMwZFqJRilryIR07RWyTdj2aBKk5L91UL+PDTtcdRyPDfSUF
DP71szP8L35xV5VkZ7HNIdFQiux0PyT3F4QzjKv9invPcmypX2V66oQ3FCIC7ePP
IUofOtgCDVVdGA+uEMNvDBGJ8WbhYxuSFTCUk6sEcCZN61dW4CGdlFYVOeCJGcjN
jDARw4kcovjLq9z0YxQBU0GOXLn09JwS0HhhkPxf8BHH7yPKsRLPAHxYkxJllFez
sA3sZ1OGthji4XjJGo2tARV8D6vQh461TMDTxbHFfVXTomFMRN1bFjPNZzDKqJwy
ALTYLPNvZAAEy9vQPBw1u9rHmw+QE/8O/SnE82o7qCh4s0n0ROCnfl7bJPZ1CuID
yud4gbbx4b4iOQlgSKtnWa6GptDYf3AqfzOENHIroI23rsLsIO29FLP0Y+Oz9L6h
Noy3YsJR6cRI9nJ2f5CckgtRwBhvABn+YuNVH0SNfEI0TOR2KngUQxR2KT5QYyYc
k9aLS3y8iqwW3ZQPaIyEOGrxxpOvklJsbXGl0N8udhaMYPO6NJaeZsdJQ+X2Cf5Y
xb4rmUYR5So6G6QDc7rNpfPV8r408gFio4jkBA5nmoz4Jz+qcGwnhoQD219HkfDY
pJXujLFbfYxEwE8mdmkZt7fEva5pB/IF6CWvAUtu11Q2rdrjSsWoiOTzGCQewjO/
e+gyeyoJz6g/ZPyaY7ehFKDraWHpaZx7ZmdUmRh9yFFWS5W5S/A15vhQ9Mhbd4YX
7SyXV89Qy/qxSi5xSjiysHsyD69AYVNrkOUT4o9syFyttlUrJFJ1v5Tmtq4SjRmi
ZTK60jKNOgFAnHjizFaDJwhqvNKtdbe1vHVDgCVRdCVjMfwRPdjugrQiYJU5T93E
yM1ZyxsSDq3cJCHwjjXA9qff4Bb3GszOeIzg+zvyvyBlABqi8iWzp9Lkclt0fXYz
2l+oOjeB0mPpabMn1HwKKLXpSXdKm0gbpt8q2qPvDo43fBoLKv2UlKikmBC4LHG4
m6LReUOtbqSndybGkXg5mBjgJX3yPfXyU8c5g1RerCCSws9hEY9WBdSFuMXvHG+S
RrO4iEYVWKksCc5gYbfa4UK+hz0IozpxRYR31P/ZjLjv9uY7iGa5c/3FLOPRnn93
o0TpCB+SMkkI+KAeIAvdCnQqidgy8KNckFS+PCj208Mp2oqHhZsM4Wlwl1Jr21vi
5DM8Dr/6bqhtHBkPWHN/X1BY3EawnLiOZzawSSQNSrchaYr4aS6AlFXBIhBPUjBJ
moj2nNF426ksjsx4WtJ18x2Ho1EUu3/TBQwEpUs8EaTXl8qvOC1xqsk8BnEYnx+o
jT308/0nrcjWbJDr0y7ACrMuE9mGrmZ9HfdccpG4hR8YLHK1TgCaArXxS9NJMl8/
FuilXEAjoy4b8GrnONzTXVTXXWQIOQBiWk6o2LTA6uJ0fkkFYuvAtCrU/El9ZknM
qDhyXyHgx33SMOPhoJ6Nl0HNzlvv8vpTTNMvSPr9P5E2saPqmoGZZa/VZjrkU/5r
FrzlQISBXehn6KBWw8ZTug9R0e1nLcLL7I2LCWobIYmcvy/wOkXjyIfC0dFNIoJx
Z5kbrzJBj37KHHwmWNZUQFxF75XkSl9XKJZ9CzNhaWNHkCsuFWkVRIhAN1Uq5aGh
RhmEIQKI+vjH2ElM1JsEoGk8gHoBkJ1VCZS0XZouTf9R1DQdopHkx4DVq1Zs25N6
POnNKuV/46li3ryVB6HovPWlbM/igaLJ0JTFzgd2PfUpNIDcvLKWG9e9NkTyMdGi
APfKaj4I2GMRDIbaHQN/OWZDlmAfMbva7phRCb0QmtyuKo2GBSMg1hbDaJb4EQTV
54/FGD6bLQxUlcv8Tp8/RraKkyTkSCl7e0/myK0NA7tIQ5bhTGmiDJAx01WcEKrv
5bfyE8aS9o+QaS8CxBx0DpX7kM21TShs0FPJJ4xSKTfqizjsATPiHiuIMUUiIwy+
fS7MGXHuqGniEOGgHrin5+o6h/ZgusDYBpmOOpEwI2lOa0oQ4CsOLbzjizquYZyk
MOk6g6Hwxmc7fCrwaDnir+Na7sES64rMPx7sOJXbxou73JHCV4xqaMSj+J8RlgUQ
UllieBWhyHHLsM75rgtvhvaHDwajSwsujOHGzoHWXNs=
--pragma protect end_data_block
--pragma protect digest_block
HSGwpt8J8yDRC9VkHbkoPFgH/vU=
--pragma protect end_digest_block
--pragma protect end_protected
