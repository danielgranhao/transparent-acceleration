-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Oo0kh+P3FV2VR4Dh+dxkxw1D3TtnayVCm87qdInv/Rb38rKBVckY8YEs/io/aYssSIY4N8PP/Gi9
S19b55CLuKIkiptWXX3wENTcDc53njZb1qIgDAaKLyyGE6FmEUnlkDj1+BKeS28cJKtWBk6viqXT
BhCk+ylaohYKD9d0bITMUh8bn3evArYgX20NBNTKdJayMj1umQyxXSA1lKp3ux6geXW3jMJruI2X
fhakAfrHGpTGfMZWFKx+oV+GMeI2jh5+uVVLuGEuthUHG4BDHVjlqq8M7rTpcxA29CfxKE+tETOl
23BNK6Q+xgNalFnwMNSp5i/8Hj8peDIYB00mEQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4224)
`protect data_block
R10v+L8ndDKG/95/yy6h3T6avJ4j7QKaxKdO34kM1qDyS8We123Ig0Y54Mz5EH3bTvt9wcyeeTVT
leyNeuXcyHqaW0OFge1dDdHQkenvdJ5cqj0rxaqn9WdlsVmupUwbpGYfg8g1cuJ44mBgMndfcUJY
Uj7FZxas7kZBGkszxwsu0kEbP6FDnFU1tSUYtIFu4WNu3RJnNQCbVXt8TqvPlqDwx4jgLqyykR1e
mZsxY624wbvF4ZK0JWP/8yniyIoQC6j0w1R82ngOdHrqL9g/ZVzrW6EAzD9NMGu2pMUzt+zgmb62
BX9Isez6L6VbK/Xv9cTs6mVs1XHYHdOwlRjQxt1p+HlF27GZcRptN+RtKLBUfQU3ktuiZBev+Mvy
pbUziRoQzHs7LJcMcY9wK6927nFvtWMIculYlZy+yXc0z5Xo+MboU8WwyaaaQt/j8v1gGBKxlEvH
rINYSYxjpJITfnSdPmQx0v/rRQBGuLhsFln0+UXgoRuiw6wt06fWt37IMWo6RKPFeLLs8VLZDlgu
cp9/791/u5S+hqDkskQZJ39Yg78TAgjE6I0VsEPi6Spz0QjLBIOLX7rzxrQNDodpuSRGVPoXfR4A
nTiIVUDf1gmhV4mwNmgoSSN9AmOd6oqR0GEloMKgkNZOHe2yGiSOvuIUGZRtKIw9l3/Df9pFlgmg
Jg5Pqu5CueMfJsm8i4qWKO3Xa/PDJzeWyrRYI549fMoGwgT4PUBC8OA1mfQ9bOPfAitWB0wVnH94
cXYZufk6iD6MiKh4sI0PCbgR1ERr8nE46b8SV/97nchgrFm0h6Qg+se1AaQAwaqdfzo/AlG/ZfYh
g1mY9IiZhMS+Mcwp/O2K1D8PUduowvc1LC/n0WYaGzRJ9DlHfTPzCd8dAwZjrkTBB17CLyhZTVHY
QsuBjmkGsXn9dLYuUxWCnaH2Oqb6G3mEwXQB4fxxKmddW1bW3iV1nRMMRMo1ZUVBOGTR7hpbTNK2
f+j9McSoX9TZcwfnisYbBlo/LDoeAJXNIIqgDVC1JNp6yyCt3NazTBok4KFYbiQ9UNp3E4ZxWnuu
0eiF6pKNUFMqnmIdxWBkz/PeJQbZ1tMAaBUXtULBX++gs6A0t0y4emt3aX4xTLF3xJujhuYUsHbz
nZH7jL7ddEToDP0U2Ss3wLc6x/2n9oNf0feKSly9IhR6w5VXOrxtAjab+8RBJlHwVGRi+foX6OMy
abq1lxxDZv0aAXib8CqECK+BSk8gGtBF7lSR8ftTml/EEWWNbhYrMa7QY7WqDHmVaYKyIUsFPBxB
s0K5pI/juHQzWal/T0bYA9TbzKF1nN0WqeYQKjoFXCi2ofk8WURc6FlwXJgyHh8D+MPfjaNwHzyu
YLcykeRpRhU196uJfa63s6VgLndqfjhgspo56F1O8igHVa/dYfc/eznYznxmT1+02XZqoBnWFGYJ
Ibh/fAlULqEGpeyGjijn4SmLDIqEXZ9GYqKKIOU/IE34uSzVzWMBc9ZKfYYgbSNDqsPQE1mhRDds
cL47tJpZ6I+FJ32A0E+/BGjioP2pMufZrefTviI93Q0lSfH0SXyexKtmDv8wJfLEOgKcbIqzCdwW
fzca7rbg0v34AAYiUJHpwOEBmM17FAVSlDjlTU49fuPR3W3H11HdQAXKY1YHTCZEXz9RdDncHYvl
seeCTshSG7LUtBaKp2c5zn6/kmGltHCibL+ehblrMqeexDHAmyoyVQtbg2M2TV+mlPSQvikIwzaZ
hamD8Ys638g/CCN/f5rN+fLFgOz+6culs3qp7aIOlVKvigQ9EnegppISee6pqgBBiCIbw/E/fL3X
Q3rd1ziRFEeDxAuNwQigoqsvQlo6Vo7VhuVtaHuXiRUcNM2Xm7Gy0lRdSWKwhfuwrY8sRjKfODTg
gl/i/x8BYxSNeFADMg4zjo8T1LhkTI/gR20qgBvdegzD7LLI3RaP8KFLB1jSaITgTaPMK8kWzi3/
Es7gisUNemF5tr/Uo2GuUxeL2Tj1NG6rw94J2XkNKTh7FCkjVkSmavVlR3aVDe9T5wbXbOK/lSug
PlMMJI60v1K/d00GKmj6T9aa6dVb823jwJDUuIEBwOxqQlO7yZ7gTnDPaljIO5AREizguJHi7/vj
wTOgf4GRHaeoDhiUQyg9gF9821NuYEOY/ljFUZqAEBWs4nxIZD5HZDQw5KI6dT+HD8W9sr8hD9AE
hSHFCBUbmUPRhGigqvj+y6pc2zG3XTY7oF+jAAr5sb3JL1m0mwPlSVlcorY/HmKfK4qzlAZEv0Yy
Hg2/08dQbiam0Db48oszwzamI7w5NzUi4lvYJw6duj3uRibduKWM7Huu/HPM7n5c6m9uouzjsbXj
5iLuy0S8SGJ6lc61Wb9SkQ4/8Hl8YXEliaSq/OcjEj/F+5RhZ7aHGUOEi3dTa86X8GzO4AaZvazw
ByCfU9Two3kr1Cx7ImWFpaS0fVQLG+5TDdwJrgLMACaXIGqIvGd7rbESKHplMzVv/D7RPJBDHrmh
7ZTkGVzlDH8yETbpisQQNjczKNOVGL/0p7A+FLAkCKs22qnOxQ+6tfN8eLNF4vuXV4WCvpZuQHK1
Gc/ZvQcseQKWw8lt5mdHoV5y/JtsVQLI664ARFNK3P13fiw697wCOrTsBjuA8dASwR4mf70uaAbw
7Yn7Gjwus+K0h1WZ4xsecKFpF1Ht8dG12XLfiaR0U9+y6KhFLCrAyFPoAzEN52Qs0TGcRc3T6675
45Bq3SQr9hSG7Lp8k7I83pXZbvBmc9wiJh85kDmFU0A8FDriWdhfquBWmtbYhmzeDbDO054wONqu
6BevyYb2QH//aRg9j2m5DOzOmkZsidwnzVcBZ1GQsyCC/mnbSg2PclYg5bob0VKLbz7gnjaEd0/+
AXbnB2a41fRtsHTU9YjY6Xt5TIwTBgMKdUfiwoRubVvXtvpQxi2zlRJ1bjh8onP8px/K/WMJ5X0z
Ildi7UzPmNRtWtv7cCOfWXHPf8j/QxDRu3MzTHtby5DpLzefj8j1QLWNSUNB8TZOKIqlTKVtyrCx
5qPNvG944yIgYjIVpICZ1Qyb4sHlYPuviC65z9k0uli+bjb3kVlTdrrzUdU2vo2xxn9GXnr8dnG0
EMxHS8lJba+ID4Zld6nmDwdUDpl+ipW5+hydQU284KwAWs/sRRdBrnAwKqut4jaQp6YW3NeON/8H
VXGhgE3vcB6Kp1Crcuc2X4nTKWhbulvydv67E/i2+5/rCmp5Gf5ZLocWowneTkcBHQM/f3oUaewJ
N06XexX4qDtTvX8HTvh5d/JROoGXlCHlPeOaFvM7eGAnzqVw4SOLqg8r1toirekL/Bu3SEBnV8sg
BC/d7OJb6qvvcQhPBIL3E36JCl/HEGv6UuIX7TWo2bcAUAm1v+Ho1hUsKuP+pzeyGLPFjorK1qXo
lH5MEGpbOJCRFYhrmbQb+r9lOUwptihrNqeQeRiyoxtql1j48XkTV12+gsSBJQDzDmxrIYN+3w7/
cYFyE02HMR/RrXpJ+Cj7Or6iciAxQGwJbQ8frZ8HHtjaIYukCXyqZ0KV18CsnuDznBpU3GR0Hp34
Q/pLoaVphI4/gyEYlVMNMySTXfpfX24Iqm3l2z0Bde/eRDo1R2K5qNc4WNf59eq8fijBkiMfpCjl
PSQvKftrAWrldbZ9VW2QZkCwlPBGoXGgYkyQdsAI7PMJxHrV2sEO37xvx6kwpvPKf8cJsPwDONzg
cuWrpoZEA8FwDloCjg6Ag15AUxOxru/BMvApxFwRpWwmr8lcchz/zE69QiEPlYEX2kxOO/F4dZzo
gOk2uHTyatE+G1ghwVN946as75s24ZU4MKJdS0mcHZgrevYE3yGJ9Rbljivsd22RWR9Nb0ccm4gH
bioz7tA7GLT5SIpAQkf6BXSU8SQN3hg4FN7XAHHKTEgdr6Kcd8JnwBrZRjQMMMQrjqTSoyxrjVD9
nTYwP9b7bcT8zDZfnM3KUwpEYaSaXhWQ6vRyHD1D4ULi9UTHqwSgHBzb6tIRD7utLt4JYCR6zXpC
KQ3inhhdhfAiV21mXsahbt1IWm4yq+9YH/qvHz8sMWqO9XQ0+RZkca4Uo+tGtwwxZUAuf8bFii2Y
eDF+J9Q5m3kGPucPLrHPBE/cdHKHRSb4phahH6dqyzICFoSYY8H2WJM6mMRpwBbuN3R6wzNqortA
YLeDLUv0pxkau+lHIyBKVI7mNcTdDGQQhi1499QApXKbd7pWmhVgq46OgfRddcy1NaJ7tPT8Gn+w
mmRHElGoU+WJ6V+wbpydp8kFfxM7b+1mZIQQ/O4kjtNm9kv9p4tXlfcE4jTuOOumpFg6ebKF8buj
xA0WcLF4Fpn+UVeCDOSqF2R7xX+mq2KnLL8YYM4lFC1Lt6ipz8SmN4wyaJLWNjhfTd627DBwbK8L
wPLpVhaRZuYqxSBM9JMXoJrgrQlicxUH/QYiUA9gCLMAivHtyXaJkd4toCcdfH9qCZkYtd8NwPP1
ZFBHvJx7W7k+3A24wdCTyZ0APn919q3rjHBmppTH4LUVut2T2fwdqwVsr3+AQq4GFhoMEiwL7G2R
Es6wZ/cfRQwwM5s9Nx+hIIPIvN5jT5kiHZVTQobXX2RXhiWb9xqeg1k5KlrFK3uQGMPaHS1pwogD
O7sSriVBhB8bgnBvRv0JxWOroDeJmcPH2YoSPB7+lSbJr4PKsv+0JKkFnkjEhJv/gwTPbdixg0sf
65vCQsRb2uxCDF2i90HX9FvL+c2oXf/qd1NtzBXDYDz5eI07c4kgaYBEBfZTNxr+2SJ6e8jhly80
fFkkR27B7zbYkTF9WQy8ttrST3ZMdOt4T20aC1ZEvxLBuCJgK4joaswzGA3FecY/jkvKwYRRMsfU
P46430RZrooa+wEDdqPtconaKFGpbCH92Q+4sDAHKPaZAlcDeZ/JeNxLz2ENi01fmww6XXngeQZI
3VLPLLDYbtkRMIHDtLisQGeFZl1qg98WiUJk6LxA8ZwY0//f3x+A1HJToki86E+n4eTi68DD1L6k
azx6GwIztkIF2l1ZeYxfuNAtN9r3IK6701oDtQfQNw8btD4J5IaZzFnXqx+Os41o3cUUs6N8hpIY
QfHeTs045hfqZpIWg4RDBt01Ao6yuZUZQgiUZ+3UOJa6Dp0ufgtynF8Ik934Wabu1hS8l5n4D8rq
oa/hpF/tKpmEtEfddrcnH7lpKEhDjMI0yNS7Z7t4lM/dAeCFU6fEy1adS9i9eFUF5mP5Bv/Veldi
/WOlnanUG85/nkTtw0ok/mowFXsPMDu19c6ux76O01xwmfYICKJxaVeIMcUZdWAF7vS+vLciBWDk
ai0Lh+Zzqmw4fL+elCkKXzi2ffNMKFZue35QxmR1lhQh1cCMF3VpdRXwEkbaRPd6dwxEVJgJfna+
1HDclV4Ytpbuzzl0p1OtZqENCpPecwdEh4nAyHlylY2ZW8/hYjOJmLdVNu/25CpQd2Hl9wwGGxDq
PUfp8cM3g5kw9ZKiZjSJQflRg+n5yvYpbrNu+wC8UbzoMxHlsaN2vlHkP8lWxwCqYcd3B1VV98Qm
UyD0FhW34t6IQTJ7MSFQqCd5UreA5EWJ1XwBGZFKQdvAsKgSu62mgBFgw6A6bPHHcipZYEyHworP
pSWrQYv0
`protect end_protected
