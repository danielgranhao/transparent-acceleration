-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
FF0YLIrG2rOa1UwWHfyBDv1ssMleAsIfdrMxtLNklItO56U/xCOXG0nq5JZRuHArnvwiMkhclTFb
U6PYnUdjiMGG5e7VCMpcIYRsYA9RMjxsq58RYVlB+9jRTkU8TYHnsB8pJuIHMrcSPEW8hBtOFyI0
paNLAsL8MNLiXBSvKlEmsRsB0r6TdVtmxTjXp8XbZtXq7FL3DXYGADI/mMO91zgD8aN3/iEbo3rG
ukRUJpP4eDyedBorxGplQBtPblPIcNPzhUi0ZUVXmHMJycXpTXC4NDiMrAii5wb6cajoxYeOd/Wh
u0jlJInQhio6RnNawVrDpQxAdQc1ZE/xdEssEg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13584)
`protect data_block
scBGPV9irJaIfDm2puwdCmWTRARkCCI1KX8NfWBXVGy4BEV/+oAs3dC9tVJcult2i2NxIUsLPetk
SveyEhelBfVuZIHzZsiKuk1cudfFhybNdGzwKmI9iHLynbp67KuzXxaK4sjG7P9G+6oU3M8Vmp3I
fdiZxebkRMzR7IoHPXifmL3a333p0Ozq8a61MI6LTtyZ0TwXA+5EiLSgNU4aC8uEMeC0OfvOPMHO
CVBeDU1rxX7q8ofhFHH5aESYITxD1oMwPKZoeAxpjVEK4CbqykSVyczkBUyukDnDT9zN8Ra/HGE5
P5PhbjW6DsSyF88LXBKKzZ3TCv+vVFOXw/4VgHrP3pFE/6lcjNNBqcJj+1QDb0BQS2KlLIn8d5ef
kfAS9x+LVrJyyIc4fQX2MGujX4fXwVZHc3tBTb6pWHpHB8uvlxuwI2TxfXOQoER/tsuX3z/3pKI9
oBAlvqjl2rjpLO74/KxAYVFiwWgkhA+SsMzg5GVRro3AHZlJTbqxH2hUSltzU95RGSXOD7BYLNPr
2ZO0FVW+UouBQ0BjLgKL7P58+7xI3LRIH4D0qqC2CbC8WJ/sTs8xkvtCa2EqQGacbCZQ4h0SQ8TT
0KMS6mp89ya+UcKAzpY7yeuNGhNHCxKzg+WYnXLGBIHemgnb04KF1ZBfJ7Ws5KE/xrfKEsg9BDCO
3A1Wh+p9+ju+hPY3U/OWRzYsR49e+Jp1T6I7lTnANVen3Jx4lwv/xuuW+hSeggcY5xD5Onyf3cGH
1wIr1gCmiol0/IaLSJYDFoGhLdJuElaDfP49+WMgkLSkgIfxCbXcklldxJPO7IF7itmEHyZsw+Jb
tb7jhrXQmv+lA9sROKJo0A+X86MUnM1VqOUgkpCQmPB0o1CphGUl8QgOBe+UONwuujjPc1WqzIpE
l+bVJjYt7nSaXTFkyT3PBF4WCVt5lOuYuzSzSyNozbkKAM15+6Pmk7C+3V9WUJrxO7lBr3Apz/jV
rDhj161Jqyd2lE/hZtqCSYSpp6fcDELaNsvY2RKtPmua15h6okqPcXyPKmrQVrqui/6ZBEavJ9hU
O0L0QgRVHAYxzaCfZ3RKDkk/hdGwZfV2NTwinCq0BUCq4LyLen6xgSsWNy6fdS6hyvcQNknPUxc1
kgX8WVnGEEig4NVy6fKNNT8pR51UKfByLm2XhkE/DeqK+xNetEIq5Xe+Xca34xmLaawfBnvBw9aw
OdID7u/3FZP0KElfqzfWjD50YdPLMB5igoKjwV9ZNivw7qdRvAZ3Xzf5Qsct0kwcozCHY4duVeJK
hvcR4zmrwmkPyLVAcu7u2C52vzzHA1GyXRUqIK02tICWo3YpY9Y3GMpX/mKEnX7VcLFDI5fHfd9q
cs+3sqGpljS0WRAEg4cWOEOXqUByCSXg5g9olI3l+gF3AMxgAvl3FYfDMQvgeiQj3pKXaYgmCiZo
WhT4OPHn31NLqz5oUeGPEtuCymaoum4kSa2GJdXWTHNflDEuq0i506+vf5qlRjvkg874r+R7Wwjo
oQLqrxBBPtkb4d9/nNrhscBgREsvv7G5jcWgpHjv03t6Dm0emCTfGd9GhGpy4WQlJwKmxUFXZ/JE
Q+YkpBd3a9qFPToPGLG00v1pFMxH3wA47ZItE8BJuerrOQIoXkTKCOetm605LAx76Pb5B4FJoIal
cPrib4Gdg6lHGUqIcC7VGCe2VDC0JZfzcmvYYQ8MQef21912rcfuGMKfZlJQzaObxMuFLD20XsT6
FM3nomSjqhr730l/gEu040Iunk1n9Gxt+lrJHk4eaIT6PAryAN2F+GT0hW4CVWEDeyUeqUfcj4hA
R/sBj1ZGgqwOqLP9CENRvyPp+3fyl8jDoUME2JpGoL7hVTPHLC4x+tOfeqkuE3JqzJCYOIka2kLx
Bpb1jWwx+NdcSmvCMqLr0RoY0Gl4cRsfdGfLUmzzmQiJ5iAcTUGtBKvkSv85O9h8Or4UAjSNloWD
GcqraEq3ONX4cg9q4NS/AxG7e62me0o4EwfJ9YqTSCzz2YSSrx+Db40wsAPwbG/ffXutAkq7yKVG
lfPw1nn4zNz50mLMsnLRc8j4tbV1rc3MvyUpZX10VL4H4Vc1K1uyYiUV1zOYostuILAcXD6c/q3O
iqGYZvWcKG+vFSjLOmjsLZJ1VncXk8gU/3oNhw+flfO4GN2wgZzQpY3BhKALx/Ef9A7j6BY/gdhj
J8/mtn/xoEc3Hzpo4W7QGy/lX1M+NM2WtxkWoC7AVVcjeT56g/zome5TVNO8QU6jp70B34Uku90Z
wkmI8U6IRMIijaMZgtl7cMh9PTXX1ndYgMkJROsbmuzpXQaMvMhZCcaAhw7dyT4um6VzJIlVhVNF
v++6OhiWcBV7j/hUWriz2PO/q11GApCxvBhlgxAsP0YVO88L+q+5URlwwAVwMp+LXxGyTu6Lej7A
ovVmOexyDM64tGhCnu3NYhDcWQQKXcVAgoO9yzj/gDPdRaNg18LAal5xNQLt9KX1Bg1C21RHUYDv
F2Zpl4UHes5a25egA7zoJGndWEn37R+en82V2h5YU46EjHq4SSnp4gGKHClmqIcp5c6KtWjtIjBy
BHOZziN/J3AoK+umQk8BUy2s7IuooAIvU0ZDmi+4OqRC60cchbAvY3oHQYw9vBGzd8k7BPDfP6ZO
NkRGN7/Hu+IFWzX1mTqZAQH3f41x39V/MDDZtmQfms8GNMqsyY9QCYMjjQHh/HI6XbIOAk+j4B4a
mgRcIHLVUjUtoFlQ4fV105+ovpXBbsCOfPVJL9Hs7w4NLcbQ4bQywNbWd9qdoljPsURAuI5+5ZHm
UQ0Fh+qhnNPQiCMM3w92gh5XR5w2CTuqhu0eklxULYuLzULFHNn5Wj5TdmGiRYQNsa/3u1JfAssi
fnFqTyYsQdVm7A5Ghj5Hm3mk5/0ek4ct83wNZqFaBJ9op1DKMLCD7mTtXCeqg8SNc77hKiPCbGX2
MI9NBad1IIHJcg/QbXL+Qe9HVgeuBAXQSRGdkHgm2Xt7dpQkEd0Cfi2U+5nMbKYqb6VlyNiIwXcG
KFNStNCGdC1mgxw2VZFrdufu41YqhtxrjVr0bpr40EGEvzsfDKtFPdcEg6DQZpbY6U2D3DdLXSgZ
W2OPoY7N9JwmopC9KxiG5uOTk9CzD8a79Ga5qnvN6v23+R6fTi1gfd+2PYZzjUGpr2BYwJZp7We5
YVXhBXc97NgWiMUYO0ALHiIANpgBvbf6hD6Py4Ecj10VpKNC+otbgRCUVd5l3ITBlnmK11KtJQrp
xVmTbSZQ3Yt/iPH4pFTQ2QDQ8FcS13xtQfuLMXmAdMRgGX4IFmgUBOo47Cm/H+9y5YmhFL+MUGqd
WVko7f6jPvqtzmeA1JaX7jpfzzLOrgl/5YGuP/X3PtXASAv8OjlIdAX0pOmAPeeAV4Qid4ctIoHM
fzRsZpT8BdbKk7I/qVGIf95OOt1Lq8GxhLV5nU1TP9r4ZAfLOMTcKIOXcJOwDlqZYrX/ximBjU7k
CTgACDMGhNnJFMGjLGu4mEr8ClnNWt53ndWvejsNO1CJMo4F5W91as5eYAbIJ/z1FclBA0xhErCm
0jjncw+8jUwiijPQHc9IUFTydbQCn9ckRQ4zbgprSKq1CA/Et7gOVBPJJH0pBUlnd7uR3AaYPJQ+
OQCxm0M2Ckv5LWjAjT8lkkhX+1bXIYWpocmqxRuIvGJ779ZelWnwa5UkA/RFodQNOhWivQ0BPeCJ
nXwpX6+fe8rTg1uml0v6NOXUI0EyTLH0eFuJdWNxaCCoyp8s+4ok2tSiYGNn0iLsjhLidDzKBVOC
Lq5I68qWcRI3EVhNWQA6IBOAVjKzC30ahUHn06g37afZesGTF9pLA6HrZvByP8DxofsPPqpRP82n
8yBK9UN6KRLft821xEwjCDog1o+wFhhmmJ7cjzwNqlTKNsJa/zewrsxYexsfo40ltsUvgdXgEjAR
ZIYiZDjQz9L5iVGvQxpsIhJRkqMjGaUl01Olv/GvoVGiWza2EkMWyS+RBrO9hC4Q601rm1bJJl4g
9PuR322K+GuZKTFq6qpz+GAVDnzTlPh83KVl3CdUnqXQrS3HU9id08MtHSUS4naqDtOiEIL+jN8k
oDh6G1cIf68wAvJLLkvQle9frt/U48ZkP/e47ZVO0CBRizZpn2KAcl0mfj1FlGAVcbEwDl8ZMmQ9
x5vz/Oylo05R9K3/HicnOEksalbXDEdX1S3u3nvth1dzopE10+hDjouOOYJr5LOtmQ7J8Fk6VjLF
L0KLLmXJDWfuHh7NI2Zj6kFDx/+xMituJFdSPEf0jvBJwh3FAxP63ttJdwlCLTdBfOppF06YQIXH
rhtlqDw6x/aP6Rc9OTECEfA0MzGe1j9dwrJe1WjGFOaeMdkp1TULkJl/FAH3PagOih8sRto0kki6
7srf+Ds/JO6dSaJyRcm+hcvXBwBP/X+440sp0VoklWCuAp9cpm2rNcbEZBW+mazI6thrBjJszkwt
yvZMGFPdtuDmpknswtXQ15tODq9182VgFx8mk+/RcC1Q7xdzeTsNGr/EhV3l9cqO/gqwz5u0DtQ4
dMUeZVv3DezHk3q3PH+TVMbN1yAWZ1iY3kXt+2FdX3Cy2mHzdEOKqtHDPdwJkhO8YRbbYjftcJoX
J7D5fx7swGzWGQkQLfqEDVkKmlURjoVzu5pGXlG3o7AXJUSzJ81k2eNzZ2m6ezkYEWdXqlS8xbNj
tyapkAU5qs8IlJ5E6/iEjq0fZJsRRWr/qJaxfVXi4En6vQFBrDcrix3lp1GevRLpgY2T3CDj7wKr
DaCdUenhpFlOqhP6tTf0Xwb4b+5EiyitgF0A2yA4rhneffJOiiwZqPidL2fFMk75guo0Q17mT5XE
4kRrmdGuF2ltesbJW2Pp36GUXzZVrn4zx/9DXWjA5abXyORnUMWQlSeQjWuQADjS7rmq22lFGBIQ
ar98pXN7VgbMr1GnTUsIwQHYnws+mhcA8opDwzbFR300eJx+TpyOgLH1iPCkK2zRv4wIm/IcChny
7s0mk8f2VKeS/QwZvsiS2PkJRO0wQoxlwp1LAm4JXhvkNy15+ZyuDpk88CGMzXPiChSuEwX/z96Q
ZB+sjuO86CJA68SZLSNK6vCkVHPFpuTWaanO03oMFfAGjio0pJXWkKfg72U4y7xtesV/pXVf4UQh
M536yjF4PyHK28TbvZRYM8M6xcCeuZyBdH8pc+1UnCwaJ6wQnAYERvu+vwc4nCMN1+i+i6adQ6XU
ciN/oywfmVPrBkRslW0D8kgYtnGxhAwP46BGkq6C8m0Auy8uYV3VvyHLQ55WJSfmUDGP4lQ/yGgz
oHvY04lgTgGWBighbE02UFnZ1ibAuyCu7+yPs/gycpIC5Yq/FHA8DH7vLBLNFLmhiN59Asde2hGQ
R8NTbtu1uBi0lIauzWOe8AeF8BYtv6u4PzTXi/XxvrHoGl9RbXTdG5rKNzqDB1LTS0sQtc1yTAap
ONIK2TZFBp3yMdzxlMksyzlHkdBeulZ+18RPbFLCh/vR6MmTfmTb7kcfRSyOiIwtpU2i0AfaTX+F
YY6sfxn9R/+B8yRX9Mn86Ek2iqTFKTgX0oXeeUuOR/oP1WKst01elwe3fuVCsCI7UpI6r6Ezuh4x
X5fQdRaYmUU3FLjLX1BmexYEvLugd1FIyjI5NgZ/ibAe2eEnNaB5KAHHFxXDmWdc64utUsazOwIP
6D00++TUWWO16qOfsG+aCAqpqByNr53Xemv29jOIifDBQfoQV1mqRW2WGTBZOBY7DmBbYVhi3OtC
kEbn33OKrCT7ut9HswnrNrecjAHhhfDrYoVaiB/c9bbWZB7d76S9zqfmg3Ikm3eSmmGPCKFs3rUw
gzBenVyGoXpM0+XJCLdrCMaV1Dt+jmb4Wp31kyXfvy4H3yXWWaZkUOPSA188ai9ynax4MajryNV7
3hYz5hQ2pRXPbCzavFSRTZmgCcMpwQQQKYGj0XYMLcRDXzMcGZO2SQMaFzNcye/qg1FbTk9hmx0l
Kapw+qvGN/vueZJR+Z2Mqop9kjQl8OELZHZ37CfRWAZnRop4kLh632oLW3QWDR/UXYuws7+aGqU/
kYFMlt0plkYYOAACJeHdfkObVwSKfbUnJC5eJ8/QfkgNJIdKPUJDjC6aImYak2dWD3Gvwal2gph5
RrvD1eHLMI4B6RAoBSLz8YfGOL/SMoDn13RGVSUVpEJ+lCykJ5APKZAiBp5qt8bSz1JTLPwDoH0p
2ioeuxjan0r7LIaJVGSOLb2sMk7fE5QsYeTcKxkB2BW1bKiDKiUIV70Fd9DOPp5pxianiDdo5qn2
v5YZMu1cdHjt8roGtd8C9QtveAIcQNNBEA9kHnzWazEr3ek0KGiMEAnqbPjftRtOk6lReAtdYUTg
xAt8hYFVZ4Su59vruFIPtgnk72EYMJlYSpJZ5nwWstlDs7tFBjM5sfxxiuvb7n4fiPauFJ/BP2N2
uHiM5E0/w3jf+deIGYMUSaXmIaNx5JF5vagSZA/n1rzX4hJiCYdkW9W0yO/VAnQCsEAxgsHvMBhg
LeO4+Jiz7gW35H28/jxv8gVqkJ6Mp4yEUnyGUXLKXLu5TKLgOGVMQmiqjpnXKhEz+Kpe8Pg2Vtfq
HC+LhI2SQNBolTZJaeDblrRwKs10gpHifjcvHsxgOFsD0tvVDz0XF47DQIRBJHpJbXpK4gSfLYjI
pPcp7T6FOONrIU9aKGKINGU31Q15ASAKmjufVzSiKrRJz50BD1sbAYhg6gHDJN5v0bfhzbxXuelC
znM1PIzksQleA30eR4J/n62oMPOZJAFYWJnjdKiotop/lqxjOR/p65Wd3cCSnzj3p7QS8DNqIt6N
H9k06/gC7CmnXiwBelddwaOriXZlrLY3ie7SAIEJPMP9smJ5OaG2id6oIP5Bn4UPhtkZe17ayjqR
RkiaW8cGjWO/enGeKRUrGMQF7U1ud7BFfv0ocQfY4ZVE16Q0g+gWRz3BfahIJ49uoWtRbM8QVnSy
WCmOV1pj2Ldy0l8wxdLw/yvnGf6cisVdEeIRqWAMMM79WMS6CVnrayS5oAhsazBQelXD7cAVll+H
hZT6u75R+MqfhWq9PpM/ifqzs0N8CLjcT9c5LUHGrqgs6qg67NLpTMc/UPbwYdCN8ZckmcTaqAdF
X/2dvrfU83kZX6slrjspu5Ue5qyYDey7W5eOpz+VV8X95cbA9RKaFyhV00CGdU60xkgoGfxp+EKY
9LRQ3mKdFqGPUqld4RaNNCqWKo9IiDrjtFYguO5N2TXIeB3OSDFPL7bRBA7XNmQM4nWw0E0Y+HlB
q4AiV1DQ4ubHKNBBrtdPMrwpW0VeMIU1swYCfL2VDcKxFbljfS8oSP2JpjDUXQxTM7wOE817KEjp
hzSkrB76Co9JwdFTY2av0iSxcmK6c4VBlJ+UEmbQ0Go/WN5yhSAzCi/hsT/AJnFqqjJh0G8I5o6n
I6NQEPxaWkj3RyhOuY9keKiE41kKZdaQihoh7dSrRucpL9HFUAL7c7mHmbqKfcd0JbPECgvDQZBS
F84mvkk6g1uzcEmeoNg/gBhs8tim2N7z2Pb6u1rT5KwiIXUoFdxQJcNm/t8aZFicmJ/1tBpQ0bmf
ire9/zbt4B1lJYsL6TvL8yjLNIetE2qGi6BQfaA6R+K7gBbI4PU2tZcE7RlgUQVjtqL9eesZG4FD
1P5YiwPC6mFxnYWjiFhARqkeLsEXO6C8RAfhuSr0f048iBiK50sl7WKvwM/mqvyMJ7iiKZTZuMf6
xx76hNQknIMei44odQFu4lB6QUenrjNxrRteMg2nrrfEhRobQ7uT6ch3DjYTOpujJWATZvtyGeHd
ZcmNkGjqi5AnXWw7fheQC32akECWGEY2ku9cqDTLw207OgC6RiBxhEwGz2md4HT3oKYKFKoNTt0N
Mv8ioaZ35A04BtjrHr3F0kalUH0OtO4wKqzA9y+q6vz6oJEOq8Dnt8sAf1L+oSJ06+GqH4Zez5Nb
GRiNpeIJTXa3J4lqwcHQb7X6kXSAwUxCh0J386DgmkinIydNeyyy+gGcpTwNZPQKHSzmoSFwIzid
LZeI+VHkgIJEVoTzdfYFOArgKae5cYFUSDCIlpquH3oA2M1L51QbV1knVFxQMc9H2pGcanGCOKcw
irtEnL4fB5qCd2fPVwEb+a4YU8T9DOo8QaGBHqAVILuuPeUuN1yjVxwYM4/13FCg9zizaOK4pAI+
kAg5p9gtVJmtMN3q9b1X7SFQnKbPTfa00VZHmx7Ia7pnIJ4pC7CGn4RziQyNs45BSF7s5X1iNyP9
n2UEvMv7uETUo5YSohoxtYPDSDxw7cdE6xLmF6a6FjvnAoiVnOGcCuC4TAu17Pa9p1XtjeiCUTqd
n6ALEv08BKZvd2ItQ7ARTvtd13x+3PI6MkGSepGICpihPLPdw0Ggmrija6IViOEEKTudHeoy1mot
ovGDH3s0Zwi8rcBBjJaYEtj3draWxInORXJbSf9RdKO7D2zyi4KkhBpjM5nKp2Nl43ros5TcEBis
+mn+saB2PUA3LanY5gxHFUUEFk6zPctyb3jxMHY1dJ7j9tUIDIiQgNvu11oviqqJWPUP2GHqezgq
kXecaxuTArzAcmf/KBhwmFEdcQdUItlLXSJirgPp+shtJSIXPofAszGkUJG4l3d8iVVhJsKwX9BP
6oRmnNmIZEiPmyec0Z1DVvuV7Be6uBeETaH+5r6M9L5mPIYVg8kBKB5bxi4i/eYrZKPKKaCDQVwr
Fguf1ETPVBIlJ5E2L8u9VEm8qnzmgJFOtCahBbHccENcWM6DWymx3rsc7MnvpwLkAyUcL9fWTd8S
Mf/if3aYVRwp6SJLAHCw0Giu6Zg3oV3dg9SS7TjZRX2ZIu4XJ17JWTNcQIPbPTG9mb6eSyPAQjEa
71IAjEvYUCF6bU42bytGV//bH+RlTEO04U7TIRGWkn0vh3a3VWKdcMis7oqobT46KojVtherjLbJ
+gs/Wob/b5WqXJSlvg5J34/j1WM+9QGOhpKZnD23VCIxsDa7UUCA3WUUejINvBa6Prs4Wt6NUgII
+Hh3OGHB85m1aL48abtEKAhzcqdHccQAAbMJEtVm9QIr3z6H0eGkmTYukLo/NpLZBvQfHvj8EAgl
xg1hV64PwkiIJeTT3v494/xZ+wip63+D3J62RVl6Mr1T3CAogRZRbz7apSeVujNW9ybVcOBOCvx1
/P0iJ+JvLr/IX6IEs9GohiRK3hQrihS5GhaE/A3EKGEaI7a5t5mYA9sCm95y8TF1jIAU2+nVuqf0
y4MYQI+Xhl116H2YkWSYb6NJV2GHJ2m/wXsyyIhJzK4q0aNrbCY0WKrkRK+Og+HfQYtLBlg+y/LK
Pz1lAKcI+bgF2ndy6UzV8/mr7pb8OkOSoFC8x95bYw4tdCaphV1JMOfyEmlCT43dyWrMwNQ7FR0p
qKeg45Z9WZ2BwqPKiyfCsS/YrHC0h82eHWjmwIMT92d2ZAMEsI4Di6JhGhYLLYfra6feW+CaOuG3
DBNYOGuNUYB2nE318IWcpDIUdFTVLHpsKyCI13FWPEVL2hx+MHZkNOMjth6mtGhFz4d4M3tDQuqI
ix7uNFBxLdsYhvqQDGq7EsMKEXNdby+jOetB1RaTSaXiSOJBIag/HNCeX7TYwj6YRwCAnFEw+u7r
e4A3p0+7FsiDYqIRp13hHvUOhuwMZlRlNAudt/tARRGPCBYknd5msOj+ywph89oyLEcin7WZ9j1W
f0yfwYeK6VWfkQ//9vGs0N/sKn5SlPCdLVyXu8gstXO3TRxNUPf4QGia8i/n0t9hVgW3CzcRwCgu
1xh8v024K2cnUlLp6NyOfWNazCFwu/5+eJWP4q7G7uZaTdVpfmoreQjJDFzeBy8XIOe2GkFYvu9H
LYZmiCFBwD1xypxE53QWN1j5eidY6zeyEPtEfXj/r3pFp7uW0EwZDjQGT7UJCF9DG7CfUv+IFDOb
DjfvIen17aAdSJhGvspBc5r4QC6FRw/h3LE6unFV+Da0gTmFgrQybQdOpKW3kRWVgBU/Fllk6s5p
dru9vIM3znYP9ti90n98RUzueOtSWGIvslZGInE/SuUShw/ZwAqF3WdFxQ3u6WGdO5qsfSUlq0cU
CaGY89+ksgU6ODTyzLiNqqS4zXlq+buTGGaMPFDiD6uD9JKv9SxFxRbw8blPXji+arfN46Z4dMxL
n6ydfzxamWGuO1C0i7SQDMg7fxwj9P460cCdbjo3zxs8cmKrlpKSqVMek3bI/Y6UBDg4bGTqa2up
FR9jTo1NqwhvWhdO7vKLaAkN/Iz4e47JezX6sVU9Pc05M/bB5lWcmLFVKJGsmm/5ZYJ/DqNO1jFj
dq/PdA6J5qOqsQRgNEs14EFGaxk6fbUoa2Yk3DvtuwZ8W4kKXAtQD3KLgX+R3IOBAAqeBlxcn3+4
sKfqYov3zANmkw/a1ISbW95/05f+7zCF1VpvtMf7n76ZrAR/3iBCvhkDtWWvr6lq9Dzp7/RPcz9z
9BAZcihvzw/PahO2WfTJON9VAVa0fsftKik9FHm4XopWbmKo1ysOkAtPW0yov5K1UMCobC40tqwH
mJQcnPEIlo6KS12kakwd4391RMgQGrkBN1qnR4f21rhI3M52IStNBRzr4KdsibsOCuQDO/+I8mpC
NSZ0qqFXsWQVo7yZwdZ4k/KeoV2BgaNZ0vUNPOjtm3zMevz3NlRj5hOMbfbzO3ovRhSNXbHyYaOc
2pTHlGZGB0Sqic17UtpFKoZyymWoSKHCrb/RyGNs5GmHRFDrYPluJ5982bsF8+uuR8zg6n8REe5I
Dcl4cfH5vq+yC7EDzinHTg1j40i8jdFl9qrHnqzaufj96BF3vinZm2SiqYQJ3p2sUBSWb+6cgiSZ
GmeYp3EHcn5ip2g6StsN9mvX4Snn7yeKOJnAC/BfIHmp4ZV+J0Iep/n6vgk9ld8que/CPNeTTCQx
Anqw8kkIiW2XRKJ8tfJ6wPeqrlpCH2kZzZkzfxhpgR7nPyLE3R5QcOcUjoGf5mNuSUneyFhB4G7d
7SnfXOCFm0WR5vOaAREknrGhwZ6gIDtKwtyUB6wWV7RW2vzLTE4U2dyHiUUj4OYYdwlyBQizoMrs
DwL7kEDOMmqjPCc8AJpnaCDoTh2T2iaEh4wKSMyGbDg1YSMweVKtJcVpRHu84frc8SJBsHdv+gG7
aeB3ca1wGtN9acXo/mHhKvMVt5kZ09LktXDRm8ff54yoNr26MnoGOXK464w8ANzMmuTUGiBxqB59
NS12WcjDh5EnYi3dG890ahnr9zu+of6Fnv2H3xR6+qM9VJb/UiLhLjpa4omicwpcn+gAzMQEWoRI
Di6A1DlXiVAsFkdWzjitBSTz+ueirq3/znSe1QyAjVfPDMhDj9yWMgZgIt8eDMU8iZiAE3fiNk6S
nnrUvvsPyiCFnpJOF8yD0w6zRJK1nn/ZCYudUEnZClncjXtWqg368/DmfxBrAolLW/xa0qYymppb
tHH8dGr8ntjZxs8qq2N3kOL+ScDE2OwkoHSN8R2sYelyRZTIkDCG3OS6nXvGSeK7tEEZpREe9i5C
AGSXtHyNWljO+UcexXzNpDsApdqi8AR8yt9EXHtzHUi8HyejRi1GNPeJ0Cy5u5yti54/wSv1YQC8
E5soWxzdBwk/3WL7R5YK9b1zmjzpkDpC20KFWkRLqWKX/mj88LjUW/EZUqGNM9XTVy10bfYcMlIs
tZ5QjSU79CLqnYYlGFT4veLwaLOYDkpN/SJqd8zBcQPq0DfO3a8XbTeDg5MA+n9nm3ApWtJv877i
rLU8KI0jb4g78SOI0oYu5mHu0XDgIwQtLMLmDC5jmgZ1B9CVaSxouHh5oRWby0MrRtBEWR2Pwc24
BvyyBjiDhRkfaJEaw6itHymO8rnuMERSZi/OGEkBcQF08cVyp4UUPLW6teomX67NJrVTu+PmONp/
P7CyG4f6beqE7guMzdB4ik3LG6lIldDOgjVkmeve+lGMnOXc36pxsT+sNLjcrLF6WzMfv0sD2rii
KxWxaGQIebcNwpOKGHsm4Tmki0P9R48SQaTXwEvnFGPbKce69Ooj9xN6h+rmCRbFKqA1BNTyU4a8
xtmP008FIFh+FNbJW4OvjgIvFnLHm+T/U6XYePPAcd0MrjHw4Jamn/tBT4urriP3JITUyL8Gxh5P
+TvBxrsT8shTI5Apx5SloqzH339E+r1IMxHOISxYBR+MZ+vE2KUDh4mDriroaiCa9CRyYUq6XHuQ
8tX6aMbLYvKJHblmtun/yUggx+6vhcr1kP5GT7iNmY8z6Cu0C4m9KuyNHqtKd3oIzhJbjiJm0dkj
1Pi0TmCZiRwflBKohjAjKiGnePObdoMGpZ55aeXhB9zBhbHSaCVuASpq7z3JaoeHKz3fWiibQqhF
868We8EHKHACiwNw3HP0RMj9jR1pt8cAvGbL2XZDP3VjDhbzjlKm1i0SRpOA81eNNGTGhObuP5wg
wjUmmraib3fwDCninfddgCgSaaqr5m+3fICPZwGHAO+mfCubRZdmO5pU46SLEfPvFJuYvEg/oESy
aW1w1QRoW1y0LrE62KudU5XIdvAFBUs0zH9glmaflDeeMcEtLJSavPyAAK9NzVSww86UWZ3UQ0Pi
0G3qBATwp6E8JiQfWljMO2aPRZVbBmNs2kLeJJuAZM2EWh5nPVECKntq31V3AZaGs+OzqV+OxLWI
sjz6oi5qjcmq2V6viq1mHcf5whcEGLR6JwFen6SC+TNp2iGt7uYWE2c3TLZv0RVhiX9WttImDH4z
7Lu2auE9Lz1t87bHy0ecOuCzCRefxIMdFZjw7Ax9mvPhSGdITll32Ze0bnNab350IotGmNDCU4Lp
sXTpiDd+QGX68yhTNvmwI6yRueXDZfo0cOgzS6e/uIkXEDLPRH+27UoFli3fziO5+7euD1AhVTn4
LbOxtW/ODBM0/Bx1WQ6FSFjXmZrOyqUPkfIdRo9spLxz0Ekz34vrX3XG7eQ0pPGA2AboLS+DpLd7
0ks6pINPvPPBZqt5YltPcWd69W9u3dFqIKZyTK8PvljwvLElHnh4O/LW7LGpPMg4CkP03i8jNNnY
gHuEoHEeqVC67qK1RpUXoK7oeu9yr2Zj5jWY6rPq62YWYhLx/YsZEPCTKAnKTqmJSVwzfF73buBn
d5XFJ0Tlm34eeutqNUUvR7PIhpyQMN+2PKhSmc/0q0+O57WHY627TLDwyYzXHLzDd7hs3Gsx1ipn
jjcMvOIy8stjenyanijnKUVIoqz6Y8WnfNra5WGC6KtYOmjS+V9oPUW3W5MI1BTSCmjAamRKP8JC
F4poJr6P56XadUByR4ktZjD1x/zsstVk0xlFaS+J5XV6RMRREi8Fpmj0468BzIliyzHZ5K1dXLbA
hYhFcZEzScFNLnqbvPbnk1b5hD79rJ0GlwNrs9IFHCR0F61eDpb1/i92m/5mO/JUmhiLK16qUhCf
T2xoO9vpsDyNNthqXGNtWHA9V59/goDbHGcfhSMh+imlJAAx7X8ZgwzS5ah8Ydjs0/XqxDCQznw/
yiOZrnL16HBp3ka6YofW07sN48p8RFI6Z0Sgv7sbdIW5JJC8J9h1Z4hiG7Z2JYAw319b5E0peese
4EDmVIBtq+6Mg8i5qxxBNkN56Qn+Kmmzu/E0AcEbpS0ILZVo87Ll5qR2xlIdDI6fBmtI3MZ83SmX
c/9ucmGnhdqRFZgaKXPX/5xijdPMrISlN0iEG4674ruZsJl8iqRpnCATvdGeM1v4QA0q+yEIwGmR
ACJs5MWVK/9GCCEa5BviHoi503iEXUOL4G8aHseWTI0kcCOAKZvkuAGDWL0lv7KdgVdn0vA1GbN1
4fyOs5rg6qlsD7S2/Slh63Xe5aWvjNPGeAqTDfvLI0K33zy/VR69TgGfbtufqpl2qbreZWUsYiYj
2tPNwgiWtWULzyCUyQJL23E0S6AmDOxDYtSp1wDoSHDBm/C97KxwMjDWmdta5RCOIxypMb9uYeIt
L7qha9yOF7ceEkvCmhB+40GCDR3C5rDiU5c8+jKIH6BGQlCPe+s3QI75RVh3bLrebKvfrZ1bqVO4
Y0M55sxT4FFOBWVjB5YDwqkvKybY0pA7WUALDh4xZpm+RqZn7oQgEV+LTlCm4vUPPpSsrMkFLDiC
zy0M4vA39iDJijnbWf6Nu22lE9C19Tj4eSjuqqyuohgqD4O2Zcn2wD1FPmM0WH+W7GsJiUMFedsO
ufxnMf1jY5GZ1DTFYqfGWHharZlVLw2WFsDx+7QNPSXtqBvcPhIIGImV4GKZd85VANY8AipEIET0
2yLFZeFIEllHIl8Pfa4qGQWa7Dg+E7FIHTOKKang9SXGhQv41tAmGp1DrHZ5rjmlyIAxCSlXFH5w
ImLnyAJeFUFRSwKJRD/iW3qQWbnWNYbzugLuXIRnoi0lC3al7n9Xo9o1RKjLuS3F9jxY/DVOQKPw
FS9XGGmZKD9P0EXPuLELiepWADK/fTVqiDnbO26dclNvez6hxJYSz5ZWJs3psRDrl6ZqmVL8wZDW
gNFe9S/GUGuosyzEKZ2iQXivbsQIERkraKcKMSCgwX1RK3qYFovyyhqEABCUqHFe1EnCkVfJf+0v
ro3lyHnt3Xn28kwld0T/XhcB5hbxKX1LZVrgtZR6YVDhCLjijaaHNro6vjVary8x1tK11iupXUDv
qDg7c584EA/LlngH755PXf7Puswwv8mRUtmiSVnxGb3vH95odb0NO+/1PqzXjgnI/ctt4DIwIpAZ
HKRUBTPiV6+zd6f2iFsVbIXmGb9DKhLqEamMcu1Cm3fTDoN9au1lzFTwJ3O0NV3tsUNdG393vcQO
PIFRvAzYe0OPbRlA4cpbEF9hpNK00iyG3EJrdj7TF6HVduPtxFbVaBS+rHNdm51ZhJp+Uv7qEakE
UO+HLYgHOly+/dUNp4MvlBm2cOofI9ouUfVcoDravU7ODua+sq+6FJZ0rNiS+vtSSGtOZlbR5VT3
rMZKC/6XvG8BTd2dkvQLl03Q3l92rxzfKctpvFhIPpDS1K2ui0BkJw6XWtx9huZ4OhGiG273IM5F
vJaMhcRM8NS+XulTVvjbx2CZ5LxKx+I2gC3Aqpppg71OIJzMlEknosClpC4gGd5XtKdS3ADSom9i
SV8L8h/V7AFx8zVhNwS0Csacx0nB0IQkSEKon434eN3MPwZuyd6D+WQ9Z1pE5QD9PPLaGGv/rRAp
uBnaxR/34kNF77XB7xl7mVJDx1JUR3dQilMutJaVfLL9XidFwJVhGIFDjuVaHnL+IBZY06wqlRls
S3lhD8zc9mKmlDsryNCRPq3inRWuPu9nVI7+byR1fhO0017Sb4T28sqNTye5g+zUxC7f/kD/Lb6l
jTCMQiIlJZ5CA/uKSd+rQK7d/DbiEwjzOzJEa0WPQGVxW4YsCMTY/ZmQti4crs09UwoSUqJypI6A
m85vBW7gsHj095mXxo8QTacE9xb35ZmNDzhnyRubrlDBIib8KpA8wr8Bb9VpV6nqkRTbrMXLlbeE
0eWFTCJKFirn0mGeoON+L2Lg9UWF8yml4Y2SGc4cVKleYUMCR+8ld4A3rNmSQg0BHrGWwinL4Ilt
+cvmtpJ/3VXb6xaDvRcbwYe4xdZoWIJmhPrsxzIBqmM1ZC6Lo7n6x++L5hpEseNbwRcoxnEgZInp
ZoKpM9CTz3uTPZW8vlmI1Y95LsFHWKe3rkBcqmpm8g5XixHEzHDCQsgDgM94VUcSVSsrsfLWzJkY
DhITg4SMJo7JL39kdJVe1Nm+PUKICzmHNWlHRvQO8hNwY0mJ1S+/1O3NZaX9eauFmSTs2wzT52Fj
jHmh34KEGPkobKFgumshSMHQK25u1fSJvVhuda24cy/m30EwcXY5jJVc3+yk5kufOi6nBuirS86G
+aRfgSNx6r9DKsRKV3AcUR7fW3UW5rrGZluYsrjcHbze0gnefMSS/Ealmkm9hUXXwwWgnDR0Gymj
CV+WxwoIaeMkjcpMPIsRiHwGC1cvS2yQ/LXNwX/QuxrPAKmhOhBEsEahkN3kZcfOmCf01I3sOI0R
CG5z0ChdreeiIapQ8wmUVqnLPcYZ1/YHiOVz2PVhwzZJaNR87T/r/2uWxW/zi+E11kHyIpQbfXSZ
akQ3DPo2QkuGV9UWqXegcEhEgdf2BePoeSDyAEU5dAsho9A0wotO0AUAlZ6wQ7AuoBWPPDJfsLdd
vJzugStWUo+mCsVwEguNo+QnNsf4c4tVKUMSLbyeZwMLvxnT+NheberbtIX8none2wB0cJvJ67OE
hxfH1f4HJGlFx8UzARDVa5OGwF5mG+Qmb1CY4pyL2OZFYtOuabn2NOT3XnVRYD1/C5uLKijXJjVq
MR0BDNCqNPc39VRMjiyoUYeDtk43TDNvyuNjg5HZtfYSYKOVixba2zRD3dcx99b+ch7RjT86sohV
yVUZYG2kXlKmx7I4SibkLt7eJrUL87YhPJsyQT8f/h5i1hKLUNfzEGSYnkEw8DivRWCmpSSvTeq6
9M6QbDFxAofPuOknfWsesQdWRdS1Rxbx3jMkkanvRzSU0irCfLSkjcdUsDeMVrf1aUnUapki4E8z
T0/80h80hExXh2wX+FAWiiQDMRb9rCBXHNawkrdlEA7FjKyXjNhpDVxmJEbvskJIeAYkq5uKRbqN
DYM40YH7zVE8eg7C/lH3LOv9MXMUg8sygTJ5OAtS7RmLleMletibZ44gYui2TKxbwbd6IqhLHedX
o+z0zosQ1orekJd37Sf1fXWZqlTBayFSO2J/gP6FhjqebbrD5Uz964Wjb1re8OBeOw36kYL45E02
QkeHzG3lBaUa6y5kffEa5XPfTRfHaF3Czh63xAAKXsvDVtVYnQKUqCKpHVAfUmRc75VARVWrWHaA
I0ohhNGsLAGLdgAmZxpA/8QvphlPi9ugoaT1ZXy2CAn337Fbfw67PWewQ2NckaXunm0LTn0CNQqD
YcEG9Oj8h09nE0l+bxsyKS7IgO2FabENo4/7X5begOxgqg9MRGfGN1KmW7+mrl/dKXKABEVY1puD
mOIg639JwP1WZRggtgONi+b30peRa1oYkZ/1tWYAWyos8qF/qOVst0MLM4b4EYWexm6sdlOfb1Xr
SzFhr7/fB8pMVhz83MRQgSV5KDarNnKXq9LdJ4plAK38YW1noexTldF62kWXNznozIXllhGsNDks
Dl706rEauf11b0/bGv0alqVwh7pX4I/H+GWpIUBOW3BLx5GZiE8zDMA9rKBi1Tx0X918x+mCfsYF
oFtyc4pho/TBmnRTmPSBQeh60TCYcYps2i7FCD9hDwUI/TKkhMUx5Xmi26oXf0vFnpgZ59igP2PY
4+2oZkfzl+Jx0U9h/qoQwZZvsGENRJ0e+xj/rn7T6mbf1a1aroqh/PMCPPQN/MT6+edctjggrmPq
yHJ82LnMs097vT0pZaP4sgtrcGnMf7K0EUiiloiZAm8Pndbamx9z3S8GLzXvAE6YoGpGMsFVyG53
YLF6pAxFLNDLk7aKGTZIoceTOnvr9l4kgP7f8quA9fBR3DXpbZo5VYu7mwTmPiN5aB7Hrr1EY9Db
O0jMZksLE0aJz/CyuySsHd4ji7OeXvSILffllysSlyFhciit53uWG/pkc6YAD82H9tYJbY4Sfc7r
EW2s37Wd13nyZR7APPpeKpFUruhbQmWcNBPZhjdL1sG4TyoB+iP8cNrTcBsvJ6se6MrBcI0i/h8d
6qQpnypIFBPHOf3E92HBQreLVlyQlvBGXcnhFIWlaAWneqmlJwMFqv81k+LmgTborvKVnY/V8t6I
crADgNLV+yeo4l3tg6mtdDtMFCBloB4GAfXilzoczMTjECloq+SKY4/wRGikYQNlX+psjkdMjMa9
e6X2LdlxB0i/xKO8BxEP2NNhnXyrDcVwpu4jwg5DkmG6MJFO53mzGFj1d/hi34gxfSd2izOQN3Rv
FEqickazZ+kb/bQ18tdn6QYTOfs4Vd7XgpEEKy+hNLwb+PqveNONryWu7wbyXTRGd6k/QATMkAeB
Unl5TTJzVWV6aW8LPXEyBnDMAaGAGLoCizzgSkase/X1YYABtrScODmZBJoIeHGMjqId3ZNmmL6t
VoETBXJ53u0HGpNw+R2FZySc
`protect end_protected
