-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uZBe4ayxec5rZ2J4s8UG/YARDdNy6GhUwUGZmkpG7ZhRGzVgMBxqfRzk/0MScBc/27iIeaua44jH
yzZOPmm2zP5wA1kfKlHmwUod/CO1caUFsifUhnN+1tTjXFAc+K6n55HqdUwmoHn98nj1uNAnCa15
dZRcNIiGTs1B0IM438D20gqUcB9kPVynk8evLQapP2FWZVSxJgxQpe0lSbvi0TAmk0Cqu+zefMSm
RaiiQk9we0BBt830qzEkUHhOjXMPHBkJI8n5evX6pOv7uNr9FvaazsidFeVlQx0EB24wq9N1Ejnz
uAbXDKPw4RP2jYiW/dAR6KpqVizBM7Lence3Aw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 8704)
`protect data_block
Wr6FH2d2kgMFihdlESexpN7HZNMmN1Aj8tkxW99qRfe58xO6uQ732qnluT857aTsbN9MDPHAFzw3
rltNLwBu3Q8IdW8vrU6qL7hjqlHMLZ7E0ETcMQ6e429ZqSkqJYTagzOgMN9vv0dkpQ/VMbQcqNyV
DGy8jEzbApcFLOuD7K8BfkAsKJIgcE8jkOHW0scxQBfiVN75noAkz2V+Zh1RevhUO9oeBN/n5Q4Q
SL/PezqyKuLW4Wmm4hZqMGu9YxHWRCFgUJgDl439g7ZbAFInIe47UHDutafFp2XVPrphTpt59+M9
7IKoCYvwclnSiElae0PZk7pyWw9PeFuud1zWP/lTz7IC6Bp6THOixZf069JHucHIEABItPsKWdMp
S60y+Qj16aZy5iJwDt/if2sPxcAJJ+UEyiyxew+ys1UiJOnsQyQmKE2MPBOQZKUNG0zpaZwcSQvC
TwTi7OkBHDZt0COe1UqeMhTK9t/O2vJS1GZp7+JEEn349oMR8O96JdvRoOQxe6+bnePXYJcRLu7N
hPGTjIdmQhvGzap5Il0Y1tH/EFnT8O4BNcc45TcN6fIgr9X+oPAdVj/GnPMhW6Q7egIGH6kskGKF
OGR/sTJyY6EaxbQXdCAVPYktDbeak1Nt1glQGum2t74nSYnhcbVeyX3/c3p4RZx4bRrSAJI7vA+U
3yPahKHACTiTHm4SyjaRXDz/+CnqjkURkkFhUJ+pchTgfN1UrqYXNxNVdqcat6e2Ap3qSGgyD5zM
RF+vryYE3CXBkNBzeNrpgHPJkrpLcCeN6t5O21HX9bbx1EYWAxaKiMcPKM7tnWQ7T0DoPXRZ6ocN
5IW9OBrg/dO033zINMdmHWcZMWJyDFy9pXg02pGUt+tVHtstPUCffk5kn02tjnk5xPId0g0eYcYm
Yzd2araQ+mczWESZlUH482AewAlEv5iLCfjJ+dFx3dQHinLwqDzZaqyDa3m1eL3+mRfg8LSFq7AY
YxhQXFcj6FiJ/z5PXw4drPbCu4AWxlT5qzRoY5iufVxYJi1qnjsOSjjjEiOQkCBRzt8DQRr9IvKt
lqPPZH/kdcOdl5F3NeF2TT66/sRapwKanW4hwWZpeIAERRT6z7nYox8kbGIpia/rJe3zqMepQG3G
usOhbaH4QG2D46j3YWlnxoS9FG6tyUJit+nhTKQ1/UWvuqPPntCdlWGhVaUXFXjIOGwgqaNjxGGB
wkWxxTozafTx9ObkQBL4/TAaNoqVCQl9x3nu9jf5DQjlhhgieC5KgGaL8SXE+mTEuqnCMsFnn9Ip
pogzHfWCY5b0FVtGlNUdWVFYwRcV44cGz1H6hgQ7ZA7DGl4tAHDDM/XaJ5psEvbuTtRJ33PN0SIW
0W0YCkMfTe2F/JyqXzbk/yNzL8ovy56Ig+S3Sr9L3UHrWJSxeDTVtJEkdyRdOrsC7VkRD2ebEx7v
lPEqQAitgfKB3mZGUD32D81JDLJstWSMXCX7exRQJpl+5ek4V8x4ykVG4sKOl5i03JVhbAAmXzqC
hcsHKR4F/toJfd9BDms9JHs6DeIQYyy+JJZwcwJ7qbIjHgXHxt2Y1faHS3VfKivwuGFZckcBtvTL
Hxh5o227XGUdZeKZYqEvzTe0lmg46hb86eDOEUHIQ719QQ6zIajMtZMmYQGcEOPsN2Eh3G/GYCGj
B484HQDoWpx+zUc7BI4lMdFP6AGechKSG461nkxjIiJ5F/zlSHu4na+XMfyv+NdET/esAF94DWwJ
XeAz5BBjFft0Vz76ShUixsdOOKHx+yR3H6tZY4+nSXu6rNTq4CC7MTI7OOS/Ugm4BmEg8OsqTjWN
WYiMKGF0lhRfakVBG8x6neWQs0pjr6anGkGjZ2CU4JEJiuL65bm1kVY4WvhqloONh9CgBD0jX+Eb
TYhSuS+3tWrFXT6su+OYXy8Tm3kbOkJRR2WK/W+3UIcXTJDJycwATPc6a+jgRKqIBBDc6ak9XfU2
RwVSdMoPf4TQ/BL2htVzZ18Lo8YFT/b5PS44zZtn3OYQsGFCC4Z4wXVpFGeGFlFFAexZuuSlC1fB
TusJA9QmDu4KpmL8pmlNMtChxmgujSNsTHezPHuxVn/2iEGiRCKDYYSeyIdogzH2qqU3s0bswI0N
8vhP97ErKIL3I9gsH9xKRfOd51X8S81nc08Ro6yvFNEzgq28BPgR17iu4ROqRPnkhNxdg56MWKqg
5sUdMb1585YqaStvSUR2e1pCTd0RYwiNkYYs0NNmx4IgT+3kAyt9ng/RCEph1BKoMPlY2gUN/isu
1fNJ56nlHkQCuo1gbLNzi52Z3vdI+bC8NeGk25jlup6EJMylQE2/njKjGVHHo8zw+Dm3nWast09f
alZ5Rgu0mcXeHwQ1IK0OnNT06mez8ppRgLkFdx4ioAXLCRHnXXUVz9oNYQrganu4eT+xURFb3LVB
YMXl/mMNxtcPVhDnT6KJkC9Wr4jJrl21jWuhzbWLcV2reAuZixyBnXrwt2u686HYbU8lGpQHnpuU
hD2ouZgVhqL7QfPhLkXwUFAfhT+BGd3fGXOR5yTVzAZKPRVuJttNuh4txRxBxyfeabVQ0Kt5v1ky
7D726V6kJrnsmySzodmTO/P0SvXZIfNnJlvIcTobwln2wu9y0R8WivfJAe+uB3zXfJB9D0yCGAFg
ziEvqQaTYS3vKqWmoXLFFt9xTt/E79VZ4oBcCy/FWKzVE4EIfItoY7kOxDu+weyZruB+fpms7zG3
PK9ffh/+kQ+hJCG8lp+F6evTv1tNgqMHpLIWJ6w0OaQbw4c9Fiw3BTZS/6HYN/PBt72y1bBbvWrv
NNXz9AMuoyNBNDRKL30nN+hP13lbHbF+lgK1Bu3OxC226tyBLOHKng001XWthntaWfLeBRU9lrKG
FG2zqoR4JFmnDy74veZ7dtHS1HWFRLl/D8Y2zGV6qUkUWqpwyY4YOJhLZO7C7QcopxxVFERwSbKj
YVv8dFpw+dit3Ja6mDlgYy69ZYC3xlsD46MK7UOCsyF9+SOstjcl1Lip9qVlHmte4cVCNWcNHobK
pdaJBIpGhOGKZvUv/ysYUmL3gE76eg6Z0daotuJUcdr0NZ4ixMCe5wy3VHjkLG2kre6p8dl0PoSi
Db6srf11vdMa09Olk1jnZnQVss9QUASK3OizXrxXQHebEsymjqXrY2VOLhU++YxIkAEVCkws3eHT
2revAZf07848kg95foTNZRv6GY42zEHdsUD73SJ1AXeub2AxA7/uTEVjzXyLE1yP+0/YFWjYX3r+
fMcAoN1HvkB8fogtgIESaoTMR3d/6MgUJYFsgmHqODnK+oDuazw//z0+rkgOiTVDNxmAB2rDITli
ukeOuMmuRoXhOaqAjZ5VlSXRseT7DeQUtBGDwryKNi03LMh3iYPC0GsHojYBkqDcjMOmD3gtQXOq
0NhpI9E+HtjV61N/XGmgTKPbBzjsi/5H6NMRTVA9wrljtkt8ft6elYjqnqVy9YZjudGBRWgO+AY6
W8Ea51IK4X7UyQsg7RFz3V5FAsbv3C5ca35TCFN5ONpLnLTluX7FqLi+yJmsnRlEDt1G3k84XBDJ
y+HixQvhSgRiC5kOi2krpyqRqsMCWV5lwYAhzcFRHXheJZ5x1Ln0Q7rFGO+VM3hcEezYQ5C7g4YT
2/E44wxCQ6/0DcAAcOOqAxqcJgRsuZbZgpkV2UXTt4wgUMA05lDfbHFuNg7wle6fio6isFpb7CAH
Te+JgjKKkF8hMoDrnyIntcs85FzjrIg+UOEKiTSOxDEosjJSMa8gZldMLJqdkdsJ5MwbnAmXqf7F
CkLt0/dtc9In6FDOjMD/YofQukxhKszw+BPv2XgBmRHdQxXP/MGSfkV8hsxWRc5f5stvecRTOQ9X
qRonGGnLcOpcgCsix+33SUjNduoRDFo+cgb6LdFbFvXq/Kfs3+bMylNDzYQvZBOFTedmdm6lngZg
+8w4ocJKrfMgCX0milOrGJmjsanBb1dupGr6Gk39q9SUihYvo7CH6m6ioHJA+NbcxSHutbEMiZ7p
gbWdC8iPQ6b034qSHiwOZLDDrH0Fi/SDAJFphy/Hitn4aNAQFKY98x4nKcuglIfX/LMfbDhnVmSu
QgKlkY5XLtPD4ZoRQlsO5oXG6Ob6WOA2Qc5nGSoLMchKY+fjk4LTA8FQN2MOZTzMa/kQgF2uqOjd
dF5AeoixtOkEE8Np404yoYrK0gwehSoONJXnmsPbAl8P2QOn/7Yo2APnL5EUscHcR+/qcOkPIwmG
gQhab07jcWrfqOJNImsDsoh5LrQcx1ndI29+FcbokJPPijbZcw7FWRDfZH0f99lqh1q34W5xppD3
Jh38IjATq01h5fRt2EEW+P9PxxAY/e8l+jI2r0HPK3rhqP16UqylLTwYCFCXFOQAUoH8fc6Xu6W1
abmoD69WzFoA1IDXt6tC66PTUkOgrXPQPRy3+m2XD1KzbLQYeDoEmLJg/AQJt2hkHWvgjk5jOj1w
+nKt93rKVPUZcZ/M3uutTtFm3u7avAqKMdc4yQwhzxToqImAKDHyNk1PuOtEUVaD2coEzwvu5Fp6
A7qa2njQlr0kRWj85P1P6FlgquVdR/aQQ4/4Gkuey/dTE8lGxWG6vbh6OPIMu1t1BHjPq4eu0YH/
jN+KWhVTtvPW3W7t4ANV0x7SVt+kYiu3L220RLA1HsfOMqTjGNLbwAj6sBFQdWqscH1kKjNYM5Q+
ULfxPUvRvNoNMewJXpbW+Wca+d4aen3huCh7YWOeuAmKoMvkU2YDwnplsFBymeN2V+lKKcRd24ny
wup6wBcjwkX1D5w2wb0f72Yc5OCV9Obbxcbid6aluuFPUyuqjUsb7dcRjrsh8QHH5fRGG0suvqQf
RseEN53eHw1C/9vD02fVEd7AQC2anoyouf1CP3+WB19t1xYYODs8sAvxmVjzAwC4jqyiusq3UaQo
oJ6wgDpqSZRE6rVF7lCkEt4slPLfpJXGuRzYnLgIt1rjqHdDErYNzfH1+JxpOEDCG5uypU1vYdRu
ezcFgmGjZhx42iSbl6Y5RAQLRQZOa77fQFyP63l5f1FQi53YRJ01A2YJFSN/AUdEKDpL3Qdvcsmw
s0Iyy2/5hCLFP+QBYLf++2cGcSXoPoxXSkJaGAzbtazYV7zT5m/8TJ4bOdAzMtostvIUbZInVQ/D
TJ7RSj4ub6AzQQ+X/XWaJRSqad45m4r0gwzKmIhMpaKrQK5QyAwAPPjlbYm9EnAssOLQts66s0BZ
Swao725iDFNtmDDIwLDTUTdy9sTkUjZUS9IS/HTahX7L7DFD0jzdciqV4f9gFBTS3166p09p6fUv
xBCa+4zICPS4k6SyN3UUsxZJVEhjhkrOZJyzguq7y5Fc88hRBvBm8tF0cJhSL9WWsCSgL8ClbpqW
6vx82RjYVD4E0vTsCZBRNQ3Xz2EPdAuWoo9z/K6ktjtUV8pkKHH1I7mdLEKfBwnD3Ll6sezrjmoL
u1Z0O79b6w4Z4IFaicSI86Eu1lvCVqDfePTVyPRUcU7szp/tz7BcAQh6kt0zLfKrdlk7qNd6kkOT
bMNd/dGRU7vZIUGmqz/tPuCXTvmltUcQbt5HoFrSy0xETDND10cBVbSl+CnF7Uz5NbFrfeWPG+UF
1kWl5hn0TNzZ20swAMK0UFtwggVIJfVepO7Pr9Ou62nH7OornbzvKR+mpzZVp9cjRqdtxkvey1E5
FWlz9nIIi1azf8ugFu5VvnpkEeeMqrE9DrNXb+Fu1F/vYi60LOy/7bZ6NpAbRTcc3x7NMzghZwu1
PrrbgkaynFGVGEcMNQkYezRdexdcWzj2W9zHlT2QcgY4QhhYT5EEpoEuuKbEO7rVSGK70UWi7oSG
+0wPvBd5NiQwhXYNKlz84c1w2gRI/zSDVsxk9/h+Po/426U7pm+RGsSgEEIk+iGOC7yV5frH1N61
1SFD4/KYE62pEqohntrbaTkJcBdCU/kRwsRAJn/7fdTuIXL8N/SvS+1ncGKrHYiepnCk7svtkbeU
mKYnK9Tn1+nWuXtWeivGeYiNSWwcl7b+kT/aPPzs9adVKGEM4+FSZooncjoPoSnm9QOx2VYCdAus
IHzIba49rWzIInRfvebDF1y12SI9usDhTkHzLV/kh1TWWCNuipX/WRc34GPVoWMz5Wpq57SVZp9W
E0BEaTZBDdvTiGAfl25diIJtIA9NILS4MmKCUgUEsE9Nh7D+9FxMwchwt2asuzjWkYBqRs9nJg4g
MSJ4t/ImbXjAYFCIGW82/EzmHOz4/6uAGJhrq3XX72gSfUfLHj5+VbJi2ZAWG19ywz4q/CBwqcT4
bCZh7u+0R36WlsRePv3FCdL2ds0RAwDS9pTMxaHQQjnsF6DYQTfrFbcZ7RvzCndbC1FM4sKCzo4V
UzkCrNsfornSCbLtAlTKLkVKvzJODf64frhNRHIpwCT9KL+UWTn6LjZJNIXvn4ON7bsEfgG7nnaP
4dBaWTiS4ocqwyuAq0LPPxa36mR/1nNzkW06ooIi7kSvhDhvT55W0t8mK91t/iwGsqgKxBhT9gla
hPnaEJDFzqLgihZgiz76PRCpixB6CJ74snxncWMT0J+60JRoeQgZSUYWXuUByH916KH+d/1OoFmL
g0LCjh/ycVA0PRe+G2Lg6IseFdU/CaIxWKqAz7h+Cf4KslZPlrIphDLFpHl5sg6MptDiuXYj78ur
jhzTwoSwasK+a3A44GMquFGMIfRk3ZPcRph3VAMIIOGGVdpnC38FAnuAFkbHJR7TSjh46rADbzAB
2DsK5siufoGyFqPSYVIbDcU/qW7kbcCZc9UZQcp3zn9lwnM5wmQKX7wJs3IC59GDZZK+fBZ1Hq1d
FbBhnrC63tWWRQeG+IotlV4y+oEdu+YCRu4Gi271u09Mp92ysMHu+1hXHilCBf4RS9jR9Bp0vDjQ
1Pde/YR3d2BekIeP1MfJLVqP5ELO8XS6445jWq+p2ABkCBHAJ02X5/0fJ3CcG90z9IeBXfv4H6GR
dVWaIXmmoSjrH+JLTjBWxtE1mGuT2c3F8vtFAewefocR1cA+R5Xft4gzxpavpldF9Ct/0bR/iCDz
L1VFh5MQF0OFDPvDDJk4NrGvQ1nkpUW1aOKZ1cWDzK1l7rLdbK9irvXZNKzQuVXE2WSQ/M6WkTGz
OJasuczhwOLfGtzxIwCwTJv54mtkDavf9HWFazLUjqrdNVrpzl4PCTlcai3IjsyZUSDdoFBjYVDq
E4AcrN1gUceEycZioRt72Z4wROSSg+QBrgsWpu8bcJqQ/VS8+9RNN31iYGRDLqWD1tdPAgrXJ9dX
DL9cdO+/xq99/UeEPvtpy5uC4IA9MUuhqUd/4ShE3cSwSzPbhICfMTWsx59ZC0Qi3AoNWlTco+VL
nlp55jnq+fKh7wQNaRLvGebILgqDPpTbJ9Ox/XGpen0df2v2fCxY6B88p6b9LrB2p7w0lnsl/BXD
DzOeQ3tt9t99bH3N/3QfjicFEuiGyQNINr51mARJB2pk1hN/hZ0jpYsG2qzaHWUFlSnU0W4nmn6D
kvjZT2oCBfKrnDWdCjVhgpxw5fnaZy+LzM26QkbNzb5CaULw6CO9MtB4vCCna4eLs0/pAyiFlRLM
rAT7BeEyt+6wfx/bNku6HMxdvSSjMAMnRZnrSBSA50gr73z00RpZLz5OTwmGB8rWQXagOjc9B61j
M4aRmT8WYW5sYMugzqg2DqxAnasEvvLQwoXJbymZL8BqXVHVjOS11nfTYyf9KSCWvCYEbNyiguGZ
nlk/yEHt6buyFCZlMhHizvQbKPafHNAXPEPeH+nU36xrxIsdf7107l8zUTIQspG97ch/ccDxzXy1
USnRr/ZI98vzNbxhFHtgz/ZDj5BxE415mWxryura+DfU9cRI07LLCWAfdeCiva43WwstcWmlqJMK
gyePQSLqVY8VWQW/Sf/BvTUttftrluge44NJu0pLw/JBpPy5JL6ePwr3UWBGVuI8UJhSjzVAHN6L
xph98aCs+9uD0Q5b/wHrqVieAP66OHWWkXQE4yBT7XV/47k54l6ewruXbdvl9SskA1Y0ueZ6zq2K
RDRgflh4VSSyteQApx97YDSQEQCJFIpdvYP9DLtgpTCTooQV+9XTHqqzzs+csRUy05U/n/lKggtn
XNNiWC6hp/JezAFiiNOgaN5JqT7Zv5wv3HtzSGVynIbMxeiEHWQmHPiFb4UkymkbSvfFhpBJ4ifv
2n88bz0VH+8ylSZlXz2AfIfnruS5GGc+lg0sxGYrieKyIjdrhOxsGx6gsfLi5hRAWnJesPv7Pk9s
3JyVMwJLRIieML1dcNKxwT6U/XdnPmGzhJoU5mxTjbIl8zuLqWnNPHvj/5bnhPUAEi6dQRl9leIU
hF2wPOCWc4I9a4udJKrlqMQDx9Yhc2blt8Txhtm3Ll1BF8qyEO7r35S/XkjkMXvgSnWdMH6WHiX4
pYeS4bR8foaL3jB0OTeOCHOtup5YJQO4AfA7ShR2utbsFl+bTDIXyEIZikKVHs+PfPCiAZVwV+3c
mIV2n3NGcM/w+6nw9qkcd5YLo7nekYuUa9CWR5a58D7HlYlccHlZUTni2HFc033eLkUDzM6X+dMC
SKMRGiUwZ35rHmnh7KGkYit49Ius/ucl/chLfsRE864PpYeyu+qxhF+6CULm1peQSLUgOkkn003T
nOmGD0+oBGkSxazIn1fslc+G5ABGMpcV80DvnzRaCA497Uaqkn5C5Qc9XiyFoN1Wm9u7lVCWaBZp
QYlpEwPbNLIrm4hERRVR7PEN/IZtAEqXhDJSdEQKalyOv1GL0T43qo1FRZJ8SgWdz8QeMdrAFanB
I1MQnyRkLo8NKtBUQvlorfavNfl5iTgBnAbOOdv1VN6NLUvd2W2tCqd7y3zWoZygvEiunogioueM
/RgVEptb0So3N7I3AT8vnjxEqWvkXh4VE2QfMPuq9MkfHNOpME5pXfIbSsEbMvMtTHyrZHZl0LnG
fK6mJvMvFkKzvsFg/3tSC235lhdOD9CCFmVEzYBM7NaKllIF+35UiJQAcUjhYRuREFXiYW9wQeJz
ITZFdF/gCIP+Rz99QqoYZcTyGxZL6ft5TLzTmBa3Z8fKE3b6vAvRFWirB4DbGtnhR8J7BEFktc88
kVQAg3KLykpPnHBGmVoLX571OZCdbELvXZ9nRk9pgefmVLnll8IRnF7eSBRDFRZ4eqwDeyBAP7+e
BS97CLNE/u8H1GRpf6iNrOqBsF9KNEqISEtV6b1spTExFBSbhNtHiuYaxyIojQKJy1pgyXCX+Svn
USOamM3fl7azc/c2U05U/Ei0L2i95nfcTgNbqKv9eocSi6/bi3PF76xnImIoXO6FzujVMuv7ie94
3vQewAt2XL44zuTpY+Vtc6xJPFgkRLvedd8sP9JFXh1ja7g5YAJiNq/FQ8S3lR+CkBQ6/xyP4GFQ
tpPh+eL14lr+kDuENmtP/FvrLgBoMfRZyIkr60a2r9qiOriqTXTdXBORgak5CpuDtlZMDDrDQe5x
1GaVBNPegiU1s/YC9qTJ1OIhlzqALGQrlVRiSmBgb4SDop/jFIoP+c3iON+xTvaKopeMuBNSCW5Y
j/mziK0CyeK4Rhwydn3KgjF7pg1Ls8iW+YIyvwCgYb2UUmG/e2PFOBLkJMMva+gYktE9EQrovFNS
JRk++TZ6/0aynwOt0GmYXMUh32+Kpq2gc4k4wbVYPEPD9wWP6V80HM4Mqi0My/ZcwPzO+L1G0nTz
vtR12FmqVcFudfsQ+qZAk/XVoP5hm35Mfd0iOq4NIdXVTrUBWoxBiaSCL4e1Wympyihhrpae9gNZ
UesaCmXby+3qw7FQbmmKiHCltz/TE7ynIkf1HTSLTJyvItEuuwR+CTxY30XxJyOEd+54q9pcEZr1
xKvdF7LKCxGsuZyEBaO0UAl8Y42KOQgp4isddET02PZKqdXtuJvw8bmDtfSTi/J9DlhojRjvXGhV
UQi/rb5SYSFAJlgo7TqxLZLMuDeXh1WlPe0Als0uTW5AWtEipppxD8FYV8N+61Kiz90cG2tyM8p0
LoD4XxmVli50HP4nstQ4waib5aJVufOAAbVP21tI9tlB5bfCZrlMxDD9zGNccTMPWf273EPsu77f
uX4luNrdYhddQft2svbCAW5iWGXaoyEcxOKhj9u7Nz3tzsLNAiNmPE9YRt2uPzVi2sImI/pPfWUF
V8S1/pkvwSbCfsiBHvgKUtwWdIPDeBPI3xK2UbiULFbehb6fPx1sAFe/M07FI1vH+1gYt+DXI8Uj
85JtMR/4Q2OB/IReT4xP3K2nkurWiljjSGSVwne0cwgz9LYolVXDc4zoibT6F4TbrmWJUOE+lXN4
me3o9NvAlMZfCMsl6Tq//CgfWbwcTglNGTQ3wSt/PjxIACggvFjqmKD848X30napDBmPfDm7r/I5
xdWziiqZAFJqR2BnxFuOXRDWHgjo8YUompGitK6ezq+v6SJugG87ytV+U48d0m1RNuc+ip5wHIuV
2MYfRy6X8uJuzKKvDoE0y+ngkTfcemY2HmJF4eIpOQGASqpCsCWhGHFzztoIxVOPCw746YEWZdr9
vs0fa4TP4ZKYS8TxnNK3NBR66c5EdBzavL4AcDE7dE7iR1Ot/cVllaif9/fK9n196RsJelzKeE0n
1FJcyggN4QN5jnzifd7oYddaTj+jCu44UWJ2sSFuVyE/K9PnYspsSv5XUaZtgKekvVwIf2WHdndM
nue/Mci+zB5BY70i9/nbOrDiQWE8xK5N5gFtYiD6r++dJGX/5vxGdR6phmSS2pZP3Esr5GihD1yN
tQj4kK5Ty5SgPYErq0+lal3dNczwSm7Ak6s0BNaCZ8q4sgXDZ1HEY2psq5JRylHGjpnb+D530crg
pirDoBz7oRzKNzd0ivbpKxKpfFXT9SzgdXfTOozs2xyuv7+IY+NscXOUn+jpcY4nIELYktnSfZAs
mg3gyCB0prLKU0cl50xacREWN6N7EvM+OdGy8hRJRN66wZLOYDFteGu1/cwSbHSLtBVQZ66IsEgz
3nO+r8FEc8ZWPQUI5NXdAA1ol4E8ccinptORZtZJ7Ox8boKrbWB4HAG4zw2PDo6rlkMI6DCft3BM
YPAViaikyHU8ZShpuQnC4tYzXfRqyUQQlJ3n+/4TG3NpaZ4IISZkz6XtF5XUj70A5Q/RAVhtKYCS
Tdz+xuK53x7SEFKCkFSOjHJHXzc2nh2At3jYMq+aCft9BP9669Vp+8RUDwyDrc+XUskdhl5AWjC+
coB8xZOODkXGkkbsTfyWxFgmAIYwWXM1b/+l/PNX6W9darkZLCYDoMIWeGLX/F6gCbeIBUem6TEY
7VzzGzlkpT+R5lVg3lgOzmr4uiuhZ56IRfDZHFFx6vtnjjh8BYHoGfi1YQXQPYnVh634IpaA5UQx
2fm6Q59+62VXdJmhRnS2M7fGbkiYR2OmsYyHWXYEggGYrwZk7mbIYPjqBDEx947SVzqfN2TQLnEo
NYkl7shRlyIUd9iuZwV4xyG3ORadXGrp0QiWFaLntjHePNXQ3+fD10g4AzkBa9mHKBI3Utzk3A+i
GI+I5MJEv7H7ojd7rF32UbdR5dW02AFRygg5U6kbkxOtgkO0/pPHXg==
`protect end_protected
