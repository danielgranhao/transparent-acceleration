-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
qGnNc6tNwR5wYjQbwjmfkoIZSswkxvIMJJfIIZ+an111GRuiCemDKgZo3/YRQ4tJPuOETxYGINek
CPS9oMtfYBDPbe7xGIuTFRD0VZXYkzY5mqXnFry4PHfDGa9I2xZRQe6CZSLDkPhTTSdkn+hVMT3Z
HPbNOHs/LHo1ouTMKEc6Tg9IV/chhY/f5ZQRMwl1PqiZFr5L7BTkyT8SEKaBHHv/Flfi9cTIzmU2
OkcaRO4EklZnLi9/Mmsjlu6doD2KS6bgRIK+WmJizHtXl8XmG8G0NmNCTQKnH3gutzmSfX16z1pn
egWv7BR/KEsYuPIkuMI+3eBLgkzZgWLSn8GX7w==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5072)
`protect data_block
Izo/3ZUgPmjOPdXOZB935MgJ0VEbyEPLQmVoZhUJqUniT7N6deeRr94SVYK20GSH/oywRqqRDDwS
zlmZQrrxUjWmswBCeEnzlQ4DU4e0M4lQVgA/KFvoFHJJnojU4b9UPDHkutcGA0EM7HQofMYpIlGo
O2JEZbrbh3eAaARQEzpj3RVW1p5EqJ26KsV8vUqetbhbQLRUVv3zsHxeW8z64hOj8Djy/SnOSrtC
gaaGHYBJADzcGA1xDn9dKSMIMgXB/nK2Bv/4UOxJIqkHAcmlOvoWIxyucZ4jr6mEXrgtV/IS1wnJ
05u2JPVNbFWG4CrhO1bGVJGf8FXTQoOlGKikZbRemk7AueDQb8DWFyQqx786RxyU1qhd8z/QhBSb
EzzB9fY/LS4VR35Zz5bLOt/kkCFaYTX4TPR88EJFjJCuP5Zwq6e8FDXlGout9xf6MIB1Q0aN/wGM
a8WS+mdu6IET5xrcVjFjoTyzAo2u0uN6hUGatZ26s68LN8HS8M+81q8xYOq3qFKzzGfYLDL3uV2m
ZtroNJ89dWcWYg0HlOHsy/WLsquubqAmS8COHLHJvqgkiT+LWNmcmzRsNhbJ5IZTEhqCie2jtAnN
3EMpRImxiss+Av4jLjtlTbTCapCQST8iMCoqIrpZuMj30jXnwTHBJio8L6JRkJRg0xNLXIg+Fepq
yv4lh5d2069+X8+gC3LiphkehgDc4N7QeN0dwigmJJk2d9Qi5DjgrsO3mlFQklwnbnj5sPtDw7FJ
4OGZFgv0Txx6o7LqEgpqz2H0Wid1QLxeej2dPggASQK6KRY7OQSvOM0FBLOSF1QV0YuW42R40tej
ycFcGO5mCTeebeQV6aoHBViDxmW6dQrg6/iaKSQoi4lXtA8gULQ5AjfXsqZRqk3SDFqiOo/fcq+t
+T5ezRl9Dd3CLPM+9ivTq0XihDsqO7cSQLMYUipNQLK/k5/lImXUDOd6kSReCQKS0wrFwoev3C7r
NKPjPXgHRvb1n/UUDpDBaeYSlIdoxiSDNafL/Lzg2YkLyIHHXHUOEEmy9m3Qpg3out033eZXmWql
lqv2lkBEobbvdVKGLdU6RvHR/JCfXK+nJRL0a7kG7Ec/7UuwvFNzrHzC4aiurPV9T+mrRlStLZSX
yqeGETk+mljiq7+RNjByGfbAfeR6x/eLKZToh8CUOtU4v+4Ahl253qY82cm4BJvcg91ARL4wUFlZ
qEChlHJx1iy4b+2O4sardKtAkp4JAiVyz78lr2hN4nTVbD6oiB8k2lW/RG2PVznvNBGNJdK1kopi
w4MZtss5VU2Kr6ZpZlGNKaAGauPS7fFHCDFMUh7KVeMPK0tiauGDlxgE7Hfrm/FQTk9rLRYaO/S/
dPwy4QYcDRDJJ6Wkm0M/GRwZerzbW+KfeejMVlouM9xuCjCt8+USSs56IX6pYshl99mtyiM2DRlE
RJPVBDGpCd/CphrS9kkb1+z4rQc1e3ixqPllgFqBg+UX8Pe1jH6Z3zldSB7xdi2WNqqx1mmne+NB
vynEd/Vqd1g+EjL+R6whSojDOenXlV4PEECE6NRVa7SAHY8rvJFzRvjTlHv8WZizklnRVxt/vAqj
E5lDJpcyA2DcmBTAiCR4K2D/Gd1Jei02/o2gQiJWn24oKFVksrX0EJ4BZzUpH0DkEV+n0o2MuYAO
/8XI8zeSOze9yXvT7lYyc3LsMQuKAmyZbezIQIktkeyk4WYuqVUlW6CHhocYCPvpTGa2rtf7m2wO
Yp5oElYUXgwH4N7P4Lhzy6XuxdTecqMkG88SRzyE+B3dQycabJAWFa56OZQm9yeyxCI5FiMTNmmM
6GJvOsJZo2/s11VJvW436KZtG5qXh9ZO11ANygtrQDx0TEnSLSgkNdKgPGtRKoQVsLNv5FJuLm0E
AelD1tRJrMMQydoAL73sBLVk19ozgNTklvdJ1q+RpOBnZxQoNhXZ2G2thMO2xqQ2AMUIVZrj0sN7
0XvrW42J4vhVhSedvQea1vAj5rWW3i4f8kjHH+xIc0OFOlu1hu9JNC5zLn48pLPJyPDZvmdhNpEQ
KNwmRKj2Hm1nJWYgg8rRKZummwnLrVPqi6dDmsil5HXjavkMDaYwHig+dpgk22SssgEMLiVURfRE
CY4fbEq8qIWSCHPpqaxN0/U1ACaoJZE7PMlpV4c+6Ty2CzjBKLeAy9oGGTk13a+CeP2S/F3eiLsE
j5saQC/gvqIGJJ/F+4bN+fyKpQsTC9a/DmsybxpOSPNZZ/kCUb41xbAY0xjw4GTLjlgKVaKlFEcS
26pIL6IVxIzWKw0ZQapavNAYyVGbHrsyVBzvXLWwJYQz0mKopbz00Ed3GYaHcUXNM7hHbXEQQZRw
bXpSVkGg1MqvCMLaXv9cHCLalf6yvBxzqXSiivSMmdRi/dsnKNOvMqMTv/OwrQSCT4et6jGvNxVM
XqtjFz1ux1bTQPSILf32+nrWIVMVtZQG2RP7UzERcZinS2V8389uYReMl1jbJnpUIg1BVR7vI6YV
p7JNim9thIr/FWwcGD5QB6EQao98nF/MXrylb3Snjfoo7zsvupGbVVT7S4LI6NKlPx/6SE9d1E32
JRa4q2Chey5L9BFeoQPg+suXI3GBDFIcpkEGBsEsyu9FGnPmpKqiYtPHNNWzMnWoTkc8VMupjayO
nt7t5y8FzgwPa8OEKQG304hA3xYsDegbx+SVKAhhosHQCDmbFL7jkV+WwK7qpGFxTVja8q/04QQK
srI2Q7RHGxbCVQlrQifZta6u7mQ9e36kC/G7P+k0yWg7lO7Tb1Ebt3LaJYS0GB0nDw4CiAByztjK
Yo+ikfJd1LQVIN5Z+EDNklB4Q9AAKyM3dm/DjEqWNNlArKFmrvpMUgIaBxOQU1x0sBpHLKYf0bK6
XNbUkhwK1nSeRpSOi89ayEYYOBtNg/ZdbH8kmLAt64e0atLoHi2m1LmKXXGvbikbK3JQDrrzbQEK
TCaHRTlNTkOf80CCEOU2zVQXCJHk2S5LIXYOFL+jSDRSWm0qX7Jxhm8sJnHu6JrFDmdf6hfxqGHH
wsTgscn8t42CIIJhmI859G4rvqQVsVAiZfPcreGiY9b5bGYM9C50UTRVz0TTr4qQRUzIfSkOwUV0
VrES8E4rnb7f7k3yuV4Ezqcc1SuI8sSY6Ef0ev70/HPCfz3rgtiYk1dh0o6+QNu7YUdqYJkYexGA
0Pf33Tysy0ednFZnG5mhKbR+lV57iiD8dBbrgdZJW/2sjchKOldYKbvE2VFJDlMRidZYAOWte3y+
48wFGbAV5QkpepvrBJz6jReG5v8LUoxdsJQ/pPgEPCt4MaLIGcIT3l3Ad0EFJHrMUWvOood+Rflx
VLNbIU9LRoiSWtN1ra34+5nx0QIS5nYamla/xzS36hqCTEa+71rv35LiDniR9Ujtm01VE75LO0p9
giDZbN6v+IdhiGlcZlAakxr58o2M5OdN4YL84XTV8hs6A97YajzpnekbfXjYnLSBIEngwAR9YQuz
8MV/jcaXEIr0kLIg60NhKfs5khCFoeb0qPCmvi9x1EXY4ZXpHrKgbxZHP3ExP0n4vFTI8pdt6dmE
CB+ohPeIsLOZCJsOrM+yr/3M/5HF/niVcUkg9swROMDptUh/Dk75SsASM2HS8EDBJgcxoQVhmuyr
0hjpSaydyyPAD1qf+4l2bYY96kwbjM331H3ZrEjwhgwrrWutEQ0waZQZfKfI9PXzduLpTvSVtrw0
rNyJovCGwmJq4XsIJhtJ8v3YO+oqSr/p5UnVTIqgz/e1z61Wzr/iztXrsp49VyKyC08QnAXCq6QA
kh7hZQL+F9kG01nU1+70aZO2lBHv6AJTtUBbNkyq8H+KxXJYP296qE80U5pwNke0FppVJ5EUc+5B
5x3n2ztclcAo7iy09dpgY1HGn/VC9yUjsv+IO55x2uNrBBq5iyeJuREYdQDzKhhzSwAWwF0TTvn5
18vkpijOuhwXgTXJCZGMGejNvsBm/kd1LYZoq09qpN3yGc6IHRwXNQd8PJM8CuYFNB6MkU09OYBS
7J1uZgJG/oP55osfSq6nxA2T+qy1I2M3ZNZXzhRCWcncsfPrOcDf/2PiAPMTwk7IPYFpelWmEocC
RRmhYAHcPSYYE97VCg1/1T94rSQofih2JzgYhKSdaUXpcqm9+XfAyDHV3FLrO1JZXCNlBExBFhF0
RE1khfCWN/hFv8RhRNMo1SLdB4ZrXhdjPEOvQbvAN88h0EbSu8di0EEVkbbLxtLRHCfaC0R6h7/R
eOQHCztadsxeWTadpENw/Cdvgg/Eqr7f9IxBvk5BCSzLneXHQD3EvALQK7LSUEIB5WMHB7ulo0H1
YYh4zEM5y3E644j/3nrIR4cU3lXaRI9hgaiM1FeUwGL14rPKceswdinkCGdY16ISLKbP4IvQB0hn
KJgvxM9WyqlKw7CU8gp4wNPgjdk0mN/nOe5UK4TnKURbPpW8PnvOL8KWfVC7a0L9XlEGUUJ9dLkH
z4DdVMqm0udZkjvuQ1We6TNnGPMTojTkU5zfWb1iVXRG7EI62vzLcClLnQwNnWYc8ipFuW1/6Q6p
RIbAMZzI0BJFMWPtQOJd4NZZJqn4X6u4G32jLKusdER1k369DLEAjrpsG9Fh3AlxAwG4dRdppGrn
7eooqLhzd7xNKeGpXyC6xKjENky9hD8uzMcSEIu3eCThe9deexYWuMJlylAOO/oK1X1BnJ0+1AUv
JJN8QFjRGLwKsc5Kkm/oYweuf1q+v8udCXEMYxZ3g3MBxyOCe0AfsYvEnA+RILPDGYKSmWX5GcNo
qirtYScpwPXjiPjrVfPODxX2mh5J8mE5CA7BrstXqvuabC5gCI6BbAgYhAxZ97TUGvLhvY/WIEvN
WfPO7N+xnbG7NWuVMEIizxB8/Zc6jFBOgt6+XdDBLp6BnJWXQy3H5Gbt/7wWrhdvHrxOYS/WQQ9j
34dVHA0UMlFvTURfmVvJbksHvGoF7TDNpxh0QCCUeY/24UnVPgzwO9XofIcK+WqkNj2z/UDaUiBN
iy8Jw89rFxBsbm2rEvmyAH6JziJExb7fSnUNP3odBYj1oZqkkAfO5LOJEUzD2rix2vSG+EmkOoik
awbEhpkKAGuVURMN2FWsKEPyXsX0iwNXQMMiILWC8NYN2AnSbUSMkTSQsCXCIH9/DQu9XZjDNm8j
kvNAlyG4X0PqktmdhKRVcIyH0HhLNDKAr2rrxrIZVnLQMNNTmjkj7Vh9rJCrRxP/EnVbm3ioyq66
FsqA9efJ470BkC7AV6PH/jap38rAHlpCKjMllm4p487K05XxjEdZ6z/b+1rGOcewzy25r+kGSYSo
091Ka2K1xG3IMKHmx94NFsnhyMOpSuCXKqTeqc78kLQcgs2AU8tyTrIc8fEfQNHHxN+24fIAY9jg
8eOj+0ykW353VE1zcNVZD0XeHdDkWYt9GOfKs9oMcV76Wgtrn29f2vdjrwT9d0q0XAJSKa985qfq
HIyLK9S1wW6aLaajvCHqoxxBXDcFmDqG0iP8mXjDkFMQ5qXQn2c5xg2IRxU4l+ZPcwGuF9zem3Aw
Ndc0Cn/LD7kmYvrfgTdZnLAeqPDKehqbos1nDRhkUYKoeVVfAFW40wiBv9mTBGhhzVDQqRsyE9TU
KONhzjRWUUayZzClIbE1C6tpjAaU/KMz3kG240/oeX7nP7YZjYZRSWcA0pskBby1BfWKIUo/2FOY
ZUGYFZB8tltvKw/csHICJPhjhcDupqDb8hQTjZh9DBldjwcq8R+Qq/e6u104fqxH90FpQbPw59cG
LauCODKKkAsZnPAaYTuF0ruK/BJymGejHn0xoAKSNkunwtmVIb+vEeO+XO0de5ch5yzys6n4WTIq
ocT3Pmh3U1vJ+cdsZwko4roXiArNsUUoS7VvincyVMKldxqPyg0jcLdP95Dfelx93H15F2iP6LPI
dqU+/YvYpUTSj5B+9MD7ZhRBV6flRMzSVxrcxnbRGFfCxPNNo3y5M0KhzqmGXJM67TF98K8nFIUm
sb7k/LGH9u7r3RVkVwTyI7zOlnsPgqpfgmGstQhNcP6LWew6h/Hyl6J2dGt+ErqZM7Pc7iz0/35k
dE46uTvcAknOu0I52WITfIOvYlNvd8bghaEmPmCDNnQE/RkehuX8/4UU0I73Z+kWM8R2gpLm119z
Z74TOmBBWNrtVzhinfDMEvoyiDXray+jRUeBrvEnshk1i5xDxsAvQDbOW/mHC7lCyLMnT9YLVjwJ
69e3NwBGbLH6raW/a/xvbKWCzfWCl++IrMvCZpO0W6O6TeqZEsBhPKAs833gGrbJF7OKOh1z+1Az
KjBsR9ckplWrFx3hWbVMP1jyu7BX4tw2Q/Mf8Wsll0VGcbLdIRPryFRwZ2iRbaZwm5W6HBeSl/AF
xgl01N3SJ9b/+h9FESCqm6e+1jjm2RbmRMA3tVT6xJdPuIPogh+X20b+ZHjdKCKNP5KOnEH1OXqx
/xJpFqVkxWJ+tPPQwPrAxWup3kjVYEKNy5zSf0VCwlVFikYstdqqxiWtnLR7GtegqaG4xFtxlg1R
FzaxfLRtu4dqKhTrnERBF64Q8mkoSnvx3oLg9/CTuxVNKtgi0YgAKlgQTq61m/Z3T52UZ3Sdg0yu
UO+geU7XPaimpZMw3I3nm3QTatd9ND4OtfsMRXSZSFrF6kYmgyB0FcbBhYrt0HYN39a1Y1MyLAiG
zKKOXNGHyXuzPz3Pp528vt0lHRx+k5/tQo3ptqp+ja8FP1fKr9I5vKR+K+/G8nt/RsMItJsxeVQ=
`protect end_protected
