-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sn3tLu7YqPICrsu2iPJxG6hpMK4Ty48RW5dKRPDjIp0OBuqj9OLSdAlQTh4gealz
8zjag5LmscrD2Byp1ahilIrM/3LRsTKAxA7yjNWrquGqGjNPXeZuN9T+qlbWtCDU
vTMKsR4nAG4QBjAINwmFlUr2d7KbGmH/jPSDV1ltp2Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9872)
`protect data_block
mm246vJQkGUma//apdGhytI4D4Ulo16C8k+Mhkdw7HBbDpiLCYANchPN2XrByllk
Ddfn80MXEKU2Dm9pkxPfLJA/nDLHREVEd5qwXSQEGtZBQnyZL9Ix5hHAkJTFg/lv
pHYu9oNh1lV9Nf6Qf80sxtkF0BuyOgnZ/O38P14+46eHnA8XduRFP7JzAEDT3BTz
NtXmeVkDKp5Arj0UGMnNkW9dS4UxVKRR8NjlK377CjHmIgAMjQJh87nxjMEhDlFM
kAjRvqqZUuSP5bVxlhIcmTQ0FMNOKPyXpkrnO/2/VqMEGpR425TqYokLh7r9dbE/
nC+8F4KCUr9FWeFwTRO1KEISGhvDukpwJm0JvuIEeHLrsLRt5+NckTgFsoYP0Vd8
uhZ6mJrzxON5iLWjpUg+wuY39njc6vURpe6FGqn51TStU0ZP5MtRoEmPZilE3Pb2
Nx+159FMtUGGbqP/FoWpAG+GYz4jsjD8QsYCN5EUHoHyDctOgKW/BQT10FfrlhVp
stEvmmYz/v9Pdbe+K7u9h8U1+BRVZ8KP38f/bx1LLETnpSd8M5vSssF7L9EdZgpC
FdU3grVjxvYwxfykN2uwp25xah46RoAc2AX1gApz/5NX9PUJntaN0RnRrisGOJOJ
4cxWhCODtqLmwHh+YDNYuhckpND8WWopi9KiC2wseEnCdStzIA1dMXBzNGGNZZeC
pJASRFGx98pFCl47jkhnp2Pu+yrc6t9kD2SKlj6phVzLvwHZXvo9Gd+C2zu/Gppm
f6LdlPba+kj37aS8gz5ly2V8tTgKiE16rpJJg8/UCj0HwECC1zK/nV3U+8HfLvKi
QmCbcBpbjpN3MecNU9zc6sFtdYf9AOa3x4pldx5ALmoEMGki0o58Kh/XgBBCcADM
SDqcNQ1l1BRaZSv4FXDK0L58/LYzBerZSBo8RaQrG2OOTbbXfnDGIAeS0vu0jTPN
pqzTEbFZuILXVCF4qUDCoph6aSz8zOrzT1yl/p2TMj8mqIM0FaZl2e7k79rmF4p2
15bVevhWBl5dmN2qI7Pfej6T5Jrl1pAzrnaBiYjH+ivr7C6L/lXZgw5Q40rADoYS
v6tGZeq4WSLjz55H+X6Vq7ozLt4gVblxBKNjS7HWKEr8KXbxA/tnHAWXfknHfvMR
e7Uv4YK8dF73/ko1wv9qaFvoAggM2kPbV4Ux1++rWWDRdgJEBWU6FpckJmxy4nNa
wZLywmYMarDDUw2nlnX+NWea4WPs9QXR8x17EbDpRzQ78TLJFik3EOO1+QDIwCFl
akGnDEZE0dLL+0aT5Bcsy2OkvOa1Lg4t5cZf005qm9E2AYPbjsqU7gGP+ff/TUWC
/2F55TbWwSL7zHBp/jaNZeWdH8idQ5MobU9zGJGLDP2B2P7agBejBsph+dQKar2z
gPQXY6iLZ98Il7THFw96iYXjzzAmDYczzfI6t5ms/4Vz+I1nQyDLJqsuk7QGuoWr
ffy5n7FVvRlIYVAFCm+iJ/txCwGbo5mz3Rekbe04jOnsySEhEqSUcwMLQuA9lSgI
imvpw1gm6v/dxhbIHvGe7du+pVFxRtNjn98tDI1Y6QRli/6eR7OHfbjmTbKkYzFL
QAC5+YrSiF7MnKaLBIImNTgGmeC2LnK7jsebebY86wHW2kVdq/Lg8uKm3XapTQfH
+nQ1BMiVa0Uxl9W9+q0vZYSeET8GEb/dgTvxmTC8cpcJ9F6yJcCa3d9IsFklmoKR
jbxjnMmXaD2op2qFz90OUnxnrSnrC6iuhjOgylnDgfwj8F+G8Ty11UfFEzGNh/Ow
ASzJeVDquEr8VIM9+OL94+h67epTEvTwoipdTLqV7SAvb+YSRIBy3tWxq3IAi4Fn
pC/6DjHU8wxqZYs2UVkDaTtSAWuwRh6rj0W+U8zRmqRIiqKOJpf/mAvYrj2O8doM
ldnK3td5oqM6SWhQrCV2AzcSQo+v/d/iJYRxpPfRA2BPDmYEsRl8mEzWgt8OtSyJ
ptN41tB6sejqv2kXD/Y2cfdqnWkTkpWn7guNGuHhmVKrN94NeSqH4utBvI1bF7nG
Sw+8k/5dJIKSLFinp3ik3sRvqZdwZOK33z65j5Xrpz6cbPcw+TRpG+gBAxbnJPFi
n13i11eti/82qj2Nm17RMzrwnTwVbVNor064OISS4RTeYFrnXo+C/iYvv5ib49Ks
GceXhOi8wuKuoRbsKC9mBOEWkU4fBRiQlEh0WElMjggJpxhUcAIu4Scjv3SkbdAD
mrgTCT25Ztn5Jl1cuGsi8NAp6XkZkNNCCUObl8TD42irNegNVrJsDlmwrx3LRXn8
8aNUr9fnB/DT9piYd9GJNqKgQlsNWr+iNGm9pQ3VtLPgj8Jkb+2t61zQCW0TMFj5
eKs+Tg5PF+ybw3aZksvuWnmjdtrl5NUDjryZwfW4haO+qyVwQt+uEAEUwoo1gvNQ
Oca4oC0eVGneHw+gYNjiB5eJQ+lQ8DWJ9QnWvbuTAwVedas/mSgYPtMoMiin1l42
yxwfQsEA6rDp03iwpkymfFFIv6xo0+cnsw/CmajYBPBRa9QAhBelEnGqv6k2Lljn
L18V9BZZ5ZSyu7AfszLJ+qk2mVBdUdAxkwK1+/+1nNnzPuDxLYwhA/99taRYsUOi
T45Is+DRlNDp8WRRFUVOEmnw3nYvkSrFGf/kpT7rZ/9z5D3ggFp9Ilfv/9OhtYL9
eVr2BAvEIXXhK1zlwmrHJ1OGHaYpFdsW3YZLNUxwc/Dz4L3H8K5tXsZODZaDx0BD
T4cH3NY1ZoKES62IpFTVXSbCKkvIUXhDJPa5Nu9yfqhiZwl9uDU/SwOtUrZwwXZc
GJjfXhzBZjqPzRejT6veolsjpXLnSk8eVGTcDVLASkyVEn0aSCd45Rf8nYPDq6Ub
vFNdS1J/d1S0R+n6era9tVIGvBy+VvNZkbw8mH1a4ciCOZLN51pJgUYym60UiZBO
8Wbu59qkThBkwndUYvtqslY12FEcYL6lbO0REAZ7x5RYXyp4amFJZrL2GNFkdabH
+NaFLHGITsNANpRyEkiO/HtLdab7/aLuhCcthlHF+3dOzZCm55lzOv4HNJbdb3+9
XZZQViC2jpiXsZxdbIJFxBBuBOcTTwPG/merweUl9+ZMG6t+domMdWF9nN0tlnvO
2LmtdGUFidOkgc0meeKiCWcEd6MR+IUs1Z1I/wVo//wN8kDIbICYSA8sNAJWYv7B
ALj7MtB9u6UaSiRn8VdilMX8KFcHO5Yy4z3x8clT7iitsvjyEoYtcXrYVCWC9Q81
2yb84mEiKsD5EJ+XrbJFLqRwexY8cJ420a7NrrjaQcz6nkzAY+6y+afixwiNy6Ka
K3/5obgx7qBrN0iqn2KhyPADIT6zyKmjJQDJ5u4Eu5o3mm7mWEII1t9FVtFZ0AgI
GsGNwpdgFJiWV5LhFhpgVvmVIuaRiQ4Uwt4swhZa+hDPpk2XDe0xr5eZiormCtnB
LNJNgO8yb2l1CBsZU6mpSHxi1wL37LVg455MA/zWDwI7Cjj7HSdo+j6yesohFLvl
Ynn8uovtPD89S18HocI4ls6Z09o7Qui0uSwVo6pIvWlLBaMzhU/KBLcYiqnAul1u
nHuaiJR/s0qzc6gJuNxRX+AldSO9EA9rGEoXm5LqTdcINRwdcu7gAZeJpSz3GHZ+
Sbc897dbQGd6aNIhv362xy6QH/yFlgHVlPt3qZ3a9GiYPt3OdfVsTCqOjgWjaBSZ
zFOe07qDAwaDC3BwJWEoaxrhM2LfVVqHp87kilbEBLyI2DxB+E0n2hK/tcG8amfh
PbaQ31XIu+4BkIMdHc5xOdbVcpasKmotwObktcyFUk0AGyw3fn+xfpTZ6gdKI9if
HNDaOsOOeHcm4PcHjBICVCgIbo/GoH/PNXC28gny/jLkruYK1pO1cQk1erBMQkrU
TYCglEpSmiT1jcGhjaV3568T1N4eHd/yKOQU7rgHgtIutjXudPWfSbFjW/Z1EI/R
RfIDhoLjdIUa2PR01Dv4V6EZSe0U0EfKMR+rhBgZSXhEDkjuq0By73u84wuGPdLc
L26L0GH7Q4PxaxUJrkDRQtPivhQs2uy1tjDnU0SYb/Q6NuNOy8nyYU8EqpTokRvC
jtlVRS6qCCcuPwN+QZzmUijA/9193VeyXAeMfsfM4VmhTmaCFW7oENNiqVxMrjCm
hLnP5i4y198Rq3pkTB5aHeCn4+SHC5/Hy2ABlHO8WF4tT+1XGqni3hOPs225pfJ1
5SRuO7lgqVemullc1mczuuoZkL/vTNOIMGVaSDGq2+CUXAfYoHaAa2MU6uzyLSg9
90ogoQ6mEd28XFCM8FYNyPUY4P4mEjm/Kaksvpq+TWFfL80g8BIb86+Efy9d3KkX
UqRyBpUZSlolIfSAMQu/UmqmRiMl6iqjv4I6S2rWt7o5ENDDBG1WRXsVhyISkdMb
ekHfJZUkeGdmT3K34jYFvzVdZWXHscp6yEDfXxmqMAryLGDlCQKryTROxjW7HNRS
l+afswJSEAC5jUUV/B94J7Ddd347p38WwBes73wawGeuDxnbJUzjSp+NLZq+xPLi
RmMuGU6C5oCLJFD0PacvVfAPahX0j7IGsuzjCzy8vFj4UEqRRK+bazAuzgaUgVbB
ytUXhvhdOM43suyarzO5yNh5RVrcm0Nd8vYEvizJwPIp7BOEIB5OsIpZfb4dnKgE
vfIG3NCqw67BQp/2zIo+cmmi+xmbvFdDNfGcxsCcRmp4daU4FoBcHGCPflOfbEwR
i2jEnLRzyqJAIZ77ZqUyexRGNxZUc6Iu0fxxFT0ShhBiTIc0RCSALCIvvgVsnpuv
TnVvX8fNMcrSyI7MsjYKfzzH8UcvfKMKlTbDJum/ueLy02lO7XfS5H/LC7x5CvZb
MWz+2qN8d7oNc5aJUvCsEB8oLKiBF3KRI9t+p9haSu79N2oElzFhhWIJtADtZ5bK
Z5YU3yhB1NhK2z4S7O2b4nSe94iDg7tEBXRO0qbElzlLDyGBQPi92iqft+Epy5dG
jegIW3Rd5pdIsXhKIktzMC2qHnJLYkWPd7PXoQ0hvsdZLNAU3ynN8GTqKKa4KHU9
Zw+CaCofaMH/E1K10TxpIt8aybfjVrB2xp8FcnUETa2KNVZfem5zbx12J+PI3Eon
QLLrOzT80woxSUWJNTjoPlihsVOyemti0NzBBHPjdb3d+K5RIr9X9P+F2R6HRNp9
4YVxf2uuFmTE193pbhz6Q07lzVlCBjNHo9D3ocbBd9VZq6QO5iv8k5R/5bz8Ynp+
mgo9KRjR+b6dFxdempx6rXkCZFjFiOy2jTtJOM/03i3lI4hdxwS9E5gjMiujss+V
dTtAoPjw7nvcLP2H0zb5OyKfQ5shZpUDilj/NaePPSe5vSrRDrEA7kj3HkhpDZl1
dRThftYl8AR9lBW35lDXfPl1Lu5EHlPKj15V6LXs/7difZHUUsTdK+RUwgfYMMQu
58ceJbDh8BLFk/f6hGMOiTFH4gtLUoZHwOv+hPBOkcm162bJuQgjoYVRk9gH6PeG
mfKxBnIdNBF0omcpXqRndpYidhrGcclJ8/kYNXjof3z4wznesTQ5pPqb+k5u5etO
eCJhv0gXNZ10hZmYpghkQCKfUe7ZHyMr6HCPD6wQ+VANILD/fyE9DjWVEp5muqLu
kR8Dy4gBTzgXf9Bx9Ue1rnyMMZQWOB2IbQpbY73rFDLmTXvqdAxVrwbG7FiKJ/Lh
UU7hoBUIuVUT5h7YzWLuUlPZvW49kciOAudUzqdwL/igbb691mfQ419fH8un4YyR
VpS/ht/ytbwRR7RO8cPdj+5ZOIiFg9wS0OOnUMXmD66FmI6qi2yiYtdUiClNYSE0
O6hjJrnLmH4jnTSPTkEh5F6dECtOS7AKdcjh/lq9jyX+OxA+1OxURkN+uDEtp7jt
91dZHZcpP0zR8mY508jysfjJPQhtNXY8kCQ25lnHYJnqRl2RxsEruZYSkJKdVotn
da+OZbdfer5p39n/I6IFXYysJKPyt6+2AXNtWyaNnYUpQZbFSfCeca5U+Ls3s8t6
MOEQCMmjaE+X3kS/zcr5Qlb/BetJMEw9A/ZBZtECZzmufBMbeumnaayMZyR/fPiK
FioxKJY4ECgdyZeLs10EgJI4cFH4BdFis+V4sHcDYZEnFhsPaKWKlCWl+U/gryob
/4AjMAoiX5/DP/kfL04+vgZM7bB7sU1QX3f4fD/Wd/LBGbPh81g1kWerDVIQGqdD
6na7nRJV64+gVSbQj/T2D8uG/O1GYGXJ0wLv0J+vm4eAYyYeEbwtpZY/oPpT8mvb
9Eql2ASlL27RQVua3rJ5a57aE/KjB5/AAgoJw3TjIf9AEWaEiiLSUDfyuh4BxPl3
xruz4lzDE8Z7XFpo0Vo7ZKOq+4p9DZVLPgDRD5jKwVYI6rCUuxWoyYREl5cZWm+A
watvu0cQ0ys81DjHY/6v9lX9qNRs0PVg/3/Av0HI4cypBA9ITCjHl3S5qIqtwhI/
s6KCQjsf9R40zpPZbfSy+U71atB+ELz+hlFmrylado4uDA+ftYpFB3a6tFENm4tn
xc02QB9d+mDL1KPygb5y2SXf/SqS3YpX8achJlJCd1wTWMMWROkkuYaRaU2zn22F
5ZUGhku49gYd2JthyQCjlC8oW9eQlrgnHQpX44pqPXA/1Y5Tn7zO3FyiEDq0FwFM
pxjUJ4apB39nMd1Dzp1JatRXawAPq6gL7XRVEw1guAPSmDpHk+I+XOV9Ynen0I3z
NdHNe5d0kVBN/R05yBoRYwm8M+eKOYeaWvf2uVwiJSCGlqoglKPsmnFOKmEh3RCL
6iAm+eW5ecUskM6fC0YlKW3Sb4YDRem+89At8JGcokhmWlHzvGXem1Vm7tUDGSjU
QwmdD8JY8b+V0qKA/hL8vLtybu+TI61PKrSKGACIMBJE3Pt7nTZt8qZ9tOSUC3OV
N5jckKCz9ezmwh+OjE2isQlGlpkxZbpDhwmG9h8uUDaQcRhqBzH5P715oEtWn7Z6
3KgMugXZhW95xAzYkw2HsR4l55bH74aKwkj0Igov0eD0usDXXtRGWdx94INGz32b
vRnlxP2MLPMrDluzBGs4gxEMBOrJ6nEb9ti4EdsTmISK7V9t2PEYRHnoqy9x3yR+
EUFQkX46HTi/7tZ7e8mNExiI7QqV3HCw8rfEwrvhtXy+fCyx0e2ZKvytFNN4Yflj
P6RKrhXVR6ICLj1Bz994Rx+4MQZ8gATypRU3LhqL7OuPwmyxVCC8q+rpnqCDrQ/A
iSJ39A7Eu9hdACqQym5h33cwL96PQAoGuALR3d1VaXW3FOl2GegLJnUIpR/AHoVR
Jq78ZjzXvPZvbWQLlokkYNlbQxoFAGLzk71cBy5OB7C/ijMLfdCVlu2I4GIpnpBz
K6+iFIXUEwflp4OnuoMYdZ3hKNVhv+PFC5zc2dmnag6530ncmDAWRAusvp8c7VFR
Rj45O4qhj6vEJvbr2fb2tQuSd3/fX6XglNvHYUDf4PpUvKYqgTWkrXw47iDtcCC5
W/2Wmky8o3JbKVToXM3wx6W/gqgfTfxbxIzX6CQ+RFG2IoP+sm6P5OXERYYngcJA
6bYp3E/zY8LWiOOA4L7hGU9pLahdBkqPi+o2Gt5jDr7gZEsizb+p8m8GunhdJvlY
HpwYc0Pp63vsEoFKAQbljtKInPUlh2ypdZorOwUUugt/AU52rQ3/Kpk5Xfz1PRo3
VQU5R5mzzxQ4+Jt77GoRgxGUhqR7iQLnwmaRD1JcTIgEcpirbpnVLzZbEhTJ4ail
Hkww4oxIYnx9jXiRwG7ZXv+EulgErejHeyFZWpUhy1fhCfamvZeuj1HxR0olhe84
EqCgJAZz9Q9WBfGmU3um4XnMbFWms4XpfQ9e71CigMWYNO8eZ9w03Xhkwmb0vfHT
cw49kc5K38I0/5VgOgA4xzuRE3Dd4x3EtvGw7hEu7YvCdOu58TgblmRdPEim0acr
GDx6LZLJ/ZY36cnZd9XNNfHTKf6txsQwGbqYb9FSxm1So+9jRB2L3VzQy99486Xj
00cGLkEtmObQsTq6TmfGwVuktWkmQk3V1HXR/0s4DZJ6ROH1re+QHZ0G3PHHlJt5
Kkkty+JOs1nVGv/3s0L0fL7VVyn4vhqSBKCcPnBQ3WSqXZq3+IeaWdb+eM88tqm4
JGYkK3qgaYroDJYAmtZU4DPfph04gENch1lz7hdKEzN86qTF+t1TvmsdYkXnbfJl
U1FqArJY9w7b8nu1UPBrFmhGHVOl2EqZal7GeO9qDU6UWFcy5+/nMlWcKr+hwQxt
ociiUOyLz7xPskpiZXlIx/I2AAkI/p8AhUqS6a+H/uZGH9aIhfqIU7eM1aiaPNQW
4uVJt/zAREqUOQPopymhbPFr5OrBKAyPrGwTLNfYpLIJwrVtqFZqsaq5Xws9faLo
GwCpDnJHNGTEXwDo7UubZkctnqPrl/+1oO452wWc0JgARBhys55q3j3eH47/OJ2n
XIo+bqYQ1DVQj8pGor7Be063IYNgVL9yoEaVyVMTUqZun32JBlFYfUQ2pmTc1+Gd
A6OvIY7rAulHP9N5mZL3JmtW68n2K7H+12Wg+WmYY7JWe1XYGd2D3VYYpL3V2axA
scrcEFbwDRdde+FuDYkAW/1TFK4pTyY/yXWOcM5TgZ6rZ3bOWwIVAoHKkQiQrY9A
6cf93vHwrcFpT5AhnSr9CD8rLs75ngAiUWacswjiZGcGw5qAf/KnP6GN1w1Jb+BA
nu9qmMMQBIIE8d+rdFPm5xkGZat4Pan1l/ofIhxQNaFyZstcdS9n+fzOYWQLfmga
H70DFqBdjRDJWKsqP8rKeAcnrn6sejFiDW8lcs9tN8ApzTs4/IhgslCSVPocQZ8Z
1m0057G4eRhp8bP/qzbSvwl+DXehsqVnprQYpvEyC+h6FKudHLLRhG6zCpueEj99
EUHTV4+VXZFJj4YVf9feD9Jg2CTgEQAp9crZTkIqguUKW7ucZiDp6dbQRvPnVAYR
fDUlO2lnzBnPjaOpAy4sZYAxo6DGZ6QbqLL9KsR0ir4PPOFQlnJjmHwFSQavToqu
GeJiu4cw1QvTDO3BmqiFvT4u2c3LXwivpV+Bth/zEdbIqgb6+1ypJFcUjdxw9653
/zx+GaqfXNu9yHcjT9Ya+yUGiyTE7ADHdJpzlgoWG0dx9XJztuzYyhyTBDmNr1u/
uORV+LLPc0DQcGOzvdD5OQZv4Z3BX2XvQYkavLhWtiWBu2w8TJZfiWZ/GJ+G5WMd
U1VafUBrtZnGFFsAZuthRno4wT7o/C9FEv9bQGML+zAVBO5zS/JMoGGeFXBJWZEV
oLXszgBLM5Dg/nUI3V0y9+2Cu29CFGXr/kXTR2Xbo5+h1reJ1B9uSojkxzBdQQQm
fb2tYoAxER7Di5CR1jg2P+IE3lv0PbMeVncwkheor0gvvANpIoQY5dFdQi/VkGkn
A5dEAIU+wWT+KUBTVqkNDu4uN/1N91VRuJAze952QUcXWRYHfh/q9m3odjzr1xTO
1CZ4lGV8cZOfsAgYvWzYAGCLQJOflxTh61YyYeNalWBN/atgvqKxrIDpT7QVuMb7
0ZmueZShiG828KWfUTiCCykXHnF3zuhjwtkRDAie4lTlrg1J8SDkgayG7A4U6acy
hoGwFavAML0FPp+qen1VUVsgr1i1iOu/woFCnBicGLOzsCGpfPLeCy1ZPiTxlaId
89Uwy6M96uadIUPRm57hfmhMTpt6bWz/jNeBg8tN5+lXpFPnkG/2QAjB/3+Sh8UR
Tyvpbf3gdRdRoAYddDkO/+z6Uvk5jtYZMVI5hlgVE7NM9xfzCgL/2HgBpspfxLU+
y5/UzYEAds0LhNdNoyQSlU3Vgup+hYKj4jX5CSjlr9eCEziPPF3+xcWQofaTQjBF
LoojyZloIqBEh1gBoSo4/HqgpLNxgox/eS9zkKlCD4ltcJ2+hbiTIHvo4IcPop14
doAfS90Yd2KdqZj5IUxC6R7Jb+JFfRFaAuNgnB4vT4pUx9BKfJfFlGqDh8YzvAfS
V/Dr9s8Z7K4gbrgWsDrGV/TsnraKim2R6YOlvmlHbkZvA3R5Lyh+T1WoyQ94qQ5y
MhbIcrCOO6PJNFHlswvHOHCDT4iSSPwUfhK9X302uRwJmc1UEgORqjtj41RcsI8A
ofFsOirYJzmE0fxuaGK6xqNccx9niusB1KdA0Ecp9P4utGd2tDtRb70zQLuE15w5
W/3rssl071fAvh6y7wdmI2hAGaha1etdjok8ru/0nWyuoBXIMVyewKTIDCvOndnw
EJNdzNjwYr2tTGNNXYqxyc2kjs7VTrphRMoP/JT0FrfBHAgDUAAAQVrnKdo02/mX
HNvOlhQRxBuL9DMS/FP2ey8GVo1wBeYTOxjKOMw9QCpyQR9JbrCMWEjzfAPJwdet
rvf91oC+h5AzPxFV0zztGgwf9TfKDTN4OR3B8mIod3Jf5ZQnprBMkNbchMT5B8kb
nEbLVaUAAIAqcL2NH4MNeWLr+elZ31/Z05pZe3vw4YPWLi/2ad8x825WjN452U/P
h6kBCYI4woYke0rGQPeVOgOIjHs/GXBj1lT5FFgdqTeHpf+RM4iU9wK2NdLoJQ5f
yvCuPMxHxAJD52HarN+2FflHFMEbt2AoejpZ+/3JXq7gdvxoroYqVx2E1tb7JeCP
mYPzPNm9Av7gFA/g9PbuDFTJsVUDg3EfilitxzVDiphVzuhVeznW2ksceEV/JDVe
ZsiOt43NJyLpmC1sNT2AREmqi1PlkgPbP/+T23f0kze7cGcsz5XZ9jPWTyXVsa6U
j4kCflI7FzbabRxWiD5qcrDfS0OzYFB4pnxmNVYQbGg5Qs7fEavfRBn1WNV44PZL
n3+ydq+nL54DdWdRkBtQz5kvQf6mYgHfm35mNNq8V9meZB6YGC6THM+K1EeatlfS
qx43ECQ8VRMhxjoWXQ93wjzwYyDA2ED3L80knvFspvR4SrelVv5SdrLJFz0Y2Rj8
kECqp6h8F/k9nv8h1ubMj3f0OP2euaYCHh8itvpdMaRK6zw+KIJ1kkezn6h4fd0k
9KHOfYzTS2DF3y0dgMcCUUv7TpFHnbrq4mC3oO63R98sjXnB3nYrCvlUNOie5MM8
S3P23j0Iuxy+SGalZh9G26rOiE6YBJsYciSCu7mLVjMimvICVP5KytWyB10J65Wt
PHVCw3czNxlh+hL4zXjfRuJGDqIBX6gTYiFtVLXA3Frwk1yQBWhI0tLqax5qL3iT
AccOeQmM9A1uK3ehIpBhHvhFIyrWUAtiOrgdIpfmGF7MKeUSZN0noYGQ9L2DYoq6
auk04qgy3TTgOMTs0QevNcUp1+BkYpbowD9NsmGayTWk5mn2jWm6BVmAxAO5RmvT
h0yn52XqOCuBVfkpdYo3/E/mzH39eKesYvx5H+v6Dz3I1gbISauGqMmL1ARs/kLt
HtlkWblu120ns8c2OkgtLD0yTvmrOT+x1AuboJc0FuJWLdKs7boF4bFMR/N/oElZ
qgKfD2Uu9dG7XNahrvZ7Vj0BMzNrE05zthqFq1P3KwZJMwJmtZx/56Fhhmta7V9W
KtOO5pcA5cW1MUZ67AMI4dcmn2bU80lD4N+0wsZwrC3o9NLW4GOksNP4UNxCB55S
mPcu1IV/3IHJxbH02JJd6ahMWs39KRiRrax9KecIQTq1ioUikQJY9jejl0Txii91
iXMonGKavlsKEdvhOmxGRty2udu3NvOt4rFIg3LXCROnHLphyOCLzNRz+rCNpjI4
M7s6KzZalHCOO4DHD/RwxzORTlurs5FiE8Pno/Bwmpe3KwZ8CWWVjdbeU7GWpXGN
KgwBKozztM6NAl69zel9nrq2S+/ulRgbHUs+WGfrL47gL2n37r1KB/J6cKlJUDRv
DL4trrCSyW7kORWBt66f3gEl6RvOKtdT9GE4PjDyPAvTT8BsFldrRq9ousoifjqL
Xw2/YqwiR87iNp4GDYd7qeP1K+9tF6d+8OSyCFvtHkYneuMWsUaJBI4zVnSUHZfP
VK2zntBhPnmvJb5SXoQzqSkjA8a0nZtqj9GWceYNAl0zfCyB+HXGe1BWSkMWo+LX
ciA6s8SM1EPuCXn4yEahQZ7JdhP9cYa7yjghXbONjQ9u5XfF/AVfb0PZQ3od/Z3w
0s+PKvQryILHPCPw1swpmcTUNKw6zPxl3vkAJ5ZxE0UJc0qT0r3yWFV+QMOuY6AJ
tl+eyg8bA2Vl0P6JMp1hpgUtW9l7NEgJLdTztx9FeicLw2HFj1ZOWsZeyBvzqAXA
ie9bYuahjD0XK4x17v9T73POoiuNypAYAprkC0+tpaPbS8r/yn+mvkHh8uNKX/Q8
bpFVj1TNzEcFXdhZXw2WB8vqPMIrhGQ0kAGuPspnzt2EBnY4v/QRQaAZpQ/FfbEm
nEbEcxoRlf3Vf79T3AsnHQ2VMZzMNYBk1MSxl/GfcN899jB5ceYPGehnDifDxJgk
GLQbDq7pQIM0PERS0Gbxvr9lzp3yL8ELQho9ka/Q/aHi/9lN4pUzCofwBSUZppe7
wb/+O9bkJTVa+xk7ROvH1PcQmaoHJScHbzjBxq3u38v+dOFnl+0VuOnFoag6Yw11
217hliF0faxs3Z5jzaVTIL2srxeywn3F1CQL/3tdHCIFFQA9JvBh6JABR6vq4nZP
9PMISbnUEI1UG08wF9yIFQWB9buPwCdgseFO05ajGh+rIayvZ40EhYqNER+5H3gg
shbPi0ebmnf+BGWMDDV7nVG5Of7sevqz4rTFkDB754t1UV9EffeijfoOJUGDM7hr
tZYHZtZrSDghWXnoujEs326X3edqPxXc3jivqCqURggct90yUIj6I4kLmHahm3Yu
Z76884GPacgxZifMWgxTK9lLfbRmKz9nMXdTRHmZVapFskPf1sFoJKTkwdpWRx8z
CfLOYTiE/ymncKz0qpezjFvVXtrM4bLFhNLh+a/rEvPG44F+JGYa7qDX5a7i1gMl
DMSLq3fZs1agd0mBLd5oLrnOxtgCYMFdgo0o5zH+2AZ3IoTZh6sws0qu+CTKAM2y
bBWQKbhC+uSvJdAlwYZVVN4eBjz5o34Bj2Z6AvZSvrh6O7Vl4rvwTfFra8GpisIy
7TGk4iPiaQI9DYws+EtMj7UQflzWtZTWFMr1q5Wmm3W3kwO4/Y9hpLLUy2jxaECn
YtZnczznP41kM2BvbSbxyFrobOCcj++bEHum3CZdkZg=
`protect end_protected
