-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Qe+kqH1t6ZdP+qdIr32kRxIOL99mP+ok/HOqWTQ1dpKTnxFvmHUodOk2AQWCBuFNHlPvbko+Sixp
NKA+KQB8VvFC25REVLTHTI82GmYDbtZwrEDyLFNItX/3vlvjxyovs6qgbO2F7XNY/qlj+5/vvxxM
qtNlDz4Ynd0MBKnWd7bYoDZQW1T+nPs0NClIwl9ieSJqymtPUOt4C/4KZkqxi4MlxGz27+GglrKa
uuKpohKp6WpM7CTNxbYdx76mdT7joNNXpJl/hFVXcqMheiYD4PoTl5drFWEVRmSRRZOT2OVcsxur
ml+2UhOZqajtHNBZhPbZszLmrApz85XPUOGSbg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6432)
`protect data_block
ZfK27fj0bBmKY1xaYhQbRthlApeoIm30pmSK9Cv0chzYcs2/GJ+2dsdL6EKzH9CWe6ICnOY7xD9D
UpSIYKUMH+2BLj2wMbmRRHg8uFY60qgM0EXiXe5wXvjVYnjFOohYIKm2LHgbbS7AAr+zGLpkLZLt
ORySWwG7cwHpOTLXZH5YwdKYJDxu+A2T8o/JdCLDK0gn4JZ0nxnljBp0y8rWDOc+RLK+QeruSbTR
+RtKGN91JBFhN4VtiBsm2yipqlb5YOInUePFCOAI9ZbmqN+pKj66erMFzIZapbNT6zk97uiQMmF9
UsVpCaFX0CnPNIAd+Qs7WgaZhCiGbx1SeQlTwlEoT8h0ev2uR6R9jafgQo27uQYEOepAji48I6Jf
zIVkBrdn0lbRZyJZzy/VZ9X4dJE17eK+7sGWzcYIDiC1bl+PB+cVM6+9sZ7vGXo6dJfjyE59rnix
AJzQvsmPv8qfrKT4Bopfh0hz7Thr5FSNrdDmJ/hjEkcadL8Pdo3UfdBmfgVKDSeHcKqkfiIWP3NE
XkGkP0bINmyYj973oX5Ak2vxPqxMRSOyZQyJ3YeW67QKnxpMBR5BTm35XXuXrOUbz9PtwfvaR3S2
rMfKt7UaWGj9KM1IRF1cfeyBwXhnekQo9gQiRvneIlF4/8cRfO6/torP4wMp6J6/yFdcRek0WwLf
glpkYq4ax4/wXlqfWhpyTGl64qhZT03I0cq78mZarzPhASBdiclVP2fSXtq+6qHSINwKBfMR+CM2
CZoby/SZDiA43ZrQcRLZ27iyy44iJDGrBnFjMAOlCFHcB9o14qOZKCrbB0XcIE7rjAyq2lOf6Pk+
EoB0+tAJ01xbo4R1Fd9meUBFrzPCgXGV7+SzkdapxGrnJYkqd0AoCbdgO+B6xpoa1Rx3k+90iHJV
4GGk+WWVmXlE7dtF/SBY+k+FG4hwWC5yYf+rVQzZ1tabWV3ZNcw8nUL2LqkEyRf8NfBgKD81vaZN
+iZq2mhV3YIF4oe14kgammThZzqi/o0bQehho4V47FHNJTK+928za6llT7yKZ17GzrlltRXOzZob
9eIsyTAA7MfzG/dk9XoQdHfxxg5khL0uMwVl73VsP7rdyCTEB7mwZ0JMuxwYZiHxdnWSEy+q+XVi
G5A0Wf6aR1qcV/Uh7/y5JPQ8C4YxIc8oSLb4jmwGuI7sJ5664NojxhD0cwdeHTKZJBKbJuZeB01R
sXqU8/wtpy9vsFdY/07OAZJsUYoaPhEoc3tr9apHaGX6wM36prnORkXMXMk/IQRvqVwJebZGh+53
owkowqCeJR1lYuQvtzcTcCL1Vsw6+A+qBXjLBBrxWDHOvnahVIPRTf9GptpjOM531ELPNF88uk34
wINm1p19aweW8dtoAL4LlXYzW1leRiV9QVPflKCO+HgMAoUgxVCWaui03TH9k89bgRHglXGJiRYx
aLy9Rr0Lf0jv2ehO9Wxa3dttqD6yQifJpwxH0ZcDEvSMyuZnkXt5IeOyQy7FR78omAOKSNPKl+Yj
IO0xWcZmBCGgbezS5P+LLmwmQfCsgqh5Q0oldI7fAC4yhW7HOxOInWo088KCPfQ1BfRyHg/2Ti7s
qqdrlmxz8EWrR0n4ZP8N7TD6IgSF32XOLjYd8cv6OFB8IfKjarb5F/x9Ac07UKc2+Rzo+Y1uJlQo
TWJWDDKFDHSwMh/6Vcma6zZmdRzckKS0/q5W/4XEh5pmNcAFxcVMvVINLNn5slzylqvsOVBiiOX7
22O8E5mJmVA3aGY3qw+fpfKlN3xvDFPnnUw+ZFy9pOG8lYywoJssWNX2BltcWfF3Wy4mTzhQ6/lB
rDfGd6KsnqW8mW/dF8ovGoo/FmbiPa9UkXGFiIUdQLFtWFAyDN5yU5vQG6REpPICOKQpl2c8ffI6
aWvWqnDQIBiLz5wg7JnwZKrY3dPIcJnUWz4RcysaFyxZEoBFwgHSxgz+yCPDcE4V1lfaoDYfkELq
sBetZirdHmNnNdG1FxIqOW7zGjfiqPR+TaZwoh6mUhxAT+v7MEo1/Eg4EPxud/KHMDh9+FxeSGep
QTElZnl67oPmHENGsqbOeOAY7V8bTS6rDOrN7r63HIykgnwT9XbZPMlh1K6BeuJC8vz6MkMCSbd+
xLr1ELlKYOnaq/iMWtpAb9KpEgXH0A1PHqNEunLjfXA8ok4iV39zK1s8jZ1KgqRvlTNQxj5VuPND
lduC07xEbiF+Hd2jZ0W3vGK3ZzswDME0SHv8yWMzQ6iZCsNfwJNeDAdrWIF/HeRBCTmCLwxQz2tX
g0XSXbTlwhcdJ8FQJgiWeBkg5yeFUj9yiSlgAngqTZirkeapq7T26A7ROtOcvOJKXuBTDbGTmVQb
k0lLXdrL6V2k9MShwD7U1et9FqhYRNaNUN89N+Nz2E3ui9x8LZ60l2fbhEMMtjI9BEthHE2JRdYp
JSq2w3XkfpNeeZJ0vOXndd/a8w3ZgO7otrC/56tiJTa252xG0GXWJbbBkLt1BuFtNlUvF8Zq5fh+
M9ZsZb1DWDARwZyrolPPafmuU+UlVZb2XQGPp5lQA6XjGQ73Ae3P55kOr1Ked40TlKS0ss23vDRX
qJuZj3UXHokvbOjnZDz/wNMDZgPI34kjVa8fiFjjGSd4d3vGCl79QQQQB+outR9Nct0Mx3FSATkc
iX8pueU4/qz8wbKdOyohPXHbmTYZ7xhbtxOKt9rCLUQXyFKmqB43Cjw2HnGR2+4hLrxAwek4vSRq
TmR3w7O6ORWHTBBzP406qUrvEm3Y1B7PTsoJNxI7JCn4mlEuX/ldziBHa3vGo/n5JCkJhLnQwXzF
+i6Sv4/tnT8+DmgYTN4AUWZfePofYDtZymqDDHxpE+DEbuElvLaJDfkJxkn5IhXcYD76j8zhataR
YpualEtgZ0ZLqHoNtzM6JO/shA9aIN+Kof7RnQFWlTOuFfNA6whyHQZEWPnoGYfSzMa7q+UJkS4o
ff+Ul4thpDKtbcQWKtntqR5JcXQDrjI73vz/93mBCTWDzgyt6SkgswCQw2Qu9Ja2IodHsbNtg1cQ
hweCwc3SSC/d9SEyPHQKTHGblNBlLCwR0UHsdLV/WDSPgnZS611LJ1aUXaVC51p7HyLooF7Ih4Fp
jmwm7yaz/SiUmBZiMVjwoyo6rFhOpBCXxPnVRTppoPVtb8o804crADjhCNvtg89dNVQn2xrRbwbV
1nc6S40//zNy/FqCuIujfHzLsLrBDyaNCrHVDogspSxu3DtHIkKzXbxDBAbyhbW22LtF+WWyI4+u
RSrH9PEXcrCBFbYyFiQY6WK1xCMBy7lQNpx/XlqcKf58QxbKx/CwRrotwW+Dwr0mZRM2TRUAo7Bp
wDtjwIKCCccL1BjccbwgKZc2PI5+KuamqWwaZu7Hb2oHseRsj1xwrr9zqa4Cs0vKfu9zw/AX/Loi
xDqQ6zV6cFRaSxayZNKm4yqqOWUQASsVQlXtrq74iLzwDs1l8roi+YmjndKn9Gjiv/n+Fhg5RnZf
9kHSQpydEAb82yYbU5yDwgbaDqboHTGUL4pdcqJfkg9UWJrhd5LkkCivjd6eLEvP2E3ASurTnQI3
HMI56Oe/lndh3vRySaAj4d4rWbIhovsxjCWd1FrBQWSdPU9hUkpgg4hUwPkEA8pL6zWhsU7yKFMX
2FGubHSRI6a4nVAMLWjUVMHUfzvPBsv9r8Qo77aemUdaJM/i/FQmQRqEwCxtkeBqtvPnfAPiShai
r8AxzmVZthn818UN5k5H309xxBPuxN4uAg2xYP3IZh4V32MAsbawbhRrlIwLcJDo8c5sU5iW5PAW
O5NuPChn2lz4lKN2JaA7O4BFDbi5Yh4K29VLuBxWkT6igQSu6U1XeCYOQ/WwZEbP4ay1M4uYeqxr
LEhIsDctkWpnIygPINWk99JKqcxrdsBTA12eaAcYaxCKjbiBI+UTBx7XcqbuujuURVHkDQp3lu+B
RuhlE2X8DHS5BE0r4wX2FXCNDLMi+aud69UU4KE8YR+YbrE2uS4Ca821soQXenUAzfUJ0ZyhuNdV
cXNVcDoWapF+a1OwsoOHcWH0d55RUrcYN5/LvNsPX3FKUmJKbUOhoKdlJrZa/7mYSlizQfbnXbWg
CZ708ZK+AMxF1QXWBaK58WfJQOCHezRLkniAW9RW7lTDLBK+lvuxL41VzhH9w6GjASpKf54rM9Jc
OvQBLyk9KL+UtvaPX2fZvPZZejXvVVpG9uES1UKyRbDRwO1C62Pzrhfpu3YmiAyb3wTwNeCJZNFR
WcUHi+t6a9FGkFRE2OcINOX2ePTQdiwsUl291m6dWt2rNvc12Lyw0AT/v6xyBLV/lMpzEW9CmT0Q
PX0LthwDziXA6KTNl3dYu67t9FKeSFeGMFyuwoHr9Ar6jI94WyMO17wr5UROoIP0U88mvMj9qAyL
YWire23jBOH/ZSqool5PQRIJayH7YUx7qwHsVw0lRGtb9yeck1xECGHWV4FOJ4JScraMi9czLERs
phdQ//FhkiKjn9nUiSxWcv/LORlLRNg3aeKdDjVwH3OylNZqIhSkQlmeNhGazL2wzh1grm3uYyRt
UYCDPVU0nslj55D98QyK0EKFxnqTZkD51IkgE5Yto/DkChblMw/ajfchpOs5HVFY05heLa9A3kj8
rmHXuj/vqMAaneEL8QYPyoYxBDPP9DTMK3OEyJPclEcS8sCZhpfCmjPxWVsPUJZC3tZuvP7UHufk
XUf0wQOlt0b8KWGmPZ/IsT5tm40HX2zbR2cDDF7kWWlCaO+pQKR+0f1lSbxqxrhvLIwiE7ILffi7
xpe5fwphO3uVE9ZZD1fl2WhlN0gB2L9eefS8OqkFG9w9yyKn6nSZifKPLYR4VbPHP94MVC3ys8IG
hl0YxP8OejzfI/Ksn/qHmb7q3+dbZk//X9pQXy5ZKNjbW+2z1TaULnYatTy6n6vkdxGc75GvoBAD
Nrxicx+rfJq8qgkzO5XedoOp7DmSlD11BhejY1HGRS0QSr1XdH8Y7Bcy2ykF/Svdtahn2Xw4ZE/h
tAQHh4NYSqSozIKjppSClcIYI0Ie8qGbGodLXCXFynpLydfSXYqAw0U+OsNY0O40vtWoDvQ71Xzc
XexPZU3oVBidNiQqaEwNk5tJFa5X60WoEoUUbFgoUbOrsgIZuwPXetZoLZ/ZAl805paY6kVT8AK8
LXspR13NCIPJ0HaI7SqFJdWgtqVyNH86Y8YkbC9qR/tlxs8nHnDksHV21SrdynrbO1PBIK9Vuv9h
oSUamH1mNB/3tSMTaXg9ABdQf1eHH+0LyRkm8HWU2cHkDRxXlhlhKPWvx847lk+GO/r2c5VKIp87
iUhhHYT8mLKtzPcSAWQB2mhpjMd69l+lr4ChR0i9aHhQwIJZy1nB3GhuA4+1yApZI80gfAJiNBSQ
v8+rZMKdnpPm6aZaAzeiIO9+2CAEa4YWVPKVx+oyo6tDQL3zjQXjHE7jhEne5CbY5JXMBmQS8pYB
UwtfKM55r1DQXROmDendViRmhd0GR1ZDYjEUsTCDbMMOoQ4wklehwzrHEHuP8wdF3YO8y3zg4dx+
p1+oocGFYt0KGUPD2URGVNJeLxqoadxSBGPFMz2kffDzwOsAy+DsENSYnQd4/v675n5ereXz7UoU
TGvT5WvqregaDJYTO9nS+D5sTv5F/RW4Xjwg6qXmLYsphmLt0PBmDXr/rRLBcZwUVFT9Qsw0wlco
oDjWZ8BI3mXuTIhPC8Qb4cPTdaFoUeZfYziZ1iifgdDu0kpkZbx8RlaNAeN0p+U5xXdPtHrSpZbs
CGWflCqMg9RWg1CEJ3VO1W1dIRczQsr1tu7mqcJHrL0I68029CO3EiDAM40O8uhm1/3D1B++WrJH
dM+mfTZ7zg+IbeSCVSc9kCqT/a7xFyg7+sleZsLYbTNhctpst4cgQzmNCpRbJKfG6iNcTfNx/xZ6
CprWfbsJXykNB0zNxr290iracD5wPsMBIsvHcCu62uQ4/WzQu8tDF1fg3N6GF8lwMrtxgtcmNki7
FvnSQSAt4gYsk2HJ9e6gCem1ZIWWbLIa9YrdlKbsh/qEOVkBnEGwQnIk03/s1zMpeRlfQDdRSsxv
WeM6qxuammmE7PsUzk6qVaF9V8AkFs6D1Zut55uGRze5y5kjsw+XfSM8yY67YegqwoewJdnNT0+z
ifAwNeIqWFswtPG4LyFf2bTdiHIS+wNfayD/f/n3YYaaQEIRL+0FtSnYH7As6LEdpJhkyZ3o8yNu
WhHePanOipKhyXS1S8IfJVXec0EwwFEabWsyHyG1oOfCey03TDS/xIsj/jhBvXWLEODZM/pgw5hq
WgyGs4rsShqnR1Q/hu/CVOL5LxrJ7Aw/VWz+v1UxUuPj6abhnOOmpvk10c75onDGTulz2izcuUVb
egItMxo05sEHmXRRX75xcXqOhC/dd2fKZQc/7GF4kmKTJtdBjzYYcV7wJ3ewQ20aoCoKyJCrjZjT
L4vFtAiGVKZ31AVQFYNbvxWYvD5S7cEp3gKX6gI/sVlahiQDM4dIFOHVRIcjElSel+LkfulxrKhE
bUTwkWv4doEQvYekYO+X2ULNhDpKbcuyM2MO1Z/K2uKQJuM3MITgDi3Uuj1KSO99cp+CgqKRwFRf
iWaFAmipYzejTT+54IRTI33p3MxMVxzOVvpv/8gHnwojoilqhT8kmeszawBTHTD3KL4aaIHfRdsl
pjjx03b21omPvYgpp2Qb8pITJMLA/TYTeYMv0nqcEGWtX7GIt8rstgiDpQXJg586k2EaiyKwtVLm
t+JWt7q4/zoNFMUTBo17nULh0vVJWt0vHA/p2+R0XAYqWFkXQdIHIvGf3PN6HpJuIEgTzHRZIrYW
BFypCVSlOqfsBOudXeOmiDPy2AE2ZZwL0QRkqANXr0c/mRlx3o+8bHoYCNPfqNuY0TVj0lCOaxf7
ORyuCpNmMaCkqs4qBFphpdG9pyOlFcPruNWClRP/40RiQR3fZQKfga2C2pUmNoOUtr0rwJtRbNZ/
rGAHpqckPBX58XtnLFqvJ7BnyGtTOY8zGlwYTVkVBWRZg85GK433O2AwJp2I7ZPHTSR7ae+MSZuh
P+slSnAVt3gcOrHTsFxti4molFd4xbsw/bO1GYoPdt9HCxjdQ1f3gPJMunSFO+NNuUdDVyB65iQs
O7tnjDvwrG7eNRQXaQ+x1hG61bM7lySNGG8MrjUfag+ZIVN77uxM/sxzGqOz7jw0useoMmwQXOEH
6f+Gfbot1+cPss/G4m8jQ0UdUvSeYCBp3oQN7fjWAvbqjMSeGYQ0aaJM+9AwBpEFdelddjNNZpqS
Pjv9a0A/amaoXEuheBv1q+v+izhzDDqyPUKAxdC9V0kPjk94puT7FQQW1HVt4ETDemBFUaehCri9
SjAFkur+3WY/jwCFjJvWIE6TbkUG73dgPegMTdibu+IhnncP37e4l+bU82u6mrXbhtXKAf+xvtfQ
x+I+hqvwDF7cSj/pthxfS+/XTe/8V4rFNLqj/YZEEjh73Ph9u7WVM8jMkDCNYpzrg4fUwXALTMhR
vNRIHMqa/gCF1/ui/8+1y3/1JqtR4V6AxOunkBn5eWreA9dLk8SLlMuHHjYfqPDayg9vR18aalYI
6cHJCqkG736VdAjQFCnp4yuQncUaSqxTzLNUl5pseUSXC+GUnqKVBGQ0nyJE0WA4qjTHfYfmqlPd
o4iZNZFZ1ypmcjzZw3CCj+/fdJ4TDITHmotdfK1dLdpSVpAwP5nPQfCbjXbDVR1ZMmrOiQkuxZDR
izrWF4NLjBnSx1dZESjjWfenQyNXvY89lMwwEJzYp7gqKW6qqenpzJ6k4WAckRuflepx3e+PZ7IC
OTL3CQBDrBpe8HtQT0MmkoDNXd9roFe5/btBK8wiUFS40DIWByDao+73Kepf40WmjD66q+6qwUUQ
aDNZ44L65k+BmCkHWclO01xQXwpZlCYE9yiyIFLpUgaQLhe+kRVLPKO08J1h2jnkZb02oIOdx8IB
a2haYCFy5PKuAs8qzzGT/drlxN7JiaCdQUBhY/W+wLO4cktdTa8U+LKIfujiiG3n1NJd6XFlnWcZ
JUeibk8HtFFdj9AIGS5xWdhFQj7g5dJjYqBkXNDkYlqmrYffLuO4xJhxWZ42jrUPhc2l8QvYTMYM
vT76wxnWZHm6U6qrX5pYSylcGPlmRMghsSNp/nHjLHr1YeXOqpFgsKBnGh67sSu6+pdohzXB9861
IMdcYg9C8g4xinpeYvfwzR95vOcDf+Ztb8QRAXNc1mZd3q3CuaR/piM4fCpWhLf5RpeIZvaVgYQx
kiwF07bGlV03CuV3AD6+ZjZkzgXyOQvddknRYiS/6AobaRXnvMamGmKUF+tv6KkHf7Bpuktkf4FX
YAdVsx7UAOYcZmxib+sI9myn7FPYIMEDYwarlPTolS2JGQ83Fp3250+RHzN9fYyKnpmrb9vN5s2L
NfpD1KcDkZDT52vVtje9J29dAF9KIeT70UKcymueKu/g+Pg8yyZoVrIo9mHTv6pw2Fo2dxE/I8uV
VeErqX0GRfGBhWD1G5GdfRYEv5MGpQtN2uXaOnN3R8VF94C6Mcs3N6XufJMfmXYU
`protect end_protected
