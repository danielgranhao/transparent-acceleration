-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CH3/DDnKoSmf35PZ6oc6TkaC7sPrEmVX110tS0YMQ2P6TpwDGamkJV9+/352aKxKuLEBDL7Zl6IT
0tc1ZzfnpGYQy2rGbDEmAEhPUeycYMaBEceMlb3oXrLiRGr5lJjyr7BDz3sC1TBlW4YNjuhoIwxL
yS1FuoKEwwwLcdFcAerqvrIaRAGC+XOqZ9EZIFLTACt9s6xehVGrT/FuUBZ5eJSV1+UMLd8KKR/O
8NNji5pHzy9+VfevBRL+NPPY1HTCS74MuVnwmB9ok26qK3b+EWJ6xqzATJ5OAnoiMqpkwPSRoayK
s3iWsVlvgCn9Qh9p75qQ1/4wY/SFuHJJF8x60g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 30000)
`protect data_block
2Jqw9EvSgijjAseo4WVvTe+FJMcYWIUtNQ/PitCMAxQdm0Ovx1vpMg4w5iTOULDUnM9DYBKVbm8Q
oJe1EuWt2mw/8YlWOCK88H2dHLt4IuvbrjBKLdJMeFq6wrNp7BflfcvHnFMjPhW2V8UvkaIwFYvO
4GXljf5khEoBzlQUkFnI305/EpdTnR0TVrJ9+qUFDkNwKmazGhZoVa3QTP5RS6JH6tNdBHBQ89PR
c5uI2RPRpeaHoxFBXWjfV03zAKW7q5kNEG5g+WZFWOCvzhssAbr2xSCuEdmdu831X73aL1beqK7z
cssW+AVQ98jOeQZwO+pxbDwHp+kwh5RPGzpqinL2928goly1l/VpKUjqEsVTDMvcKrfckqP7ZWot
NL+zdaFUuiJMfodpjxdulqbjC3ZVZBWX4YtSOai7EmnlAei93XE8WSO8tOHCIO39qqVrG2ke7iYL
hsT2kM9zPUYHToUWYncf26tb7kq3kOSVdZMsAKTpaqoc268w21aZhqssMcmfIvapcZwTU5Dx98XQ
/y/2nFnT4W6bhVKEfD4rcemDf0MwK1N0bxotbhW2ETR6qr4wcWTqzGqmZ5a5sdgfDC9ydnchRAqf
Z6gFIa3uwd30o+M2GS+HlqMptsq3wwz5pROj2JQOt0AhAmtuEAXg/6dgFY4KHOv37dpMDX+2nBir
/ijYyMSMrjqq4yjCziVrMKCJwEloNsbH3ybRVxdiuhR+KUmL1SBWoOLxiLvN9mGej5ZxuXh1SRKS
ecaGoYGIa5csqE1t/k4lsUzR/0QBchNjK6ygpDd+FCJ2UkwWv44Pokb9sBkUXws0NGvsWxN67D4J
U9onZZwHiYMfiaUoUXShiXL9XT3JxoSMBxKn1ZNdrSOQql/7GIj0EHTsagVrn60SzTknQCZFKeS/
Sg/VuPBMwi0ees74S3m+gZWtta142BmdSSoA7LQqRiAUnX/TsvhZwC4APJU+dSM07vuX/zif9+xE
Vwft1RNq0yTnmb706FjVb8tDYqg+hpRNT7ACEtoIKXjEEJAYi0/BYlUHLdCbK4yHlGvZEPjIA0xk
+l0lfMvwgC2lBGbGcFIB5reUWqUlt5MdKSY9G6/Ru2Kc9wBa0tNSvVEMeooTeCbUCY3Jc87CPdPh
uroPrW4stvtXFMvjLaahp69NhRpviIxCwxoeQfAc7Na6mqoeyVr2Lum4I95d2KVX8B/JOt3GGzNC
FI+wJ0CwIDWPFSwSiCYZZPn0cFUDDyq4vDbowCOAOwbwwlbiJ19wecNxYAl4soVoDljBaECaUooB
Sz+dlM0E/XcVpvx5TBRxiW7T/XMwjECcjsvLEQf2kRabkLEKGqItOUaXdRo0H7+xR4zongOQxlX7
oFi19C9nrVjETLpGxdK+copN35fnVxbSY+G3dd31tqIRjcTtODWnEJWV42avt8X0/ym7RpQWiT4n
DU3gUX0ycEXAdJjbdH4Zu6QgLXxa7s3o9wBeMArHhaYlNi/3EeFr5LkdMk9TjDB3kzKLk9eJI7Id
eE43iihJ8Aw+KouylPzvYMTX5jLfvNEBAqQt1/sBQ1nm2uxDdDaTHbBUGTowNELF6kCh9JR73PhA
DiYT7ACuDQg82pT6DcI4fe7nau5foS5XNmG+kJY4T/VUshobBgTJpawiI1o/YCkjWf88T6W9qkO5
Fu+6jMBE1+ztJavloc/6Uk+ew5LIhzzOXnXC2la8QWMH0NnHZOFR6W1bVt5rQS73rmpbQjvBphPG
FdSrOkisrkzy+YCEPsKeEzC+VXuN+/f9+Iysl1YTHmmpLjcAl+FDaD5rFupzvjPDDCPDFWG3Gz9L
AR2dO8kHLE6LXsJSNDxi7QgqfxgLt1E6KO3PQX/ZbsVEloIi5Y1I5TUEgDnpmywDmUQO0kxO8zIw
Vpb9REZm0Gf8WV3zqAFL11fCeF2smNJMy+Qyh0JmlCX66I9TzlRIGXPnIDUR4xaya5LqviT1HrDF
B31aDHZp9xSQ+VIx8tbsXWW2qYAmzZhAk2vfUM8J1qn+wcybu0lx95rgPAeXIdgB4/Fpsfld4iwN
2AXU9HOv+nhl1Yge7RmGGs1Eg9Xrjo2r5mjPvvODunmXeWUQzk/ZWbsNB4DnCcG6+RIc7WozdWbV
ip3Kx+xCwhecTtwa+AMPGhCLIuGygRkcH29WrwvTAUtpbMyScSS/lFg/lvwXQMYqpUN9WadeoS6/
+jQtVwyYbJ/blg/wIUrvuHGMM/dJUprnHO/j8Yh6dlRERTzp7e6ZEDIRs+bHCl/rzuJXppd5Xurk
VHROiDz9r/9OSo0UvemsfsOELVuYFyqVTVYYikhkKab3PH5P+rDOKEYTwTPN04ZuIX/U6n0Wr0Rm
6j9EE7KUKxod2v2X71T3d29duwAefF7CX3QTjiZSLppqDjXoeNy9Ugmy1/14p5fQRYysxVgo6SET
vmS3AF5NCtEtQ5vCarTmPTO0La1I+oaPZNYjm6OmTmGiBROPM5AcUTB32RmnuVnhizY/VPFni0BG
FDYccPaiDYCmpIZqQZ1G3Fymupfq7Auhug7azRBfRm6gSFyvrwzjbTMjKm1xmDFOCo/exyekVoWD
6uMeZuAEGtuYMtNvwyetAt7BJMFbD3EagGr6knVG20RswQGKXANBtAIEuzKVatbG3voNK7hbcQ4L
aElNU08hipsnWlhJN4m00dnfRDXi39w14sYJdqp7AIpIpq/JuhmbyzLAbobYqzFQvespf6o4ouAl
10czw7oWCGcXLJYNx5wD4ReYP7auDczoBcgyLL/TbDtFVk3LGa5PZTNsUzqfx0LFsoIddQNMHQxZ
kOle4xyYf2blrr+YwzXX5BahLi3v5q9OwGlQinuDHUF/GeQRB2cgX7hG6aSqPqoMDxTa/qOGmu0/
e+RzZoHEawFh3rD7Jy5zDxBnOGUKWCKQWsJwoAiPbjgpb3eh35O3QdSF8U+cieZ4EVy+A5G0uAEm
DvDKkva80tZPdelflTzTJdF+GcnZ/iD1+LuIee2FuePiJNuFg53KBhf+bV8hpsmxS/47wgpOpsnG
UDYCXkKhvNGwSsKTSGFwH4VUItBQnHJwP2J2tlDItdTE8loe3aySRW/D7K9AQhJNBYXP8ya4PqCm
QsYxf0p5n9rk+TdKXw5Zt1dQy09M/c9LvPZPJuejQou55N0YE6qmXgLZHkxBGRNpxKO+lEDnU2Vh
gs9RSf4hJ1uyf/LWTHluTnJwSZdr5StUHmjWj6gwMP6kdyNvCM4hS2VcZ1Ys5KThvEMrO+/8vX2t
vKMIZo7hFxSEqfKH27GfSvPvOmbBovQCw3nYF+eJSF4i8zWc61QYw9jj/B7V8oCv4Rmh54f6fN82
6oksP0JyxzYCLoop3Z7fn1nsnsxAIXZrjMsIsSQ3sHaH7XLNBcoAiqgPOPAsLA0n6seIpCfRRMSM
k7iI/NkAE/RKy81glE4yiiMPdrEwlCVNA1YWAgVRtpARHm1KBuHeARJ1L1MTaWcZNplDnnT3KboM
WeDufq7aRjigGTFQK3oNPgv0X2050c76iCwij+hr0iXjM0kHcjqjgSS7b3AExJSW5KqzS2B1m2/v
7UvwN2unB4bMw7xJO8Qv7eqjPNcqTTnxE+R4jXAPphLvL3KOzhnaj09AgHuciQqo1fPLWOUF22/8
KJJXELYo0lEO1+LCOsooWGCHL+J6RGKC4uG+1i5kaaKA1jQXFOlhMLTb1WG/iBufVgNrRf5Z4JyI
Acvn58OmZB2m1pasPsn/Ryr/YGB0z1yCvsGUOLl7xKXwS7yGqImNrLQTX+TARfdK7FOnC1VOp3Ma
N0IgIYEKedHjaCtRDRuxp/mCZbSu7PgisqARlP421Zv5oPld1oH2z9YIZQHcxnk1JVz3MnAhJcqZ
rhpVZCuyyHkzvHaEz0eyiGaP6PBouRB0d1CdG6uU4Rji9ClD9rrH0sBqQhS/teLW+IML42FE/bGL
Y9pSmoIfE+zQ8ww0o+9TIYTtkjx9XwSaNK5Br/vf9LdOV49Pz/qViyK02t4JAVwUMlD6ikRXwat3
AQKGc0KMMxa4uTDnXWbRxaiYxR160NYxSP98fjqt3Oujc4k4jf6qqpNywGIMlKWIheIngZ8YznU3
AcOSq6lRb9iC94DM4bOEFA6YIKK3oHVxlEEkHfURi16if0I76DgcdVRm/eoSnAcoehhE6xsamqsu
nN9J//JZuDflOMg5+UC3Ov1QKir8uurIpqhBqAE2JrOGkrf+tQVJKraYjVRWe+uMXmfqHt2vuZlH
Ns6tLVr6mHnGbeLFgGMFpiLIFmnOOgY/mBdHxcFkP98lg591Ov19sWRayOLuqgkf1zM0XKmYP8Xx
B6cj4GoFwENyFUFtL6Casa9V+o1dY47TS4Zou1m3Gh7OUcd32nFRKatFdNI0ktYLhszuGGG9VUt6
sn7cIm2vLhadWEQrqzmW9Butk1S7fwYynLefXVdZtlwbHj/bLr4yuk9zYRq231ZmKvFZyValB5qI
tIaOUHWTEEzkU6V4nMft1ZteYQaOQTcPeMdRfH+IHyeLEH0sTPd3Y6IKw6td2GEJO1Stdfg8cLSw
KPgUqJrEcCq5xh6QNBdTy0tC45V3jSesrMkhYa0QaPTKbmQvyex43S/8kmWHEvwFPTFba4aKVrX7
MlCZ7B0LTsrhxolQkFEhnEOUYjoXkE0eNs1Wjc/L0k2XLc0LaG1frj/fRejLrAqzYp78M+vDRtHY
39xTP7UJywa9nJxpXb6cWFBGPbtiR6t4AATsDOeBD8Q191RoUZ1UcjASuRVmXcXpmlbb+g0QF+BK
3i0MDBwNI4S4zGtwCz4AIF6jT5bQiDXs/CIOytrYEehvj5d+K24e7+RqqcepQKujkbsZ+Vru/XKv
hlfuVpVxmjkrTIrvfNXuXsuTpeZjG/fjz1auop86WCidSANeFa92QsSgXLXNt4wf2NFOgEjzpXjT
CXJyPnlVGvx+TcXgWhAPKPxyBFdhBLwx6Z3f7d4MumOeDO/fWPairtQHHF9BDe1S4U/eYUoy2T4o
qB9g8TXH8y4w0OuP+O0z0OWmMoyNcHNleEGyTAQHk8ulTKw9nWwUxzoScPdVjU2LB9PuJ6Smv6dY
cQx8NnoRDnzgomKyBuBYAQg2jhjxzDGs+uEbhUhP+NTihTdvH9YUoeKh5nRjSFQ1Nj3/v7+YKOGr
kil4sbw8kYTwi5yXYF5Kk5gYNgc9eAK1PvCDBjFPxFnjF0COMLWoq2qiWEa+/+dDmlw4YuBa44tT
1+7LGQqAJviM9encCQpwy62I4Bk5CNgxk6PWs0e5C2aQYbUHXU1tqJHclrojb0D7Q3uLWLPySPpm
pIyjzu/tzrVyf00owjT6d8K6Xw/57XvjpiHVvHHPsvNy58eZn6haUZhzQj814Zl4bzJoj1P1739O
pg8zDjEsvCyYOClZZ/v9r351I48CqQpmb+njUecT5DgOFK693y//VuUzmsX1IW5pLVNjPLdbfGyw
CH3pWKkuEvaSzy8yn1/gJSBbZOdkDuzIvWsI4R+lq4Itplaw0yB4ys9G1rDrkuOd6UPQPbt3JgaF
dSWVB82xmpnppIcslQXqnKf+jw1pJz7GSN3T85KuEDSGAjASwaB9GCROvzOsrlF5Kfx9/VMLTVoZ
pzRfWdNdb4oD4e0t4otZtAGklmqKwhpZxZqjfxDPUhe9EbeWoinicEcWRdmWcI0nsTj1n5TeqiBE
WsPBomxCR3V0CytqUvVVTDizessdqiEP97EF0BBSARiC5FnkbfF4hhQSmQfe5nOGBgeS95dKAdob
6xt2hb+G/aVJBOw7FcCq09mKyW4jubUyUrkwKC+STxOVyP2rH1sf+JinwDE+YKZhgesHcabj0lWC
D13stvXQ29PCNrtMCF5O4WfhkVEa7MzZBDYL1CZFsIOwWGixbrM722OxUaS2pfCykmjtt8E1SRB/
tX4NxEocRzBWDKOOo4fZFLQQJD9o/QtyCzkTxSMGRi+SwmWF68MHwf2DrLPIGl2DQHzYAJ7khbwH
3wAgMCH16+paQGodJ/ScyFurA1HmKfjxfzqLpzuAbF5VneZ91SH+9DpXV3aQlqRyhuS+yhWDf8rF
zv4TKQ1Jxd4XZN5Mw9K5Yim3AgSmBYkXcFdeMVxYX5VvoVnvpMEsFFi61zJLnKsgY22rVPQHQwOq
zw1mQuEbgeGKrToDMG28maRD6YMV2Jw1otB+vaSh4kQF1jWJmaI8XRR0GFBc8TCjsspNzXLNMU1Z
vvK8SO0XL3OvOtZWpRTb4UZG6gRSyPKrMVZMvisW3FKwePbICHRabgxh7vZ5tFLAFEczADPK+a9F
S31kgyQD2CvzNwz08rrOQBG4HryFf4d6vq0Ueqw1zYJs+ZHot52tfSh0OlWaeTKFewBA9wb1oMIZ
SemutBNduFVC+BnNm5skRk8htd8O0uzyq1ipcrOxfg5/oMUeQiio+m6uqDGu9y02PgNo0vbwNJUx
SNz1TZypSBsIcl/KbZ/X+At3SNeXdDk5LkpYs5/G3nIC+US/C5nI8Nc/R5iMhDlg1GVTQ8GfofIX
5+mi9iDBVDP1mJxj1TO8ugkgKtHqhYfaKAN+3WTMff9wk1+tFyTw5YOoHHCUh5GuNWjXGa6sbTF9
V9SuuwAOkGtCZd5fdi5mkkRQnM2UPTYqvK3MfOuGzsATc+AvuSdM+nsBmeWannsIJrjSM8p0HHkU
9rnCb+wd87Mb25YGAtKsdG0wITBlWYRxHrd3r+v3+4IrRJqbBdjFP8mnVOUEu0MNKpqgG7kWAIT9
Av0O66R10FoX9LT8g42VScLPNGE7zHiU/GWIZL/EWB/WyIAB+9Gz5zqMLprccigjaXlhXOADfCIQ
VnwmUTCfOGrytiB3B8pDtQu6lyaYNurSuC+YV1FyIkKCJEynu2nYyVVniFtFWr+tkTilrQcXIMvG
rMK51+2MTSjoCo2ON53/scQ2Zjr5+JFaJG1R95PYX7BuFbCZuEn1E7SDQN27cPIvQ2IKEO28H2ER
qwtjB7wdYYqKRBcg++43D+ChxyXBf6PxN60bU5tI99mLjCblVu5ctxLy8amBOoCmMXEqQj8LiXVR
3bgPZgFXptw7SQSzl81FbBfEtL8a7VBcPvsIFaQXOkyiUINc2sfXSgsOvarnDt283aBzillZ+wJO
uOfmVBPf3qF6/dZ3dPeOVzj5o0CBnP8ICS360sP1yp+EPtFI2XEolLZ2dVs3wBAPF69nQ47/n5yi
U1bEhUqqLo/TfgoH3AmIAefF1C8bPPd2kLi0JwwAEfrjB2KAW429F8kHWF2GDQivKuwe37HHQ9cY
pW7Ags7iYr7+5Hxn4Ilm5uxC+vaEWpsFn8f7LPzfB5rOwk9xY0vnQdaC7KTPXlQdteZfDIXh2C88
dXSaKYZOsndFtig3FWeQdogkF3XL9/dsZI20BF7MfCLzGsfG5LRN+wqAQPBl8MqtlpdsTiYaa++J
jiIo5uI2yIzQdmcx/5OC/S0NJW/xRcKG3RPXftzgCDym2fRkCJxLgQLrCP5RSd9Xz154gZmmM9Uf
pIIG1GNvjcdZGA+aqLxh/C2YeuBKIbHLES4cqiR3cT7X/LLiBMfQrfrhZgjDSW4mXYLYtoCrIsMP
+ZFkxvJNAfUo3ZXrmFlxGzICNrXMLEZFl8GtM/0zy1BmwmuQeHwKZK5H2d2XJRpzpwVX2caw+ZQr
QH3bNRIcPOjNd9lS//gTUxyX6vCiX9mfS8Douu3QYJQ3M9FR1xr5QlH2Hvy2nq5m/BJ+G3Aou4Om
+oZkERWg5v3RqeEmjuo4jU3P9Lf7K3ChJgDxPadC2IQE915AVIHV2EDasy+vFLPa/ICiApBQznzG
LE2HU35QKRFcSS47XAmfeS6i2BwLLEgxfI5KghDPCNMy3g9juAEu8/KdCg7OEviJ2lobBJX9wmZh
nrgXO2WTAlcPYMkscOQOh/Eg1oCzgOWIzkXYsnXm0M8a9jYTLCUkIoJbslf226xu4flo2XbuM5II
ycekREv2d5z2O2ZXJIZSazYm7PgT407czbJbVeNc6WPfYgeIPA49DMXQN7uWRm3tE8YvpnkGbZtS
sYxVm7b0qK5LluaD1uvdlhB5sxFFc+kQ2YUWuLl6hKWInua0mHe7souVs2g6sir2wp4wJSv9KlZr
lTtYQ8cZLOFeG2K9HdsKHssdktP37EStPIYjBeNRQjKg/adkN5OQ367mgjg7JRUJGnt24ogqsczM
hTEJjkXmstyaqLHVsJbYxTKmxnK+FxU/fZ77p+laddIVaLH1AMwVb7WDScbH2hBCQEaC1Wm+qw0T
X28QaIixKowtm4r3Ze7RA+CFCFRFZDOw/Gf066i8chJisgr90lgxW7abFWVF19aSIvNAtltJedDP
7zMQSptlZ00BuEShmN/lSdVyl3L0enPCn4DKBwZ1935BjE/QmtwAccYT5FK19WU7S1GQnf2v1iHp
BzIhuKA95AiCPSmqWLQQOk+wyP02VGobv8Er7Ct01+Umr0UHQywnnF8IMN9P8VTaS+gJRxhoRpTo
pFSiizB9YMQ3DSeh9YnLsXmVDl1tpEr7kWlkz44ZrqW81lwctT10kCwp0j1R8fWlrjqsZzKKsPDm
URESr0kRNPXF/SgWHMcAmY4jtNmCcEqz4qcDdONwdSopDz/8GUt5lZ8tz6F/7njKJNpgNrIrvUjB
xBCiufer6fO5YLf3ozBB6+eM6cXCK3+z8CLZOIG0Ofe2CTL48jws7sO2j3fX7ffBgTQppO+opF+n
vFLNUYUrNK6XZM0flYVZp1xEtP5XQGwzLNStlAdAUm1hZG694lLQspcQT5w6xplKC4ny/0OtZ+lW
rJ1GdNJk86xhh8g5ii8DSvI2E4IuVcCcK+PL/eq9SQpX7s9zzlV7Sr2cvAH8Ac/S1/coPMhFCFhq
Yah97ioShJ2Uva7JCA+vKhspdB4dR/BtExtg8B/CvLQRctoHqCp1VuHuvR+AfAC/QzkpdFxJ/xjZ
afOqgXWousHM5DTFClvNMXlaYCOUsuFESt/nZjitaPd4l03yGFMSqFADASxPytmR+x1Y+VYQvJnn
hQt8YfHpff8GqA6StosWeQQEJyV977XOO2fT+Fg5RiDKpOxO97Cuk6fpPBIruqMBINjea0L7+3UE
vSdJh8H/dtnwSxZ7enO1CKxc7uxHSMPJXiJVEzBEmCFF6KxUUHG3eI11HBqsT21XzXfcf4GL5bS1
UZsaw2qvQ/How46xOtIyzJhKayI+dFzNEE2iyYHJAWLkbb5dUsdI40DOlxpeh9mReCzsnXQ/qDUz
hgdo8BGS4SsHJW9b+pTfwoTIXXVpHlmDY/1gIJFp1U5LuXIuh5LWXz7DqPupZYV9RFdVBu0fo5pV
XOikMNvWXQYgvG6GWoIPbRID4i9WF9k/Me3ENclLlSpK8f5pbyfeDhRgFJ41byZPS/Ar5EzSt9h1
NHK2hMlx4t04ladc0726mX4Jtzbzbbp5GkF9YL7llKnIqTUS/Usc/vvn9YgIx6q9azq1XDBUYpLi
hbnZIlUccIlhnSuxWw7OYJE2jXgnBvU5WXRQPiWSger2M6lQgmYIXBk44JXXhoUZMbla1FeUQSGa
flzcHjA2DHSvW9Wwadqml/YZdOtK86he5i3ANHSqDHgBdtnTJenHQKT7feaiw0ZmpBOQmOWYdZt8
5gVqjdSb7hIO8/+UPEZ3tQxP6IB2CAxC3VyA1z86VVdEBz7kniNf0WC+lihf3k5wtnUb1x4vgaMl
GPQjW2pRbiahlVp/vkZfSRqsZ6HkTo87Tqn2z4R0HLwuiENismUlYW5FUjUE5IiAnBTQEZ7SuvAT
PsxqHI9NEfH4s3yS/CitHVid9K5HJPFt8FLQKNr0oj8PE91Nn+dBADF0GjW53wGtAcHVmUR6ceVV
6cSgIfUhI46K0RG+wyGiI3AbwKqn3DTOxQf80E3DRvO9VwMw3p7IhjPgoGnLEDupJAxtlpCwEjNQ
XSu/0v0QF29xxtAe+yFQDxX3lf4iaY2gMxGMKw0y+OlYxGLIUYuSxybYfzoDUJtBXX9ahkP4O/7j
227VvMPlC5CtKp3WoUpt3hgBf0krrpP03ynqttICITRs6LVEpsa5oMhFF2m/aY8sK2Sr1eTILbn8
KrLp507LxF2iYv57t1bAGAUPZ/fGi/BQPZNjIpjDhW6rF8OY7A8tslH9EkFFCVYiynb/wUJeqmdd
lmmLC/iadg3qQ4iBz7wlgs38jlonz4uS/GD/cCs4fwZ+SNKN35AOlYm64jCCyznSw8H3o/pQcOh6
ZB7/xxiLDAU3cHqRuUgXVnwhfK+ZN3tvFZ/Sw0dv5TTdNXAUa0bDXh9gvUptFSyS+RzKU6zKcP6Q
DND/nE3h2RIDk0QJmS+lvwErlue1JVoQxDTi9sB5oGaoVvNu5j0016BsGIinnSVorJhPFPx/hVan
N7E9iTSMoX1GxiluEKKT6LE/RApW69MQ6ZQ4W72q/nV4BCrjQSx4XRI7G1vfEwIxVbrMTbRUeBMa
7e+7HZyoiYuzZGIbj78r5YzJShwGa88v7OcjfxirMyLo/K0MBA4JRWNaAaSjVD+GlZiJpX0kB70D
B1SnmeCGLJhYe4lBuZMq0nTsXacsVV3h6orYIF/mDE2/Icm4r9CrdgaHAUJ5jODz8SBZIRr1VYN9
pWnVj1X4/69RprnecjMiVIGMbUDeDJVfXctnzpZUo5yxSvqZa/nYekENTKdAH1W8G1ny+ZECJko/
iGMVatFF+zKOLUXOX1Mpl6nSnJhDkr0bW2uVkTYCL28XUN8nbFhbAhlpD5WXF3sXXvSxEmzkyquZ
UF8iJoxOuP7O6xLBO8AR2bjtaOu6I9YDg0p1BpzZgQxAThOQph2WF6M0LXggXiKmHw7vY8zsc8t+
Pse98uzMDCTruLltbHi4l0PU3Rjt5Clhy04CD/jan3Iy+IES4R8Ke7RGMsMdU18Q7bkXnjijk2W5
r46kqLGG+KkCKz16WiS2cptqi9FmlFeA5crBbx+f6fp44ylHc9hC7H76M+wj6h+A8Du/1hU28XDq
ZRXmLMk1EsUy9bJkb00IMy4PAZTfmZ0xzcoZfvA3wx8Ebcyv3RvWlv9hZFIBBvldwyNmakZ3VKJm
keiwIPN0TzZNzJYUDyqhRW5BmzmHmUtr+Q9KfE372i+XU+a/efmO+qR030A2+bWqcH5F7OOhS2tN
DZWBJ9fIOsRWVc+QSpE2LRSFy3xptJ3DUnCptdpNBTwnELVbC/CWKDq2gfxPq9QYp7/C8kUxYv1B
buvVGQ1pWn72opqrhSYwIoNbZ55OWjdlvXSBTKRwA9RwofrP6hFGFFKI/ogpzW7x7f6luKFrLr+Z
zaClojcxUMLUN8OBPFcq4N6VSOOmc5hBpTK5I5xJfMK6PmimDgwfzj+NPG28QmCSPy8NQT5cYlnE
MRvG2mXW5RaFDf6gs2wD+b0IoxIM6brg4pnaisuQwaBPNXYgEpwTqfItWO8A6GmC7YWwGwNTf0tO
EilYR2Cbf/lLgaBhpdklahD9cRmLq05M7nMQ3Zofj+1SbW9FZnu99/1f3f1zprBMVcl4tyz0ItzT
uyOue7vyydNLc2cLvO99WaflnWWtpizZK+P5oEtmd6IeKL0OypJ5aBD3oouKGFWHv8DbDUiids8T
RS4j+TqBDbuHCU5uuF6+/jXtDZ0+rj9Eae4Dc93oslolPOv86iUJfscc5cWRqWKn3wlPieOYe2Cx
pkcSq0rVH45SJB43kozvLdKJhYt+zlqhXGXi/+ii2HXcadp/0mSTkkKu29fwTFyE8V40LHQ42oEr
LUNvHl47XOA6MM4eLCZFqcR/FxTJ74f6ulvbmEsKMy8FsMBe8MYV7j/R11nZVe4sEZ8zOzA6lrSr
KkwvqKq6hJaaONxtog24NtFExLV9S08WH2LLC5o5sX43h4iabflEvzTOF6gGl/XU1ceE5jGMlYnK
wURAECKFYUiqhxj33qd59oAIYvLJTAalyM++4h8MePTnGb7PcuSsK1wvAPLa8QP2JBUsGNGIsiFy
CpyoIcmxa9rFuq+ichKrctP+KHWPs4Irj63z0pi+aQRd3KKnXDGXsOe95388ugJff59SwrVMElWU
g/ZCpiWGEDndR/qm1IQ1w7HiHH8/i8HyrURwKt8+8FrT3xcykervLOrDZISc0HzH/BGkiop6KmUE
PE4n9eh4TCZ7tGG75sahI4ofKNWYBnhO3CyDLNgInJkhts1i8rK0I+N4EIefYtBAoQwi+PR2fku9
uqi93lsZwIHTi2SeaiSWNBVv83sq9etPbVOPEuFMP/4DgOrr1afYzB0TOP5bG0hM0QcZ+z83OCSu
yB/RrqZ7TKKQrBH8+XCMBAAZAqji31xzDL18NBsZWp0UihmuLAdL9LP6fNEyr3nuKjTjWCP2BHat
8vsfBCxfOHf9tloh8vFrxOLNnlVyPcM/t82gP6ps52JBSmV84cqwoComieSfQIQ5WxvaRhMjZwDI
4IPwDDTfPaEOIuPvThVKG03WkIq4pCluxY8TmQhIkPHXlkl5OiK+Lii94PCpRoQwNpyKwYh+bed2
e7Fq60MnRfpHDIc9yH9qz1Ymu5uApH7wVVRiB8FKyhrDo2N2V5iCxMyIzcl5tImqsLTxGMve40uR
F90MY/gsK8Eh7HAt/M1jsDbhn+dJZA84EqVDH0PRUHuXsi6vX9+TnEmrx2yzR5MRTs/M3fqL/gPk
iJ6MVuURp6cG3IjEQViTyEkq/UGoZhXU2tSPZILOdIksnMkIJ7/EaduvFchgz4IEMiRemRtDj2te
tY+84S2Jw4dmr3HpIDEU8c2A1ZeH+mSk9cGbR7sLQTG2jG6J4ecGNBW+t4N6nA698CI5onJfW9q/
7HyTZxRBkFOjdixVDYBU8fZRAli9IqOVzvlXYCLd/x/X7nNEA4N/pEAaYvoS14rqV6mp9DjQ8TgJ
OTcuEa9kFu5cfHf5LG6aSZdSy4VEggyYjxJL40gZaCFOoTW/a4tzRLRjPgFljdV90QQw81p8WWc2
9K8J6sOjIxmMWHyqnDf7JeN1sf1i43QqSad0OktLa02c1AvbqZuV5JpjTns6gsxsShqLi89RjARe
sQOsyW9CfXpE4/9bGQKAbpNEm5JCx1wLXhKZ2cVhwqaKWGuAvSZYeacRHm6oqZw6orF8B+IFjCYy
z5ftbbpqscQwAFgPZjkGbBmYaYsyv4bz+r2QAe4JkHUng/uhc879+1qs8oLZ3jfbnIPKsdxVToeZ
zhCUqTzanByFH1gU0To5A9GPACh3hLzX1VUZS20TsesVW9KOQCzAg45XhQZL1C9QL0JrUV/a81a2
3ot4vYL5cf2eRzfrmfNOKfXw41tNYh6DOOIEcNUgL1cxnEQbLond7qr9GdSAxO4/oa+SiI/w9xcv
plzhtOr8ue7JkJuHxss2hU64Oa6B+i9vKWRpcDOn8zjHYCYBaJS245IQqX15NI01+9BE4775naxV
IBS+MV7Cb8bUPeIJaYxORFtenIw2A6zrgehbLIstNTN3AHg2tRxSx4ZWWffX4B+fy4NndwMtm19Z
oJEL2FNo4OXVjniswBFUdedd43D0UkOJCwu8VQCqoHK1i+LiLnE5ZxApkkPqUiwNHA+CZOLZS4Uw
+yaYBDd07bhWj+zJujS638/IflVQofVJXihGgNqP07bZ4CADgqaZJWhsA6ESvqRjHyBaWpM5EOC5
BQytP49vce5KHlGB0t5XNIJkxHOSLighmZjadjthXKlw554H17WZyBp07GEObFAs3Lz12oi1kHVx
1zpmt1aajdqgGMq3hKjKLr+4id7XucboPhu8b8zJRQRGzGgxjuA2+9pBRBPNba1M7imCY70/1SNC
I/qKRiz9xf2txWPQ9ZMq7JjwpSY+nXfaRe0NI60Dle1EpPqpm1xl4i//JDkb9v2V31tUFjpzseLY
wBWIbMYhTZ9e3IBRp1RsqtTi2+P3z47V0NgxGJG9WpsIZ+dSQOuGblyo0Y9R9lhZniF6DmIiwNZq
9m5i8gU0KvAPkf5cXpjCffcjY342BOx7jRMILAyCc6V1XLLxpfvLxXAqsdzIZ6ZJETOOTgxalm8m
VTEeXTNBN2luseTW5rQyMfSEeQIpe+IHtkjFafeOtxcZ0Q2niCsbDorOz3SsSHNEAHfWfNCUKYt3
iENKAKasneo3IGLAFkrI4qNUZnFvqRM8bzD6dqckGVLMh9bt+8D8yukUD3YJju59XIJrnc0VsqCl
VEI8t+HZFgXbxZgpl3REmcVKz9gIsbTHf3Md9qaZX1yCACRG8oCrQVoFmhafQXIWYy4QUnsemSzN
nkk67kaxFhEPCExIu7g0fLntbOG/vnoRpP7YQDDJlg2azWFB6i+uq8gcFFD9kyWRO+uJtCJU2uR3
DO6Vqx+vRwWiJMfMtEW8vZHC/HWyfctGc0tmWOZp5ohQv5m17PYZdVhUtKq9aKDk1/6zdiCITNUj
L6z0s8SV7+ToHo8SghVe+TncYaNnq4vQ+PUcRJwEWLg9wEe70t5AZCWe9+fPpWbnsZkpRim/4BkJ
pfk5UQY88u77z5hKXlmmdqbP4Inrw9vbkhJLwVKiQAG3kDxyirvtGwDQ7YrCqx+oB7IFxMjY0fRq
s5t+RFouSXJyxIF6MpCbqqory3RfH+tRzygu9RI8Zn13TqebUsWxPIPScDl9rBc6N6fIspX4uxJw
z1VAq7MuV+doBLaCC52dKqIPhWwBbgtN47BjS0uBdyEFx3mCv7aKmjrsvMKbpeZ1XVVnc9bQRr+F
BJAquUnSm5hBVlmrfU5Lsqd5+W3vdihk4WRse79bxbZw/6SfiSAEODlUjiQgGqZ3i/hXQg/G5gCv
IrzbnWTShnqbBFSeGK31AowpJKh6m+trjiumwsEsCz7gooUpiXH4N0WidHlc/+6fshHexQ2E4Clt
bvlhrgDsk2hixe6AAt0WylfGwYzVR+DGxTZOJr0E+PfDHYhmAc9kCArtL+DMANPeKoQFnCRcM1HU
lCkSRi0SK9VY4VkZAQfQauq/zcIguq/nO/Uzoddu/NfqCfc4heO24Hyrh/aecFNSanHTZtg7HwV7
5lCAm/typthchmi2RDMSv7nGA+R10fMXQ+cQnpmntHBrlSli6uv0EB+UGMBHeY1z8OeZ01Y4UrgD
vRQ8l1Tf49kIwVFtm8hP2vOD2BwQIohhb5V56WTcjUyhhX94P2rPJRowLQGYQo4J0BtiGELrp35e
PBe1a2bmF3yBvVt7/z+is1f1e5PXHsuGYHCMgTNjOg9pni9fnkIOKHkUhLlJl8zgM5EeUREixCcE
Z4vFEA4qEXSwyq83ueyaa/m6h71/xdhGQ80UmbjMupIRF+AV3C3tgN2DioQnMz2Q1pzr4bQsVJIM
XTpOPYSdTAujz+VsY5uZ4fCcV/ZoUUGiv7Dpe2sqdd6k8BvOEvNquUXCnoshMG0SzwUoQLqJfC3r
kveVaMsrmTQHcOJ7UwsiNmEjEDAv9snv7TZRbjhI3vfgNnz9Pox+DTSmiMigvly8ahvQY8Hm1vdM
miKTFgvMY1Vy38HEqAghHuQybsSgypd1yXl54TFYIkThs55MlEW43svwu2vsUvnj5Wi9FGiuwGzb
8QU/ZXaCxTfRlyE7oYpKsklUqu8N8Eq7g/byxc921AzSRKoEHdEPWk4uY24JibT0pctpyJ8C7Ruq
BK3MPYQ6HVgQtxO50HuLwFHienHxODKEkPVGbht/AOpoK/s1lOGOoMHkJNScUtmaXZzNnVZOEEi6
GdRWFnrj3+1RuT45jGq2ZFesRcGNHQfE1I6G0Tq4u0ENYtswKmFxel66lXxAvxffWCfawnICatLK
+VAnwaGYGxuDxGmPAnJOob7P59goAN9m+S7zyuKMkUsVFobDEgpnSn0zpXFBvoCFkU2+RgWH95Sk
nIn8CCBcs2O63SCnOEnPuNZ19cvAgNHv+vvdUdVgFAVL9oXCVcUKNIbIU3RTxZUGjozHsirh9GOg
fgrq+KYzSxAkv6FxXDxTLnwO0lTGEkpSXR885u4zBRY41+i5ePb83nw6gAQelJFfKbAPgBMj58eY
3Wy29UOtJZRiTnjSXxvlsNe5GWYOaM4MiveoZdGScandWMx3pg6C216M4VOQQQVoEOuZUcixip3q
sU1ZYYrdanIu36C4FsNP+rtyWMPmPySAN8G2jiZA+AUzdxoZ1RQ041tMJO5aquibjgPvLmqaCLVJ
WG+sCMG/rGirxoCVWwTUZ6LoXUJCvkYBPQDRvJO/lkZs+ipkxK5b28ZY5Me6N3eXucpVbOfRxi1P
UH0J239M+0TBO1nF5sGhKGNzjyDnO4olTd84pwLBOKzF0H/X/HqGsZ5h1gkv0O03hcoIPve8CZyJ
ZRzW8+AZBEF3hA4tVAZ35Y2rn+XC+kkE41qOLW0FbI1C8OYhMM3L35sy1/I4oAkG/cItxKFewE5K
x9lWt1vx6p2s5D5yB9Q46/EUmbFCP4UXihg+//HPmSzSqLta+yJRNpkjaQtfe14E6ZO5Gn9pJA4l
HI+SevCGMLsJ8ZsJLQ0clcPyozi1zk0LBlmzanWlf34tb9Ze3yfxfsojnNKB7vvtkGa7o5Zk0XLP
J41MhDmcetUM4V5a+caGw/wfRUnxHg1zbkVt4ikYhxj+yZyC4Nw7/Vfa0DACY8pcrrE92Xbry3YI
PflZz27OuGFNM3hQVqpbgTjHbBUQT0vtL3wBltyBUE7yffncsNd/0o5+cHyUkmqC9m9IVkgzFsf4
EzWMebIlheGWjKIJAIAjcVdnpSwdqiHUSbMw4CIQn1luMy9Z2wkAmoUR4WWCVO62w1AC5U8rDhXN
T+lE2EGOE8KtcbTvD0lm6uB6VywtXtEFeqkPQhKeV9nE3ro/Ku6JPl1WCFvJf2IjGyFlcktME/k7
8YV+H8tLNg9/gsZrNrg7jBZeLM6P1Wx4e6zvjaIvLF9VnwC1YJ9si80GnY2EMrmjLAJRyXRs7DOM
X1ExmtgLMZ9sltFXZ97KU1xMLnFkh6XF2d+280f2evypGMH9KvB7f9kg3o/nK1FgUqT9iqExtqHI
fvDMWCKz2gs9MKKDKiuc34Xc+O2o1KDtVjtbOou6/fMmiZJrlCnJZI4+IE4pHt6VTzPVe4laUzU7
dY9nVfw0S3m7YeuZWP6wq2riQvPP3Xd65gV4JDPYi/C3AF8EShlQA1czyn7jxnh9XFWSa7Uj/zHd
7lTrmpdAr9A1htcz1ZN5A9ZHfLKGsIO3zyPQIIGY7cAKy7EJGWuAweI5dnR5WNdFCgkTtZjepFcD
EoPzEnIixIgZOlVuafTq1dYWyOvTMGE2yRGNqYr1YTHgkjZUe1MOcqilFhQI5A18Qnv3axOUbl5T
Oo+WyBgQbP8l7ELI2zv1AhqJAiVjUEVU9Ad7yL5CEqU8tTXPl8sag0F9JSWNixoQkElUco/CSSQG
8SnteS5M4esAaTrJMAvuPfhO3Xtj+WHYhtRrFlxx+j7n3XNEUPQ+L5489Z7CPQEnOb94G51o9OME
OYaKqgnDq2FZ7injIum3SjknW89yjrwqLA4s6h5YUcSIKBZaMfIbZ8hca0MmA5wQbFH3jZZztbFv
cJ+uuIqiUESbzlCMYpL1D4+Bj+dOvOH3YYGdzH90NiDZyVtCjME5yWxTKD55C6tIXS+OK/kNu0eU
y1W/u6+ZD22Xv2itcUBDboRxP58TnwaNcM8jW8swPrale1uwy5EC5TbBBf1fQ7LQMTN3aXHieVaZ
6QCcEL4jt3QycuoS2qTiGzjk/De0FBRw+aeWzrGUt7PGH2tJlztI208AowyRqwj4L9GnMChL12R6
dXdIwLqQMBF5b/+n7qbtkISHxnc0ga+IEx1KShArm+hWK07XRwr4f/sq5/DqnzikxhSNZwWR1WC6
nO1dr/YGA9TSWuPSTrPvAKdXCbzSe/I/cvXmHZalrWqMEEcJ9rI/VRc0o9mW8x3wDhdFRg6eOW1v
5SkR0oqtLcnYPUXiMjHyt8m+XdZ0U/UCVW8DwrKjhaXA7rUogMHVSktK9lvVNaQJo7CdIAPk25dt
kYxdCL7VAhHppdOuCbk/0/FDqQTYgyiYzZ6jaGk67bco7dhOvbHkOTDed9lR5Sb5hUPRiRTaR302
MC1oIb1HGDDVF/nvMSLMW4BF8v2b84JzlITqLy1w7Dey1DUlss/tY6KwBeA3BXTMI5zhQUPbolya
/fIyqV/falNlqcO06YIq4HHKEXSTZ6sM3XSdyee+TLD3IaIrpzb3O0cbQY3efszvkGjcvCKOFZVg
flw68WuzXfN5Z+N8asyBHKV1dRaUqSVtpV0zOXsdzOiD+/ste+RbH3/th7XViIPDZiDLts7EDPUn
DEPg1Q04qgFggcXqGM/W9+vh7Z44jXiKJdyq7wvnueV81mfv8xinOh2s3fJmKEii4YNi0qbmGf9f
xRV/WVDA8/hdd9SBDyNBd4ZgPT7FkUogRjyy/fT55Lvpr0+v3G22xf/7ZQU2tkYyrtQsA20PEyU/
Q1rxoz/6lLmMaCD+PX787bawylHHK5ye2keQxjI+RkqU/RLOLaVTPuOsRoRnr0POTJIamDSUK+Pk
+zcJxU8reL8dlzM2APjd8jqP6cCLG3wG1JK1WbplSpLkQEHRXmEif7/WkLddTQ8OYDzREotWkQ3E
EybF22WQ5byK/2KS+MwjyhWpp2AZr/jNqNe4HqzUJXchD8VF8UaUhdoc5uG/KXMHgEZZIWhnGm4/
0lvVRr0tEl5eC145x9Q3l4PCpytF2AMgvVV/Iji+oeqVi2xAAORKBFMuiZA+Iit8R0glwyzVoHVY
YwShcKuyIrAFTB9mZCe+1pRcO9bjoC3l+bOgbXM+8+ngHHroJnXIRV2az7kSpkALl5WXWhpL2iyc
MnHUpv7ValdnhyTA+M5WmnAstHBe9RvjWVzkD4a07PlXTDawI59bvCTNOlx7AwWVAwor715FIng3
ZWCP4DeQ6g+BDrrAfiVLTIJzMRMIHRa3wHMsb63tF2ghtWSimo/RJO/tij7dhT+h71wfxdivsO9L
MycUxIxrJ9OzB1/69ORL37UTas+YkODTFSI0t6FClQQ9HVOjyg6eEArZ7ie2i2CLw49QyYcA1GgP
6ie93MHNYbGRBnLWeqrwS1XSJyeFdFRDHRNiGuW0qa/mRktjuweRUkBn6rx+WPnFVFZ/VQHPL8+X
JRwIHP09+RtolvK7tphMxqdZBfD8KAE1YZg5UV9mBWqYQjlKrXliQs1DozeWh7g5u5XFAAcozlPQ
1evPOuyy3X9DvRpq04fBLE4RMTdAODJO7grqnDrkK/Rjs8uT6NIVZRd6HG6IdFMOAxCA3Yr77dCK
ECgj/jEBwqB/vjlqVSkuiBnzRo9q0IgKSdF2HD7rbbeQktC8zaxSBdlpSVdVrPUkAZhzrzELBd9s
mXmY1P1ou4y8oH92Znl3IWuAL7WOh90Yeas3QgzvUeWUYAcF87dEuIr7si2i1g2vMUrTqtdgRY/w
EnyH0DxWe8ZbyxoAvvMYGkHDoJuiCxOHCQvaTAMWedgqAKmqJLF7+FcEJky1Cd91cdMbU7PlIMKO
P/zWoCgJ6D7oWqCTvJs5VwgPD7cOiRE90kbrb66cngFK2o65gGgvMhaqGs3uVtnR489InoE8KNrN
CP31+MokJBBv36iqcCqsWaA46IW6i2ENDEa7rjqBzJqqt3PsPSsxfaZTGkWYoP0R+kaqFeaygy3E
NkjI7iZlqfFiMEruhZwnV/WG7KQpAkYDX2QGfLEzksIhMRPiD7YxfqE3xlkvK82VUYTUfkCrYZFs
YGNAMqsa2Y1DKjvwYr49RJ6vW7+XHtqF03G9WZiPnmQl/p81G9IMKqER21xlE1ZY8IHvoxn1D0ZD
HDQFt+P8B8KwY3pEVyNPVe9p83sf7jIZGT6i03kmVvOkP6PA7DBJE8RMpCoiAiME1qWno3zEYPQU
8uu81SXUngxYMD68mz2BSUMuwpjIlcUTkBeg0u1qNLzSbDfiGsJv3BOfCJEGDGDZj8X3LaAjlmjJ
5Qs7hh9T6bqm9qF2A8tj4BzTu5bmcrykQ1u5vlAZ0F+4KgmmfiXcSz1ZmPTZtCfmrN1DnMRgUxJU
Xni++xSq12u83ShoG7nla63roHy3+eGkLWmJSBbBA78Og9NP9HHZ/pYj6YnKa2T+ZD0QdRnOOjuq
ASseeqw3as62FXXfAXqkwBsX+OAFaizSFEWVXsVHVmk09tk/y7j9q4682OfNrR21k1xWB8YAri+e
l9fKFsbTGsd1SpBOVEk/UUlbaKMDMTwHH7T8dthHJ7ctznV7dIfXJ+Ww6wM1HVCm0IYYGFgge87f
3+4SA0WHwud50AMdCpVntpxDBPCrLk2ZWAxnDqIvffoNJXurBWgejnqgogYC6XivjVy/HATpbtg0
l8VaBHm3y8iLLKAxt3xlVG2VKUbp8rhEDapuYx5ZSqdkpePkySMcAW3iUyQUYWKKystcOLo7+qr2
D6FGU9WjVPi7HeQ6OQN+KX/kAJhcpJJEQ+yof5J3svlafD8w/Q3UdurEIphaeuShRJSh+3bS3hle
1rVDTAPz/4aIiER0GBE6j1OC1t0D5yb4mCP8P+s+21M72AxlGd298Th2ahBBAcYqI3W/dCxfMF8u
/qlQIKIJ8bGHvIpO4GV8MuIse/SNjbwXNLeHXWnH6OmXiNOpmnG456k4bIcyy690zy+f1Sb+sVHi
iKVuZqdkh48kjDPrcN/5J3GdbxEMinh6qNi0cLX/YtPmUE8FrUkqdSfeXrzm4aKOgCinkFIk5Mr0
LGqXZV3Wm9dtKOPkRuJiEC7mZNztJVHXOB2yIUZkUAvWO3MzVPkoWCtliPYBzjAvdPIDeilGkKkD
0hJrJ3H8lUvmXKXPGIh2iGl5QQPgq1/9Ahr+xDfEa0geRpw58+F/ZtHcVbBmYbBqpgKODjJsSLAl
/kuK2xULu13CDJ1M8guqz7quJ7IQeGPz/5Ra9AYT2j8oy04/zDNTaq1yNsuIhjrqQP9Ilk+q1/3E
PTeliVeYlYiWBOe18dnCXIoAox9XELJVKRujAa/E1UH2Q+OoHhH6MSpfyFaZIvAc0mus8MM2RXtJ
2S41/VcjhjsIRU9tE1wFArN5llkIJCgBoEchIRhHVXrGJJru38Z8b4XZJ8Lw1sTcgj3gIZaYzMfP
jvukds33naPWGAXcewtkKlCPQYuhq9UprLRWaaLruco6n54RyDJWsQK9xGblJrOLqls75famjIec
zxKcu9bFt8Q1qY7x5c3+S7ryrNGf+owr8R+isJBNo1a44dPmuGp8x3JWsQpDxg+dPrWBzD+NzJdf
ceOPKFhIwxqz3gMs/Gja7RoTAteJo5I6/4ul0B0d7WwkkBdHB3t6YhzY3sPWqP3htRjhS2Orxz4S
BBfFMBrt+l16muBxVTh1EvxTXU+WeS84xO3/nWGF8RXaVDxN9v8XuITAIMl3ECBk9uq+sy9aEwQT
XpyLX7Nney+XS9Sb3ERlH/CVv1d2w2LlQpwYYgsGKBLk8nznzEdaADfmhLozRyGQsqnuSLftktRb
qQExbfyHpi1C/pFrk9WeN7t+tRYdO+wfEtCDPMbKVsYcf6s92WVy3J23BUUUc0pv1rGEVdtxoY5U
ib+Ub4ebKpU/vUaILiyGwmVApU6zHHyW86F/FkQMqOgOTcaxMxg3lgycz3c0v9w2Fkim6pu7Z4M5
DzxUlHAstuMO7ScO2BW67NTiUoRgYQo8iN/TUIue3q2kdmha0t8/cIz7cgbAfDBvs5v14xoqIS3x
Z9tKWHSH40IURta4T0GwOpDWxkc5/OBlVdsTl8AMljag6K1INiGPylxuBXVyyvTh/KAwuPX28eOG
fV5+i8ewSwfh58KOs8uRvKXtN/xn68UvB9mTRWrYE842UPm2jNd1iuBNcobHrHI5ydUpxMjwrinI
dKSIj55tFPaCMpx7HfXUS3yjyZLzH4182a7mo6+BtihWV8be7e6H8Qp/wrRH4nJpBTDAFfBz0xiF
QG27l9CMqbORqStcgJkXd86/SPNJqfqBgO/9tqTisFmwbWIoOcUc/ETeeA/4U+azrTysTvVxU8pb
SReZBNGGaEcmN3RjzBuKjaB83vLkeYNySKr0By8oArVeEjavSi2rE/fEFwMo0hHIdNanwVZcHVLg
hz1w726pclYmVMJvmKhNn15CXxYca5ZzFjTSmol7lLyTBuca+FhBIltjB1aaflOIRDCAKQ4WokdU
g6jCKY0M2tzp5cftohOKwnGs9iDxvjfOBCi0ipwiOabyBQkzAUWlLzvzkTVBZ8BzA9waVV3j7Tv0
aPgua4N435h+L7n2Bmv1CluJBQ//CaJUf6xt/qlYb+JzVepkls44hSkiz6K9IzNy4PoS583zk8bU
heymdjlI6Dq5jGbBoorU68scDkqk/YsVg3wTmUDPpG2tCI+SqiGngsandbwRW0dLQHIdonTwdlfY
Be83V0WqE4C8OBwpTRTFMvCfQVik/SV0iWD6H3lYvR39GwF3Lnm6eKbdxOdQD1kJmM2kmZdgz72P
EAx/IJ3j1H3wVRD/ucjqr1NSnO0f0FNff0Jza7A41Q11n8H9Ek5FzeVtUDC8zOmOX1JG5ZI6Kyb7
HdJ6x3UyV/CuMDJGXJ2LCSuu+6vsBLWR5yt4IEITN0S7UKmN0snT14NXRa5UeTSR6x2J6hSUK3Sw
JUycOhSDGbUNBOfDAiZJ6eGgUim8dYdlI6Ge365uqyPMXYdZ9ScdMgXhIvaKQu8X9h03doKhWaM3
NL9VlZbV/bqPLWJyhLzMn3JbrAbYvL+mrTQ6gxqNDA+0egPy9NlOYR4qUwX/zTsW6digJSKoNLDt
Ownxj+ieOg0dCsqi1MOmY1gSgBuGZXfogfe9AyWu50zlInmgBmJEewojserRnyJzUbSCamOmkrx9
0+QLiqWMexiTZmjzDpSIBYeviTgUUOZnadZOBMZnRRH/lxiAkTe1xilxxHJQKxwbowyOU7fsoH+i
3OP2SG1E8R7h/eSyP15xi2gXgn7Vd4E33/KS8GjBuRpQXfDEnlWttbttU8Mh6cS+6kBKMJpMsmuH
WkWnnzZGLKYmMuSP6553Wvnxf9/uEohL5idK4u+hV/NzhAKXaoNmHPIXN/BKcsFn0kl7rRsIbKBz
3DKj2+wv9uVRJ56p3aNK+tjMW/D17sOFPiU5B18wI1cxYgJXBf3zSkVLQKswQbGG26nagjtshwAS
x9HXwfFAcweZnQOd1+d+9JkfCHePfKCP0GYiLv+aMxEp5UpKU5s8LI2oAuOI/a7XssoanwsSe/ZA
KRViVeQFJiotBLpbRSjCh8bUNg309cnRRUCDpmIHg2dbQiOelGPX4gLEcNoFRA3HeQYx0vlGAc3w
AEoWnIttXa4lIG7Y48IbLiZj1gPn2bFAkE9tj2DNw/henNqr6/xJXb2tr2DSZ/lrwfVxOmtT73C+
GEYHBopn7zEvoofWvWodFolJ4L7Xtxt2l+l3FYFt7kLgdoYdyw6bIDERbz0uzCfIpewbe8SKIImb
Y5wSl/4GQDNllTu1k54dAl1mfR9E5hBHCOYMtQrB8Jek2mHiIZ10sadnmuQm0vgvgVgZlIuyhdHP
mURmCdT35/17p+5GNWTzJh4bNzf8aQPzt5+l7DLEy6c65F625aMeCkBZGAGV6VdxE/VlmfCyr59Z
RJOOrC3GI4Ml0uaOPP+XYlwQh4oaTtrbaB9W3K0RkgUoL/Q/1CbeeNtSaGJw2hxIH6rvYNntg5DV
F2Bi0ecWCAg2flyG7Uptb8VfSPXXHh6rg0yCQ2n+ol862ZQRkGdW/siEKxJC6H844D2elqwwI+7d
KnuUxEOv4/lXLzi7wrq07K6riVyfmg+20moDZgGCmYqtHet6iQ1/uvQqVlJLkrBApcI+b6o7wY9e
QYdgt0qc47JCeoG/j8elUC/yUh1wgCiH6rdAb550BlpomxrB5yLDzK2T5blv3jKxBSW49xwDKUU+
qtq9+nypz4tAhIrYvhv2yc+42XKwtBI44JpxQjH8mLEklDwihGliYf6B1FnLKF8CbbNZVBvI2WhI
7Jq4Q5fGkKUw7Gtw7gV2sWpoSc5LeO1Cl3MRk1pkLhCE7k3kpViRNxqDH8ECHIz3bvftLMuVB760
FGwezpNcsxtSXRpbOUfefNJrZTiRjPRBb9hWzuA/AaIJMc2vAND+jU2jI7hMQdV2KO//QRKnyfkR
HMslHc1FT3rYMO7s2fmFZbWhuiYjPqyyQtnCncojHe1Q80XqqZTYcwqUZGAFPWewBfJLvavEnG2C
EeU/z7atpQ16jRqBLA5ev+XBqnLLb4BLUWxUEqY0MQAA/opORkSgMQGGUiR25AsvpN21NC61E4ym
Soyq8cyJdrJKZxv8zxCyMUejFDTk2yrp5yWgXKmLhUtaayHMzVqUsHdFgl1iluPq7IP12qCYWfVo
iAEtom8ADns3THbauEFTqfAsCleKE0Tx2XRbCNCYJbTcbAGKBNkMTAQAABTY18+0WB4C66JKLxAf
CRO9jfB5pIe0Kry3enLWj9MH3/HmJjRyZD2ROjF6uC4msJCQ3AAZ9RJlm2q4N5C88NHkXQlVySHi
fELxWgU6U9J7QPQc6yuY9jkFKBOgbOBfsOSJksgarHPsizRZZsNXFpRn+1ylkYKcV23BwgjN7qhR
prmtsx+BFYeFwygdWjQnnpDXvYobnVoeOqtn2F8P8g8OLV+WLqt/X6Vb6VJ28bJN2D5/60oU8uly
rovD5/f7EHhVS0LZ7MHavdU4Xp8KdpXU/s+yczDMNzh1Jj4uYZHH3Ud0tK+Ro/xiZ7k4RrsNxRjm
ohM+k81Ajvs8BXb2D9P8pWFHzOOUXwTMgqpjbzrEUQSa26mWgaMKpZRa6X0OZZjdJNTzXzV1qupU
0MoQEzlLtPjRgLOgMZtJDpZ8sY1Nb0p//OliVsObRSPyBpFIiz3kUVHJmmYT/YGF926TWUfR3wli
yVkBtCaB9F0HqQAWijHyq0Eukq+z41hU+XJbd22bYunr/eDoL7fU+Masl1PgpVI+b4LgcCh/Fdfq
1q56WAJlxZtqVOyCn6vyRK/7v2nOak7R/6D1j46X4tRZtLjrvKShY85YKgoqHvw8gh1K819ge7Ni
3EcR9NQAWwqgoRTqdm4jCQZquFPg9cOjA46nICD9LvFEh6rcJrXMleM+MlQM/+52Z3IlymU+4mcs
7aNsRc8uYojIVh1Pupmhi+vUEj/lqqELIy2M9OApRV0Tgb9LmdtDTQkj2/pk6j51flsLLoAKpcav
qwiKqnG+uWar0FZJ1SkxuuPaxHZaadNlGTYD3FV0QXdmICDRohhDY5ZUuZcUHUGSetaHkx7QThdR
7WEMLq8KaVLeUlYAGCYX9CY2By9eAKQCGyF9guZwLmdl/6HqJoK8jrkmYn4BFXK9Bw2tnJwkZ3tR
zo/kK48YCmRuP1Quc2lCteIV+gyRKSGK/UYfsgcibPzJzw1BsdgUcR0XeNsI78Iryxfo3pH+W4/4
h9aNdlOtuyng6HCoAlXdQKNMVsjQqccIuc5DEeriReaQ8WIe9Cqf/0f8NdYXB4kmS6DOCNefloZ8
BiSy8udUzVtjiROSR+mmQ2LugiwhwEwvad/JZZf9e94vzymybWdV8PgAk21ItgNK+v2J5I407pr2
ualjz+bxgjb779hbeleWWhyHPlHhCzYCzhcylqOBMDt0vVsr/ytFhFMGSz86RSQOc6PG75S7F+0i
QkSURYoHzBjpDOURwx9upTiMDB7T/8+LP5BZhh4dWgwBolI7ZFFbysQQqLZm9vRFDg9A0VVFAV2b
c94FsSgvsYkM/CwsH06X833+/O4prkzKAlB0OfJ/kioI+1TPAdAiy0Yn0MgtvUoAOvN1iwJThSB1
zLpQWV3fPSDLGSkRwVZ7waFG4ZQ8KOVqzR1CDLcuXPJaGmOvddgEdFwBFWPkCbzynos0WKxd0rYG
70thxL2QX0yLwFGiubUfQRmyQ3TC8Nje9f5gFsINPtTvEBqDoDJFbtPYhUkIhhAl/GTLYoc0Jyxt
UfKDEAklDw+nWaqsGLg5inwbU5GUr1ct2smtrsFLXBJkvhxKccyrgIZcZNN0EeBT9Do70Jx1rtCD
hx6Qy6UxGPijbkIJWtE289mJQATzIrvOd6YqWTaAlBafUkIe7Rp8kBah+7pK7HCG/tyAnaufld47
mOMiOY+WD/fri1GnBIK1CCBB4fX/+FJb2VW4AgYW6y5IXxcuKIfgR8gUE8KqLYk/xHvLJbJa5of9
A7MgYDqmECOHNFxVujSn8EosBRmvnavBt9BsnKxUf6vsQC18Sr3MC3B56myPvNZl0VBIe1bZ7CS6
arIuq75B+Aj2xItXKLU4f2McahQsaGj/oUPQ13lTsuTpA3VEAxplksNEzE8gZ66gHUSPiEVd6NM9
/GPewlTIbNqveVNCzriVPNjfaVFs77LFGTeFtnekDpVgFP3+BA3RHvbCENmvNnP9n3ITUZoCQwob
8U5VLCbD2K8RjXxjQxMftzTE5iB/AMXKGsAMAvNc/lS3+88Oc4NnYS9uZ4Uu/fdeGEpPuH2fAXr0
/ViN+d35xriI/uUZYtygkEae/jRMEHi4oFQTG6d0LJxxREVeWmRtCsgQ+eMaPknonVpNpVI5zwg8
EQDVi7/tsN7XQaKcqWcdCJ6JP8S4ubqQWIUf76LtCcDou32Thb2xbnWovNM+0pQt0EX9BG4RvSxy
PPRh81ijqcEKFr8cs1e7gTU5h9eHTePp3Vtv1m/DhLN9GCaiDclYsWYzMihNXedQLs7U472FVDcF
D4N39GAJSXVKuw4/KuXdX1NVGZ6P6BU+wqDReSzAqJAkzImwu3Ou0yL0aHFqljreE5S4t9++Q681
/iDYXr4ItYNcADDCl9xoe+zy5DKmwb8nB8JmD76E72WkmKCd6ZIgHJflUSPQhpG0gNwA0Vmdp4AC
/VAJZZcovJ3WLvyqkVJz5jbzhpoo6c9VkyMY6ykBPqItLQYEujZcyqP8fRG6aztnX0QRBdMqHbeX
jxGA6jNedvsI8fXs9aVjU9GjLLe+BRZ2aVCMtKgt+8SKCOtDiNp3iPuNwmr9JMqZLl44baX+fFKD
lq63bLOENQLqwOS7m1Z9x0SI6hBr2A2xuH2cHZmS6q7TjDPwzi/M2jKAWGQUXsLH6ZWCYBq1Igar
Q4qzftmcR9BXd6vPYrnsNFtsOcpPR9B9Ugd5VruAuz0CUaWbiXk6zqc2YTiwEtxSLQLCdN7QC02p
Oc643JXlKaLVc2+fA51vNGXDaZUeWIk6+eZtv9e+ZsdUsLnIGKQKpJiLD/EBc9yj6BEKhjQynhWS
DocANLjN+nngrkCmlk71lvANHRD10tpG2jmHQoyI+H+MZ59alrGFACHFr5wiSfb5VX14YqdITKxD
Rfc5ihyeXfShd82DH4eoUOA4tGstNeloPVjnaTn37ELhsf81djXE0X2jNVesunPJr99aficZsmP0
jnnEanO+XtnfhBGQonIPXir6BdRWGryENKc5c3YYQ+4sZsORWXzx1J1wwR0DxstU6Qlaw53Wb9qA
AuaPAPXilDYn/t/jwqAfMec277sJbR5VBu2ryFyayguuYrxI1JYzBw+/YpfDf/KGengovFmEUZl8
7vC3rh1NjYwfRXsf9cCwFWHJokLulDKEsltIAIVmmbcDEWUx52jzUyypkPz2B/pJPtUdO2tLCZd9
nETzCy0OkDadSCTkZsWBkCDFb9NKjQsqeSVZxle0IqD5dTimELPh61KpWNjgQQ8+n0mSWM8uR2GG
Uc4zNy9Z7KgqKYtRxstHMwpn4G3bc6PTx/k1G7+MrdsDbVaQANmOjXyHPcfu4uNySp/JxpRJSOyu
I5ovjGF9BaOwNTm9/uUW5Z9LivEsfojRL/C18OVPbzmNawAdw2fWbWZ5x/WAXYxrOVAN2Cbs7hgD
BO/iEK9zfGatSDVmEYtm8jN1DTstFxLQi3OuteGeFDHjAzO0vcJKvADtjrzXWfimqAxSAcF/9lwL
Oz9KgwHnJ16VgzZZ+iH+yuXLgYkxd4eEo+rKw4ADfTFM2BwE9Mks7FmuxWn59pF4geBvDNg/mz4h
zaeJ+629X+W2y93JdCJIkd5TN5gs0mwxMoWGyxkchNBBxkHcpbg6Lfw/0o45P8D/vItBy9dnC2EB
C/AyFsA+/q0UBLhIzg30+3p6nK+hRIw0KXFtFK6MsN4SG2WCLFIee6u04dLc0s1+f60bIUnovkoJ
BnG5+XYTNL9IwuDuJmcXsKxyKMboRKYE9kfax54+LPlOpY0A4jYQCDhdWKz9L5hdCkpqgdhnD1Iy
VgJ3awGuIt28j6sbnKsWJoqI6vF3WN1/m0R3RvTFwLG4TAOR4RUP+15RFGRbKLuM7g7gK0s0B1Rd
RONH5238i84jYJ5X3/4v5uS0o+7IGr2UKXlMgm89igeK2xpcenmu2JsZOoc+VxGxhnFZt2/0t4g2
Qno7c7Yx7JuDI95wijcYkFNxKAv9eLllV21jihJN+Amf2YwYL4BaMp1VWpQNbzQ4j2bDjMVFw0U7
pD+HKKPxu5t9LuqrQbwTmg2aL/KbUiBALIqrMwcd63tkRUQAW2mkwHCVrIukf6sYGkWLhSd4uikZ
03+sedKYR5Ekyxl202k7zPmWBcIzydeI4MYetbMY1B/1frOSNLAG81BO2oxlLvR0t1+epjF17tR5
UT++++SGt0tE5nLBv1kuzjMAammVRSCemreJpoD6lNv+okn7usyhaXu0YOFbdgbi3r+kbsN8D7VY
GytnxyObHLbvr8gCjbfF4u76gfEf9y1FXFN3l5QKzzBHY+9eQng92FWsan/rNMSeySMhpT2iJPNx
AoN5w1bLH/+/6O64TOjJ07DyBtBBllGyZj8AzU8admcK/uiQV+u/6Xpse6pvV4W1aAYUQjPa9NcF
b1AibAGIc3V/am93XpBUd7ccnqPAO96Ohs1bzBUtjFnNdoVtMTFiRRQB2H1nqhN7s4H6D4/LEKSC
kYb3BJh5veuz8ipEx6l7NPL5ZobBwkXkQSqJnmDcuEae9exGytNjZDiEj5GLf70kxmkvAAUJJ168
V1RnPSv/3v0++Kd3fXoEVTP9ibJmeow73ZnSyFF7ADruosVxZcStnTslqkQkq0Zam2QGSlYMRMnW
5S5cjEoOWrKWG6jdDsJSDIplV2VWUJsReoJ5WkPqvFib4xV1v9nKR0fi0n8nCR1LjyhPrHb6dQ2D
PTY4jhv6wGxURepbab1YlXrG52lJ5gIFrbHBRr/NJHOcG/FvPtUZ702jWW4wBKSmQJ+6rygjGSnP
tzbPlAIhFpZ1KkY+xpBeiptxNwItK0URsapUyXHoVI0DGvWED4gkkJsNJoRtuzig/4+NQFPSpx6g
oQJzVUNPrQ5Z/rocsl3uhGIhyWkBlurpDNydOLSKrl/TGf+6YWemVOexT8QlxTc8sQDrUM8cSd1R
WioF2gZb7w/jELRTh2QHW7j3csasmPNX71FrbirFjUBeXIALKwi0M40U3jnHVl2pyz9bYPJCCzme
hZ881V3SzK6NiTUp4JlGkpH81BMZK4GQiIXCZMwUgcwnLtElD3bv3jL4MyZ2XwlcFW2q7sxz7bPy
x7DX6cpyFwXPbqQeIyoQgVlIHawlK7cUzPcxxAUUT1gIjU+2zcc7kK1fkCmF7R6dhukUCl7Oz7cy
EtZGGLIiIE0CjlM1xmYuM1NC7Qhcb4rQOMhUiQOgQc8J30XiqyeUYYwDzz1IiG1WUmzPJgYMTe7R
6Y8eZj0NIqlXse/s1GB/RSSsD2OR7L/qDvJRFS078ira3L/+XgO+PtDGrpVW/Exii3/51oN7kiYf
cW1B2dabQXSk5xZEuFaJ01rixpUVc0Nxlwex4HewuF4/K/0bDDKIongKxP6u2sXTrYmrGzJ2TD7/
mgEWgILhU04Dw+pg6Rot9PTYEq0w52kRMpYAV9u7hYy+SqwrzX+rm1xiCShAgGxXGbFidEA7yKFh
mbA0ZWzuX3/XC3r9vsGazzMgRLXOOGJsYLEW1besEPoFv+yVpK9FFMPW/hNIXi46SbQePEm+x+35
wkgvZYG3gpg9GcBrGbj9IXtcmJ2+HdPXUUV3rx7REeKTnic4gyFlakW1DODMKiXNXMhtIXR8UVWw
yVg+h6GwVtMJcVCgGWCjNNKc8Yako/Z79inb97GkI4wN+NeevcTIEXuY3WVjpJBugeWLtWBRMIYk
SF16rvamv7A/Hy4IRw00pXdX661sbAqwc9VBywr1GfuEpo/4whp8JGNrjun3kJR8sI/Bi+v5XuKV
LTTXFaTv8WzUw3Nn2wFlpwYiGHuHyxwEQBF2O75hr4TveqHnAc8QEohLv+7bk3CkeO/3Bkiyo0MI
SEzj7Q64LPZ6NOIk6VrhAFQOt8+MtDdXzrwiGs6krYaiLoWa9yeNaXv5YWwSTAE49+cirG4YLrd+
lGZ4w+cSVxQkrCzJytSLRepAI7DM+NnrNa79z3rVjaaEWt09CbETd/fWTZV/+3fDhWS3c8ooN6Ex
m8t+7MXHgOS0n+RvaWgzjwfHMx7MyqgtyagO7GGRDCZbaQl0WY3PHW5P1xvXjf7vu2BxDGrxy3O/
9v4JKm3Y/pTBzP42p05+SV9I+jEbWTgdk3l/Ys7VroHxTffE3r/K70FlGBCgGLBJdW48A7OeBIlU
rI3uvLS28+rAcZ3SzRZHAq9UnYHvIlXI8F+/LP+ccOxx/4n9lmtEMK8XR65lrNYMwccxrD9E7LTd
CmnA7tPZP7CbbM+WYbZTGDjoLTGpyRfGQ8CwHahnGyLLip8LH7kmHvQwmSKQUvG6dgp4zg9yjJ5P
PZbwemLJmDsFcKwbeADdfTns4Nybm5jVT9ls67Zq8PefalH+smJqV7h17KhJruZzJjvM0b/725/c
OCkzV/IJN4t0MtZO94lOtRrKyz4Bi/y39i16WDTUDXC71DrUIzHBedqJoKsoW8jcotEoTAtSJy4l
eiwZTgL/M558cxoEc/T6gDeEKmw8ijdIr+T9cmAI3vTW9CoyccnTRxCaELL6xzyBW2E37UPKZtNd
2kka50ay6Xn3gF2Nbly8ycZoV75ebL+5bsiUPHHHpSA01FRGH7mBaoyAXjoMltgFL2Qud4GeoPVq
h8Cz3nTRQ1Wv63zxeOgANbwtM7ZKuM2lh5eUeyzGGjcwhG3q4jleQ32xt3LYatQViOcjBL47CsqO
rQ17P29FOoawMJLMfhdqwjJaxztyqM9/ntXLBXIpu4h7LKpldldjs3lXf6E923laj8HHw4Z0tWL9
KTGBzTSwAGbJDLokrtDj5S3lxSKR57YLMQCKVixsYUYdoWhl56+m1LzMPsS2WPJ1coGFv38vVOO9
HZ7cCBH+PcsE2RPztkb+vctJvErMonx9AIFf+1F6bQ/Gs+1c84Fw8hFBJOFqIhtjXiZejS5L1+GJ
QbB7198f8eSn1EaGc2PABy7yY8PuEaAKl7zZONzj+N90sRzPdAru+SRqJhXk6L3irs4EC7G1xAdP
zgoFlVJFc+e4R4JsWGDR9wq+o7ZI+8cRoo27ipVZifKcXwP5c5L2HPtY8BF8BHpyeX/JHYK+wsyG
jGn3EF7nzANFbu83DYJmxruMOKY4KxM6xyP++vdc97t3KNlnqcHa5mha8dN67gTnXhgE8i+pOEtc
mW0DvoDFq2bdcHGUy3k9S+hfbimAqztTG/U864PjUENkCNNXmm2PEZPMDqqxqN9hbKjhWDroF26W
5NroMi9RbxUhgimrBoeMidFZQRrv0pvqlMN/hVAk/A3ejdDM2g9/7PVEg/FneoT09a6zAF/U4fEG
ONNL2qg43aalZEoEwa8Gx+Yo6JampjnUPCtiNeOIkt52aFnkUw6qNBgRi6Qc+bBdv4rqn2cKIYOn
R0YwAkhMKk6BUv8dshjbr7ogs2hEjqKNrTkCP1lTBdx2HfkZ5mdlExlcAaJyb3TCvTS/iZ3N7lp7
pZP7xEdo2PRgtIziB3AS4IM6qnyV57HZ+AvPnHNm/Fwr1A4tfWD4toIL9nogfFhUrYhtdlfZIxH0
8orgbu4UY6DH69rcFXMiTCXc73wKcIkwhiukanJlpxb1nvLl3tXjUTCunLkOqnikI7VqoRJqlVFv
v/AI4DcareyREhSiv5H2QBRU6PoFbngXHrJNjZv9X88mS7DAja4Fj07/CBZOT450TrwY4rlJd7Se
IDLUs/v40h+3tND6vJeB/5fRpMVjLV2fwqFVZdkTeP6LTcwsIrCidZQQ4HkfKSRGzvo28YiYBMtP
QAHWPC7cV2CHDu6nMAXD+jZe7ASdU2+QMADmCSW+2aNpXpiO418dkatLjAhPcfvk8s8JI27cO/0u
+ZjsX+cDDuTInKUCrgDGSrYUdWOnjv13HldTC/mykR7LxrkRT25tIfmGLDembNMwgU+/BBMd9ao6
IgtyPGP4Hu57jFDnoWOK0ywduEHFn7MPmfIJNortSduNtiMMKmSgxeQ/baxBxh2hzP5tyxZRthkY
2YyRxNTTaR6eY6gyG/Ij5fH7YFDFoglHLWS495bzlVJiKUl3t40YlleWgbiCqi6HL4IOeN7YEY+8
W4p6Il2Vr4ZfdkC72fbDxywkoHJnlGO4OuvrvBbaZT8lF7GTuyzHbQXAMXv7mdkMrAPH+rxgmQcB
TjBcKH9WdogqbDeNcPWONyYiuZ24dvrkJ2nF2ak2zI+qsOmF61+W9jyhd9TBFFT7jk4QOAGDIekR
DlYXjv++evjNJCM3aOTMiTKjGEVQMNNRn2434u2gGyn5RMdym/rk6qabiAeAp30g18zPo5NpNJ4X
tXEo1Fn9knDlUS1fMyh32Axzr0YUh7ZZNQczHaOSIqwT5ccdloUWN9tIZvfeIrsMreb64XSDpLQa
NXWFytMy4Qf+Pi1Y+2vvwc2PUDLjf7Z+DZ5/LZIUCy3oxYtcfOgfhqO8ztDOFM5KfLl7z9RMRa8U
rZysmCrPYSyOMtYDeuLvmCTEPGtKWWirHZlYfLeMOtkXAu/Wr5H6ZjSiw1oU7oRvhJuEf8qV8pJm
/5C6IFTIJ6VnOQbA66tXOvpq/aceZX/rovJbOlDytDuPcKleklg/3FKPrwoUctfTPLubyQnBu2zZ
o5RVFC17ikNJOJvG5xcnvj6ZUojiHYbkkiLR9EUZKQWTgjrJErJZRkxEM6ZoT3EGvm0ZZtizVDeJ
LxBkGBhvHBUsg7UH4g9NKlTrUF6Rlq5L45G2W33tuBGkFpFZZHx+dga9ssO2I1dxEbTAdraikJwW
xnQwvWhmrFXRAU5OUMr0BzNm1MMnKIOE6QqQZfBnwyit/aWqvEV0blgXtrRy1KBpPzJGvO3jQFrO
Yk4owwnZMu3YMBxO6HGYgyP06bHUjD+01q0new+GsLN5xMHE2/qw9GxO16/W4w3jQdP52mgZL4tL
b+P2oXcM7iUSRp9FWTNSwBHRfwRS41EXDmIXRvffWhhh7Glr+HQeh5GEPfS+Jf07Rx9/xtTp3GJO
WAKVh2QNrsvm6zadMkD6XtOHbLYGZonr20GbLGiCDEoj0qJ9U0ki3RqHQh+u6xfVTZ/gTFpfcVkc
jRTLQdoMPisaACnwjMVJTO0L/6Z3tnAuafYPDTV/vYavt7KeMV8lS3vvQccs+DPGi9pMuNMOxxyc
ZGqieyviTH1h5Apgegm1qX90IGWtgyu2zqj7l/zkV5vt8ExZxOzfqL8yV1d8J7HFzMHVgd/Hrgke
KMErmmqQRlD+F1zBhvs96ifssNfJfCO61vu4b7WionWuYnvPiz6CY69imc9FHnX5NzBvVU2zc5vR
UqCGgsPHl50BQ2jEVkqmpl6YAhJUj1STg2ycgOTud3AVKiIEQNQfMORsNZ1XCBf9661O0hjaQBIF
Rf/393PvSkm1UXr1BZFhdjRrQn1Bq4gsX5UN6VZqhgYRgxwRd9rqoiYYOPBygW0nF8FV75Mzrwrj
8YfXmAKHWzy6dMJ/myTibAmd1PcJVAzMfhbKJ8PejYDXVLfBIJvoGtXi+x38mu3U/rGnY9vBbbsO
3qIaPtQ0MtLcgNGR+99ZIViNuondWPGunNZEh5f9eLDYjfX4WKeDZEVfyLjN1Mb5dOO/AX1W4pmS
IlA+d6veeUHkZNvNZopfnz2AEPzdODt/NC56bsnmiliMf7HUiagJcGZuZ2idIGH4VEOMeBb8YjaA
EIXkTrR9C+kwWWXkvfVzdCWv1J7eCRMiPUGbiLjks0vmKe0jn1ytJCTAfQQkZfdDMQsqsJUvyarA
/gVTbZtCpdpF+5Xkv6kKa+IdY3+1S1jFI8PgHhYzlfUhl3aZNG1lkKBzQJ6wM/cifAezwjKNXnHA
gy7i6/lhq6ZJtFhh2JCFcV+6PsM7unMc4TqEj9weTKo/1DlLAxgNPmH5xN5IgpY4mfZfPR7AHxXo
pOXtoGrTQvlOWGLEgzF3Zy4s5VuIPZittd15ieY0HUvbfHG3y1/XTK3r2CkPr6+yDLCf2vLG66Sa
UF++4ox6ZwF63IZRRHUc5UxzQyWlymcAHOWNVgl8VJMywDn0sWn5Ip72u9qFuA2L2D+PwtdfTbPN
v9rYWsekBWlvqjIiBhNt/LeqAbLOVc/OHPQQDUI5BPiff+r2FZGtnwpI5Gnej9sYREP0a2mwypVt
xTF1pdIKmkuX0iD1wBGAdIM/pCoBxAHJKsNdPfMKWKPqP+NrXNKqlFEaCDFCp+zU1xuTtmvG5BK/
3uoiLcAxhuNm3dq+0fxb47TkNKUVtIJ18H0LFWiMj44RBuO7sYkPkaU041ncUZnMh3lgQR2wbQ3x
l9FadYjDBX0eTLq8SAh1ywSpIjIbkLokjFz2LIHKYYP5B9M3c9Kvil5vVHJ7OdVdycPK1lpPuQ9I
E0jz0pPnPjbbRCXrm9U/fw82ikMIVY69MO0GBCYZa340BSsj9VKwDq3K/y3/dUarO9pDg4nNoTRI
abk+PdJLoUylvGeE7AGkQmUPZO0zuFPEw2XX1t5T9bkTlgp+fx6mlz+q8CIs9vVHMs4ekadlgHy/
b9kbF1yLgi555DkAkdw26lZY0mbGJ8PucO7HmwlofFrOUs50/0ylqvLe83veW22b2jT8AIiIfikn
E4wMvTY+Aj98vSjmbAbvUSw/mOkLJA/hpSH67Scqk2yacy17yVg7RZX0haiqxzI4jd1pLEIcDvWZ
Yn/lgxrPqQhDe9F2iXAeSq5G4uAZNvl97Ag8B0BRJUha/VB2N/7s7HoXOLqa2fKUvHR7cbr92ML5
clZxhLFmqxbazNpUXQDznPTvB7H8PsHjGLPVEjBTKusctb7wW9+S96L2OV38CEV21oTUPnplib20
mnfAXTstGisJIRRggAxIo37xfX34VQjYEuUPPR2KI6ZUZopytx0qNKXkOEuvP40Tk3OhHqozdEDx
C08eNlrh0brU4/PdPzDSebqVdh1YBt2aju0zN9Av4C3QCgSF6bToqTuMvaQ0atw78oAYAZBEZepS
LttwUvhxf0/0OO2ZBt29mDI4U/Hv6k+BotS1XQM68K31u9+hLT3vPbT5G9EJdf0oTvkAf5w1diJR
WxhazHCsSfTrT2wPkpVPbImjQRf8/SnanIYV2CrH+EchNYwRbaGLxWJg4Jbi/R1IUC2OP55POHas
bg9dfKFui6udakcjJXXww9bP2fvJ+KKIHuXkfsmaa2xK6S8HdBS/f+qABSO9PflX7nvoElz20jSv
MhSr4obOXUBz9H6CxLBLDpHXPiTikuoftfu2pVWx7CvOuYuKZy58jXIIpoyCbbXVLqn1R4ri3eCi
TMRXHUpbWFoR98cGgXZ7SKp+rGom3PrWVUBlVh9toGUNbdFri5YrzzLBmAHM/dUE9gKCGR7vILMX
P/eJneIYiw8/FjGW2suPHlL0dixBOANMmZLtD53aNA1z1co0t+Jci7HhCxqTQuTrKqylnPd4bAzE
3r1W1k11uhv1ikmi2aThif7zRHAXeJfC7eSKYRjidZO3/UO5sbTuKa5V7rFqqHeSqGGpWPPZCYu0
9su5Iitj9pc17GfTkCkHkuZ3ggHIIef1+twn+1dGB0SpUiuSCjhZBn11f7jf39md7BEzG+znNRlJ
vjnHvtSA1kUirUwWlwbqyCDWSM63PxYgABekGZN5Y8Bz6ooWczsED6tfbgdld/2EvfuL1tKD/Sq1
hQ7kl8H/MVa1ejxFubmP/ZeCgRL4cQd8Gbn7nHchCUPrO9CY0cBnJ6TjhAq7EThlo+T2eLrpFtLo
luTN/FKn3iCDOsG28hkVqP/gsZfZQYwwfqcE5lhLiKjyZRr3BmbTwiwHCXO6noXoxllvU1ATdsYz
70kxyE/cVxO7pmmZgGyFvZJJrIWDm2//1+9SeuxFY+I4Yh4iSYQoDyT9wJeHiqtCp4bgYqB3pBSz
Aj2yGIq4SkvDoffTopk23DYMzANwi7Wjh2kmBL85Yhdj1NenDfGmx+csHlZO5CTBvvVw1BW9kQkT
mlrDhXrdTMrTNUMc/ebftuDQvut/UPtfdUfVBcMY1iNQGVYKotUCQp3WhWQMLjJMOv5HLHG8AQ9X
nmIQG7Kf+nlcbazEVHQ89B3UtY6j6Ba/G1wUQbY8Vg3hisRbIIyPzULdTzaI0am2LiR/N7QwKpQP
cWv5S+fAPI8vnpAIssececp1jiytUANWXXd3s4hbk/LmtehpOaAocrWRFG/7b9S0CVghjzK9Z2Lm
cqmKTLIRPpCstjaCuNA1MfUvH1UX9zYxSm60ZszCWPU56m3Gm7NGI5TR/hu2u2jsy3cdr3zyobmX
SDgSytTvuOLcMRjNksJhfjCE/yFsVDVRVBdU39pVAX5lyhS1ySp7pfU4HGqtGSPAIxkV51KfXvmE
8F52J0xOwC6u02fG/bwR8HKLKtdLWVv/KC/2/tRBHErEKeI6hF+oUYPMi9NTHg+CmEFGPmf4M7Z/
hI7+yX0M7569qAtK7aH1S5Amn4H7dTwdAeoRfTe48GBZ1UE/bxwYp2jZ4MKlO1wEo5mOVT/RsWKO
xNS5UBxTHg+vo9pxg0tc8rAV2sBagvfW7JKjZ1AAM45SsVQ06AmeRxRNsnOOtqKsnR1mg9XoMLwV
exD2ds592elTDTTSKYoGIL9K1EO51L5NH2id4Q7Kehzr4M2NtQCA0KBA80s6UYBdjMWGgdrdPfDv
LYmHY9rzOryLCRY0rnMdasWkxfARU1C/nWZL/z3dSCsXhQp7eXYdRxY3wkuj/EZzKkpyBzCJHku9
vdwUNnWC8m8ACSxLNdXejxZqnxOIslsJTyaCxXYh+PplT9mYl3UnUjS6DlApc7eXLd8e8ijZJPqG
ZAcfQHqjV8ka84sJRH3ze4kj9wWseeJ91GT4oQQ6PHs0GzlKJiC0Exw4YdF0gzfqjbeQ9h5M3llB
nwKqHaI1b47N0KBnf8DQdEDz22cRiVoin3fq+0A6Gha16MSKHKkzhk9qeJfsBEiyNbpchcyu0Mi1
1+gD+kmyNImXrD00PlYsTQZTdUwklzTDCq2+SJahZSOiFwzWtGRxmjwS/VJA00qc/0H0n/oFeimh
WjquWUNZRYBc3aZRWvAGi747O1iNtybLiacKW9AMqnkLPX9Oc4GAT+6AIDfulsck0FRQWwsNop4l
Rf4OgLvcmIAJjOjUyvW7gtBw2NeH2qbTIiv8eTjYgapB/ivWrPEstw+hN18qYSRbzsxUKVueEX0a
Dg38M6wqsP9JTbvD4GeAVZEc1YzCE+LAgNNF4kFVsNYx5NFGEc+rkuNR/oPW5O6oQSlaMHW4WG0e
/8gjaoD2eXibdKs0Ivw8A1mH5+QPXTYqCMsBUHr27okxYqT18GuBDhQ38kGd0eqT6uyHnB3YoQcC
0XlV8bCZSDYjbl0+EJ8mAFXJe54z1Ym/kTu/NVnMhlDuZrKyiMQT1KyKTCLkI9q3rD1ydkczlRQe
fF9w/YQtMXF/5HWKXv1T91qgLIigDVtg5ShemutUjrG5HJvAL/p71b0yDXKa6L3B48qP2oIoYeW0
7K6O6YLKBj4qB/Hhl33E8PV53HXm7s/zsjMcCQ+YzAEByBsphdUNQndWMRJkj2VfH1B7rXbFYChA
1WWD6RpqIT99ASkSZvsz0TT0rVG26WO3QD9s4aaOLpkUa760yvb/d7O4dx+Bjgr2aupYf0jImBZM
B+x8+DLrqvdUhhznA6jHhDVnfXoaTnnPGFeD4LzHlqqqV3gKbYYIyXfJFXD9zKySOSzBMuL9TbvU
agDQXaJ0g+rMq394r8Q5Hz1wZnVIQ9xAYRNd3qWCkX/aOKM4p7eJh6opvJTHmd0eXR+9DoFSkprZ
R73ftcj65m30uccZieZci9NY+8o/jl8t3qmBAJHnnL5N+TnG+ivjAh/JIyhELZ1fdYHKJyC13vCc
U0Yk11LkF2Q5re/zgqrLr4OQ7nXuiAdv7KZxUOwAmBFsvzCWlC/JwHRffjaiKHRsyg+Kq4osOWGB
KAVGC6Ln7LXecdUL28QTS2K4cGWKynuDBS5AOaVXBEld7HovxRB+3fm8hH+EjKRw7+RfWMDlfpDv
+erR5vwum6GKy2eL3QfXmn7UhZ8SKVjYglNp+kWNXKgFGLQWJdYPtMicxjhhx5r1edtF3n1R/FBg
9QZY9cOnUab0TNT5TJ6EbVOPQKocmNaK2sTlNFFpuOg/pGDgd+uuVrt0x9rbOoSP7HpAWjhg9nWy
xv5YPWBaj/VS8zw5Nn6wYok6wscQEJqTCnIuZ4qCRsV7JvP1FVPS2ReNVaB4/Vp6z17hR1k0R2Zj
WVcNt+Vmrql3tD8xwN4NokSpa7SH4tybm8/fahGJ4ANF4e7/uYSJP016qRzsoYGjIPuag28xxmAv
bHCWUOFNomG/5v8dHACYQLJ6xLnT15iXvwXdAUtQp1xTpFkpOmlMUWq9TIjrt4TExgV8CmnN08TU
ZaWRBIKko4RleWSrJ2ylGv4FQHFXfOuyySiwy2wb4b2XQAokcdAGUZxawRM7ona1pqoRqDzed/gg
uJYeqpMzdmwtnt6T200r1cTCyi6ND6mqJSnI3E4RcQ7jcjHvZC9Xormqb4K/uN2BS9UWBsoJljG7
KqXW+gCRR++xfKb5+FT3kW66rgVnNlfqVXaboMzUgAkDyO3mZy89+YqJKsWyAeXv+mnTfaAr6UHk
KsSwimcbVo0nQfw+QvmDzYSs4eGMhEFQjpnHMSaAUpI7z/RAmNBXj/Ynmv+9X044MbJ837yhp8qP
KYfRA60fVOi8S+p8YR8lzsQ2rkB521udwDy4KWveKh4dHl5mguvT/jTwz4xkirVY/A6crGvfOSoo
uCVRS0nWOX1lBEeN0mul89ejHZQC+uBFMtxLf37GiEzLc4+vp6peMPFTAc1PoiqROFoPoDlpseih
rGnYTH3PprgVvYD7xWPwcEq4QnCRS7Iz+w6r9XlthnRvlwqW7jBwjQ4ZGFhIvrxNpBvredS7lhOk
ZNHa935jROI5ZaodvmX1SAPIhd3NevR4MpXLoqYb5hSqGD7EJq8SsdHSm8DVqDa8T6dyRO4mT3iw
nyWL2+Fbb2w1WYkry5u5TLoKTDqK2fxcQFsZaDBfdvSxAjtDhbf7nuM9/5WvllozRFLOJ0VS3850
70vLr6yqYj1OyS+fNPaiG9BlY1YvpYnVdsM+TRJWVcFDt0zzoIlGa/RHg794OThNlobZMo9QnQpe
gmXFDBW739Gn7a7YPnkLe/VBSOf58P/eL7J7znjJ5/We/ntv2yxumlyd7q3Gij5bjqLTChcYafnb
usZv/027ns6sirZsKmE9OTPR72iCSXD28ne0SIRVSUQM+SWZFdNk+ckHXUMPvTefon0sCoZ58ldO
7wFbExdcUUfSGlRR4Npn+wvDYp4Qs33TELluUi/uumTihXWk8+prr5Fb77Jd2TrdDTdt6CUfW6SY
DNbM+cFF7OjRXwdNNK6EGljG0/5otRGZhQB3ccv+MKlRuh3t6qjMn0+zORN8ukCPxYjK4nc098yU
5GeeByMb2w3u6Iopk7rR3YX1uURWCLA/fDl8YQX+S/1Re3Va8dzzFJ0YvEkxchvumMuwkEi5Dk16
cPdJXpVSDllPisvJEjefBe6D
`protect end_protected
