-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
fS0EnneWFqOG3K77LhJsqa1ubzyj76IkeHT3rh5UVj2L5A4e7KcItvPuLDsN71IA
YYQk6UVNOWvmVfH4LQc7IhgfHlyr0fsucPzYhUqeHObDtsHuK0N0I8+ca9TFdeMP
lhG4U/Nx4RRARhTx1EgWHxs+rj+phFlhcJsMh+SgvDXy4Tjd48rHFw==
--pragma protect end_key_block
--pragma protect digest_block
Gfw/BxbVmdGb5BEPb2Xrxjwifjg=
--pragma protect end_digest_block
--pragma protect data_block
E5rWTMBsLsR4coQEi9kjmyMZE/RGyeAHjbQdIIvAaMKp4o7we3oV+55Q2TBazVOc
eXl5an8vgsjjFPh/qOf3GdRQIplFUtsHE5jVIW20AJ4/f/H5lACKjXu47F8lpJsS
eYoQPEuchpPZsgmHCbMnjz8pODlL99QpqlWGO++drdfQioLPwJzWpmJf7XvsC/Bk
YcLgDdl80p1AcQR96kmBToCd5M0xX56RkMwx2qJZC8LfJ0LPxNtFchcMTlRCUBzN
O/cIsw6fBlsYqAvTNjEcrNee0WzqUtieIfJDGikXp3LnY4J2qjyUNX5RQf7y6JTe
GhRQf0STrEXEf/fo/m3clUb3SmE/kbYvSQfxcSex4CG85fcIl7BFqZYO0Jj6lcmi
/BgL/Kn9iAO0NHOl+XrRJs8EpBAy7cZRR6tEFN3OfLuz7lCjSqOKhUM3ppqndap1
XBwppwLfuCbKSHtlLL1Efa9GCOyIzlzRWvj59q7KgEIEztgye/4xzDoe7JqeM7fM
OK0xnfNQZ1UxJTnoxW89Mw3UqdUyAPyG7JCTD8ngjTUu1FZjz42W1u9KHXeBqes6
eJLjX0uWk82zhSlfA1twVnXP+w7fS/sPW03oX8YsJJg5ngNbqaOduewOEniQ1WBC
NvnI02wjED9HnvROObf8U/afXFW8nShaITKIBRF9j+p4E9oI5Fn2Gt8MF6S5tsQ6
VBYdEqMl6BqoPh3al+UIr3OEQIaRXtR6lpZBqq6KBU9G4kvoLf07U8bqc6wt9b5v
wo4+c84ZW7kiZSwMwUmH20lintR5FUzOgILUmbAAWMSsfTpf3WF4RK4gxUdoxNip
kgPY2IqxyrACh/hBoMNzoG4e6/S/f6988xI/tjR9Sg/9IY6Nlv7jsJDMrES033xl
S2d3rFvYsfGNgBRe8KH4zFYfTToVN0/+ix/1oSdaHd4FQJPzmmSpbjtkICGUT3zo
WtVve0pGdM1Lx9ukRP05Ff00djOTGJ2M+921t+ziDihpyLqKo2pc46n6cEbn+FZF
M9kWXyxYvXPaviSeEwoaSP0XfvJcmijNHcD5jvTrmDOGhC5URhAaFGh1GqhQoqbG
wleQOzSgaq0ku6tO4pNsTOlRaiZJXV/0uMCHTe8knTCvmR6kIPJzLwCytlQQB9yD
uEaiOdmkSmLEd/umzGUviwxMlOOxNY9hsUF1b5mMZOp4lGaP3oQpfyJQEmlMiLAM
8RJoBs1QJOSusw24vnQCbfgvI9L/bBaCfPZX6/6926Zfq/PJZ7arB7VMqCrCUc0L
3BamiBAa3XUIxbgCcMVpeooyS93lp2rG01nVYn/BKcAg0MGgPLokJWy9/a3rxuSn
fvhHA0r3NZ5TnA9JRuaDmBv6sqq8RuAIV3uy8qVNWCLQWSnB88SpzAfdsGbAKCQY
CnbgiK49wJKFSLn2W/hDYENNU2FC5mvnDOcBLfB6W10m+lWZgh1EJ3OwWpa5x2zn
u2+AcCFTtS7/WUEE4GKNYyB4COHV6AW3jkMT7JjIJGY0EBhAGICUfw01lvKIGm6G
BT976Ha52Ju1IRHU/frgLU/sWfx1Uj2Lf7qRIAdc77U2im0gmNE3OLYL8k0j3T8B
0Jh3e6tyNyjjo8gRRr62CFGZwxCjOLz/f6nd2V3m78mKAKMg1JbBKTgy9hxYO+Xg
O6lC+BDYapKhnx5Otol2EeTfrCN4H+4YxNmV8nMld2MUIYbEVe1owWkBczfcTgt4
2kHZQ9dAy3N64avTwb3xA6dVyx0LuqGP7Jz86qyWm3HKbyPkh2Bn8YRkhrVHJJ1V
o9ysrhzVPQojYE+DHUZliIZBgEgEBPjrf6SgzGW6YdFH2jJGAyJdN3ciioZuceIr
kVoTv7oRQg3OLewNIYlUqvZ399Wvu7pt1H+hMlW4IYrsj1zKYOyh+Obs1vZFX5/d
42bqxm2GJmFaw8zldJKFw1iDO62kSCJcqQMh5FFrRqmgFaqgLE0LIHZkID7/C+nG
WPJOBMX020Kgxra1/XidEjEV7fh+TTiGgm9j5YzDTGMVKAAcwok4ofhxw0WDwkeK
OVnNzgoIaSoUJ6pCLCAlCzDtNZ+QKTYny6Hn0xrlXpVpgDjFl83HN6lVtd6aKy0e
yriy9TNuKNNzmNVgLvt3xHUwvGGROorSXFun4CArXyuchP2XqZAwRwW49LcfDwmp
/ToA74D5oQlHVJTbRLE469EIkAY474DmPKYq1AG84oYrEETzxH8vQsCbbRahKDUn
aWtDATjSueeL2iAdVxK2ldVun4f0THkSiZ1w6O3aOZIlakkp1sUCS7xFOTIt99yb
nHTJglHpWZejMmLg57CG9c7JaCrxaR5DO5nnirqw87pCWE2jEZLFp9yUw+zPMiH1
Vs2nqBNG30lAn4jQWyHvj+zf8XzYltoOh+btc50/jqGZ9qAS+CeukvybTTYY7Bud
uB9BbFMCg4sNaBp9aX2onn4SpsMDKlTZjyW+PFLXlvMnSWjpzNTCmoK0UVUsaiv0
W6lRZbScpa9e6ri9tXr61xHw7P8FaajO1RR490J2YEeNKm0JeGQ2f5pGuyE+Fpld
YZ0S4DjamySDdr0RzFZSX9t0naG022yk+kg8i+hiRm1eoBkY1IAOigargyvbirfE
a7k/TtMZ60xCpgdMuAF5Iuj1M6qpEWm8JK3FmIaXHI8mFgaGbRxR8fOm2aDxJS7O
ceZDDwHlZeyuwYq/136hR98b+haMpAeXJcs7rmAky8l+x+CXomptTD7phsusWGB4
o79G3+CxEutZUMUSUC8kb/o6bJdMawvl3oXK6UAOeY49d6nLETTLrG/jrhjPRmay
E2axxWCRtaeGXP9k6AwUnGjFxI7LfoBJdbQCUsC3ooWyRSrtykQ4ClqIf3B3YIRL
cNSOcO0VAxFCHgbThaSwvLDHI6g8wxUTHFYapiB1egTT9hCY4+98BHO8mOinm+9x
0U9FF4TPzQo1TeyUKNK9etyZ/q7Tf1zshetUmC+5bb2bzGZ/urX02HaclSEXgSYx
I4QrPGmjtNVpoz5Zx3GYjZ9sSxKVf8MYkVPcYHyI/cl4RPv/ipnanCqMaa511S2c
yS1DE8o2ZPTBAiWfv17SiuxCPnNvl7lSXDl/g8Xv7wL3YxDKmlxSwL3m/epwlGxa
pY5WTE8et9AqUoCUysWyjbFJ3qrH8D8iVjBWUHC1JEGUacPu7b/lfISptaAgzOSY
+oLbqNNstIn7WJdxrg0HnEuaN2kWUiDzDD4W++lEi8sWmw7AC6YDvXniSdaOz2pj
g+v8T1cqcwaW06TfIvjlzmA+IZfia2D47CDXBO75md/dQG9JTuSf3GM6oPCLNn7R
25eBpYuWSC5ZxAmqgy5iFSXxrniw5npzhFMzy3lFux4igNzys9TndV+IZNTP17kl
wgwgIouMWveazrp+rwiwCXwIXmGo4SipYDlTWYse3KQ5iu1erQ9MtCdbfPlH3xl6
WmB8TtLZF+9Bv+ZVUbqVBAasFeLzFcWP5jDzU8VRnIpIkohtuuGjGXCWq8HgI3Wd
dgZsyHWLBIZ08PpSMXVIv7Q+zZImyM0PiN6OKjwtBtjwtW2frYtrdz8nvNZe2PYn
9NlGs7fLmI8ZjWRW170pkrO39jYLdQvO0Df2g4dUF42zgSv+6cfQB8t0CVyPbvYL
w4DtTA7+6UjhC9L8TOIj/bOM0H+Tc27+2uN4x8wyrMXjA7vzRnNJcNVCmfZEKjDA
evFqwXPg1iWVbjXzpkDHX+4UjgMKDUsgvYpopkflytt2Ppzv4j5615YmGbDPHZJq
I4QfUXBny8QjCn9TI5OKFj+V5a1+ukiSOhKk2kOYsUL/x7YEC/F+Hh84QXFO3+Od
rXBXD6/IaAfXa4fzHfcmWl5IlVNam+1G4qLwz5qPBUPmuo4bwnPt6cKvwdxiXMu5
Pe2aYcHRD5qn4+ksx6Zm4qzKffhc4+ehtZFQWy11vydJ6E7ToRtkGb/QKG6pROpP
l006MFyD9H+fQzYQaFpcziylzKvrZDnqqmiXuts7W23q8qdKn+ceLxpZHZUL6dvf
ZKY5puHI7bDkQ39XOSGunMlIVWhwT0c0OOpeqvmkCVB0DIW2QIzaEOiEqO2Tubrj
vtnXLWTm8jUTBiOzKZT3psUezyITmcdL7og/lJcDEiJjNLZAuiGzhUyjxY6raq18
G8HHwM59P2u6S+lAwvbTUMeyFju5d5S4S05zkdXalbNumF/iRDooid37+sskCKi9
47a01vauhLhHK2GNc+ibqBJOgQ366rbGMPYOJ7foT5xtlwYsI63QPQJZ8R3sSdCr
Q5ZYxmIwAJSSUtR4S/G/SlwD323ABoILPUOyIQEwiUn9XDvmekHUFAvllp2W8lN4
QxG5mXPtqcYVHTHX2/K8S3AHxsw6GrRYfHJB/7DIacx0PcWV6sRAIqdzzPNX/kxb
98G6BsEHCu8FoWUm15v3Pp2JrFLlGeKSzh89jiVTyEzmFBhKaDUiVfZ45/4Rb5uZ
ssCKndJPgOiKMrxsLk0ksSs+Mm6BmMO8lPBebOobNcddWYcYxzl+tGGGxQBKKmIg
YnI9xsemZsHoIkr3W2kxsPhWAX9dUS20yft2lRKcqEtFdXbuB0GKRfpvLX7SZZhr
KYvsBdlpQI0YZapBM0T0ahyjS0vYM/9b6RaT9PUdDgArKs7NpJwWkgPimS0lVSjT
n+vJ68xjwqzYQCzaUKp8NwJrfDJs27Vm6BFf1/HzOAC9kva68NkD3zW9QITsHyqm
dR/q+l/KW182cYb7scq6/7rfpDd1d3daSXnG/ovVzALcSMUKsOeABJXZTpajbpwo
Dt5Nnt/Ki+ezLGHOfPn/j0YhtlqXA+qhDfyPPjck+MzCJsuP47Znfz7qqcd5HJWn
jM83QIvTguP5yngWG1OiJZKYK+Q6vTr474YcNddJFQtPeXP0z995JyT7em5Vx6z6
wtj5mIJtB5foFd8t4lgdPjy0JBpqZPqNFLuv/1cx6teTWlNefuvBhlYQR1vGMj7z
+hlwzy09PAPNi6EQpouQN9rmvyjBnx0njHq3CfZKeNa/Au5mxEFa+tnkFlnOgibK
PeIQ+gSrsd077mGYfonVMpsjUNesS+ZIh7D0XbK/K/xYQdprE2j8gM6t8lhQzUoD
zwhMHPStpZfAqH4iH1otLLlbdxw0J3bWnsqIOlNbj7oam09nYeNjlfHUfkG7jlAX
/VzgNEdrEKVImInpHJhxIJtr2qH8d9u38Xyl1/mngeI/f4XDyuiI9N4i8lASZd8g
ENYxhRd4Rw3NCvvQ/6tflFoKpEmFv7fXZnTB6a3hFBfTWAXrCr3mbHSjb8aeN6mH
BerYDlY3BV91V7NJvD1WUb3csvBoDB/6Xkh83tP/X/Dl2NJKlCl3zBz98XNHrg5s
SWaBpgtaOmlldGFhzCF5Sbr1XaAc8v5HtD6mz5mR4Xe3v6bJW8IYAGPjCGr6CZN3
SWjdStfx69FWW3FY4K9XWq2RbI/a/lDKepQ1a1UfUzjclwodXQfoTMMMMtLbqt1z
RqEdrmSot2HKIKcIazmVqQI2aDFnO/uAwXR45WTPqArBKF38tQOmXdF8X6XRtFa2
S8uDQw5LAiAfr05TFkw+kKlB5VVBGfqQrzLWIgyoRRSGjHSxzPNtvRvuED2wjrUK
PsAgpCEM2c6fUqWt53dTIiRAoW/NpD9D+FsYI5PMBId1GQg+kMH+4zy1Tbzss9XY
i69jxBaBsU4zKfbd3JqAuYYV6fRqW3tVnA8HcUMshHOejeAGhHHoBkr0eUS8iiRh
7vWIrnHikJugfIq2MBNmxiJH0ll7SLafG2VDTSi31crIcCjZCAMEyHS0kBWtuOZ7
gtklPYG+GJ/x90m+nmmePK4q+KZUaYXk23ExljuU3QcZm2o9PbKsIn7yoCSY56wd
ezwxP1JpOFmAfzrkld35Xy25t8eStvAC3ZjH+tnf/ub3uRpwWLo4ZILoUoz8j1v4
4RxrTaTQJwXugtQno3oIMiU4degU24elaHrWR1dsDehPOuye7k+mwJ/13b+1VbS7
/yQT+FntKBZIJ6YIboKXMCcevxdmOnM9IjR7lKrOBA1cqkkHTerJY0TRoft8zTq+
bcyg5Zjq1Sk8I9E88j/oki+zHBk/TPOAx5Aw1arNRHor7P3jqjU3oowqDdi+Gugx
Rh+bz+4Xx5oo44DZJBmmvjGEVJ8lNzNILdwH1Z0XzlsHeSq7/VZ7WLxx3Z4CsR/8
uNC8eXl/Apub9RrBD/olpJNF4HebCXXKCuUG66Wb0pHrs9ciiPblEb3M4qiXXtt3
EAKa7yD3AF1BFxQ8uCU8wKLIA8fwpxMgdMuYHuocXZtEvmaacms5FTbTn/9nfnm7
WOzhoa/E/i1l1Hd3/NHYKVfMgFMF3dAVZEeuVdSqHO+qXV4nb1THXIKTixnVbxNA
flDppIm9iJ4IBvo9suaWopTGMQzbVp8geOYYrwH6ie5f9dtls+k1kYidKZ2XiSEE
my/QKYLn83NuKPc6Zh6NMZGt7AW24PEQp4W1kTmbiU3hIP89b50kz9fnyvbgSrrA
CyA/umxPWstGkuAteVW7odhmStE/js+grdS2GVA/wuSVvU7s60vpklf4FsNoN6R4
IW4C1WQF5MhmuJL0diWc2ZRUrXPMkJZRdt84Tzc3HgCg9l+TmipS/rRC9GRfRtHh
zagUOl8NtE5wE8kbbUvPRGivNq29MSiu9z8JE12gHe7xjx58HL2mGxnQaZKlmjhh
NRaCe6zqD1s4im7mj2VfpwKSAK/uTiIruumcc0sTq3XgL7CGKqkUiqZge2quthWi
WhfqZqnmKweGKc2BqhEM+VKrQJaA7+dCTDPQm3+//+FpmvRNyMv174q+d74EXuIA
kIePZyvKVBMJHYl4lSZEJuNTHcp54608bhNiBj3GTv8TXZmPZ733qVXxKYcIjcPk
tgBY54sDWVrgCu+siebm71hebqXpELC18eg0hcJGD5w15XpXrQpx06kKNnZ99yJd
ayzRl2fZ4dK7wrYZsarUooZHULLiIwDfAs1m7uZf3kUpgTEDBJkAEpDl8affPizC
fAgkE6gPMm19Vuz8QKj8ym4tGaDpXMxTMxl0vsaYTT5P0jpDLuPt1OzYVh/26a4o
2gMjxGCkXRBCoWM4RRlVvug/MYcnfWHK34xCZ5UV9qsy6+zy/Je3CcVvHeBgDk0V
CGAyQHRxKSgW0lq9pnzUbu28F1nm4dlUnQpQnsewm25BxLZLFdeSA0QNjKsKAGP9
PPYbGZgp8cBG3QjDr/WkVhmQv0k7JjrvlRmI6bR4jbX1MZdwE4EKWqoQc7Y+JVHl
9QgwS2+SD9g73Gtea3dAaGuDXB7778fTbuNZJLhsHOvhIf5IAh6qpikp51MJAGCX
XXAR/XMjV8Z8Cvd3mWznA1rz6v1gxF3k0PRW/DWaUZSZ0xEqmK0E4gyDmef0K6Lp
yIPPFYtGykLIQ8YfU3BTJ1QWFuQn2mGI6Q48hR3pEpGTMo3gfh2S9H0D5daABlRx
PxEvpzzxcvXqGGi8G2doyV5HQ1fIYFaHNsA7PKcE4N8jHUB5SJIOy54LIdoMMEpP
HUjWjwXRz41l2ZIslkikn8xuYcDMAPL95y5fEX72HHJtaxKGt0iSwNaU+ZAUWhw1
scCtch4QKgVp13AW5J2AhZRWNE7Cf8zBQTlAPlwmdXj3c9SgWiGsKA0fo4g73QgL
xAFXvFO1Oy2cxViROCJZmCd/aW7Z4yXi7kWFXPiVka1UT1r8cESKvgThPDjbeEmu
mGuwgp+Y/yxfZOCuWIL0DJmsM+gSuzm2lT8+WUGKZNbbkXdLM8GoNf3wAk4Goi8P
8RLD+hvdyrFzZcueBbPjMc7Nu/3omrThnQKIiIoRtNFH52PJ8VM6Pq6xlqiqrUI/
sRxe2IfnAaPMJfwDmJC/KYdDiSYn8KUFgoBGilBO1GBwy6VfHaKJuzyltOv4Da9K
HoIRD+EFtQqmyzj6aCCJnD7fyPE7KWLvLcULSPg/42sjKeZuXCDgkCaLr/YU4GA/
uqpQBsjnQKmy50QkifRDExyJuTDx1CVg3wc8r5aq3aqR2Kl0THvXvWdpakUz6yC6
FbtowcQIS16uP0anSL+ge6mH3p1tfElEgxikFj97RoYqHvxWj9tPOPHmRiFRG+xa
ZBOrHkKHpr7Xg1H5L4LEFF+jcxbMObaFIsl49NKE0CAuGkX8YItydvlzA8SQwX9A
0GtFRgOZefrnQH3tVXAPdRQ0+MLBvaXAy8gxS0mlqwkCySXm0Y3PgAFJfxRGTq4K
6oVUzE5Dj9DBvA6aSSyo38UIg4HZi0xvnNZisBnJHnFy6gJljk4nuh89pK/u6x9x
nLrYILmSj7OvSO/szD7OGs1OE2LA8FhSuEn6eSrChyabMI0en3pyN+v8By/HeQ7t
suJySYONOJmpXQ5jPJiCyLTmqzOMQvXgsfGgxZ6Zl+45a3FLuWmnln52rUjg7lrE
63w3m1dJvm/TyX/1PKZ6bqjj6QNoBSC+d4AAvxfDw590i99lwD6/Juoz9qtHf93H
eyQycITe3jbV6Kb76eBl3vJCVyNEZYOEV3qtgiazO5scli75+PQUt0TFkzBhXloZ
lkK8oTRy1XUltEgcNQa6XBBSqmSfSD7oRZPIrv+Nbpvah6JUJLu/O2p5cMebf6ID
jFOggJQ5jI3aKC8QpY+feAWibZoEz+byn+hnsuTr2t++Vdxrr5Mosgt8Hp9ZT0mA
RERQWWfwORfUeWmuSks69xY5RDpiz4R4hrhJDkozAlYyu+4H2ehnHHUOwxF1j8ED
Pf2TOWz/+ZaReyBj0Vd9hsYBD7qf23kDRMAVW2T+T9oYnPbc4t7ul5RUcihf94Xm
nYxKHk4ohe6VprswipYBRB4uY8QsugnJZvTC1TJ9w0nGqcS45twYGPFQeAQJPjav
xDUZlYCOQCjIYymauJVfY9JLsZPf/dVAlz5JOUP5EUeI2I6fZexDIWn/Pf56lyqK
zmqdfHPmlfenNWTS0Rfkpysq082PyV0Gfboyjt7gmw5VjBGuBmK+bdA3sj7YaphM
hOsEmsJZcHTbZRgExY+Fdtkxyr0CfAQZhkxbauULyyYW/izFSt46PGvkDM+YCdp9
aHxxFEHfxddVsPiMBExY6BaboITaIDu/C1OACGos5AUS6awJFXxVylu5SDDT6t3K
Aq3helP8kcgneMLXnhv9Q2VyF7Sa5z5AnPdlBoSM+vEDPM8EROpdkgv8X9cED/VG
ZT2VwygtT7xzwxUrOMxEeAtqd+UfZPwEd9xzCilJj2/q5IONZCLsUL8QdemCrQ5/
Wkf1zEKrzS2Ir3jZbnvS+l0wtPUygjj9/nh7ceOSidcqYRNLB7DvFh4zHXBx1drs
GCa+FupToUX/NSjS2a00PXXvbbA1BsZWIFVHRJAFWqbQEt7YbzlclDfHgZTj36oi
KLB/OiqEFd2HITZEkI3SxEEOS8gy4nmK2s3wT7+9tl0hCH4E5X/T2xuyzImL99+E
AaHlKaN4AKn3DqJ2ALTD4Xwi7NTC45AQPMRf47VRLUvy72JA8fc85jK4+k8ELeFP
+irg90w5Qtzmx+FhOH/xZdDGT11JD2TXtgHVvxZmLe71UYpIwz6a4BzDBV8g/Hd4
Bhv0L0kLpAob9ziSnqtl63SwwUps/wXm/BAkgekPyDQi71EBboxz1bG+O5Y0xBhr
+bgOlMYvfoJD1qTuSz3ZYyaO1zDCRxwepUYW0YNgA2tw1r+Vl/xfHzQaatboaHse
K8ZtngnooeoUCf7FJbYExOsJOrzs6tXueeyC9dHt7TSN2ST5WlsevVGaqSghwfiO
270Cf3pwLoOAFqBjJ6WJ7LzFvSP5lA0CkvLWeFXIOj2g6ZC7q4IYwbbOZZyadJXb
Wfeou709lmDHQCqqUxpZ1DuBiaBTwmzs5AawVvPCKQsDJuiVXdzwd6HhRq69mOiU
FUVVvnfz7RAUOHep+gUETPNW9ojugrvofx/8EeFYCEVJwxKatVQr2RrnZA2h6m4l
rCEaNmc31DeO8dSUIfUr/1k7DYrgpWDVlV+r/nCTNSVrrMR0umFBmawzhClN1177
G4sAUgGeVv6Ay47b36YvD28vh9sUsD2GNA3Rh6bu2+OqsYXJgcTiXnToid75V1tQ
6xwKqFwvmUXsENFcnY+JOJMl0NDykOfAZb++w91Y+fV57Zxb/0lKSx8aY+MCbjvc
Kin0PED7QULiuSGsYm9LfOFqfSFYY/PygeMH5MJpmThqdrYOEBEQ2JSvYY1wkHCO
KqEK3Eo206Y3JOdNhvkGaFL8SZKz6BjkPmJR1//eAAiGhNLJfgrrWLPITfKcDn6H
CsnSIfTroOBbr+lqrvYbGgqGwHXBCzCVNNLh/R8SFioMaq2qLgC82LOYSUOfNOEx
ThBRpJVpofZMmyxIiE0w8sXbKE0XxCPBh8NelrqDGUer94e+M6CfD75Pc/JhGeG0
B1QRkJspZwF5casrraj6NRksPPFY6u7wTSlfbz4d9rWAkuTa6BihAGS1UNdaGH9w
gKAJo05WRh3gOG6Kt8hREj2DewXtyNphIFY+bWitiN5Ao2M5Z0LIJlrP0cmH+Swx
alMfbrHnBaqkx6qi1F/UAVmSbGT6pjBivAihLhukp7pg3UAlYqwKSGRvxOdX0o+2
ZRxgxuBn3P5KdNjiTY+bKqAAGwpMp2NfVyAYXgcrCZ1vbWyYa3dxt+WdjesoogzD
CwaXd0DPmzDWOf3jTjlynFTyWp3GY6OgTAX9ThafUC7DXrtUdrw1NRcpFnv35np8
KhjU/FohKmeWmIytcGUQQO/bFeg1D9M+sTb7RNJNwtHGOik3mn1TAiZ5HrAHIeqI
LKap6CcHphiYcUNoaRYDkBmgL7Q6Owe6Dis9Vm1VAG8fyyTxFiRga6++09DC81HS
pxkJeFJ0kEn7jTDFKOJ74FvYH7LsNU+jP9G1B/iUWKkux62X43+TbiGibsC5UBpp
6xt+jRwva8U3H4jF5EXH1SrcqEDQ5HPiM878tN69fJL5lse2lLYEjIMT2bGmC87U
50DqDuP9AYxpG/PU9JWc/TCt4hSwKpnAuGWiTKOFhjMKp/5s2eEpzOkOOAmOn3+X
LBDrqdIWA2H6AjUdL247yxjDkSZCwxjsX+ks4nId6a8moH987Hg9yh65qZF1hzF7
vS8veW1LGUQii5DCFadQI7YAEAsFfns66la8ccsm01e0yycp+NKWcv98MCkD4qXo
MaFePrOtGVb4dOpjX5k4sRn80tJQSj913lDfj8paDpmFcEeqqo6a467oZmeStLm7
8KA/Ej1uSWmPjZP0viVC2Sqbvx3HIIl0DUc5fMK/EkeKaywDiBtv7fitLLntHhRW
5DWLwxLLsu1zfyVlhuQPZttALVh5yXqW7+tTqqkf5mbZ+XIcxg/wgWRoZRBG9rU7
h15fE9+y8J2fN7Q9QOBf0smjv1vn9KNPpLPUqJQEkefgXaxs8ac/ThHi0QsXDLy2
pTdQBioXlSf0Sae9kmgtJllQfHNMYNnJ56gTg3mEKJiMP5Xuv1dg5IIyo3+VeTzl
mNe0ytxWLVsW2GzeDsgzWhHcG6CNS4j+e4ghc24+4nqVbgtaCq+ECsbDQigMJ9J1
PGrsx7tkKmXnXIusPTcG9DvXcdmQyeyWbz5sLEUxMkIg3Xvug2ZyY1iL+m2bQ8di
BDKG3WHXDINnzSrE5GUWR7MRKkAKI94/mdZWJaA9mM2xnmnhQLEJa9AB0WLbvg0F
17IxVAukWWj6aCUeHXmyhYDtxZb0Zkq3k0fUMM1Ii5ixBiIBMuicAHMSbyWvseXW
RQb9fzClbAHCwRzVKwtjMmdOVmg4CuFUKH3js+32Wy4PKXbM7UryLcL/yLqigv34
zlIetRm3uwC4Ojn8Pvkno7Tbkz31+z9Sv9JxBjKC7VoCK80F61ugaTzlE1lPlgQ1
mpAX9HeLpQa81YrWIaWc3lx6UgYr0QzkVMXC21us5AEElr0IX4t1XXQz1RyvnyLe
1qvo44tvTBCgCiFbUzOF+JHbjQUIjf0fuimFly5+2ZkgNeKai/SEKLlDLCv48Spm
/LI5L1ZN7jyU2u1vTU+IEfzX8sekXPJWEbNUgtdvQy28Js2qlYoKqMEyPCgIwrvO
1ZZ1vnNiQz0ggO2EKcK1ZrXPn53dgZZ/kh5E4znIarFHoIznYVUazmvKPhr8DmtZ
oVHD3wn3bdWrnUzNLQWSugOV8p4/BRc81lcn2yMms4h0aG0n8Wt//fNFRYNAz1jP
uHKBcLlW83LpvCW3Bn2LLM7+SuvDYINrDWE7mayusp2nI4ew0RdLkLsnlgtLHRLt
cPTM3IRucRIuj148X1UYnZgGsPW5W4lHZdtAVxPSyXAjGka/bu/h64ZUWLiuI9np
QyD8dn9J6J7oCLVQLf2wpr2wNpZ2/ImQq0cRy9b5vBwYjDrriZ/PXzHFfQACZ77Y
TBJ4fIwNwvS/V6dAMC40UBoVvDFTJvCaz03DhHJe/3Fsqi5cEApXE1gvtRmLdey6
iMrJvauYoJXGDxxkOTq2vRLVHxiUCi3OOMtpQodhKWlckZq+vg3Q14eZvsKeSiao
hhrOZU6ZzpeU22mRKzpIJGm9nYgyQw3NCTpzf5wmxfR8eKX0reL4Hlq2+Rslak5b
NY5UzylFSWWT74PbRzBtggkDJKjk3cR7lKjLgOhXLRwZU/7NKpF/6+wQ6gp4vHOD
Khcd8hAR++FxIiZHuYZKMKY3OAEUXKf1RewgbclnVMm7i/aJQBdZgO3D5nD33KcQ
ucMvTfIiox8sY/gElole0PMzysG6anShIqBOh7xegRzOCGyw2Gi5IAfOBUYdhIMB
w3Xg/b3K/pv+VbrkFHpWplliSQaUpqppifpuEyRDzAKQ+f28Wz6yom9spDef9Cou
8IykE7U4Z69e7Gncdj2WWOJxrLYCAyJP+gIb30Vvnsa6ACx5zdvcYCRn3hkvXzrF
Wfl5NY65zS6fd6ZHdxF0u3MvzonMs92DAX+CfIqPQX3jMJknDR5neNH1JtBCGglQ
wnY8WKosCVXGg2I23KUgM0EQ/WATZRvwppUTxKPiC7gxVb0WDWv6+iGGCCcf9xUB
aRLvBLQlgqeCYu9ykeUgDyoJxonxjRzod0envpENwjHECHjPWtOx1FcIUeS0r1CO
tdod5EJicWg9/D7VRYkqQKuihpz4zn03QxiGL1XFRPuKSxZsuHnVnF7OmL+FU7Sg
Hcdnp+FZ1EpzCnImnZCCge4goTGaXoTMyvXgUAs0OA9slghNYQOj7AwyyulwFJsl
tgkqhXkX1ZgsAR+tTjkCvnadiheiEiBr9QM8KSwfTif9YoAbj0rvkykkZCJIbTFb
jnqwnzILmtd3f0iM1uJ2ZrZ4mlsiKwaDHZUU7fl7XkAQLBSB62sw/joEYj9pFH4a
U5S/RwPNS2at+b4f+UJuKl0yOvt/oK4WFbAC8y/UUsVY3tiVTA1q1q8ebzcyib5/
lLVoIxYlK+tTv9Pi/AalhQt68mYDYqZS/AGBgAp0oteSIqE0ZS+6+6uPkca2xc+I
vAlgTYoUMvq85CshcE0sXSndVGsvZrVxLvf40CZP11CqwmuprFqnm/vhWzHi3ej3
qNcoQsarFR5JAXVGNt/5GMoGz0QTKX42/UMibWw4VLOnGsFImqhQUwrE+qBxLmTu
sst+MRo0RX9WAAK/79YbMInMsp30W+HCTsKIYGSHyKpCBMKnkhBFIo50z6T+403I
L3wxBQpFlIuFYWhDlkMwyml1srieGJhBsn6EraAOaf2CQ5pMyqIn2uCT5Ak4CDPi
H89LFv8EYbmmeJGysOyDQOB0ziXL/AMmHQTqLT0RuMF6s0XDqMtFq1NIy7DNMduF
z4taXQWZ3/p8a8ZHnuKn3nlVeXIRLphw7+JdLpv9k4n8XpFU8CikPCZvzfaKGlr/
Fbj41YVPEUO6gljPOx57wEMM74C7L0xn1SbKtdTVtCDOWjrUSDJG26pJeL04J4Ki
pXOgECcTIEkuiW2KpZEM57V06sUnaPShEK/Aol0ac5pguMtEXzjHoRNyETujkGiL
3gcmjDySZlAYbwp521AOeB+LsANXXic9qHQdeYEJ+6WRl/59zWFAS463Rwzm4FPj
BLO8gqfOtQJFSl8+sNcIKNPOro4NWQsGWdSamqZ7VJi7a5LT9vk0aVLlXY+cdyUl
wSY/KompNlWyYGK0Qozaq7IqIBDIjkaGJvoEhYEueAjM5dJWEkyDbqdk4t5zfGY6
/+J63ppkGdEs6oulKoe/Es0Pt9QgeeTSKGGASTweYUT2Xx2FJAdzIO+s5UM9AYCs
NERIvkT7ttBk93DJMw8E87ML0e10cAysWilz1fRmL2LiVihH1Rn4vFJn2UO2IFr9
dO0xeea02LrQ3Z7YN0tLohd9jEly86I/LvEWZ6fJEcAM+UlTUWIiUxnR+6pAmAC3
K3U/WHu1vJHx+FFzxXxdmNWqxKTJMdTW5N17YHvW5f4AQ8NtRys0Pnt9NhsFdUud
hjb4ndVI3xul5Sd4HKEX0gxs4tQw+KvOsrx0m1BuW8pxMrJOlf7Ct//FhqeUB8yd
ZHDUNWDSUDkySGVA8I2Bq/VPrH/SPoZLovRbR3480w7O4OtSzuyggYn/GXLHuCGS
K/vy/fDfBd3uSsrxnLrzSW6JZq3tFYz8vpry3LKaqaZIUgvhJTnesMo1oPf9Y+vs
lM2TO/Fhr2WOtWWY/v8lInVfAmiOWCM2PIW5wt9wbMnd4wrVesAFeUYg2rPGo8Vj
JLep0jYVKK/VdaY238Ut2R3ytIFiUMUACkqDLSPH5T/G6o0YNpGTLRShJHq7mbx7
6KiAixOd/2WXyWFx9c/qKpDyFZuSsqKDCXPL44wec5+Xozg5tRusSuDuRm+cHvA4
g710oL0ger9YiBsvlsB489x2oECR9riffENRuTzWbMyuTSKv+p8QWJ5Tie/f0DEK
1I2t35XL60b/4mW1jemD0gMvPtz0W77CEeGUuCltFiRpmAf5K1/AVfm5bweHKe2j
JM1qE+qALPWLxOO6YSHxh5GhS1gyVXK6oQM4atok4I4QaP9UoMt+82tipipXz7XB
XIJBqYc/NsOK0reexd/QJqg7O2pXPHboxyrokoWyRgiT3cd1uMMyU3qLfndaA87k
aWbOYcXLslbITchfluHZ9cfnGf3dX+1hzo7koybjAIxLDGaCDx9xxr5KKOQKiry6
4vOaMMp9UoWWrrOaJKspgxtcgB+O4uBpKkGS6Yd0gl8DmbXlufuFN74wcmp7b6kA
Br6nUpTry6BTQ3aDsJsqlO7nNBKqAa3Gk3OZux/rQINjKyKUiqpcaAjw/1blkl0z
R260q0VYdSSHlDgYugEKksMe4iRXciEdFDwls8lAWjIqkMZeoZPgLvU8S87zx6yU
RyYIbnni8+Q3wpD40a3lG0oHgR1yJEHbv8zlY0dOtPmkmPDXUvOioVDtGOzX6RQD
H9UxoQQoIvG6S9e1y0JlPrXHfPi/HoV4zAOZMGDLUp+eNwQc0mBhLyHhayyCKkY8
FgmnJqdxlgiwfZE0sCKVhH60MIh3gD4SHJbXVb99F0i/YOmdZFT1P32UNOOYgfR+
rc7TpuR4Mm0ddUKSOo0aNyRt1YuaIWVm2Oz1mJd4aU+Fv/LnSzk4U2gbMNmVJDwf
k5Sd11di12nYCH7DtQQH8ywt5fFhnunviqk+n6FKwH9PHI71JC+kvAMuatkSna7b
xI0HPm/m06pMZrlReRdJEMjtsTd5qzmE/TW/ONVWEtHpaJDZ3wt9ftxtn1T/cT+5
KjEFcpivLJtOPXMkUHEEm7NPj86bBBPmE+pRKWMWSCO4b85LXYpm7etBv/QVKrkj
OV19VR15NDUCb1JneTS8EUSuvA6CGNN39UvD3Se+PRsoiWGT5jkezdHUw7vuWVLt
FKvXZX3WY0M2GBlZ9oueRLGv5XDZd14cGPddLcGAI5q7riN0DcMulgeG6Cd6BXJf
sbVva+kgp9ozfOb9bNISUku/kt9IoaIVl4jOcqZyDuSsfQdcNWwXupfTr7TBrNKB
zw07NfhdhYRleWC5ARelKfjpuTfpbEDJRrMnansPHpKStZOm78JxZX0oXtY4oyVB
yBEKTc6BFlF0V6iH/4huWZoobH/kMkEalmsbRfYUo6yKjD/1DoCNrSIy4LiinxPd
Mvh3h4T5SIy6va4g5CepV0Kcfcl6Mz7n0L2MFn+G4VBvk7p8kZGm/TqHly1RbFkF
8IgclHPL6GY+JtASLI+D7Xcie4M76duiaFTVnlJDxlank8qPqBfkXR29zZJHJP/Y
AYZCKnI81536JDaqOWyqqbfOKmJdGeIH82dfeavR5uIr8l0ojKjVHb1daVKHFjTs
4s7/SXKmzzjWERnpNmVTjnexJF8c1/QV8blWcKuv91fiC5BXXuORzepRsXkmniW3
k5LxA2cVCjS61jvVR5/gUuqf0T5CRbvA5qtNI4FQCQUug4Ti4mrlwZDEJkbV+JRP
+x2BIWWswGzJ07jLDWFmnrw06huwRmQRMS6oe6LRsCUdZzdz9FkiVKiA7oB+uwuZ
h28NvCRF4ELK48P+ZmjaTpPxbncvwQsRr+5gCAynTZBqX7y10Ax0qM2gDPTk+VDc
+IehasJDSP8GG4pR4t+op7WxZyTwTk+t4ZVJpVjMsqrDk3mySnHI1fN2lFeW7KTV
fMIKNXmAe4cbEexcve5bcIfVQ+zmJ00wq6n7iy+pfuYzeWgkMNjkCAWy2zMcXZum
VjJFQcOelBOAE2DwgqwBEMmZKiiRZyvdv5rSjHHknbKo0FH8xWvcV6oSMO5vhRi7
V5FTb8dS8Dny4MVRjYN7HLh4ExUKKqaewa94UOAFF/PRvdBt0IMOY9WdEQL28WMY
FEpC/a3DhxQ7MJq9JZbPnVhc5QpNLADF0tR09dWVpKvOdzQGCRF/1r1vbAh8+cCK
1U/UkNs8oP11DUhz5GoLBv8URkYQksmYL2edaEgeYgies93Vvh0Wbr8LVkyAANQx
1UyMP7I5ULfn+ecdgELgIyrLNGiZU2xFk/gqK3x5glx2pBv5p0O9kQG4E7dcCUPF
Q4jTX1KQg8VYhRdzN4Ho4YoiB/r2cjfOFi2TUSBd7fDN8aWiosBoY15xSpkJl7w9
WQptTHHZW68StRXe4ET+8DIRRZChbmfyOiliYmpc6qGMlyjSAS8Xfy/TUXuFPdTs
DmFiPm9729odOD1PxPp4aqmJCjxPnRGKULEZeS2H8hLUAY0DjpToEGp2QpWB4lYF
3kKK79arR+EqmE+uI/xZ4sl3vI2zzBJspxtc8qd8xX5oyGQ16BBkx2AddDX0obBf
af/S3lV+xUFT1D6idUqFhvVy6tH2deI2xwoOwWjNOzz/M/KsL/u3+6Ozqd75feKb
13zdXNJAJzvHxI6mDCD6wCPskTPSlhcA9DOu0acL53GJTe39PTSJEeEL/t0AvZri
RyVyyizzQGEsRdu9Bt0k1RDRppfyhIwc4WNtjw08xlqwVmA00ZofoNtehGYjPuek
R5Cwu3/PsnzkKRTZUCyFE+by/7SAwfQZcuxKQzLvtRnORl8L/q64ZVYkLmGVUL6+
fVtgIch7/Jfh0PvSBd/hobSRKrHSTVZcfyIEk428xM4qtrbclCnYkEuGUe8Obju8
SmXtSCWHCM9CV33hd/KAQl94nscTGv6tqjRog5aQLJ69oQzysc4Cb5tJBGaUrxAd
ENUSDzXw0M92KfswaEiL6QFX9h8RyPxpje3N8Maxa3HitCyT1PVRX0vnGnFFPSon
GxlPJlet3WQlyig+uRG/a9Z25qh8Lrhmp2JMK5kHrUTxAh7Qf/XUCnJYUxhK0iKa
iqfDF7EYXH7/BQFIvZnfVc3ENBwp0V1BCkw+yP2IoqzrczQxQj1ibjzGuT4aNIN+
opACrY99E+T+fBDxz6kF5mEtaRn/JWBUbNurTwnbxr2lN6DswtP5Zw5IvL/gN9ku
yjzpBfGr7hwWAay502Fhmyz82hPuNb47bYywpQRoObxBFZ7HBcxJQNLQd2DQX3t5
jkPW0KSBwEQP9+Z1jnQHsoV1ShG/hWMLnYYA0Qg1UrYDUteuoC8OgO0OBjD0QqXI
Xf6CMLv23Gniu1GjdAzKvw4IZKLJuoIx/JAK2iceZSjH/jLnT1aF9PdlhrCFzgia
0Hf7BtLEcElGoc+wbG6eav8CqnWgoumDZUFtmMB7kbprQRctqw/F3tui2T/1S7rn
yVQazwA2mIV9g7vQToBI3MMnJaKhJ40C8ULnUEsxHzDxQjLK+PD4ZgbzMW3b9GLG
jyFQH1pSF+JPlAsOWPWFO9kO+W0u/RCu3XghJznIQdvxgAk+i3Zl8V89Gt45tnjA
Lp61luejF2/7UftMgC//VJOKPdOl0aIXHIi17oUcOJq4pitdGWnWYJqzntn+k+gr
7qL3P/E06R/gFZi9CSRP5SVmlk5t6O6lXBPrHdpLX9lxw4nW2J/+ATQEcPrem6wj
GheHML+L105cxckv0F1wdQ7noudKQ03Fdk5UgFYjtDBgvt0v0NKdK5eNFQ7nsbKS
a+7TvYhJOTOxs68l0my4aY0kAfOOhbCPf+hhdBfbeFjjIMmmkjnNH+2ITiStbmen
Tw8pbbm/IXbJgJK6xD5S+sK+3jpgm0grQ/gqYn9U9OWfgtY8/BEChwEzjrNyrkLw
rVKM8DobrpYJT1KqyS5YKV4B8FPj39on8JTgq9E4vDEJn7AhIBX0AD7fL5m3WoJw
iHaqLEoJwkyN8vb2q5iylY1W72gfqMdjW8x+YHU/oksYOC+QEAJIJ2kBGr0e6FQe
jqxktJ4dhsWNLoUHxTUUzXEaEN6ym8wvDM5oHEpfutbTSVz0Fvt61I4ei0Ed7jP7
d1rY5ptnUijTsBmCvH9OFMDnKTd4qgFX6crkFiEMYHeX8C9XHmTxA1yLig+TbYyD
ATBJLngG4cMJG3q27CTtuHHSTV5VQ8d0RwQyWoiJqmFdwLe5+sS9UI4ZpZGrz1W4
OaDQsmatpWKICF+lKLxiW65J0xaG8eMi7Okqdma+jkfx9tnJMSkHBdnUGY6D5S00
9VqUieusZbvPLyDYxyJwhtNQYfdN3VbnhmkfSi5VOX7ApSaywJwmazVJ2PiefEFb
UiaN0M1mcdhmXAL1a0UVqoLzIqRE4PCYatRCj9XmYqhczyxUcuJIe8fQPphnq8LB
VX5Fp9BeN2p4r08dj9QaXzZdzNlnTna4aSNX77mxBAMYCZc2R7bLM7HiqSmrx2oQ
gXSgCkaxQ4P1V4xpo+B5DlLH7RZOhySiMEYET3zSQu8gjYd1H9xY97ztjrOy0tfW
AaVOYAyjFxgUptTA6UZ5EjKC659cCa+njJ0N+tzrpTAw696hP7vJPnc/Dwoc7Fp/
MXT5QsesZnCDzUUluyidBgqrWUpycxC1z8vY3DPzSgmKZcQgr128LfvW+iP2HzXK
lcWpXWXj5PJxjdv44JqeIGrwtnSyB0NxuLlyx9KigNulL9U3ydv+ng+7aCRak8Qi
P1LxdeXgNJ4WHRtr4mIDyzlEIIqBqRSV5xKVANSY5swTiAf+4jwg2CbE5LMVCXYh
4vvEwKcS8W1ZvL8RSzKp/Ha1RvS/VzUKgh8NpMrOyXcFYhXY4JwO6/+RII0IvHRY
PFllO8UAqRjsgNq5ek2K4OfqCtAHH5Bi4NCKEYLsHaN0Ewf75EivWBJHrDlxDtF3
TRj11JYHTTOPtCpcACsK+WwVC5B7ph+hcXk2tJMwwoG/cBTwtjwCzM6h43ya8Jn/
UX7aDKrcn7yTeX8jfNZS6llIEI0L/j5jjw+ozaB4aJkhzDkheQgl9yNUqauSuAmZ
iZVOnBsldp0EiXDRGpMuvZzz4IMJ+XvD2QKo3YohFjEDSSZVSwtnDbMS6/xc4opI
M0qAtlME5ieNrZedi4h3CBIdn1gIwn5WwGDLUWqKkLlrUtP3KYWbdmx3MDK+gaJP
fGhfyibDOzWX4RrPBSrqGoNjKLcRKqoP+o2SZXak+XFA4rNMDCrw22w9CS/i3OwY
W9nqnRBmkIuvuHjE36xPbYQXOW1Wyw+oVRiFFP4LpO1VbEOHWoqheWmGllcBIwMS
cmRXOnogELDl7qna4UCZLw1h59gxw6I7iPA28lelsgTCFP80491SjY12XUmjQfPt
whIGpDBSnG1OR5aVdCyJPT4HVPiQvDKffeFi9i3TGAFlE4G+DD0NoVMC9Gqzj4xN
vuu6zqfevQrVyT+DYN8AFkPRVyoHfOUB/g2+tqF0csEr9xM6ywAD2jq7n+tFp6XJ
A5mPWyPbmlt8+qpjcbslgJuGNs9V3xXCq6I0uA/Oa9cQ3THSq1p1bQ1NGWMtKDZ1
hzzNwohdFXjGY2jG1cWLhCXTz32FM9LZQIP7+SAjbybEBra2Gg4Hwwa4JdyeYKfy
PrES61gtzKg9H5fSDes8Bm7CF8UnG2BGqsAhOy2WseMeRU6UClQUer+BfXpW5Wc6
DQ9FEukpLygwrY8+yvwMuDESbRs/Lrl8LwQrqt1evlp3uCq8p0zG5S+I/iJHxLPc
60vfBv9J7bvSkw63C+8C1BdAw+fPglJvhWtW/kTOOQSPmIpXB54re1AZq0e1LYSD
7EXsRFicqJBZ7qEwMpciYdrAkhnDme/RRky5R8z1iq2O9GUecalyoABMyPdAiUrL
aNg26JoXcjaZ9iRoCJsBk/fkBwiqKevDSHSJCY6OKcfnQnyewd1RyFyI/mZ+440U
mDJtB6XBh0q5Gq0KKqt+l4Ex0uWtiTWgeWpSK+eZh9fgVXuu24HwHPPm8bXmpNSd
0RcnOBnWWgzFhQdlTyEIbuBHkDCkMH6DEnlnOgTqcUBGGqW7BXv5CNm6SeyVyFpn
Q7SiPOEWCTuXBkGP7yRYx3fWmuUnuSAjNiP5VlpjJeBZ28S+XlCy33VxZ3Shpyvb
IwQxIgd6AStew5Joy9U9ryhTWo/VWTaakqQ/k1xhgumOJxB8HJvHcM+66bED6lXq
D8wmujS90NtafaRAeW9VuJk74D9wm3y2sadD8OwfF2j+/wmijJajWbBNfCwT46PK
VNok8wFzroMs9ZYxQCF/tGBBO4GFuZMfv1pRULx/hTpkbcGq+1kE1uJKIqiHudOB
0zdQUpDMZcs9XXjSmPlI+QscunCdSRtlMqKvzKFXLOXsc4HlEvVZPPN7dHJvDViV
octWfxQMbBNiBbEaRBxE3AFgBrqWBje5N/oVad4zeN+f5iCCabYcCx2dGdbLOoeL
9NYb/ZIIR6badV6HnNqbkgyk0oqA4LUMczClsMgiduxITBleNNBq5WVLRpaeq8Fn
m6hHjqey4+zVHr+i+IJVvEZ32yAQ8+3VRH9T6SbiqriG2/sgHjf3bJeQS90armUG
o9//WGByo9tWrD4eVdJcRAqKJSpXkaEwYGxr4ZymZeHPeSwVtK/bUIKWPIY70ler
4/HKZITJ43Vz76A8l7O90cCxTMj6BEg4pMDaJS601VHk1JbbQR+tjJqE4berUoYf
RU4DBEuhsl3J6QBWaYBNvQ2p/aT1woho9aaR3bb2PzAPCxgZa8Urf/BFgYyemcS/
1ADFMdq9nR4917gY4vHgefJfL60GFLXKaqwt4EIpGRag35anG73WGQB5jO3l4WY6
eNgWpp5qkTY/cZNHVuxzcl50wjBkaQ5wU4m4PULQjy7KtY3mP1s0wxlrymVI5htG
LPW6T+0RQpyPbGHI1uxq/WE+19nOw+v3N/AVpxvjQgDirE4/xpjMuTgzHemeQITe
11PV0KsvZhB7MZ7ewkvC/DgCtrXPT6XmVOq6vQX371c7G6xFwv9JAGf/MDptoD9G
OaE3AuAsRCAEw2DhQSgm9AkpBM6nEUrfv7h9dgNWP8MZeVne2erEV4dZKOu5ZUvU
M25bjiaihFQKr71SzOEvikMC8NdRC+KkKaN5KOFO3kKimc7KdCwiXilRXLFhUn8G
LOudYkuTXkAba3QZGoC6bCKO864pjl+CeY2EOGj4i5MaJO4GaR5Vl2iOskvDtuvx
7gHSgielO67Jb3za1OhknLXHh8+ePtJoMOVekzgwJaK2NTdDK74juEFl+hTMlMcS
ZjtyeQmrpcLLFLae06YxiCG80+2h+9IChOvI00KFmpEwE3qKEDs5cEFvNRwx5awr
1fav9ssyNdBzxylCSNurfZ8u0jdYm+J3JYLvMPePk6oN59JwAdOtr2N5RpcbLwlM
vXDvpdNJkAoONCWjWp43Oymj+HS2UzyKqDFRFO6BSJ4FEfnogX68vjOX9xoR+YXb
zUSXIu9HOkxQy9+uje8AFvDxZtRcOWQQApA/m5Vfz3dWi4d4uUe1e5i7DUAVa/UK
rFrrYNNfY3hVX9hBtu8ENsGAC5W7hvsPq3cr2XtqoTjkx7wZXjgGnWLKp37H1SZ8
maHJyKFTpiS0GJNu0YBTQ77b72Ol9+xPsI2Q/k7ODz9DOlHRt17Rjur4CL4fIn/w
JHoJDAxluWqylQauOMJ3L8oMC2sDIRWgCoDrtr7Kfgd//oih8Adw4YooS8nMZw9r
5x+10aTiaAb92vOoib4TkJ6WfKAy2sxf3sOU/ycezR51pPyel1O8nRugk4kG/NvW
NqnC2ygUDdOMt4QEYWayyCdX3q/h2YQEVzce566V1grf+np2TWK2LsF5IB8fBR/X
ECwhaPKE37htkoQovaVYwwIOUQMnE/oPwYwnSHIGMewVB07kOCQ+gR3+pK6S4qHP
gw03qjzUEIwECCucFXnbvLJD3wx6tcQUdNe81QuTUjE/iDGnYpPBrGtc7RSEEE0b
ZO68wYO/8sDlQti1/7z1/+6CNJ6zlHBKZHG3TPsXYdJJwnM9BJ3jMiTR5rqGMmcg
udTIc1X+hBJQNjNUumP84sX+VCXHkZSjixBtaaf81bn/CMiRLe2iROxZS0kjrzZd
+lrxX1JSfspUvh0lGs/iLiM2kgL53avLSpokrEnj9UVBAfgYzgS/p66LZyhNeXnQ
TInZfaaDSkzEB4LXMYOISuw/kCxgYYuiEwhwbJ2c5jZyKLOZw+KLDN5PF9vUYa6q
GU4yzCXyv01dUTzWwrfAC1twxjCrxKO9w8BUQNPvK/rMKI24f/uxO5l/fvB+e8Cu
9JJMAo2SHnvnFrT6J5Yy3M9o7TiqoSImYds2+puuejuc8noj7TySa5x9fyy763YR
hG7VDlx8NJuA0ZuT97sf4Ix/S1agKdGSH+gQmn+td8m3svtltBrqMT4Hhtwgqotm
4gSc45TyN67ctX64OncwEpf0lkVDzLmLo11KkpdCyVtV8ejMUHID2QL2g1+2DWdL
KFyfbc6rPLznsNEMdGWWv6hu0mhZp+8hRWpZKR3Mpb8MnbWrJgSSlaPJB0D2VnjO
WAEVzZFBqWFP/S4qj6jFBAltP0jDxR8MRxsFfHDoDPhc72J8R9pGhTNO+YTas8iU
N8DBJEsOEgAkb9b0TlSPxK4VrvZJtgCQ2MlmWjO2gE1xO+NkP98IpiabQALmidsl
rDswpXnsHxZYNQGUbOcFRPEPxCkRn7NBa1ezF+MylQCw0tq/QDDQ4VfrElP5uZSw
pqaEPAX8soo28eXPtoXPh51zkAHYB8g3v2cEi3OdfYEDkitBX/np2fpWF/YjIL4P
RM/AtgtuTTPEsJexInR0iHsf0NSjiLZcZQWOllj+ZrChBGSSMLewwFV0v2sNrYC7
Tv9seT6xAWGzor3+Kon28w+aMVmctnYMRutnx/sXZmqvATtKWXituvVD00kb0tXJ
34CMbkB0zXKg2ALjcuNAMjjJkfTlvBzZdDk7+thRbIkKi5hl/+S+R9nMhuE2m1V0
+l0I9OIi2xoEjKsUsKTO7mqEc3reSku6kYnJC/8wIzB8HnwqYVwG7psPI1jLCMSq
5va/aQTiTHjIsdl0SmOsN/H987eJ1HH52uAPLMLdWx2Cu/GFKSHZ34tSDObLvWaz
QrPBzxrpn0jn+3ECSYS+XEByPuYWaGGR+ma9bCPgtcR21DHp2zM8NM4Ioyn2ySlH
7yRzl+rssF8PS7srjPgxoCLg0+8KKmpNUqnwVIAUt95GVUms9eKBBMPAB54uB+je
6Dul9FjKDCG3LlohYgVIyxEAcwmpVK089W+wvaJYuqOmZX3HMMe8Z1VH9Cnp+iNa
DDg/rKW7f7EO9XZSvytBOe6P4NdCJXKwehI6pL26EZrHZIGhW4zEL5jgm1wkM5sY
+diPj1+twzhlx1AenIaObpqNZx+X++bO/DKQST/2u6DSHnXT2f5CVR/EiSSCKBCr
9vRnc8NeaguRTy2gfOIfD1JnOwQ+8InpTnzsPWcqpxg9ED9+b8bhFnMhYHrUmFIp
2dIsUHRsXslvWcT3zEzCFMeHjnMGNCx6sK/N66ZBVpXDCqLwMer60w2uC7VEwN9y
D/1qTJmcAqVcDbiEnu72E7ZDior21xB2lAWcwyc5lxwq8Wa78Tk4EUAnqJ9ltGRD
KlSHQlwAKNNfCUGEKN5AQJBp1Ij0FC2ds4WgMqfydy7PZE81L46DvKGLiHPlOYF+
SbN7KEYfvYP+IIpBqzVA66fQniY2nLGTekYH6OaN+ec7dT2KmJiX9qGJuG0Bhv6x
yiqvDU24kCEW9I5mu7nDsFgjOsGhMlFU95n95QGAaIYqG+7B3z3zwJ19i14FpQDE
sjrDOwHDLr2Qfbi4J+vqjVGdIvXespx4jlb87iEhaM/o0YP5lI38bNe+OeXhr2qG
EGO66cFezcoMa6+96eLVtVoFD6v63VdMb/IczV/d0T1TFsc+EU1qM7z1U4jUk3K1
mH9/gu4vvP1/8YrmI9TM+3GHSWtXAHkUH0CrLLbFPmPHwZ48opYa0kR4qzfIdiWG
zVt5kqHhlmS5KcS1Gq71lKGVfrBYJeob+VHWt22sQbZJVLXNcfD/drv6l6EiW5kj
i2gc9cl6KIo7AfZfy5VIHLRWqV4lD9mTckrMa54Pvj7Z+R4NWtuFrXQBoInU3pyl
2JeIo73g53QX/dG0qgMJy+yPDixRmM2t2RSGIktFXJKKVbHJoPBamcYJAf/3wPUn
EDYzuv11XKXt1yKiYbUYlRXsYpUxhy58D/iMukEPQusFKwz2bXLQjg8LalNCetox
JsgrK71AIgBEphLf4qL+cuCqPIdNxaBtMdo2Ol+nPRCbBtoFIyxdMg1+WweEpLE/
upfl2ix8aRiY5GPriT2nkjE6sLU0qiPk45W+EibeyAJTHsjW4b214ILGSdmcWr0r
QvTDgFonwWt0IGe+aCZr+k+pqSZ5fZDiKteV71ddf+2rcSjZFoQy8K1T3IRBEWFu
873tp38T+sD8siNRokpltwNNPVD5uQ4K46PvFkbdX4t5wNWDAcOXs5UH37PH3b21
lO5ZpG4q3Gz4mo6HEI6dYvOD4pkyZfBwHQq6ChhPtjDx6hsqg9wfYqTxNPJpaO1d
p5T1KhNdS2u+MV8LKgr7xI8vnovf5HJHBzxAh65HC9s4NJpjMtX5vekdXc2zVQ+L
en+zPOBRvZc6lZwJ1sWhtHYEDWiBKyGthIiAKXrAa7swvRluhsqaX+lNvCjNasFn
Ek/XgJ44n6ZJp+SzYD4R1tDR0paa4rxOigz/pxt26WUeyhZ1xVvHFb+DzPCzFCrz
2o65GDqa8SPMQlQg0evedpHFNynEO1zJqgDRZsjB99CPrUubvjqspMBx/Ax5kGB9
G+O26fSQSHhdcaQxJQga0mx8l245G6fh35AfVyuF5momnHEB1ykkB/xkn92hV6kr
HGehA4Vs4XQsPMFuxxlo+E1UeZMUrSUQkTUNhxFlR1fLGm/bm027CV5i+l3coaFN
MCUFeMbR7dEU9xVZtVKo299aoBZkDbunoPGJ1q1dsFDiEvBh068t7DN+jW9CylAv
VppiUyHMTDGo5G/XqbJXTGaswRSnVX0dqAXADQ9vW73Cxjg2C9Z5Tkb5t+GbTWJ3
ZplxBPz3dLuMzef8wSTqZZhVhBPNfva3Jfil3lDRdT1SCnRGajJexavyZ2HzS+B8
N9dIlmqqag1m7Dk8XQzC5GgdK41bUE5M0DTUQSvVoUVJQ0jzag0+9fKA2uTeU9d9
k0iFIamG5HX3GuvfMFGKTK1+/tcNwMIAmNymUkx2VCCJudbZRaNBjR/oC9EOPaM8
gAeFijO3JB1oQKUAl/HzhaKL0g5Z/NLpzS62awVJ49RTG9HbvcTV3uHUChcHv42x
hMLsyvoJXtP5TOe7STaQuBlN21CTXaZwp4e7Y02EolL9+JyV9lrpwqrvAD5qjrgB
SuAw2LaTjmUAQzDZ11RbkMFhWFuuQc3uQYMCus67e/JrIEvP+L0uBDIA7WpW5gr0
V6u9fHKjX0DXU6VmaMBqLwE6/a6rjmQbSQnDJCwOS2I+zohRkVWazt9lqjjdl2Cw
VLWEEwMh+fphzwjlpCEQB66xZWyDoMADfZlTxP/CiIAgckSzpQmBmvsvGe5dV71d
klKZKfmKde2tdNLydN7zQB0o2m5HgAW0EBwWnsuy/ZmcnAdQ5ciPCaiMw4tqiZN0
OK2uWV+B7KhfvSekyEcMeNvgm8Vqq5560dhg0dWqnMzbWkEqJ9jSMYGDuayXbUhg
aFfRZJ1TVmBxz0yNCFggvKpofnu7Z9YYAwy98TAljcOR3k9o9SwJI+VetTf2wIMx
YtP95STCHtlScCrEISQ4I0h1YzlnhiKF5ugoV+ptmXGmLQ5Cvx6LOWsPyf2SzoQG
1bp5n1lXbGORFX5mK3mYytTy6fcxlW96a9AoZ2WkEZwnre3L7oo28oIKvAPSXeIL
52k8G1JIaMn1WDZj9OPellqEH4IuM7ckQNsvOcdcSgwYIAUQ9fbUr6Oen04R99lo
Nouq82svlUFIsoCNnSDVRq7F0ujJD3ST0kcRM7bIzK94Sbi4Hqs328nvoHnx1zRh
1sOAScZ85S+ZTFmOVBRIU3SpJMe1FPRlXXm8j2gfnH/66BizQNc+pmJ5JMoK7m8j
lpqBWOsN4HsnLQ2nYkzCZPZgQNxeRuoVkJvnbbwSecSUzhLe5ZqUNE9Ryo0Mn0hq
KBf5DYx5uvriZ40eV+eFislNP1aftC1tW3iTqHgukBycQz4i7ZNSJmtsmzqxr5Ic
5lntPFgrjb2bSYh2wHsXNH7uvgSPvb/Zoh0zRqTm4efBn6sxSW1UFBdrRBe9de7B
Qx8q9tGK5ITFO+GVzvCAl6pRhAQNB/TBI3HicVTO6ELNSZiyPT3IL4GHndnGRVr4
FjGaNoNpDtzg/AxNGg7JoU/vA7e9fVz+aPdlfmy7mL1fYaxFGsVegbEoZJBoiMYt
WcoMnA64gRwO3Fn5G1yWv79wFYiPOu24F99Aw7RW6VzF/qa35V5HguaEyKUJKSzt
2pEsjyRIH7Em4+UtPwSNQyoYt9pldzXvGhyXME1VFLG7+zBoQf6GwJYbIf3BNhUI
r/rGLil7MGzwlKPbyr8zg2ODHG6VU0KoSx70JwOgzlSbvl5SmR0819ufRr1lOFI7
F1ZzmaxcTBi6VGVXBsjoIyDNHmHnmUp2GAcKs+e9Gv8GZ48GuDE7LcgfjGIv/osS
JQTF6yv4iBfJVWkaeJJDYn04f7MmvgWN8qxRNSuGirATCz+1rivbRQ7GDzkMSlUe
UTXBvTS76ZBj7yg+FCK2N8PnelcomupcP6JPbHu4ESPeTin6ZGVNKdrCQqztekrJ
MgbIqpD3wb56KT/1pJBPzAamqqhrr5sI50+sRTq/GOf0bUL1Hsqnj1u4iLNjTMoU
XHPMdr82ah5yaldF0fo9zZ3jqGhk8njhOHv5mFvKB0D1iWffbhGhcuHsAgBumM2p
MXAquBiwOWMh3w86yhf4yMGmkPryUXmyqe568MdjYFd9tUffMlnKZVLnrUy0cAxG
kHwGmpNk0QTZQzC7c/X5iJI5aMgQNifka4pcGqGBnHBMKZnzDAFHwHQ59KPwwAcX
Qc82Z6MBFcBD/Y3bGvYOFLucX5uGlUoUo4G2Ac3bPoXOsbI1a5GcAaF5uZ6j4dZi
HfgnWOc7Y+2FqYIXfShClAjd8SySxPvSmgdXK9XjM1p2MmWqdzqHbkZnhlfQmIMk
Ells+go5lG2j30f5yHDTzcPUEXPPGeukj07b1BzSl5q5QT9aeu6z6tbi3+YTfzBv
m1ObdkPq2CsoqCHgiTqznRMGSwi7gPTtTaIOsq9E9LMcvObhPW/kRQU/eQcFjJ0/
42Rx0DflmC5tyB3aFtaW0N346SaFOOAi7oniZQMpUPplI717vCfIFsJtUyV9uMIl
WMvF4Ltx2OChLz2GTM59etN1xLlAFyipc2RVqRiABVV9qcAeAYVRqw6Ggzkm7TPn
suRk7B1iZdR9MbLISFRUidKMlErDDmqYunmrRIaOQtcAZKsbmcvPwh1VwuUQ1U61
gvlMNiBOpI7D/VfRJN0JXevoa/b6dvScORxqLtPNM7UVSymhbg6bx3bNHHXRrxwy
lfJkXyYSslHbhI2tzQAijabAam76Z+hppFl0iaYzgB0t6avzNiZAEoMcqa/XMxLl
q/6hCu3qjOUXrxAjcGqrakAlmMGwAPH4C7ZwmbGmUGUG2tdrphdYHFCf4Mqm4Jkb
3rEymIU/xrvRiu1846ywqCmxrp9pmYi4A18nEXn+Kw1d47/k7DTTZspL9/uoTDki
21l1ayJ4o/p3kqgZkt/C1xCgqOqbPY2ZKcoFGsQEq2atVCN4U3Cp3vuy07AtJ3D2
B8OzgFP8pNdBrQ8wQaqaf3pTrl3JT1ifcGrajM9lIhbo6t08VR4MDfQdUSP7Fk+g
Un0AgdtQ41/4/SXYmoa2vWUtyHW1j5zXHR2wZTFetF94g6XmS2HF3On4K0m1Q2S0
QwnwUGHPlknpLeNbMV6WLWXgeTxnLgCPrmU/vH9SVJjPxrjDxFXz98VK3GRAc25c
SdsfN/THMLVNB2XonTP5DIup6UUF0emqs0qxGC3t8iTj5f82uNyLfeXu0DJHSlUH
fpq0ntd47Gay2uuZEyx2gnvt9jTMVKsTWbJpSFzyqudzQdN2cxpvmCDZdEtCU9st
fp7/UEPli1YDum88s2bQbe9MFO2YCAVtlLNJMShfwVTJHeCrwQ4I8LYawEPqxVSg
6bDVmfuowGChuN/QFCkgyILbjnCR0DTY0Z60QP8n4LKQxtDp2qtXL5HMtuzGf1jo
OcN9LU3fht2vBVs91Pnk5MEiyRMJQBIj75KKFSk7152g7xQP9R7vLgPRJseON/S4
48644AhZ+QND6ycsSByMidMPy30uMex/fjA3mb1oPw8T2I1GLw95PcyWpwYyWEMG
JEWiclRkQxdPWObH3l6sLXA5coggT7dqZogmSK9NeDNyfH3UulMSRby0ksn/OgTf
SDmeXoGoFDEPDxcp5jPUJMhn4r6yDsPf8JurFVGQF/s2ppEqRrvaVuUKC76ScYYh
pXBEdPd0ul8hSKEDKrMcN8Z2adm+DEHYduKYKSujJDvyKyW6ag+f/l4SaPN3g1s8
S26P5vd+7T8zPmvZt8/ccBLSp1F6AQ28AiJ9JV8gXAIfObSp0WYSjTKHrtRTxyI8
rJzPn1itxCM9zpWdCgFojs1fprHoTVooBQuqhsxrH5IIAs0d3OR/vud2wbUnqvkU
TcYnosCRJAgdncYZ6atL6Q06nIqBmCyw/51WL9YN8F4iSLLk8nI6eCu2z1M71lHC
dfhWZblAK+VUWvU8GUPBBps1pbc27ruAD20tA/QSnYNKFD1W/NAT6VCZOsE1h8sc
u6dHJ4XXtJIfo+Pm8+RMOqHQlkt75i8461gaj8Pm6+gZfNcrpI1ees+aK+66e1XW
vZYjkevEVoWUB5nAb4ECt6kPVwxLqhHitx1Al1ZxC/kebqkf2ZTAHcJy5dW5P/1u
1dBwU0DOg4Cgok3uy+muPtgLuA9A1A+wEXdaYUXkPklrC5lvrJU9kx63sQDaLFlT
TWqSO9Ie1zdKihAAKog+ZmM2GobHCPgaWp3f2xb6g0Jg3PA0n+DAQ37JOGqPqY8o
w/QTe8/k7XX4c2W54K4c+g9EolHbovtzYdPJo5aEWQWOg5iR+7waac0WXD5K6ZHM
DThtmSDeNUZOOKCUmR3d30dTGpTq3ZM9s+oCFmRpKAZ2uZjrMJ12rlzIWp/qPPZy
DI5EGYuglhxapUWr0Ki22GIyLrDho8BFywh/hS4DYtnCU7HtztxNENmnWUtOlrLC
20uiuJ23t72CUQrM8R5Lv19cbOhGwDCkCeiQPZqZguZZrRcPoOAL1iZMaG5qpyc8
GeU+ghBzowLP9D++1Q3e2m1Lu/RWqSUeqeTHpXyP9chY4Du2pggYPMiOl/M50/Ky
SuyD0o/J8PybV7c1Atalq3ufQL+h0usco4nUFRXJPw6xOp+iV4BgkoPjqLfateY6
75YZlM7w/DO2NiV/qRVZvxBfis9xlTYVLjiUANALjRpMfW7INq7KyNohNiSNEEip
9qwcvpyPunyB4RuXvlqiXJga1rXGJlph8LSzgi4Obv0iS/LxxDYIye7g3vByOLAD
YUqNwQTlmUKvm7xlZGINrw71LoCzgce3p2zaxcKf9r/fyr0oduoEcWbzuWQtstxn
CdIVFXsWCTowvn6+55fFc69EdsJWC01UG/w79+i2+Xy7SV4D7L/gRQhaHSDVz5S7
aAh2ew4vYG+gaz8FfI/DHbefkBtfJcNrXcMmWbSMGx6+6x3Xinsu8ssQ0Bi9plXr
vQ4dfw5p5IHVGS6qlPaPZ+BDeDFfapLa8FeXBMZcSP4U3GPoEHBxoIgaX78ljcMg
8Mwxyn92XnNMUIwfl32nkWhzPPb0LFF3XFvIZ6BiyFWCikxOmx5U1sCtXaeReNQo
jRaU/MY7/0a7gORHAblTJ1fDDpcyXf7YgWpJ20lhoUKV9tMPk/m84G83qnF/gYUF
2PYi+e+rtH3NDF/XKItm7UwbZFrjPG9GKPtISDTUwbGPTVsRid+AsLuDf0ySRQJr
GkzEe3b1hxALuwBWc6FZAVscE6MzU/ApDQC05FFQ3pUWDmJoA8eN1uNKSXHBLkMR
A+2OZvZqIsHhHPknBPtnxrIN56NFpP3wsKEhG8E6sorxxwWELqQMNXmlWwSTWahl
ncYGJ/kl7u1PULUhf+8cQird/ouA/uEbjBTkOA8fUKtSz2tOay6MibXm4q/WKDxV
inCeeq2+VsgZwISC2QVW1gdR5SYtLTXsCaQutY6Z+YNEYsEJdA4hpwXsByxsKPsN
NAR3pJJ79TqxpNjtmOEEVBz7G/So/Vr9LjeEMUptVL2EMtSte1aEww20jrDlxG0/
Xdx7XMwGzvSuekxbEbvX6O4R4y34WpNdQRmJumfV6M1zPgvqpTfBk52j7Q5ANXm2
w+WU7Z5HMTTr7rie8dZz1ls8UAikU8rR1AR7Rk1+xG84wgkjU67+y/pG7QtiNANI
2OXB9tibFS6KvDN5sSyzVlUNYN1dMnthU7bpoS6QGa+7UO9hQn0uszLTwBDDPxLq
sdzXbp+fYLOX74gEAEfaD/cAPCDhXQ7KAKS3ruiKNcOnboi6MRuOkGzn9w1agrBX
plGxKVsqOo14f4iIe9CAbBEhQFTfDYcZuOJpLijJkRu3eDBYSPQPYa1mTSFXacMn
xbHDa4O/w5ypzZ932ytq9atq1ZidrS58lmnJa1XpGbB3vuAVkBux4+Cbkhi7UYru
Nt3ECZSJyf5VO71I70lRYYrtpDMIZFKSoB2LTaebYu1Vr+OPbMem5Eq6KCeFH3EO
PuyH0t7HNppLQ44On3H2kDCIjOi3vaSuypROc4R81N8dzvANHiMYIq709yM1p+Ai
h6YnArCQ2o8onV7eyirMJlSdGDIl1Xv5m53Evz302c0RcvT3FxI19XZ0iOdcBB8a
qVMSxpzG+J9kaglV5LbW2IlP6spOXq9J0bKWRF8J02/pti5xbqZmtNnbwYWH0nC2
o4cIKyUSiB6LScIYmQo1WREj87yxJJ9RVqxCTEtRLviJlu0kUAEL6wXyhliIfexX
8hGwMAKljnhXpIgWKejshEzHl15JzkAvu+YxT/XMN0tXO5rXv17J1bSxK77HdCqu
VLpk3ZP1X5UDW5/rzbB52mGd3+3nAAIdd+p9abjfZ9ibbh/53aO7d9yLY6s/iav8
teD6Z+2tgdIknw7dHiIr4pVr60NXW6UNsrarwDtBVmgqwsLQOfpWxfQhxvXopUWE
1wDyKdzRc3YxixuN2efUavEi/3JuLi2Fy9HO6JmU1BU8eUirdWVYLpTbWH7Bdpdf
d6okSkb2Aa6mv6SydWNTxgMDvIgK2M07BrBlOVymQ3ZKzejZO06BGqKOogXcj96R
FrhBPCu3n0QNFCg697lKUgzcS5GdMCCf6Tm06RSmQKfyKJBWGcQsTSEpb45mPt56
KjewhpksCJqhrJkzPfWwS7cT55tywpmbjflm6F3sR9leGtyEzWOTPkhJR6CORcvk
wDHtsIShtvKIB8DL1EryKyyIpwCZKUt6sOKIUvQXNDsjQwVYufCx8mQmv6Li9j9f
/Ead3X+Hh+wg+UMg2WHjMwaad88b7b52bj3DyrrEtTWLlysGaGi7TF1af5t1KK84
0GuKx4olcgbofpheJEShmTiSZV3oaAH0UecOARfEH7eQEeXsid4vTUsPR5Xl+Jue
iyZiaLj65YIqil073+3ye005aNbgKaFxaDjvucCJBXOJQ1T30lJ29iHFmP/0SHHv
ii37DsH9AxbjI6ZOROqG1i3fHNdXyMfglLoHnyfIsxRK2PlnmSMf+JfA0lcPv9cZ
5ry8twZarNoy7OFdftKujg5UAhitoh9n/sQ5klZ52HpXi7tOBExJeQagh7OR4PKG
NuhlqS8ntWA9dk562hx410IM6PKnJhoUqTCQwQ2B32upbuDFJ8UCqPOpprKjsJ5j
naAmT/BidUsWozyy1DPnrQWxrqI017zd+rroH9/dLeC930YhDBslDx3IxS5bAgKG
IMT3UxWWLyT+h9GzZCwuZFrjMbnbdMAN5aQBE+nyr1+BqgT0ifOw1Fj5Q3I/yDxz
9a2Qm3fvQzYIOq+UZePDVrdPk7FsPCZp8UQM2pPray4+Ibt86k7279rubtWfAhp7
n6lKIPQtWL/os2/CRsCkjZQhyR+Z3eSkW3TfvbjN04Gy5RqyvnGcHZ7SX5WJEUOb
y41Dme2fLhAK65+drGBcs9l/ehmIOZXg7NhoCyUyhjIs6qqJpvvaHY8lPCOg2Rgt
wr/Wdy/F73s/ykBvupIjTh5YDnOhv/aNqQcqY7Jx+ZJXipOATRjH5MVuBJGcf5fn
+Y6ieLh2ZwU1VOnk8VnelKL4C5nEmBgR/obA9NmN4PjZbMb9D1K2Nl2ew4K5fmTn
vXx7IGr9BqTFvq+KWwCrqR3ePbpR6Zi+AWyHZIkVbhVTh/JMdQ/dDPcK9DlknZfp
mb27MQ3XkiREoKFpaFZBN90h8euvjw6VF9UXMmWUYAHEpUZLRDEQpCKt0YVdk2zS
/LsS1WEZ/anZoAHv//TPow6Zvz/WSCTeAa5xHL/9h/znAKEdb/c/wu/4LIFbBTSP
nwY2cVchXAH/1VAkoyTs7exEOFkgQ1+kuEI5DPPL8ytkUeEz1P/xRs4Wig8eBuxS
XCq7b0Pq6M+1Yyd2+uH8o2cqP28lkTUGe77htXo6Gy9oZPGM9NMDgYZZaGROS9Uo
woWZ8Xj9egbwlDtKY3zluy8jKqWcMhAuJT5dpKDXoX3snsS8me1W4H2ET0P3RGFU
0ZYKcaiBZutwsx6xUSAk51aOhpLJCDhV0XsoSd5Hmw+JQlIDdo4BcCL4mlkSdDPg
SEw3RDGp3C2sLctA0FIw5O+EC5oWssL+3/I7vGjtDHotzqyY4FaG3r9vREPZbHJS
F7g7IUM203AYkYazaT/s9mmXyB/Um/K7VR2bcmGozwYAjFESRIr+YCqI7AdMeeur
4x/1OwNzpA1EwHsBs5NQs7KV1LeFMydVkPpTXHdUMuGPiYWv8qCSqupua0pa1EXG
CHnVIEyqLS56s4IF6ojkbxgzV1WDpL7mOHo5dP0E0bzlr5Ly1XGhAwduQQ8E3aDE
/lQIC1y9APIUfVYaPHoW4S1d+XRJFfh2DsrPcqJPLiVWKe5TX7tIDL2Gfi2Ma+Am
9hJkDOk+4ZNLPx26nvRc20HtVpiIu94iePiYtl+/bhjvPdGYSoa5ytQDpND7uJj7
v6fxhGfCFuu/2o33N5WrVifWlRQG+un/6P94My0k4Ne4VSf7ylMdzlwvzOsKsSxy
Cs0y12ybUx/i1Spld30gWc8er7L2rabv9anh5rvHWqlPmxBel2JDrS1nGrQfq7Br
atqj3aMClpEfpUkqgXzGqy2ZQPd5kxswZoBuuaCNlZH1Y+EMEyfM8nMWgX0AXT/G
z5/B2vktB5eDgMXlcchrlQLfJ/1KUrjcVZWOC3eYDY9kHc7NrAFikB2Cl7W1zv9i
O62CNfoYv1/CiZEjSc5E4+40aB28QP9OGscxO6AzP3Eyw1NuL+V828us4W//QyvK
5btLL9//foknuVi35wLOTPIJFlUwoRjPc+nuaVUqPtusYif2v9/6WTGqgNCqXhYI
VfnHXBaRdca6rCig5AiS7kWX2h2lgyAHyGVtI9A22cfCcCjTSagq3p4ui0lc4uRe
qvlytBLBtHlITE/fmEnVUKh+5xorjNO4Dr8EUbbrWhQQodNEcTjJwAELZoEqrUYf
CYMyVe6rzvjVPQFPPiuvIPHlaBQF4c9MgC4dOM4FXx26wXBNXEkIgZj3EYd708z2
TrF6f0aKtOiULzQPH0wA0qrV5lvEMGRAwCmqA5sUGYWr/2N9q5+D5MkczfuGIyjE
PSYydzTWoFjkphtD9CoYc6Vwg8RYVRW1+m3Wa50bVR3ZrDay3HmHXYsv4vyN4R3F
W33RNpcY4kAMaDXXDnOJVrHORgBc8VkeCFrlwJ6jpRxMDmUJ/1DocM84pSznTwXD
bEEkwa7jN2XRlY/57ktpediry4hDXJId8TozN6bAVvP1UOcHBacbY5ZusS5VrAve
ZHLwoj5IIjHUtTs5ZHvpThmPA/C+ASNs3tZ18I8YOeK+WW2gjtlv4qYu/L3LyX+O
tlGv+/bpW7yjAXwhh8LOckKaWyuiP1jb/glyhP+KcjlvEhIg0SOytWUmEpsjsNig
g+He17iMfYuG2B/T4pRdFcpGJQTV7uZFkg+I4bj8zUJ33OzWm/Swzu+/gxCoNpJ2
jlpIauK5FrCYpdN10WXtFozUMEeExgUXtLgPoOWpl5awnHpgQxx7MMfY9rFzGi1q
+Lwbs+Kjd/8f7NDH+uEZZwukx82nJekxExrAENRE9TVW//yeha+DPtmIKqIGkcWS
Foz3MtiGjH21sxVhRIHBocEQl3JloOTLu4DWEfnN9InzBrnLafLFGDFJotfF286E
xtCupE7OKWvzn9tilkhrf9a8Ah40KTJxjJd29vlgUXe/okNDN+ut2VpOV3u/zKWM
MVlfT9ZHa8Tbb7Ka2sotMpNeTxOBQQsF8+CwlY5C03KD7PzUEuBU4DwEjlJdv/0W
YsTnpvSqrkF4Y/gnIEKSIugz1xODj9EoGleLUEhlewTGlRBK/qz31IsUCVumz6WQ
8LRNx95ChvIbc6Pc7shI3csX7EsmlkY6F2lr4NkH8sIV/5Fw6B/DofqWf7aYwo9o
epfsrOundlM/qbxE5Wkn4OudZCTNZrfFRUbT4BjCQBvs4T/OUiO/W0/neavEAqJf
3FHQHa0TsJ4oJJbJcVwIZWKsR0HJt5gRJrdKXtpP+wsdaO+MJT7M5fugNceiw1UG
itkhKMvBKVwnk7k2jPSYPcE1oRSblTrzNgDYBspZebnqZo4uugmh/WiJiEe3u1zB
a9D7mMZ0KDDOCJkFy0ya5+8C0TXmE/S8fUKaRnamSqHxmVuwxsy0FnF2TNSc+hmH
4fzRbg0sPKUnNbWg7lJW5qwEv7WauLkcWVJ3jd9Y15CyKDP0grB2nv088AA8i/vc
W/xnm7qoxiEUyBuw5Vfk9Pt4igueP6rwUx6ikCXYyxjevPjV9eINiFYcZXzUsGlY
DrH3DrasHWDQFADBAFniFwMrgBKIG8MTBngLTZZME3FGphNFJgrKPX3FgNO3nu3H
aPXNJfHms+6WWGlH06mh0QYcoKB+pligj62cM51XapnrZcWHdatrGW6CB7/lVPPw
Sd2VzwRriGoWTp6xBSJQBwmZmcy7GrCkszSTf9YLI8lqhExekxcJSEW2K5NAmR8c
/pS+RYdusrFkyam6xtpOLsZx1W1U3bhue/ZL4feOIo7sABZL42rh3ISzDaMWGUA8
ZYx+muTd1qV5c49b7jpnqtJEH126yLrZqpgB/svUQ8AghXYRjYYCtAKpl7ynLTwf
E5arfT8iQw7FCdhDpAZQSSzfaS5dmZa1LBP2waHsNwlgTXzMZhPuMZJyOOwXBAUx
oP1F+c83tzH+QKTbLTrVHRQfj+gGlQQHDW0UmYoOjSVv82j308biOk6bkShb5PA+
TuX84akMAyJMEnGeCfhG3SCZyOPysYVvkvHOMV1v2Swt/+0WrZhDV5RNp03Uo9cL
Wkk4peHPCMtZT2bV6b63YlKdRXfgi7ac+r4Ecu4reveYjuu9LB4Jax3iX372E7ry
v25Xk8GVRUGt3ITzsOTw846pUj6yPR4qZEDfDVKDyhzCSEa8KPv712ZUKBLVoEWt
Bk/nxCgSJAhtnLFrnSNEauE7lJdMvVFYyke+3F4tZ1zxyl2HV0QlUZKRODH+ksDt
+uMZMtLAHbUAprmUfIdVcnYy3RlDNXi6NHIJkllSC8q0WCZ8m7AwWr4j6b55kORT
epiXrrGfGJ0vxlKmqCY4qZ2dxurMivYi4PmqrVAKHFjtqON57VHQDU/0E75rJXif
tGA6k92m90OeCbK2U0tHMyYvrY33DCGR/H1ysSVRSxmW7vOEnB96JEkEqjLsELX8
54+DYELKwWwrHuxC+4uCdJJVLzSG0o5SqldiMvX7Bx0Hv8dOSrdrggI+fLdaQfy8
xyRUmpap/+K3eC/ZPYoNVEwhmkefyyYKu4GHalklFXXAEZ6nr8Yf0UfzpM0vYrO9
djfd2gKkw6gk42X0w+DxgC2XQO0Q21LtU5fvuAWANEndbpJsJGgNUQpp3rY7NExa
aYSKj3zT/wryg6dgykmCNlR7RWNbb+HmrnILE5YxoZl2WqT42T26/OECwUohQSSz
giQuLHcki7WkHqxDdYICnjzlpcDaT7nBbia1GZ025uGl97DiSHswhhJCRMYA6W18
xjcDA2HibNvnqHB9yjxy6VTAIxp/K+HznTBytP0oLdoCS4hjj77RSGyXzae0Kv+H
eKg6xMSmJ5qj+RjHnWiimpYS++YzJcatMi3+tu4/wWWsBj4vYWOGks9dbQoJNFGB
50usm2RDtFl69+gihf98Gq5yMoyCZTXFYRaw2vqsv3q0oxPgOmHQVlV5veQSQAYZ
wmQiGe53g23ZWvffGp+iwluA6pHd+edz1/LKzp9qQC19tWXIsKp61QPpUq++4GIh
q83dq5bHssBu4o0W711gRC72zKxrxUZb/zw+c0BuL0XjLgP0BVVNX/tqpC0CJsZd
mzpJPBZIsI6xlCWw4tFZAvzrtZkVnR7zmSBmwFlIOAieZY1/lWZYH9rshjFWEvos
x7LUg4BF3/LjEWsvaK5VFWOFlV967UAzrlnqYs8q1Nf19aMyHIQyaeckXODNN7lS
6VnJbX4ExVs8sAyrXjjRvvB+tn8gFMfQm1fiXYAS9eEExthi65UiFIZFI5fHIcSp
XxXoOY+r00lj8XzTnZqkxRgRqLJXoS/0VbrA6AvcbthTdHy89rdtaQPsAn8tRMA+
5KgPVUj/pLM9sLg+GMmGlLBKgqhVELwcTEmevD50l/VkAcIS6GrJ5VbygIaL9qam
+2JBLZu86mreUYRfC/lazlBG71u+pvuU4L16WsGxE0TU6+3Yj8Tn2C3+aXDXmEQP
WDdR75toEHiqLS4Hn29t1eVew98X8Xq5VrHoRF3Rt9r6D+a2D58oegOLxQQkHnYn
BNUBibYIWPHNZHVJ028KWKaJeVIjbF8iqnfTYyC6+AVRdhZb6kNTU2YcKj681N46
2+5vVrySFqiF8o3eg1fW7ZNeVRVYCrtya4bSHeAhBBdiOTaWTvJbp/CEJF4v6RQc
537dksxXxc6h00KwuTRXN1LDc/CbVzpCO3AjC4WxTpNrD3JsP6SP2Tsrr2li9ViT
rynlmYaGjTgxW07MT4sGneG00AmtcALnyVAGFP7k/FNkcKYc0YdLo+N0ctCeC/tD
dnqdAL7lD9kdwGeack7cje3OnfLV2h2W0VqkMO36S1N3b8X00SfDUIdpGsEz5F48
8HXGvYnZqS4CagNeXFL9W+788JpOXo+ge5m0oNCAjjW/73Nr3Zcmnb1zzZVPYvZD
DsZPdE0QoZAJbT5Ojw7Y0LML1hn1HGpnXUrKGYCn/ZgEHtHWpT/uak1WWK7pZLRD
kniPaN7Tmii4rqRPvL5Nlt0jeq+ob4NALqRrzhzaBVbgkLCA9NPrs3FvUws5G2mU
ppVWDsCVaa/+D0nLL6weXZLtaEXjf78oEzKXEiN1EAg77bxS3aRCvCpz/jtLe9py
eRYqYS2q0XpGrXhzpgDU10+RftlqRcx3RGsg57Nrs8dYV8noS/UuJcOB5rOMvdbD
u+9swULQEaQD+wNB7kEa9f+nTxCOslrsx3qDckxmiqgV3r1WGFdOvDeXfqqLpZdD
oxRaLu9ec5jBByWBCEcdQ8lMXwytF8uBamCBbnHJqmWrzX8jUkGTLt5z02+A2oPs
/MCkZYOa0nsHEYVQ5WeKlzEU62vWqPbJB4AN2EzZrOEJRS1WXlwlSTUBpTk9Pj7W
32MWpM37d4w+x/UBOpyRan6fCvIJAO/hqSmZuzve7wCH1eoq4DdOXz2ZXqqNMqy7
R0Uqtp0vcw4n2KTn1vEkcFoWjDdioVNCEvn4yb1xBFQxxqO5y4RWLGj81EVLAhvy
03xQEtRfbAkwG3Gk1I81vBx0KyXR4zHB+EvU5oIMnu8b0jmP9E3Klbbw0sIWXpvi
IDweRuMU1SHuVC1S4SyMaFFmRlawLD7aVMR+xkegZYKsrAEO2a0r02vRSWp5Skxj
4c8/4e7rGrHg5kOXliUrTxltpICCYDFRwTCa70bDyG5T04qiUPmIBeHodKIXNrU4
24h5hcCcms24LAmYhYWCelkCiywK/hHxHzjIy2PHOtMTe+miHgCRB4QTK+BHyZbH
NPeBMy+ze7anljTp8lhZaNW2hq06jQqAnuFRknB3JF1VK0CbE0pbnAmxD/Pw5rGj
+2EYCI12ul61t54FUgdL+spM0kLoSI0WAI9mlTSiYDSYDVg8Hk30/04KORWo/w+c
GgPh9ejvwfUeIeleIJPeoqCJT1ryAxxt2k69qOG9q00g0g2zR550hb8Re+Zl8W6D
KL0cjegR+yvMoFQpfpbXRcMue/TXwEq2PHeuGZjziwuCj+XdxVSQvraGHyU1YC5I
0UeH6wJGgxm4wkVIeowx62hDzW2rJDOLrYyVNpoQojsd0PVUWMFFi36+CrWbkjM5
WYywu/Q1DBnyJIulYO/XR64LWNZQ3zrw7IjliU1FTxvicwwLjU3nN5cF72PG0ZmF
l6BJNo2swfwCMmEANqVG2oz6zhtar4cQp0UdBfe9HuT3/6nZko0+bn0DQkz9hD7U
lj1llxKppfAVCIP8SXJXtkuVp9wiUoPvZwMiiigj76xn36LNYNal2NSlAeRlkNcn
+r+nDhp3JTHr+t+MzvrQJrr7ZRvxw2HHuceZkLLdqdGcNATxdhacUU+63AepouuK
JrUm3riWURk8h/EkDFHri1StBkSf7HSVdvtIMs0VUedWONEc1f0ci9wnVJPmWcwo
ErvGwQLFagUDgF4ItrjUsH4FSw5lxPsaBMNSEi5cQxl01V4vVbP8ETfmXjkOVwkf
2Xxeo+qLso1WdjXgtwFuXkwAJfeS7vsjMjLpTjcfYnrWP1Oe7es0aCklF9QtUTvI
soaxU01gXO1wtDaLj2R5l6ay0Jj/gE6x/h0BcyhFbuBfsyrL+OKYW8Ae7ZwvkfP3
ZxpxsG8s1NtQQs4yeI58VoQpHD6z+Zg1lHIsP1eqYb/Lq6BokpHu+D+eIFjr7CZJ
M5y4M2WoWcX9oZOTkwwqZt031ESfaLJjmzqKkYRe5ulGlwhN75zt4QdV6T8evqh2
BD767eYPNS+u7G3GNNPA7h72ATZ2z8/1fOWczQlN0b7gzZ4AnznS0CR4sueX7+ZO
Rbj+k15HDPCNC6AC6TNCkn0KIc1u7HCrNSIrVuJlWlhS04jvYx44HuC5DdR9drb8
bLrqk74l+IxNm/KVREcb/POD+OQVWHDk9rYqV8I5xIA7ma44m/1Qmd1+arbb83Py
6DnF4GVmqZZK08dmi8/RS1p5TNInNSGvcIYJ9KcJxl0=
--pragma protect end_data_block
--pragma protect digest_block
WxZHcGafHfkANdvm+o234rKjq9g=
--pragma protect end_digest_block
--pragma protect end_protected
