-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
4LF1eLcIQcI91Ru2MkPGDfnLE8kmb/1pLhxlHojk28Xje9j40thrPaJTLheyFAyP
OWt4QCIKaV4VQeVByP4sE9JRbePRm9VtXlEGobN0nhLH27iokpDI+QW7huRdCfV4
D5eK4dTxg0Kuv4l9qstuQnJwKbk8ZTmUdoFjydtkVf4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 30000)
`protect data_block
mW7bYflDIHWldSlKBNpkhl+v6ed7U5UGus0rbvv09OdWaWsUHXnaENxPoznOt56Q
VP5NX09+rHbpI9wc4yWCIgqT34j0Hz2o0Ya3He7KCHFoKw8ckXyuDuGABqudvmZW
FNs5wPFryZsBgnbzeOKPZEZ7DKCuKlVI+sCxhLw4Oy6lkNHl2gw1gXOdDG8oGvVE
OCEYztDRjS3s+NTJ7ZTxq9K6FUCnnWYf/lwhaNY4i/ktiKVGZGL912qeJvie5Lay
dBysJmiM8MwgwijXNwmkkGDJ3LXqgZij9w7PZ9/9omBTZNalE7+vC70YdGB0KUax
6/ziQqbOq6Lw/tQ18bEviDTZ7uQHE46OJ0uFFKU38NhLeUO3NMeainDV7pac8N2s
/fBZJOoNuc6o0iHRML/PPlPrK8ANp6YeyWYsN4JWIgEaYLQ3WljsyTGzQBgi+pAb
poMOvxTXaKWXhg9alt4Hs1clSS+KO8NbNFc55J10F7bgnZWsavtVZLf9tMlzecqe
8enLyt2KDgIG5R0G4CTOfADTXf62BI7i/ykpJaWygH/ekhO+/YSy40hWGszQt3G6
emrzlT6+7Qrd4HNMO9x2FznEhl2BzQamL7yuzsrZsFmu6ObsWUujJF9G2eVx4VEC
1zCPan94sl4hVvVEKu/Nm09eeQPPqp6vLNaFjBcIzz5hocHOeH7lS2h8kpmDfpma
Ah91SLytipR4Nc3hwrcHEA+3x7F/OuGvAMBdPT8j+YehApYuVyKui+au65GXsweL
T0sp66Jj4B2WmpIhMLqs7lByx/fqshUGfI6AnVOOSaqLNalOYKu1tIpMnbsk0NQN
NQjnZLZFMgzRWIVDvsnIn3lRvYSZ+DmNSgKUv5I60Yuou6BkLPZ8q45mCM8yNcny
E2xw4mFKukK6xtNeVMH8nCBqiIkU8nUOUwN/ChXPsJPjaUleweuuvj3kD6qQwY/J
ikXQfjDhAAj55R/aN4gVcxIQ/HrIO5TIHjMV5jx30+PJUgStA0XCO6b1MCeSRnzE
pg9xU33/oddQq13SHarcSIztmcVxeEvHGQXd8W37YaYLiWU1ApGIhT3b8qpSJurw
TfHjwy8pTZJrOCvwYcG82UgOU7RErGGPWLznK6yOv3kPdhu3Cebh2HI20neeeGW0
UrSes5HPZnElrEEtQ617x/dMmXIFQl/dTxtIK2396RHyeSjekwMkRm+cmKZwwwzu
4szOuM0N6PS2uZ3EqOb2TWX+i4cGySxfrGd9Tv6VOadu9FxvzvxkqkmOTxYbpTWC
GdmGLVrLszUMEbktlbQQ6sVCj9AMZUywqld5Xwf4XFpHy7p5/VcL0+FJ/0jLhMrI
ZV8SAtCLPbQ/31epKbGrWD+6AMnIxfGwgXbZgXKcWaz9kGOufJEBumraUSWyaVbM
VIwsBUVjXso3KMcFc7d0bvj9G6Hb3kgPt9SOhe4+jVUGM0XMlMtmN8Ud+GHYH4qR
GFBxQnqzp+52qgzuZj73KEJ21RjaYdevPnLaG6/1Wm0RZsif18cqqRpybiFDISWj
Yt0b10/G2H0R8LjI8Ss9XoxLIX853vk3JfF8pwf98/ogelQ9PyWwOMMCh1NiNYr2
ketkxXmfGcVq8FvrhDo7nwTEe6Ke/0hYwdAlG2eXfYGLLy1+6ZqCa/gXP0HNwkCz
lNvcwLsBO6YWiib0ebXsl2mJGvUy4RmU/jYDIaqgDzvT1AueWJ0ynoXubQc57TjV
WZeqDJsDBYLnaBw+LyD4V6GoFv406WyPjZvE56d3bAc7JJ+h1cf9OaVRFzsDYwQd
RiC213/0YC0aa2zw7XCkRRNs4n+csRyNQ3kz9kmIDv33Pz2OmK0TnxjoFOM/ag2p
8ownZhq5M8cWzMpuzjE1ztG7tpn5sw5gZYtWnUAV8DT+0ZN/bwWKx/FL5yd4ZZJ5
JLTTtXMDYTAnxQYphgdE7+KjVo3MwG5rD95IdpclKxPGeZW+ebbQHZF0hql/fwdR
yIoNOEuxtw07dGdKIvoq8+MniOY+qez3Tlgfrb1+ZYb7+MUBWXMXGa7wZK3NiHM4
M23k3hFWcM45OwPgxWkjWH0khZafCleDEdn+OxkuBFnGXyxfI3eYZ1A07ITsHezC
CloYEjpek8R+REcfdxRnlbPvHn0r38vh9kZ1R8D07CqkVqAO0JDQ9Cn2EIXMYJiy
74Y7G1fwteAW7WqMMwBan70ko650rkcngcvbIeeupZKbapi6lQ9MVXEo6wDhKC9R
OVZ9ktdiZ/EbTog23XbLCpHVGH49mj57bS5nlUOJBN8Mhr11bV2qRsrFpT6wxF9t
zmO9nq4LxXfo02coWt+dIwWAsyEbH9F3TkJuO48APQTyDCN5QHlMgkallEGeU3Jg
3XEBy49bvOXxpOuCqxirciDkwKBPK/yu53BVkhWQx312KhUPPklVIdiofd4pIav2
wajNJj0vERjGGLT8iFFCT285tWgZ+6I8Z+F6gkAMlNDqdkntV7rOUUGF0q/5Im4N
PFdjf4rkFS9JrdYJIZLiECBXFRt/FhJlnRvA0//MkclVSlC2BKAMd5h3m9bMqXwr
ZGAupRAPFoUCSFs2M4JX+i0jUiZfItXK8aSpUulRDZyHhYtzpg08KPbgOk7TT1oY
Rfiky4FbfEx9kExN53XujvkgOf+DeX1jcffAdGPVnfJE+chp39Pki0ewg0Xdzr3v
eozZ+YYkgbuq2BT5yEoYPlasJZDAjwFSQMbzzH1AmMztDJQDXhkqQzSmlC6mlkAU
72U4/S/J1yFqQsp5dQwlOdTPkhomsx2k1EsPwueGlV08p5zVCQc4ggEGi3ewVGjA
jPwYg7ESYX7Ia7MRZlcxkyRWnLaUoKdqpfI12i14mVoYd+Ceqc5/5/qXGMlLT+5E
C24Vn//TWK2ionrryOv0A87BTwaoTeg6lmhgjU1/KZN9qFkXTgcIxMFIarCwQ0jV
aeIsRtXmunN6Ns7zQykzp15nIUvfoJ9Ae4WaGsfsbIwksxbVAXXGIycZsGDakAqH
xCc3d8g/TcWuVUXaoRkzWmfMozj0vyufoFOHoCJ8Q/Egkze5Xgq8wO3wHG9qHx6F
GuXhEBxD1rh872ATqLz11Q4lNzGfBM1uG5PpIiYnT6wR0WIVwnQc2xi0FErKhEw7
U+Un2XOV/laGG9IBvFcNVlHt6Cgc4gc2zz7901wVJVJ+0pCzHgu+QnlzP0t3iZEp
RF6eRD99AInz5uVn0d1CHjkPg3zIFzeS6ZHBHej1NKhY4BbZBeU4ZjA4kEFbjOd5
XKi/28Y3LN1naKyMGO5LAXo1gx6Klg64xk+ms5THeV9rVeRxHuU4+bsg+lZj3gs5
kxbRPLu4dfmH/iW2KOuiWBKggQ8KEDfsxga2Q4oIOX3HcXQp+crkubMbFMyE8OmY
VqRxlF48rZSGpE8c0w2BMMtIyII4JP4xqX9GKNqX4nGNxc+2bqB9vvsMUGqnYQXg
bRL6lYYcWVUtdaL5l/P2NOIhjLr3E6MMQzPgV9Q7W43Gby1a2/iEb2FDkG198j0I
PhLOSD+NkPVjH7kbyqiXmZ6XpcB/WzI+PZF1RPTGhFzJxNdHNb3I3/dWYGm7ckRk
71gX4nO/XncLNpBz5iH204hZk3+wQarrKPd3exw1JgJx9e4vAX1EPBeskuU16X5q
IhMkWOjYbqXqlxvsCNnEEh+VY3IqVQ0+im2RgWvTe+eesIxr7NTPiQqN2h8O/Etd
sxgwJYEgpUuzVsPMP6PAuR1uBzRZBspluHxCEiVSmDAQgVn1lfALW2iROD35MS9b
s75O5E2GHV6puDBYpYAtArk9J5aqAFfMJrfbAVVpPu1/wG9rgeGSt3mq++usLrh0
ckmZt78OAGIjC6scRlrcpyDvSTkaC8OlYpPRch5WSz31oNTA281WUHuNsoNMPRVW
JmQKp/EM5T3by48VnN9DkJzFW89xTAnZPpkJHr+QwlQc5TA1ylZr0fdgYQ7KRjes
cRuHtTYuXOy1e+CjFkC9ZmetORUgfoWz7AD7DUXYlq2sXdjdqTjT+BlTUbOxu+N5
dfLU5Id3Sa5x2OlR+p4dRqnY67KUII6ojmCQsgvuow/ZUGF/e210JJJ521qTb8FL
wRebEoNfiynxG5Si0HrWNRDACvrqXcov85bc3jr6IS06MmKopcPtSDt82lOS0zMi
GSKcdXZqs+GROj3/nnlOg3zyImPJSqYWW0H1kRBA9CXNAK09S8+FNgM30rxgFf10
rle3VthBpCz5L5X8spHaaprKwxTHyYf2uy4EsiXdTFPOFDnM3LcaQMWAeRQWI/N9
tOiCng/p3hN99TbRdTxUHfyu3Fj+fgtwDN4lYrkllRNvTX5tcYo9+GjOTxJiHmBH
29QsT+8zfYIaXCq2voGHlC2Pv16NU+ySVprF4W4USPr0/n4j83lbIMjzM1doPxon
zi4ZY0CTmfXWthFoHadEYLJIN7Af6bDkCkoNBbO5MV5HSlVkamvNFgdllYYH2hCL
XfapE+Ru23ZV5Y2tFw4HO7vsgg3l3dEI0F1yzkb7KfkTV/NhgrqdDU56Klot1CMn
M280dJ5uQnNUY6GV3yIlTkX4OB05GIglfP2HPQ5lS8BZvSPx/UTnorCAjkMUhF+F
CdtQkHxxknXAiVseop4wYOXAbbpH3Czc7VknEVTOT2gdpktMG8IGTzrv4W8+HyhG
lFAZJNui7AGgSVDjd26OMlTjpZGW+NnVRqdIWL7H8rsrz4ZhXvZgRoREeunNky6t
fzeWrLLiDIefmxvs4f/kg6J6I1mpTiemrr6AFK4N72SJKqDjXYRzkXa1PTL3gHuX
QpKbbft8EJ1Xg2L9Kloq8e8BWad9V0TnH1dWW77dASt7Ys7ea16ifZ1JAYA1MKBF
wHA2R49uMWE5hKkzq++zZkpKfkADN++cAFmVlJ72WvFibEJUsF3jDzrhjuyti+fR
qISpMvfJ3iBEuuqWv0qdNgd0Kt0jRXhyyDklqyUzRRqr2UpMF4iYA3RFO7FEohI2
eHyWsdkhywWcxiZt5AbNw8wHYaCc9VUzYtoZZGoX0UfZtxGlt2tKncGjS9mDI9+o
wb+dYJm5XQaQhfp98u6tgU1ghjl+dKWdFCYmXLfwdbR0uCR/7rCBSENGFxjmQ2Xn
w6mMITDan4JKhTA9lhvcO0ZmOkqYGScQ0Oh+BDvYAiszOlbZDWNpGajVgjPOZ9Is
mmbe998kueezl0gWoQ/V+VaQvd5Q74yp/np4q0DHGlQmtw7AzFqxdasM1HUk0LDZ
nUsgV3/rh5H5Z/qBE9qbvouZDNkXBPsDnsulXOA1TZbmUKeyJGBcWy544VCHhhGm
KtMhb97m/kcbN1omVg71acyPswkTbPnxfdkx+1ASjaQOHwc2GUq7WvXp+OAEsc66
tHOBxAkKun52nVlzFRfnUwjRKom+eaaEPjT8/Xxo7Zd918tDYa+ke31ZcNFBsHWO
wX+f/YnB0LBQ+kH+eIGVMC9DKOGnoM5hdRNuH/ocYlkqnxr/V8ii1ywTm3JSEpiT
hp1GhmnrbLnXCSRTZz2IjQ30UoKpk+EdEBdPC71msr4TZf1gwBaTMtrAgJTfG71H
GhuB30fHzJ5Ys1RENzWTjVoYeTFzI++BuKL0Aq5zat20k6IddcDq4CkbvIZRplS6
ZH967KXuFnz0bYE6EvVU9bzX6gX8d+2XO2ZpAbbKRonzcxpjV8uF+NMQUucJs7NV
LZ4aFmjxAMyOj3ovR+xkvqDrLUl+VoNo2gg9fncER9tSHNBdyWqcUHBjmnPDhPKv
ayq2Hglk0BcCFBZIpJLF7PZbTd6M+1nskVL6Y8hUM4g6EDWEJ0X7tOGFzzb4jzE7
VuVUJ42bOehiEDxahgngUh9Gwu3uZezG2M28VWc7470KRE7ufpD6se5P6VDdRVnj
KaZeOjQiQoD7XB2/YDEYKiV4LuWS4wiBXypycs/dK8HeW5Huv9ph6JPy9fGIRrb2
gblS+Ngc+iCX1ek7VP1TJhxmQUoO+oLPQg3ZH2LelGyIm1a6nMXxGe46D4eEjqWT
/G31XSkpWLI7MCwBp3VGPa8MaQ4S9e4TjpOQ3HLYMIfHIeguf9T2FsYqr3Knm8Ll
fuD1UEjDcg+9uhm4QSifwS5wLzDR6o8gLNMwnAAEL4VWp2B+Jrs81jHVCaWmI45G
Q71Dqy9t+ygK97gXAQRVz+29QWXj9Ec8WWhncTxEI4oTnICA5nB0NodYhJy1XWjF
jAsX3+89rrasfqvc4F7q8zRL4txWb70/1ScGOr2eF0/dLh0dYJqDYFKmUB9js98Y
auaxZb1BEjkfumZboCxXuhXOu3Awh4C64WN4zsjx55kQX81xW6YvNwZKLk1pYqSs
OSbieAgwnzgvWWH8VkhY4G0/QSTODJIWArkWj9gK6+gz8W2IenKvYi2CJBCjD5Fz
d+3Bj0IVbtuppHz0xbN/zsOufxfhfuY+zy05DgeeAi3mE2yWFv9Tm/SV6zFr3s7V
kTzvBNMC0YGlNO4TEnWUrHgFQZkXh8XBqdJ6x1Di6iBZtpTd/UxJe+Uk429L6dkE
UtrjCLTX7dg354y/yjuQgf4BW3jwT3ZgCDV2jCdnn8SwK3Cjeqji25xQdIoA7tX/
e897DJ1ClgPI+HP13rtlWRW4zZK4SORrNzwI47LHcuh1tG6q57clSbmcQG//HTK0
+v4ShhGJgHBmxRE3/yXcSOo4UL3HDWIK8pk7X24GE0q2H/cHoRiBp0PaM8ptXSmm
tdS0AhwBFuhPfO39Pp6/RtF1FJIty1hgtmmoQ8xhRd8Nqgq/gBntuPiLwYKQCSGK
e9B3lZFOEMSInK/kSxJjK9+r6GWnGEXQNWfsHCeBaor2EXCDi4xB6dQnvsDi+MPt
u5OsfYQoyp1jqubHVBjsqCm5We2tOzmbToeKTAzs42QIVaYXmrTUfl2pt7ksoLcc
CviCLVmKeURoY0MgI6rdJU8c+8SS6xVz58WutcMfst/5jxHDac1Pi3dNI9GJbu2i
KIvvo8lgoxub310jD4Bvb/qoV8PD/pbK7VhwC+pV85niSoZ44BQ9siQYPzoSINg5
umQHGfccthpbbBTSM6iUDpQ6VXRFu4fsVET+Ujjpb5BN38RSiU3pxAvnHhdLeQM1
QXOqKsBDffpr6USZoKW1NUp6QiD5IHLXM4JPZip6EtyWg8PQouqROwiqfK1KUoR7
NfZuszWH2uJ+RNMJMtAwrv4rpt6OLfDMtRycgm4wBtZQcx4FUsAFSm+XZrV8Su2G
A6tULhVg2GVNNb5N53V6zyrMrGYMLlVXI+GlhkG8VxF/sb3JCx0jKCm2luDO5NAc
XHqiW1SUy4NqfRJ/enNRSTxVaVMDtUJJXEONkw8XZniPLCtDtvJBHuBjjUNvu92N
+ixq2ExHRb6rdSun5xXkvbo19OF2IbPY9UD+oEnu6ZRZEeueuX/WufnYG5DQtJqj
lpZ3HB6wM1mo/vlS2Ug9b9if1E2v+1obxKMxNs2GsvYV3B2BMkWLrHusxoEu7XEj
L76aIJ0k3lpX7F1bQywQMsP4ropa6/q9eEIY9H4pxqHno8Y/EsuLiw2FTbn2kxog
0yjfJwH1VDxh0k9JibMumQ9H6nUB4qLKwExh1tNnZvnIZN+9dOupc/y3fhnz9azk
LG+Q+XHKeOGZYnjAzC5pWBsTP5TfuQQ9zycs3TwOctME/Laa3SPTlSLEjDLYzoVJ
AMVRBMUSYgE6g5a1m2ytq3H0FbAnyudFK5xQh3JslhJDy8ngxpwwzr90UJPkvA0N
mW23hcXWb3b1BcOvkH0yjPzCAR15b9ovDqn6t8xRrOr+9Mj5JiXFNhn7kKEtlN48
O+xkUFaYjMCOb33gBhJm12qoHihHQRM+Z3Oa0F/cGFlojKf15n73zBnWy8VVdUMl
CiFzjNvVPhpCyaMrFnm7dz5Q6Xf06B9hxWI8trs03gAafxfyupUrqknxa8xBcoTL
tgrqpQDyMsALKEA+Bdjm/k39Jc7NrA4/Rh7VJlB8JTOzVhFMDBW8NGC1hZNBuZAv
t100XrBpvzy13CvgTWMj5nBhBrtzMSkWMLaCMO28eB510IfEQI2onSJhWxGhObFn
K1hYxy/eKFZ8sdna/LWz4aIb2FjF+L1ArCp6+l4xa1bnR0pB7zCHjH74b03OuJNm
0RyKe62CGZX2mehSFxm1So/7vdZU4QrSRuyC+vzzLeHXkWNaQr3asM4xZdZlOTX8
Tg7tCE4oRRKcONHVPyhbuNiLIUz8rAz96zRioVjAQ4mYlRDMG261IcidwjqeTY9a
GCAq7TnY4vboyIf7FKixApWUGr1J3JvNC0uobUIrPutdAuVOqGkbQwxAH/DGi16A
5/mhVoLqdlIGDSqQk8s78KYWWLSquqfYLfmX2ew/zaesRhctTj+CyxTLsPkO7SbA
H76Sb9PQfS/CIPoOMN7lPQ8M0V/Vk998OUFj9koy3oCYtaS30SN4u2I9wmPNO7Jt
pSfhORcbd87obphXfnncnO8ykXSmX8vjSjKv7qGNkfcl+t8IVkziNZ4CAp/9zUQD
IcJXaBI2/uS4g1zEi+q5oSP2aWVIu5we+L4QkNNqwFaYWCJGFu4gQyaXI3iiuEQQ
FHUZZmvEzaQ9DchvAAzCBLetaXDT8IYSkrOXpOZR4LJt9e2SbkTFu5pUmIKjPV2b
sA9XMAXOFviPJb4LQKlZhCiCUYy3Iiv6YZGVkxSVA8fZtDNRBoPes4Y4o+QS7E6v
N/nEpePCwanyj5J3A3DIHlXi5n1sxh0DsVyKYwz42rJDTQNTYEgHouc0Qqz9JmH4
cCiS+/LqsL7pc1vVNjVAilOYtgfi0s+ECVnRnnGFeVa9VPbpmVpY/MxYNorBlXRZ
CUNT24UNLDffLDfI6XrTCjjJT92NUECGIANVkZml6rHPK/zTutHFRYMhoyq+c3wp
172E03oBoFjW6clR4g2Rl4MtxLgLWLZYOUZ3nHS8kFRmUz0N2mjsODAlk/Bchu6j
+oJlfvSdgjJNSHBcEUq/tNajO2g0Lggwil5MQrWyr8TdLHiSTL/tKcA7yaIVqFBq
5exbU8rzVsQI61YUk2wKdShICgiF9WDrIRYISdpuicn+CuY6m9y3Ime7+a1h5Wya
OKFvZyxFD6vj14t0rSLQUdbItRvXrP4LIjl9dTJugtDpf9D/RL1+g9JxdHEFodb6
dCGYkn+GHrl7Df6TK8PhkNntRq0T2zEVxq7mvLP5w3XMcMsjSE9Mxosf30KFAZKu
hPvD94xmrXrVEhgBWeHsGQXna06X68EgPOKnpYpUNG1P/GuKZIrJHml2cTklmtCi
SrhsO2XgfyYohh5WtEc/UDZmtfyRj+QRr5WTv64jO19RBRuyT+OLzdKRYQDWX4wH
aMfd3Vz/zsAggbXY2JhPAQfPLWHkt0UhyHMBMtpdnt6/wPTywMpdUTGbDiWtptSL
oAbQ9KAUqBKgBLeL7Gqb4RdY8wI/liBo2wjYIq4gK8tSFB6sK8GCdqFkBfzjpZEe
/4YsJ0OdSr4AWLnLvahMhiqpfZ63jbAUDdEi/HS9o0jEBKLyX4I9/jNRLrKktI+L
ruGvOVn55ZJ+GKMzbkbBOvDbBa5we31/n/EjpkgsByWL/XXQI6M4n22yjI8VxoTm
CfQb74ZSz1I4Bqtj1oft+vljlFztRMuupX2E7KsZbbZEQ1FUg1m8fVGpgtoCF17M
41cUaAS0LNW6U8MjsxPg8ZREtV7DLeGBXsJcoKW5QT6cdzawKLhEICFXmBJcIK35
6agEqk1V4l+hghCh7TM/u1GnNonUkeXfFeTgnbwGstlVYrkKnDnmEzvr84MExL6k
02gbaSdRgJVI6eFtgaF1WiyjTTwQ/ZNcdmrCT68WuE6V8mUn32J6/oU1sYuoJKDh
nSghKgnSVGdbngbYdHTYODw+L8UG/ET2/rQUmrxGMZwnS3NJXpWfyvsJOCxcogJT
Bs3rYX5OgUOKp523LBe6ld+D6uRiHGHRM8mexyRT42b+FungZrtaTyUSzfteWThY
4oVSWH6Nr2g5IkrBvFOeT3su9d19xlgXH51RUWbcNeT2bH7e+Ak1Tw0mT28JZExw
z6pkWKlXxpyf4FOv/ppYg5iHvKwKLiPwu77rBkjK1uOQ3nqTcmqO4HC2JreUuO8P
Fd9dl9PRrRKhe/I9840TMKcJSDD18WYcK4USlSDxSR+v3zr/qCs2DzDnMP52biCI
14K65yVNScTu+coSA06ZiChuOrjGqJio8yGo5go+4Bj1M3ovy9h8QwH/VnIThaMt
0zgmq6JhJoP7TRg9K5UDt+88Oi6SDU2aqUV0SPG6BO8M3ESWTOq7U457b+pItep5
Iw3wQ8xuBBl8PJxRchUezxsJKhsB0cVMozjy04PlcIAzi7eb/xm6o6is5ZrllCZY
LkfFL4ystzyv/2qL6jSP0s79n5LNWE2YPnjDgshTE7sJ9ia98qJAfe6QFOV+YUaU
Qt0YTFnK1fbCsTcpQ9cw9mLQtHBhLBtJ1EsHSAfiIXtm8v1QCSslnvpn8V0BE94d
ARoyBVTOuw1tdY1DItRWwYE5eYoZhrpoH7aD+DwPGlVhkCAH7teEfiB4GJTOQBMe
LHs6tHWDu+yTTfXplAxeAXO50Oncf0wWFxZCpL6B3ZN6D2aShooxYWAqAzmPWeM4
evPnUr1GnN5KSgKkYx2dvsXPMe3fXsr05HoEOR5QAJisxTpBM4qbd/m70FDVqWuv
q2Ar3wC6dMnglJnLq9GVaaJ+/BqO7kmhcHKfPiijbiukWeiijAminiXuSHlllbQw
IsNUjg5disw5uejJM6vkBw1z5oiQ1WYfjv1LfveGTkXlA/OZ7mWcIxMhL3xbDAdL
25J9yuxUYlqZuVt4hSPr2zGs3cVvihC/AALnuTMsGcrB+qxBd22fy5liBarIZlwB
pz81HkGgMOzj0vq0Fh+LOiLXB8mpM0un10VKWA1nTo7bJZ8+wh3ekjMncbc+OO9H
2XobHRpc2ZIuCu684ICUoCstKhoTKWfUjk6svQsaVptp9gisfti4ivoI1nnuLY2H
OucwDF3b65JUh2Vp09uaHmyev2bX/sv04DzCDN+fHGgOoEAPXcEROHy1o+6VSi8N
ermdLH53R54AGXOSWjfhG2oAg8qUX4cc9BJG+KAOb37NeAOnW9XPd9uTvLa3tScR
5WwT4CisUbuKxet/oiKTNU1tnzpnwnzIOZ2+1iMUMsXP/h1ihY/4T21n/mF+kreC
coNlsSblD5+GEVeZLQA9I22RnVWPcA7T6RNPlTSB9y1grc28IqSITWLmRDclmCw7
3zKEUVyQsgAJlOJRLKGnmhB5l3zLwY9vQ7EAtT0SxzUI5oaG0rQwncXISY5hwQjc
NXPvSC4hS+/oH+t3zQT9GX/DCIKlVw2t6z1t7dlelPX/m0TC7OisumLkhJEX9BBY
5AT8SzhHAt9OdFhkTYzT5Zlz5KUzphxEARr1rmmdwmRcsND5J1fB+/lOjB9BYff/
+WvbBDfQHZi2phzMEAyRxztYgfWfZG5dVN8dxIupzeVlDOUnfFYOcv5JIYx8T410
ycvYhdTlcOsitNkG5oVxqXmKeKtPwZEWVqs7zyZhMG8PqjfsuoTl7oFMNpL/FoBH
saE5cmjGPv8VazFFqBPuzdqXJx3lzh2hkVC3BySyJTeKZwaUcKgQoFrNoja2zLYM
OimrUmcQo9Fdhn7lR3hmhVzoznyYm8oDlq3PugcMAZWYLSXZ/hrWK6V7j7EbwFLJ
NdSGrvBButMjWvhH3D3RYHaKvMb4lFx7X42nSUYX6dGwS2BTXG6YSkLrBwK3H7Fe
NmIMvR0vw8q4gNqfmblxZdBfkBFjTcv8MWpqdDpNHDlt+k0nu2JKz7jdpBZqJgA1
hZW1osz0J2gOiwycI7o3RPucMdclXvvMfhV/zgdNtXc5BxvfdJvYId287VtRqfYI
LX3F7uQ+K5XTZhXHRToK7HhocRMDsgUqpcH+uCrYgUWk3YDLmO6V80ORHigIu8vI
vLLY4UUW0KK1+DEYNlkTHA28Ik8OWJVRGs0ZKWaKoQPF/aOU1qJJjJOyBJg9v6xa
3+zIx2sRmJHYqeGz85wfZElN9nXRMctllWWtg35qQ7piHYh+WHndDF6ezmctUzvL
S2ThObX8+1RKDhYwHRBMqxK3xV35Y1+e71pZQixyCLskk5t6gvhZDZZhPJftbb18
4eIK22VMrnrqxbLDn0140cVHfnr+ChgT0n/tSLdWH1rykKHb6xkK1fkVOdBmmNBS
MgY+fl162HUJtjZXFE0IfhqwsMllB01681lULiO6I+ep3p8AYqo7lF8fdl/YrWHp
OaT9eApOWeBFxDNZ6nGkx95E6StkOKrUpMj3Qy2uy+ndSTWcP6EkSB3yWwgrc+CW
QU1dy327ygcDQJkVZ1rAS0lQtCw6lMXfoVGIsNQXxu6nGJm/N2dLq3pb6UhCwRwP
QOrxGe0Pkl7y32FKlygmpWdjyum2r3cdC7Whejk1etCDEVejWQ9zOg5rJIXLDHrB
RzkaJN1z0jPWFkSiDLv+TO8vUkOcRNWvZg9dVQ3AEhQhsU143fMZ890j8qw3uvk4
KBn5Uz52dXXFqiaTiljb1e+RDNt+NwO/XxPLRpwX5bkUk8KWQBBJmPXOZUZpbRLE
f14EcB/K8s4oXYOI6klznPqrV5wGb2PxhO6TmWS4FLosLEj66PTD77W+iNN80QI+
cJQe2bKYqbLxnSqFsdQcIhuW/f0ZFCKHZhmEBIo6cTe80vSsUNjYOKUnn0I2KPyO
n2wdETmldDsGoS9pGsjrOQoiP2yHJ3Avd4fNikAEyJvpDjsVvZczMFeoCXuVOw6D
tuGRSqYktMVd4sAk08zmXD0dyVGUoMHT4Fm452MPNqEtpSiv32zHauztwDCYHoJ6
FnEQob/PpekV/5YoiMR62btMrPs+b5B/4TBz9/Y6OdfoalMyVaoScZla1Dmi9WCd
ThI/xgM6s9KpAdyIB3CQAK1RqIRahj1aW9Wxp3ehQfT4Jq2YEZAbfMo2UD+Fzp47
z0tD9uu8P0eBjsLHU4glWK7mmap1MGDSBm4DMAYMRNhL4Yuy753BsbQu6CfIAxnF
sm5SNniPDg5ENe863oq0wqJK12+bc1ceBvxs/5fSyeYW8JVdDwoI1Dw6J0z6YuPt
9Kx9+JzZ+kGa+ilJdaLAuxcSnzLgIXm6jTXueQxW2yjbxGoPjMPfRrqW74W+jd0v
8ZxxlsIdmZvvIPhCLzdXltVPqLbrC3coCMfu2Wx/E7Qz00SrOpmRe+hCGrtGMuLo
2xOGyCsw/WXwkneYHtEe5ZJjv1oxlSUDBmNkPALhz7oGKROJheg5s9OKHGJizI/r
P0RED2L2crgY6OAG8KXlbKbfmd1NcREPSSdLgcw1Onz8Yc6qOO7Bo7xjArnXZ+l8
Q2JuI3Y0nuGG2aahacK3vIZh4gl5cjDsc8tcLgBpDjeEwH7Kq9D+qrPT4QP7uvcg
590k2CA7uvSLqTZG18HfeuJKAnG8hYfDzBUn22B13w4cKaTljjMQ46w6N3wAYYAd
FLFDQTCawXTNYCpany7JZkn1SQ/726cxyGeRFmNngyC4hzIgNyZGyv1RW8o9tnG+
FJ6oqVmi7oVchq9jIeLH8usfM8QYrXb2NEE+/4kDR+ER08l7Kc/9nu+p5gmaDI+D
+R9nQ9yB5khaq33YZoYBLGkxWr3vydgNPfGD05WHU3SS+5pZK+D/0UdIE3ypyBBR
A/hqM1kEVvbclG11+HdwUEK4VqZ9HSkX9diT9aqsYReTWoYBU2OEvkIomsiB4HPd
q+GS+Hyudu1l7/SErwYbqzh9DmbB2NKqeiB9My603/Ly42AcbXTpMT4YsuAy4tOM
47M7hQz1rYW7GldToK39/xHG8KDsgJRRgniQ7LAK1DLckSsXFpcVrvrqqXs1h7cA
im6FqC51NL2yH3i/7F1LAjSSRFbUmldm8nYBfbWiDKeNVOGhd+b0j6u3gEd0Hs2v
c0kkhUaqL/rTcKDAy6dnytwSMUSZEPEIGmE8uwmf/CZgzUIEgfVNYcuR1df00yUh
4SAV4lhww7kLVOG6AEePczhe0cVwo7Bj5INMInZK9J3oPlm4cbwK4z8AvChDFEBc
CLyo8hNhFchHI1uVIfzMacqMylE4hdJce26RNKSMpHCEusg87brTc2Jt19v/hWW8
OAj533Vexw0cwdx9Xycxmsg6LIYGwEZC2VdEhe+LBE8LJYdG26agOfOtTZAghlta
z61mCNkRvs1Zg0Ta6RgPp04d2sWCc+hcyzzRq+QT2+n9BYP4/9OIaBc94DAtwYfJ
yfmp9iYA7Xo0Baksxvr6wVUtJflUuOIEJ2z2FoydbbCn4Dv4zU74OiaMoRce0Pkh
I3eOEL46j08MvpvUHP3C19ElxdkPJkcHIbL1FevrZifM5F2i+zkvzLCmH+y+Tplq
V+NlA/AbB1QV7OmeIdm7X/f8My0FBLi5lj00mpLwUgzjJ4XYlOkvU5+zTnw2lmUo
kI1NdBot1V9+T3aXRuh0xWn22FT59V4ORAXaaR1V161V71Z2/euyt+OShCotnF//
qgJ02CTSAQWc6mzXUSI0EAItMhzTBShAnrdoRhYlG0J8s6Q3svf4afoPuWoS4yCj
SH0zK+Ac3+2ZKS5rb0QDRIvGVrIPlScKacXirOubhX0I8Xb9Jc4e7pdu9f7Btl/O
kk/woOYmJBkOB6eNWA+HizsbljRuMoHETMvj6dwF6MguR4i4x5BhwhDaAvDj9RYx
lSkXYx6WZs2QNRDPiMqmS/7uuubuJB71gzPk81sZJaIcmSrPns9fus7sfisIFgAv
5G3jKYK/nrpVUhhW7rB311rr4ZlE3488/yvhBDX9WHahpn7KWDl5Nzf7k8Z2wnka
wLnrTaCo5UwDgwJ5r5FHWu5QNu+Oq3+/5eqExbugHI1U1VoVj9o9CwesfusHiK+V
HlAmodsd2eyU2OAas1cpc7BJUHAHYKLT/Ik6pskkPxMPBy8USxPV670q5CHIIozd
fx3yJstiiOMRSpdIaGTGxFm4rrhWuX7L7kKfGZQRD0CR6YUZ0Kc1xlGcwFZlVLxh
ocFAK4CWuRs+Sn7L3kzMhgkNNCalxHNHlsuUV5R9VxRoBifb3Hyr5YNTKrCCylxF
6N5XEmiQm5Ao8E+RWrYHh0pw+uYj3KRqeuFDm3HBEbQSZsA5xAsOX+LLcTnyRUOo
oSSAwnuTy4L4kaBWNfsh2gNhPccFyw8o0LJmTuEHXlz3Th1yaK9+nW5dyzmk8CQe
BTSadxBuagqbkTzeZ6w5VvTCoD4ucJMfSrkOi1fUpk9SLU20AHDmM7hMrcl2LT+S
Vliuz8uXDMuIdLvKHfURaeCyZlQeBsON2idmHp+GvvNfMQOlwso8pmJ+cnPHxW24
C+K2h4iX/AvgllU4ohHLRWVJbpcZ8FT4xi0s0bEPYuB/dR/Fy3/c+nydiaJ2Y7Y7
Wg7hOKkD5EFSqh0bIpMOC8PoXDsPmN+/zOoe2xz7290wcyu9W1PESnPbHU0cqlgH
6xAHsc4GOxHfzdU2dGYitM7I3sYzgBadTBvyVv8qc3BmpbNOAtKNUuGen0JKd9Ao
J1hVC1k4TclvaNXzNFeloln5bEySVKe9Xtbnpl8h6fzRt+u2z0zyNj1NZuofsn/t
CHmoxtDYmY8tO1znXVUyY7KhORSwWe/XmeHwzTGZ8eAjljHqPmuZLF+Ql4S2qdca
uCFDdJf5bbDafrnXDvBcUVL2aexEF5LtLRTBWa6WC4DelD6yLw+vPMta2YKX71Od
CK7PkjyPbnE3pp6xzZZGwCHwBZn40XU1HKdcCuc7RJXpq4aSCm2QGNaAGzod9Mc9
7//b0Oh6eRK7KyZBKhpw8mf87SQSIiZXeBsd3CJFNaejBn4UvA9Oqy2NmQf6lq/Q
VNxePBb6R/0X2FOVo6BDdNV2JvwFYVnARN2NHGkV3aUWIc67K9Ft6c0iRQzY6j9V
HABHWA/FI2Lv+HeGprBOHJDVgnw7EuFmz3rIEK1l6pK2JETYxLpo58yO25RcFoR3
MyfPCGjLPdV6rjgJRerYQct7PvtCF48UfBdUTGhwELcVXf6d0VPVUwOeHhoPZSgc
hXwmoI6WLMGF8qaarXI6kiREHkLubMP91oL08GtGf+N9p6HWpd0HUmxv3+mMdAjM
HpMNk+3Plj8qB/EsuMV4SQTz0tnKHfetRHBd2DS1RiRbofA8PAuGqbZp1MQxm4Ot
Cfv8GGQ/Pbb8mPVOrgXKeTfu9c5Oj3AGayggTu7ovW970Ntc50+r2ott+Yhfnqzt
y1HtyoYNM1AuGwzozs5MfTfKWGMzl5vZjcwi8GQUEB6iWcdv8Pj4FiQf5AFJeEN/
2UCeWcWfzGF08gIRupkVq1l/sDMhahKHWoRLfmXGNXv0BBYegwq4ifp+y3HR76Ed
7b5o8XSKUy6LJgsA0GRBiLepg0ditv8w9MjEeXO1QiYrn4iDWEFN0nEtgGhMzUVu
Hc0nItK+IEX8HsP1odQS0LNbqYk6k4vbna7Z5n1EhdwKB9MndilZhnVmPbHByDg1
2edVI9ehfctLiZpUyxxkRDCChDItn5gW58+MQYzpmcQ7N5/WdxAhAkDACyZR/sEF
dSUx3cThtV6VyLwTVIzkKWdPduyKZv1Dy7BhmUZzQg8zMcL+GUl+YsmrGNb5BQ3n
7KzV7PwdHlaCkPdGSyqegGVtjYx5vmYA1vmQ7oeQrpUK/nQT6vuGlLQZgNpBPmpG
p+HzMttsIf3eq+oYMmhLZYxdiS27nu6rZFLw5wle6FEmMRsjmnGkqj2Fs5btE00C
HvLkIVGCxmyZwf8ilcjXTSAEPPmVpGkNWycxHq4c2DobgyDf4R0DgEk54HtY1KRm
o6KWiLYr1d25m+fO8ECruc/jpomPXXnN9t8u3MLqXYbicjQxhgIQ7B9Q2Nd78vH/
H3xniC5gxs/nXy585RfzywrUSFB1hsO75Sv7e5VQjKh6miWiwzfGfjDkGGqgcdnA
vhlrTsp5P02UzsRDyRkDGPFZDZKs37WAjEB+Yl+XBAl+hrzMn7Wdl7Qvt3TjEt8O
VD4sWSxoNN0l74UjEoRtU+Qp5oXDPKB3r4zwHrBkCLcLocgNVko9O0MktT+lCP42
OWa8Dr+PsHUdfkbc8aqsqZQNTURxbaKPQs3wTatTW9AbrHOZb4YMTgQZztC/LGYQ
16cxXRGj+tlyfE22fWFrXwDaZg5hWIGJpGSFrjsWjX9T41T2OehjnPq7FQNfGfIR
a2Ff2dZKxaR3ga4zG/rP8CH2rg5WdFfN2pp5mc9shuO5bKQAI2Tk5UR1gHvlqKK7
zfrBnmrj9Xsw7l80B8vZ257M4SUMJE5X2F8LXanmQ+H6xfNFEA1E3tO71rurpwgm
fHBV22WhMilkHABoe8qjeLeh986A59ikys4iHpkXuKkRlwxQzjuRPytxZ4pYl8hT
a7I//vwpIikB01DTD40iOE9OIZ8S/XbP51IIWoiBnVbHyWtmIMEriiHcidloqQfv
1EqkVcmzoLOaEuQGKrqHrB3x927SW4asgPk9iziaDwzlDlLea822KtGzsHAg2YGQ
oDOkmJ4voqnz+Uk6/oPdpo4QBYNE8EcHOQ+AMzGdUMRMU77Tl5y5aH33Z3JFkIuX
27zgn76fjUf9np71tasPTejZHFtHayALvcm2AjvpM60DeFDXDLdfFvnmiGo2Kz7c
qTgJZhGzZviAmUaS4/PuS0R853flVe0y6G2Jxi/VEVfVNRNAKTxD9xhcdpl8YvQn
i0i2tBDR6qv2K/m78lR1rblqG9trPU0ij1c4+opRRqhkekg2KTH11sPzQVrI2sbz
Cu35nK1X6/Y27s3yTxvlugcEg09HIB0bcTyiW476ihukl6MK+oVg6Mb7XJKopxag
+oVt21I1MKR3Ud7iUNOjwqYCCWLBgsYMvQaUhkAcDW4mLwhvr10OTR2+4OYtF/SQ
pwpSCXL5F9ixTO2N3IQLMmtRtaJgBghCB1slXwpYI+NrasuzDkb5uk6fb/SRTT0R
V9KkwHT62y+bBqfUq2UQdapjHNzMLWk6cIrHKYbk1E4QimR2IBwp+NzFoYn4CRQ7
LWHbYfRycl0NcXH5/fd/QTLPEKMruVOY34OuBfb4JAuKjPadl0VMeQbJmkbm1q4f
R+XtEKZ/Z9+S5RGuOyAv0AcrU4sAc1uyuk1XyW6HtJOJTULwBn/8hZmDzW4IoT3W
w/Nt2dcVmgGSvrl7m0UIrW8qWR7wAxfRuHk1twTnsROIGUyaWv0eE1uIux7/eUkI
ybyGUuAbAVfplchAg32721Taf/kS3CwRbA9d/1EPI5rrHR4iTZLBoCOr2uO+xpI5
KFXGidBayK4AA2OC+CuZeR8eECbWx+uZe8iCZ3nZ2WahBdfnJljWf93QFLGqKMgm
DXFpHQ78L+x1K9cmXAOvN1zqTk48bYt8yGfzTbmmAlPVV0htkPTNP0PwpqgQg3f8
xYotCeyzQ+qfkJg2VZYYtEc1REMT0GhjSlrfjg+RR6bL0g+7LHiOUwfPy8oC1Ym5
O1/epkDV4xoRjEWmhJwKyjlX62dtHmmz8quy6W9q16AghnVCKNO5Tz26k8mhNzDh
QIjfKCEHGVX8bcWWqyS7dr/MYQNwypT1pl1W0oquTm5ZYRvpIi8Mz3scZ4XDjMQU
xwVlb2EvAuXAQQU/dbDeHEK3bSHjLBqXa2NsV1NUvUg/u38rffIVHmLVeGrsGt2w
HFhkoMkNSFPV3jxk1Le92cde3JyKiC4c9LCcamVIyUv2DNT4vTXkP8GRvZPjc2m0
TNb4Pm9QLZwtHOFeFWwkt3LeJ/aHvfmwBQ+oQ4sLMmYUTQdin2SZGBld+LCPJsJ6
w/bHL+Y9Z7+1SbSXFiHOKDeaiLH15PwJLdFtApCRLa0C+qfyo9RuAoudSJx9TYKd
h+tungevENz0qtC7ruMcmQ4GpIvu4uandodnHaety0qtD/M4Xn3+Drkfs2EJF+ed
U003XcSJqHbAs+Eq2olCNleBkcvpP4Mw7cdUyV/ARLgJdv/EVzMbHk53sIR0I0py
exn4FyaaE01adhCscvDedQFhDBNCKXIQiAvqQr9pqTsQCGzISv9YvaDDQ2AJBAnC
YzBTVmgoTpEabNU0BsCPNElxWfTGRwqIeMOgbMUeHmUObeuoXijxxgu/zaUl/GFK
yOjmDWLpw2mAFsqAa1zKQ3+VrAoxU+bGBur/tEyThM8B6+P03AU/OaC1VKDjVb+s
wyd3+hMwth1EqfRdwE51PuE7bVcMO+EMSFiIFmsMuujzlyKhooXd9r2hPekPyld6
OOW2rZABgYVbUIj82V6wzYUNURLBEc7qCX9Wn4cIjaakLeIVm39OxhbHoLNh2LYT
0frJoxHiBSi6IFdgWyWE5/AbIu+xnt3hH8ukaVk97iSkGYtA2hrzC8Nch3tiOIHE
9OhD+TceE7iLOrXeTj2JL7fKAuESxvnwxNl9f3mc9Zyikm4XI0sMeA3jP/1GBkmQ
HWFDk4grV1yOqHo6sv76DgpTS4PJAlKaq9jmNnYtjqeUmb+OcldIV1k496Z+5Dn/
IG+lC3nLwp8F60A+/iqlM9D1uCLDRLurnyIlBXC1siAXp4nLCMsgFYq3nIi8jB03
JQ/ZaqNAEwzPzVGZtCMKWEWq8GCRdsxSU/dCyiPHBTmWVtIO6eNEHKvO2PuEdDsd
0NYLa6a2k+SdQ5zJgdF6tEMaZgjTK4MFrZDOStrVQAB8gnm0FZm1m36sIwbeXrYp
bmvEKfbv0U4gIeVD9rOJyzMuzgtzBSHuIjJBF9UmTrZpKhCTbXQ0eU2fJXFbH5ZL
rrmTMZSFlc9KxzczI8xugb5mGLsRjWzrxb+B1tN4+M9sgLeR1BrFjcjcdPKINIBF
oxJy5LNEiE9UxJf9Qz+PUmZ3bjJAacVnn01TkAc7l9RzDVSmXVpAoEt3XFNooJG9
HhdpCzdTWOqfMQ/huNaYjsEmzrFBvV4PhQ8TlLe/+ysk5CfTlmf6bDjCOBSPGcYw
HB3MCORlQggJBTn7kMnv327jlaquS4/DdiZ5/G5aXp081LLEeREYCaEqnV4cEi09
qyVd3+Msfxj03AhFy2EZ4q6ji8Pim70Yh+ZQ112not9Sz3IrbwagwToZYthmMQUh
5lxm0TS9sgpzTDaDe9mt+oQrlIIfizRITFPugCzT7I4VSo90bW1LNpWDk5PDYhdv
azGNkmwo2mrAoUhWFXZIf71VcApTCkIFwUVAYecbmQYYzeM0G5xRcK9yyKdKvSst
8IY5KuM8q7VSrkhYdvUocpiC76gcTuP7GZmfyoGsPYvCB4rDI/Fo3RckUoHFzTED
zuuKyxXKARnOktW+V3w648BWBAbJQPDy7+eH5XPqacB1qIO3oq61Fz2x4ByRaKMk
ngOvLxEOoeSgL9VMdmZSNvmq+yNgADA0qk5SUOLIwCot5GsuSRsJWFaWnWjVRBYq
W/3qKYQTZkM0SmF8hU0cRYjdQbUIiyRorDwY/63hsuY4NmeM/5p+SVGZjc72eOt9
8kAwc7vVRCslZL26x++peDsdQFxH/MO5ybvOGa/339iH2h2d7KOwTPvGrWFsn0FZ
KlpY3pNiN5roC+BXd2z+rOIn9z3ryh44JsBLRYwl9/HWoCOL3Sfl0wvFzP0Nso34
LfjQpjIpCaeH+uMPoQfrx7UbM9ReY/9mhoDWEjA7WK3iR7hfMcsyfzifqwr/UPKy
M1MSX3BeTO1VkA1WFyzZypPTLWu9C2Gjk17lMT1zUyT0w//qIAGzSXJNDX5M9vZa
GFKx2BLhoLe2paYHFE3hxfu3Y7YD2RbX0lpcI0dRPnZMh19Jthcj/rJi9YySxfqH
+SZk4WaFsCfN/0j3U4oGn2qzmUnCafn+zFma96d/aW2Xh97QOpYStzGi1JWvK0gE
NsVBFrioClSxEygrPvdUZOFL2tt8XC76+qTVzpPOJFU3im+rfEZlXikGHnoihu12
7l+wK2xPZlftrfl1l+S7yACohiNkdv9TQBw8QORknhHmRZKXoii/d/mYLJ2CFgBS
hjND2BNXj7oA05x3O5ghU8v9k8ddVIFFiMqebZEp++bSGrl2+FoHftnKXF4Ldj6U
1XmlDwuuG0+MMBrW1opzBWa5XQNM4V0uCTtc4SsIvnG4blhuh7E715WN5PAxOry8
gYmL8B4ypSbZUCjQG/UHzMsJhP1Ss94gYN8v2oa/JrXgymPZEzrmZgnGEoxHK52Y
RuDJ1LyEzc8yOIFPYTvk1Rz9M3CjNhbq8ArbmFNxg4/95K2m1vEayXWRGaBi7NrY
525mdOyVcHlt9Yxyfgrx88qJ2544OHfA57MmFplAXVnewml0CydzkF2cJZjrplo1
mZTwAv5hVTWgzZB9YzBXdK2Ipx/ieRfveM316LZUZTvr7ngfolqiiDzHBhPf45SL
7AoCPBTxis6h3qScqKLgvyj/RnkTh/SE1FY6Lfv+WKFSkC5LFevM2z4CULjqaUJD
nBxCBv+Zy/cst/E3/9xLaSTA4bzLPobhnjc3/JEjSMccHW6Gg00dCIuEGnEbDe1L
ZP/oNK+4/vAKOLsPW8p1fbweXfjQ7Sx9D3reDSuA6sVXU51JqjRlZFkgO1AGc32j
NpU+J4WjfERXHCEB2Q3XsXT2KFl64YOUFzwRJpHN+BQJ76z3Od0+aTE8xTjmPNph
KsZZgxQpD0LvLshex7wbhg46RVil4xcmOJAycGflIZLoqyr+OUZC+F4adUaTvKjl
RW63DmtfNmHBujdJckDarAUVH3eAOAMIqvZYh44qwvOLMTyc8plWxfkvgyWDnyIm
FW3u/JxwhGpHg/vjkruQ5j0P3aj20Fqjx8ASiBxaUQrivg5hwVy13W/ZdXsyPXPM
je0J8NdkVR/++2Da59kEG716O5o4RvrQekZRbvAXCFbrbTl3eM9IOIOEshNQW60p
uGVydaDgncWilQ9ARFQMR94oaxJqgWQBUREgYmMxTz9JoRmFDWhQDUl4jILD1l9T
ahvogZDFQ4iM7LkiI23CDv3vcYVVvFWv+/zkesd3J+BW0WNNgraw5KWXhGN3EyDV
gUUfeb6fK3lh6SgvFSyDOfSp/tAHcn+ARSWnI0mwL8ACxdlP3cQT+jbeLKaY/xvn
tiYuJWdLKVKbs/R+cmvmUMcMWEabZnitgRe/gJnEGId5BqiFRqaJmyaM8IJ1nIS1
KqJCXKZdO0J/HJMBCnHrAdMwpyfbAv2jZ9gRMSiPOtTw3xqiOurz3ok8sK5upBOM
N+iIJwGd0BIA4PLWdXN38Co4BtSTlRZTzNl8SH2GwVK/9/gPlZ1sbRJwtf8xIkyA
ndA9tp+u1UnWaZvJsYsO8LccA3ADhBx+e3+oYPyHA1Ef086XALbo/stChbrdaIEM
oIA+QDgsg16TItnqw/7YfZ9FTakp81Uo+n3kpTPH5zeGDEVjdPwyvr44OEvnIjcP
Lr86Tf5hYqzH9unvr/S7GvBnF+VGjTzIB42bsviN7GIoVCi4SdKomhQB+T9HSmxi
hsoN9tzm5WIYNXI4LMfdJAK3lI8NkcEdhVog5TG6YUSuTbKDty3NG7q8RvX2PNLW
RvfnNrcrtkq7uMdGh+g37U6ZjYaQ6A+TZrNWzaRh/HA7sH8g4pqUUJdPU3v4eMVq
o9WonO/gqtLTujpD3mBumYb+IcUC/cpGKwvM2AZ6/5gRtD/mYyf9wcg1Ybc4dbY+
9DLsqXFEPlZcVUhHNjtMtvbrNPZ8wd4b2KWESZrcUG5zxQxWgrUMjrsCfgGpMpBM
vpf3s8OGv8io1BRXJyacJqpxy6M0JzwdOQtsED0OGwYfNiI8JoutPul3ov90HDxS
Mez8VONsCmwYBHAEtqC0eKgG2Za2etB+KWM5vEXEI9jmdJGgPI3xVPCA9kXsPPrm
9yZOlciAJ5piS11E/lSzisOCEDkI/Q6ZSAc+THmDrAT7fhnT/PKA8BdxwZh9FCwa
ZZlNYgJ+AYoYP8Rt4B9Z7qQ9RQSoghFafD5VIMpivqGBmRlDnlzlrCXCmwB0oUyx
19BzUnjyDap8QB683zIXIi5g7/USa6fQxUDD82h0iQquJLu831jHD/C/v8sSeoNo
0II9bhPzjc3GGO0kbwf/ThZb4Jo3bfWJgWs5D8Qod6i8aXbMpmjbWIv2nCRkB45D
GWI6iec8KMPXYblyPKJyHBTtyomjB2AuKdOUNsCizlBGJdYpyXbyaX+L8bxtCIDi
kIZvp1bMLSex2tA2dB+1vWDZWMh6A8AEWl7YuDz/T+W3+GwBbPcUDWnYqKuBLJze
+ims/X637hYfCJwOjLj78RLRljK+ITbMUuyHGW2ii4NfF2A3wiPY65DV/h5Ix7FE
xacEmMENL6HQBPbRMzsKLnRHaPXnvIsDzNdgKVnovRJNMWxmcJTtsXTc6muUqhbb
RHdtbiaU7fc3wjlO2HVtsQHpiYCfrLulSFtG0bPpxjK2leCdw9Nzv6ub66CxhnhE
CGTk0KNKpElefVKPx3pPptqD8XiQ92TlPFMTGZpWKdDL33bCLHW+gl8KNhrFBrLO
J+sHxS6MP9JrfqVhjepncbxR33QAQIKm2pT9dl2kYvbA2Nvt/l5TjYZBjQ/+Yp/6
/VAXP/B+RxQkMg15xLfwpfbo0eN1L34tc3oR2Tp51Nx8eInFa3xVrdpgDwheU0cu
pSmNAA8LUeN52tv5NCOJp5Xcbv6nywmZBeK9Fgo3Tquk/keUWfrBiu6BIMrC1kSs
hi4dHv90uBwESsnZ7zF6H/cot3Rzb5kmzHArrSgZx+QpmT2eDs4ahCtWzdSJ+/fO
vBO7ZjRDUl/0L0ZwgL6tBmEWTrAWETgeRm1Uq1RrjlsgclaTrTqRTcRg+VbxMxwU
wq8Ac1V3JLrB8AluigdbohjSBMnGt7nCmYjoOAaRdKH6c+PY82sSLw8TocATkslB
fA8F3DvRhai8o8MWilzKjYNJOvVsdGs2KJOCSQxmWpEOLmAP1t8O8JVIKkDAgLfB
BANzKF7aFQYBsnqWPCBcI4cmL+y75NNFkld0FO3ldtoWJu/W5i7F0x/ba0D6TVJl
VvUybrWl8ja/2SPV4pVo8utmjj4uFkJnbpDV9rZtlcQ9zvG/7ut+brLIT5rlj1YY
MKvUHAaugucDSLd8sDalHYm7hsAMg0u6XN52AY1R7eMPQZslV7IyVFwXRwUSELXx
h3iRwH4GEX0nRgLGgl/5AyO0qjsL6Hf0ImvUefG9xkAbj0C6u/vKfNVJzIJCyF3c
JBkAtryOSzN3chI3FKfPCIPtfGNXNwXCOnjnuC2s+V/ueu8koqetlusyV+5bqgji
NM7Ir7gLQ2jfKBxjNVZMoDRaQuii3Q8dJBhWMb1k60MI4PrTkGMlr123V0EHvK07
cRJd7hObR5/j4BmPciw1g8RMPM+vGzWmd3NY9dFdpTF7T9Olm8ZmYnufCnqCMi6p
UjZn/e97z60TcI4DTx6/9fsrq1X9IiVWO0XCqYicDqttrsFn3BgVoGlhtECt4QFZ
cZtyB86QqgWg11Zc4UfQzsu9UjFURXVCTU9mn91LAUcTh5Ttw5BsygZm03MRgAum
9R0GnvOPwJCQ8GJ10VNBNeLrBLXZ7inU3QpSNYStbFhMxFv1vNpBX/vEt0SRTU77
yYJppY/4WeVSTLuyApdeqN0Sf6QRPuBuW5xVWUp8+dRmS2tck8wI+dcvMI7z/gg9
YtZk1EMER1ikR5/1IfawUFSJz1jKG47NZVYGYUGPoa0aeWyjW3rSpZniMQ2vWVmj
EBLhRs9OPkrTo70fJGO/63siKPj7x0COu7wljvf75AZqsqeq1QCrgrJNJ21jNxXY
uTya4jz4kUBzSAHregzjdfPQeeGsYQRg46gHEbndWx1JhVct1rQtG826o6z01x0r
GDFDFRQUEy6OleuBxoXfKPNSFaHSKpJNx8HPbfHlDI8+EsXCirXVpI3SSabNHI4a
MF/6Va4h7Qhe/3Bybaskfh+peoRlN2nduCEPVn74Egk38+5XLaj+NUorcpRPT8zn
S/IOj0FkjWhxoFB/fc3aibMi98maFEyXNKXV39bC6nrWrZUADlVrgSqz9S2/cNkL
YceUZmj6uC0HlwYEM02Dgsgq9eVwvZo+5covIrzofjdfOiH6L0m8t7OJOKcRqXR1
h4nhLhfXA+AYIzSirQvHp/v1xdspi4phYjPFphhKx3wAWQQXm3RZQ4pDi++4qRwr
P7EUDkusc1YsdD+7Gpaqk6WAo+Bhs+QdQNLfyjOUfzEoRZTNVeSZYNrqwY4RDrtK
bWdZ+8S1fkPJTjNiwnw6l9Y7VbUv+9CFnu+y0XWj/XN3M/YJpIOqpvenieBzaqNk
aLte0LJU4LSLp/j3S3ZI7VX8yC/Cl5KT0x+wePFwG0EqeMlRtVdAZgazr3AzE7zq
9F1XS79jwLrYvfXeSS1BGiXWbveYW6aDdt5PKs7cOYRz5281QQxBPNGxD18wm2r8
nbT655CKBwtDsFfrXV9NdgGSPRa/J6eCMLdaapqDEe/3h7g2RV/anjujuuc0zjeD
kVPyftnySoGkv9t2/cyCZdhyowHnaLDUYi4j/VWGH8iR8GqTJNrYPrIn2xEhDPob
E18H0sQ0OpE8K49R6btuLnRrQkAtatsg6/tXPilRiiqbVpOUFq8ou6hz5PMtV46l
UWUqp/mofctyV05PwAPFS2qK3hoBvCNpUCNpeJrXvmHOhf6XmWNw24rLj8jCYUEM
fuiB8pZehUEbon9N43vLVAWovdlAA9OwMuL3zCAr9VPvA7yRKBjB+zSpaYkygv0k
ri3nahkt3LX85Mta2fX02Bad0n0cu1pc4gcOrRKzUsYoyIwmZOsRLDztanAC9Z1s
7gCC0Py8Vpa1jBn3cVO67WChQt7rXmvTDXITwFHhHfeIPTTrq38ToFEadzEGAhzs
sQdRrAYfNznjSIlPG9jAR5iltGy1K7OlbTzf1m1knsK6lQNWoXukPdoVAuBHbWXQ
AuUhMTX8Xymwlkw3YBi171owV4zuJbmNcl+T7iqRzSD+VPYerCgQAOmkR8ixqKCM
FmlUm0e+TtJVPCrkDEfgT36+kpr5fRffGkGaYqRFu7qg44CutooO2pbb9r0S8zpr
JZikWEc+oADL8RqNSEgFN2ABqAnJDlseTtAZ7eXQTm2JvPhjUNZ3Zi5PxkZ1mamT
xI+gIC+9YhwUSKfw5t/fDYKAVgdWYl5BJgjueZKHSfdwdlkS/biex+tkbW/+3LZH
EbiPAWeKIJCJZpTMV9NOoiW1wLx9LV07RoS7XhvB50qj0n0juFOJ0PCosP17EUGv
HzOD2XL1OFkWzzZjrU+34FyAtTbhuUhoMcthYKW/KQmZQlbmr359VDPQSLD5NNHV
vbPmZUaxATNk9HgXOcqdtEIEWdeVcrdD4xYdRH2CwPCnCOA01X4q8S95M3ocxgTN
h46v74D6BYv/5aAjbX9xPog7rPcaIDN6xwuHHBTE0+KVTjQ3ZN8MmEROgLLXCK06
5SlqKJDmXTBZb6GC8QnfQYNWydlkCxY56jUVY62c+bB/IuHSRhR+lIReRskhgNnN
o0NOJQDGOuJQ/qOswj9Jhc8jklqtQK1Bmcfc1fpMlVBFAoSTMFF5evUpyD7lP1Vp
Z4wgiU35oaBpW3wme53HokuIvQDejcjuUh8ZUgHGqbYdbfzYAt9PxLh3nl6BowdO
8Xhk201Wv3G1D6PxmanrYzAlzNb6lP8gB1MzSzgAf1mTNN8Fg18VOb24bYaJBMop
LxiHJkzpwQ4QbuMIVujEmhK0Dw0uhza5g4i5IeU+DMaf4p5U0F6x0BaGsmNshmru
+GMUUoskyIo2DB+YEkeaz5XmmAoj4fSR4Z1GB8oak21uCcejhD6Fu2H44ibrDd0k
3eq2jzgpeHF+784Cly/J2vUjSscY1UU5bKAF/CezB/yWnjFVdmGdWV8OzE2t6zQ/
BF1/QffxKMlzPW79oXyRAeHUNPz6YSzspIgEPvJNDjsqe2wXnwGV/x62qakt327U
Q9ZM+jKmCmeyaXyj5E8ZItwMhDVhfyWsghKcjh0EP3wFas0UmSklP2TJ9c6tDDfm
X4ZVhO3OCBJsi1C88089wZBEWuM1GM1q/TENDfPqYQkZXtvXoUL4b7N5LcpL1bZy
KXkxoGJofqc6h3sSR4iXMQhRqPXE8PG0rWRQgsUdTZNEDxqRhmkaQbp6snc0AyVf
Jx1KP6+5dc2SaG+TGYqBMnWOjI9k3Qc3NdU1i14c4EXX6UkcLkWRBV0ibs+yGa2n
Qc+GwPCnncOdjFRAPZqILz1k4d5TEgc21SCbjJObI6HB6Hdlay4dYvtmomsjJCbh
hbhP6g9QtBROsUw+Qk0hgMEbX6rmoxOa4uFGBALMDMLFqayc9mQc0pFONU5B3q0h
kSoAsLoZJ2oEuhHwYuXlBKiPVfoOoIfWg9OGUblMgyfZkWezP2tOKTUPexjL15VB
x/5x3tki+1ZNVSTfvg9FKM5C2/jw8Uax/YPqOQ90t1E+906EBa62sJNPK55me8lu
13x2a8qUY0xSAqdwAgBc0CuYXYpgCpwaUqMjxCyN0aYmdjuy7Zdp5vdazTFvmd20
RgOfXIGOP4hWoUnpwtWWUgQSmbJC/xCFDA/WUgQ1icsikOYIf9hKvGxUp8OmvK1k
yqVK0W1j4qROh43gxvb7SBglBhoxSVlW9QKvQXFC8sODryaA2EWK7Wqbhonsew/T
9giDN9ZN+6aVLDwIGRsao70TQWzmgHMHozXKonvYT+zgJqsIBUKb5eOSjsM0uG/U
bjH45ywU0/gRgwvCXCwew7KEKHa7QSKpR82FTQuOw/vlvBho78wiMdFTdZBciO4N
VudBUgpR/CFILGslYlJUujIaXPPOt8eeJBzjLoJT9xwsBAklbOP5qBVjcn/AtIO/
/12MnGTfQh3hGjd48uRkdSuks9N3kePmt3x0jypCyoLDPOq/RX//Mehi9gh7Rvqn
0+zbh1Cz9ux1sA0In8fPj6KQKY22a2RAcGGvW5aXI/1oUh2cZm5fwgYOXijzk8em
UaXdezOSU6iYPTUtH0QL80cxXtKcD4Xk/8nj2VR1LWX3JKZfgJGez7RL0fbm+5kU
aB93V5mrdRWnc5mjlNCpKSVZJyR4LLamRhjof284jrzBrXtOzVcJwlE4OEqEbRxa
YdmIfeWIYh4eGyzh27LHx2MUZiJXa9bOjBArl4SnPtsmC6D65eZ3YcFRqKeBcJ8R
NZSduS9tNbGv0qG/6j049K8JRO6m4H4Kv5CDUu7JSmAWgnYxfMTBig/LVysIOvJv
qDB/aJwkr5sSbExj5HnSNDzsVTC0bltKHGLeqi9D3j5YaaF7XQ2eJZ7MLf0xYRdd
5GD0VjhFZcAhptFpX1oC8gniigfNUp4QL7su8rGIuPCyGk81XjMmw+RUAqkI58WJ
uby9EwxRG/AVj7nyMr3c7M6buqYKE0Z3+zK5VmmBzx+T982F4njg3m6jH8WLVfoY
5zJ0c7VPoxKBntecDUHIi7bTud0KVDVfSlXSLN3KgvtCAa13YehSISXoi3kKYRlC
6YVQBFz8Uud6CCABTLYsD/cptsGwLMPMHufTBo3s7IWLpE4Hy92cRiUEGWpAI8I4
4CsuJ8WkZrUyUDHScyj+ALWxSCLFxNg2xhFcKZwgu3x5h2Sxinq8YCE2ju2NVV1M
WXEcrRHhntQceGEnBKDziTLgFmqy9FAH57qkHUSYaKj/FS4cTrintTHaoT+5EHKm
GhV08IVkWtujuOErstCetFt3OoiI6itfTrpt7b+uUYyukcch3fZYRcR+Q0HWnMB2
uCUYeLvJkes6FODEVqVHXtTtSFVFKeHEkSB5yh4pec2viqNtbB12VvbglJXj27KY
xb6zCXe8mFuF8rBVNyTgD+BawDBTIrwZPqdhsFwg8uoQIx2XIBc8Ph79wPFspNpT
SnLvutWVUdNM+Ro9aNu080WzT9nZhuYfxmu+dGITSk3LTfpbY0HsrbkqvW60Wltb
SgOLD9c3bauQC2i3ZFQSixlBsW0kKAa8zlC3rYBdowxCPZSo35LajKeCrydiNqw4
oVqFBPwtK8F1iksjR9jYVdGb9ycZAHgmadtNNfy68TfjwAPupU88/Bfll2hAt/ZL
xzcbBXDps/9QOX0Y0rS4cYaY0cXOwJk2abGaia5K/5yUcvhLZa1EbgC3alqs1VRi
Z18FtEf1L+crfyPqjm6k3c/vc9WXDwWDh4SS4NcmWTqkovBlRrCf5VFgGmVILGaz
ozNDHoD8SCx6iJVFl7BTdfVhFFdsfFBejYUIa5dcTp82UhNieTO1DAkWkLR/ENnk
9GpK14acvx78Mv5N4UKzmJR/oDXZ4n5xLlzhGqUG67SboioWY1NGm6KNNZLsMjlF
EsF1AaHhGSRtZ9lY+wArx+hfvEI4Dj7+v90AhUkg98dE2TySM/kyd6ZkXqoM4GMr
oomt3E/j0OzKc4QrN6Bqzxvb2u6se220JsshHhMnAOAVlXjxhup/Xd/gJAus52YC
RYhMiLgpGtvS7K/C6ccr0klkz84znTA6JuXiX+jKBkddl5jvW0DGukcF4D8ir6dx
VeEMO3VxFuwW7mi93x5sTn+Z6sOT2pgWVH7eZIvoG16YSp4eD6q60+Y4nFIKczus
WvganCuS9SqjwT2RgfjE5hH+FupPro6LqHHA9G6QeLamjIPHhVak9ydQK6vteUmv
H7aiF4eCUZltNsaNApKZ7graBZ8JV3/6oRxZGCCCivwTJ14APRi8KthL/dX6ygby
4rNOwhWoukDfG1tfp6udLigdYkvR+Gl7kaOgTVnXMkp4uPcFIrhY2AgZjJC4e2l6
A0w1WnyiBf+9XW1HxGWqqZ72I3/5J4xBR/fRHZBm0ZbtbEcf9BX/9fUZEhtpTkZY
jHhZzwwjPoEw5ecE9AOp8FspH8ULtP0WNTPiBe56OGgirOq8phv3oyGXvzO4OrgB
B01NoSf7bp9XoQI/M9aDn4oh8gvUSBKXxngCziVPAi642NPvfYjVxcV4mKkIRSG+
MomgbkRbLme84vplXOrBLv1RyH/L1ObhtxoZko592O2jRTSLkV/Ol6eAzJeWUlkU
+yjlEDXjOUN8IxYj7H0NBHH0X5eR/d7eAU7p0brIuGtGbwEKhlVyV+sc+Zvn/8RL
lxJIpZCQRbN9lfdKvvNYmCElsEIDDjDhLD123tUsraLVujpjMHq1c/K18l/0DGUN
NBqZBizrVnVgZIPzjV8kgOhS1reFvp+B2rh/XZXgwu73qiHZxDj4CDZEs0Ir3YvP
dGRjkIX6Q9jB5NGgJqjfVApXZ3VGu4flM/GNdPYgCq0RijMwUW4iGby7dr5mFm7s
2dO85zHztHmbj6FCkYKQiBwDqnOY4EOPXxQhlBllJH289trKdzDBYUYJDWxjmFi0
EgXVipfj9uZGenU/xsu7g2U3QjnZli2lrHcAIG1pqd6FmZocoRH94yZBkgVQ3FmV
aqfti5BdUd5drXT5F8RVSmmZj2t9ouv/g6rclyy9biAB9smSW6uBvHjF4DD0BagI
QlFs8MPtBmtSCmalV45dypWYdlMkb8ZWLPpr5A35Tc20/Ncd8ENWCqs7hioylLYB
jZJheUrI4D97rQ1tX9lwagj9tQOw0naQXS3ZKUk8H6Y1uVr5w++JJ83GHf3aPkxq
RtNWnFm2U6T2mWIo6bTiF6Q/I9JMl93O0LRW5422HV7T7dxhgwEpG9fx0uSWSBRH
K5Gmf5boG9n3imIMj+DworV8qPEsqNs7l4nyObfitxJOKCWkEeqH3ocVcrGtQfvb
iT5Og38GtSTHhdrOobhFqQ21I+vvIrjNgB5Nh1Kutg6IA8lVH6BGYcCipRXgpfGX
hfcfFRpumhk+Uw6SVSW2y6FgH1yZy+y1G43L12MS8RaM7OHwieBG6AGAn11prj7J
3YKOXjU6EbWnxoPRxIb6oy2IRmhTlW6O27ZkHOOa9VVP4/MCGFgKytLbIIQOj+0a
VJh10MnYy/PblPeHqThE5E1k7AWR5aC9iBAHfgdZ+O3bOACKM9Gsh9h/Bo8u+EKq
vmGv7Ggz9DovdVgY1QaOgCLdKSI+tdH7ZuEGE5hsKoArPQWqKx0xRsebqWFuHP5m
AnJQVO1ZmWyODYEQpIFEkO4iq8+1AzxY4LSiHgF1+xExZayd7v5S/7GSWlVKUYYX
cdlPsUeCeoRmlviYzmfjcQ20mZlnm2rRyw8YDhw0bdtJn+TQ7GdBwDQaSI23PdkN
zugjV8e8sJKq9y8V+9lPY5YlFTTk+ieFevLpgbITVw7/CVTCZJ8WyfNygLqzmDau
v6uBeO0vSUt/LkRJWt1tWCIY8QALsUDf06ipuRmAVZ6Y6PnnYCiPETLTNe0DWXCZ
NR0O0+VkntzhkU5LvTdSTIQ5yDBLB1pFAQc+dGjWtIczUPufxm7AYVivqvmUhF5t
Xhb0Nbl9nHifN157uiQ1nutpF+KUSC99jC0bZGUaqLi7wahULTwN0FJcpU9PBTFi
ftjcEQxCAdJKUkBa7vStXsldozUR+o5OoR4jiBFKdUhkPhk4c9rX1p4EJk4IW/85
TC4Uo8TAbMB2Oz3MNf+9KJozJieVuFxboeCEkiS+HmMdokKrsjO9xl51rXiSDJlf
4cARvbAYTltS1ae1W8RXP3WTxsiO8bFnyPDBrQBM5So/a/U4y0DddFO6jflvo/eh
8SBEXFwqJVV1B/4dpizxtiAyIN2eb30z+yATg9Ch7FXAMC2Nk1JbfDAwOKp2koMP
sSoCctoUcoMPnaF7P+I+cDPnyoWK8WlE/Dxj3UTuBmW2qVDd30RSfwFmsDzKnHwF
rkU3WCdbS1UBN2RJDobYEiSKi0lYBhnjc56+gzrwiMDemln6NbelhzxhWwu9OvfF
3p6+BtWrc7GhlRX3iJDJ1lNH2f8hfF0G8D5KmY6K515L7zryeszbXblqY2U1FaFI
vVPYR+v1XunTl5Cm6IqjcUWbVRIumuvcZlNC8hpLO3s5gPmpUYz5AETbNQYKS8fd
XUJtbrIZGUm2rQ0dZUueh21GDme9bwWchgrKZ6KBskda91+LSuOijFOq6zNPgLj9
zhRQdJl185qduQhRVc9hXn/jpXxZ5Nd2dPoLgiDzyM9i5HxX5os8ce5zUp7nwpG8
vsBcZxV7Z1CCkzIwg/6QY4I0mbmWsZqeBAoEXCH6AKLFVNMcigKNPBjk2bN0Tvb1
Zr8rNCBPCbuFiFhATnqaddcNQlPzmKRAOjkajCW5Vts3pRLcghNHN4n8CLiKWrfx
pocuiiQ7BjCpfZl1tWiXCiB1rYxBo9FUnpYv9+Bbx7tx0TfG+OUO3ibYNZ2wrpxJ
n1p9MThiLJEBl6JSd00v95s/tt6Rlc0NzNkgMMyEPUeAjrZ2mbo9L/L8pOZZx91c
yHoU1ci/aoAIYBuvxAgPav+n6+Sp7Nx5dhuRZF6pm2mVSexO8Z9KOdz5npSDPOvG
LX0hzAawZazKF/5Bik6NVxpgxfHh6SiN4FknkSmj0FD8fwMtsRbxwbKZDqsNyx8H
u8c919+N9my9Yc5Ocg3EwCDwUCMHy4yz1RfgeFtM/vmPKomvcVDOV4JaOwxjJC9g
SrlzPDBkAdC4wanJHlj/mu/K6Q6q5iEAYVckGwuFO8RhfFKc7b+dLGGk/Z9yDWyE
6rF5BYCgeZMhLuhfdi0wFRlwF5pvki0sn655eoFX9K9xWLN0DX8tutbj1zNfQZgd
OJ+wDMaaxHTbfF4E1HDI8TzGrQF2FXivbPtVMoSb7CcZiy9CsO/mdGVZiN47t5uT
H9lRTxaXhlrp+OKMqfvYRLcKNkNbXvHusCAYn+kYEKEqP4rKlz7WHiyB37+GHLtQ
slTs/Yqae6g4eVDEzw5aVx5v4wOtH9oykV0nChrxStXtTQTZghpRZ7xbbiOh3xDr
HAITozRNzVGNbz6emgmu8GeOXTuuO1Eo6x9Pd5N5BYwknhSmBkr8ypGorgMGI3Y5
nJHyIR9Qubk0vwEJtH9znvcVqFK236EPv7uKE5Cc7OXC3PukN/ygiRXhpE9qyyz2
ftxgAZ1kTelgFU3LEUJxZKixqxNcTPMge8dUKRUV4R9REdQ9u3ICe5AO0onf+kjw
W5780xnhVCXiTh7NvgxMA+FnysZklTKyqX94agUVt6bYxdiSsONYXkBkao8K3kw6
CZFhC/Jlu+eBDw3CdiQ5G3ewvO7jxRwcJoIivm9E9uXo9vLHRFVx5zoqM1GM774a
8bo0EuM/dzZ0OaWDuejOJ43NA/wYLaj6zkyyaKExnbslKix0ACL/aZOHi7PeqInu
8cSnIx9JII/8MvPqS7uzF388sbPTuAL8UuSmawYhCIUJ33jmYWe0TH4UcQmMFAjF
E17BsyVO56idsybtlGtkZw2EE765LBPYsNFg7uWRJKESXnjo8F632zWQ2k4s5+td
mjCKRut27RGoDI/m0imLC0h0cO5weFcGtT1mV+LV17lFlsnTUL7ZcRfgN4P7RWyd
j8aEDvQN7WYX8qaEGtiazfEslcI1lJUbpLC+3cPtyPMMPWoh6L//46mYnHQW2ZmR
DlOygd0AFzVIom0onknKNo1EkT1VYLiWGh9YjHAO6PxbD2Xf0VbaNjFpPc33L461
U5HI3mLGr6bEXaqHL5lzLmZuQJTaIW+jKnU0P/kJwfuFlGrygVXLj5aeXEy0+1sT
1HtJsp6i7V8ffgojPXlmE+t5QYM+Z8qI9p4CovXBlBxMWtluga0MOueGvWMtKhMe
qCnDuWktaqAcqkZCc4OFb9pfOKClqBaHLEKl8JwhVDn+rpnbE6VMB2NDl7V2HTF8
4AArRv0MQ5pvyF7D9mnNlCmNaUdePCj5TR4ChMh9Ub8IT36gy7ij2TvpcZJ03Thr
ldCZ8b9K1jt+X3p3+qQdGZDw51F9i0WWvVH26Ij+iJUvNfbMkr2madlkjcCvXbvJ
IHuZLrecfkjLjYYSCQqe1kxq5/wmSgGyCpiA1ZM6PlMbebm9z7XtMCfhKhywTFOF
/5z7MXjMou/1CaHcwRnBAkS1fZShZwq11vZtGfjO17KBABG1YFnRuifokdNzkfM/
Vk7BjHmnXjbP6vOy+Gx19EbU+EaHeIoYw4R/of9tctvY4OwQOlZgMsH/QNpSJsQV
HWg56K9c8PGxnySzxbWard9VHuP/OM92sKR++2f5EA3Okov+/E9RmGC/fMjtiUMb
0aRFOrrWmsgSkG2IihHyyDghoCsSN+iJzJ86L96W1qo4yGQPqx7QGB8MwyOm2vnL
m6ZUxZC6rKMQzfC9znhSKDyLa3BqyE+P/jORnHO4OYxGTyPAyp9vqCG4OOC7vSCZ
EWmPkOoXAqUff+Oj9w2Ck8wKkNWeehXilwc/3GRQoocVaS0MgwuCjDHv6tV08mR4
AABhf3D3Q7yuSzP4vhgCQGyR5z0I9nnMgSvfg1L0OFrifZfmjG/LSyMZhv8NxzPP
uI05m6FCXCtWK/wvFl6prs/kpHRBUNE4eJSLAv1FnW3nuu9AVs3dh2/3SgV4CHvu
fhkNZO9gPfPPYLjP5P5VI/264Hz4BwHaCSyjM7Jk+bP+3EGhKeR/xirm3BAzsjw6
AZ6ZVA6rd+tV+7acEh42bZ1eOwkIb+jcVH6yMOBNEQwZyHCAotdthK1h91/FaSWn
nHUnHHvW+vxK3fL1Loj7DaNMxyjD2oQq9HGBQKLdCoyGWRGc0TrOc6vqEbK7wOZ6
0IVC9Htp+xPyedwk/iIINjuueB+kIM8AiVxUK0UcRO1+UcutUTnCH6GIVu6uIh7e
CmLSIwk4jNgAmNzqrrc4k5z7aLW2jN6NAWUyR09ufouJDLvETyaDr9kExWaWD24+
fRc2eFQErBJIAQ3cnKk5L7DTQN1WN4hLkubH2GP29ZhOw/h2eStd7F69vMaIwJVu
DDhSA70rVvgNf1Liz71u9WXHMBIbwfTN8LiXHHpjW2yf7o08pHWumnBXc5bz7fYT
bi26ifrVW5dPwLzLMMxvdDAA+6WGIi5NZ7z19ny/TXYwtw5CizBSPyICuqeBvYq3
eDpbyrv5TH2Z1lpJ3ZoiEhKm0YdB9qOBxA1hkIljnkF5OtZdDSxTwsZxnzFUdPwI
2Q240dyTyOB+eJ7ExMrOsow9QA3TvSZhylmHOHGUtcrMn3vBtEUdj0ITP4nS5tpY
TB/0cfTSPb743v+d7JUmJRBQT7CfJ8RmR5B71pcsgCZ0ls6ZpZmJ7bwTDyFoaaWK
pma/3y8iL1/8NpQs011FAFr+iUndzqMcrUUQC+U3DVvXoOq0naOOTi1KzaHSr52f
b9Dg5qymn2IqQ9ynuHvrcJEjf6JIUds1xBHlQscANTW2lSZShnVa9bE24MpEHgOR
UvUovZSKgpt65WHIJrXSnORu8IMyh764neVMAlu8pvkQuC6RX7abqn4tvdivz8sm
fTr+0eCb1YRCVfxmJEyy6Adpg9ItUQyECPz02GSmg1op8nR5IlCf2NwqVbyK34OG
7zTu22eHu2GNxeTecMUByr4Est7qHzffxHVtSxnuCu+MD3CXOVJDtJKKnVfWyeJH
1NXD05gKGVDsrlpgayf1YBnz9qIC5uELgWabLWMIbQRo3H/XL4RboP8jaXr4LZ+Y
YDO8qCvib2jCh592WwVFbMDpIQAPUzj6y/4LNMYgwuGaLuDnZ0G1otmhVQuRR8sx
cp4enummVLVNpbdI+FVb/k3QPf8NCLKr9pDBBeSHsqqCHWlsIKoybdQJsgG8iJca
uTldh2EoJ8FWfbLDJp5+CgvU+wLPMvzw4UEP7KJHo/p8TIe0mvxtifHu9iqxcgwB
1dPLgbFo8RIA8Ks4qjDKtGPkv/qUwETmpW76rua1h9QgWV8GYEgXoI91fqQ+JekO
VuKdk3k/OjY88nSORi9mOrPDGTrzlnBYqQXd8gch1D66qxhX2jzqcPRVxhndj9Ka
65LJ6vvjmthmrnK3tvgw0DDrwhvQ7gKZX+20ORX+FQMI0XJOeZjAJ29ItR+ZX8Xz
Lmv2Z51IfPUh6dfZ5+I3RLfcTxwnhKThG54fzdox8n3ireWY0LZE00bbEEGnenwq
7Dc/gO4K99sgeYaxSFaUEfwG4mrE2WyfulKOE+61WzMSU8bOvBy6r2Lh7LLbmguo
MKK7ol/HPY9+iXJfgA+B+VupWwvyP+p5YCW2pJnlKzoNzllK1l3ipNl4Ac/fsEPL
HnGDTiXGiJJjkdYvxjOS/n+P4axVeJv2jwxsk4nwiihm+QDqQ5dy5Q0bEHcMxhJf
0iVYP8EXx8k1ymg84X4COW6o2qPWDUCJ/8wl0f4a3229cUGfss0kHvdtSIdeeeTF
Kge1ZHfnfO7NttZ7R06HUY9jcdoGuhXGUIJy9+x4CCd3hgpAp0SJUbKpp6OBncfg
7S+wYrCjKegFxVbchZnEvgBYgWjKpLaMOE0jrLs9uiw4srVYiBzybHuMRUuWfAaS
8cA/WTBmMh029ZjjUBx9CyT76O/YifJ+9AzKVMdWfFDRf1Cel1yeXhXgOSYKb06y
+9IZRFLUWeGE56XgvgaZIjA2bMGZenWT3Q57vR8krodk4SHe2qz4GAByHuL+4j2v
eO4qF4CbHA+a4o/kJDOm3Y8eHlVuwHVYetuEfNfqPrT8J1yazVYoXJaMF+8kNEsF
SfvD5x0aDaFs/dluEmE/v3rYyC1Xxe27rI96/Pi44HJFpsRN8qwImb/XcGmLUHZd
y6uXMGGd8ZILLybaa6SDg8iIFIXYqJSe93MpBnWGWZpgQlocD9dqHsKx9sxA7YWP
uzQ0PN4vmLSoXB6TBWkrFI0mYjUsioIyWLsr6YCmrcB3lwOFcXXHw8IV2jMduFbJ
gR10yncyxFfV8aN/4sAmVKDE1PNuZJrLjuwlCHc5EA7nj7hOz87nnXeT3msGRFdC
LCljc+dce45yHkjLFeBSsscSEXn0l+K+u17Q/yuaWBoHbUvqFgGQIiF6N5ou2mOq
PTmyTd4hxlbkVZcLSQxM5M78mVgWySCriltAfiA8xtXFKlDl/VPdFmN8FtP028/b
l3ubgegB9tEfUD6d5Q2PBlMPkY8gsChVYvpR4vzZB+guWYF21OhkMl+sqcONvfDB
BpXaphH1wcb5T6oF+XwFjP+re5oVxLb9nFwn2RXRzDPSyxMPrTuJpIfiBIa+IH8c
P9X94Ydj1h40K0Ol82X+kgL126D+8GF/m9Ro6j2n9G9n9+zejQuwLXRlsuSebPxl
hd1k8eBW+gBMtbbnnXrdHIbpGxN00z5ZN42CXhfk2Z5t0zt8mbVVca+7y75275f/
UWq5/Q2b4DlMKpbW2oUFr+HuwNK/bg79QheCpXVmmZ/f6WuUZJpkkqnJ/U3boaiU
8ebesOpYDj7kLkdmvLrIJF1GKz7GwjyvQi80JFQZ8dEWOibj6rgX2v8AKyHz1UiB
CWGUj9kdRuK4QDZobraRUFoWvXfWDxYcY6XTFIpAHSfB2qWURNslaPzVPwWzmKbA
1adRrvdV5p+BcB6kMa2mtx5hqf94TkJccdwC4/jtR7DZYjf7dqGszk5PPLirCa7s
Q//EIvOM4ujeRGjyLhx1j1EUcOz/Xx2khqHiKnSz+JDhCqiW8M39E/Urn9MiRbLc
rVml6ir6hzPNwxGRMNjdL+iDaOavDbFQheBs4sf0RuLC9qkNCv025/q0BsKHtZbF
cQfMj+uRmx+VItOhv5odCcqudKt1/406fIzRDk9bIdcuC3BoSlnL1lNcCp5WmJWM
zQCjvIKW3MYl3VyIEFO8qkyodGCzUZXWrmi9a1EnSrgTA1MmD2w5aEcN8hdXTLoY
bnRDfDtIlgvvJBjldbtlkex/ACWxe1yfvpjy1DsKvlO16H7P00YQ5W0CHWAuJn+a
a2AI3B75htbGHVhbpaiCy9WoAWmAjhRJhpbqKOIYOD04+oA9mW58Xto1H+y+k5Au
d4YTFFb00RB6kHcGSq1ojsQ5vgnvdt2Xgtiex60dtA/vYcTThF6F+0l1CnBVcSRx
UlFD/G++GkpAMBQ38Kl7a3FD8iJrKumjozvwrTc+s16zIk4WqhDeUm1Ws+4dn8+s
6F/3HCQFSGWRPbRDiO4pvcpsC7M6e5QopNP2Z1Njro883At1yrKkka26t+g+KFJL
meBlAF92v/hrgtmz72xd+hYWpfdFM1xVUIwfOylshxyxJ5qIdSrF6oHn3ubbx9uh
fpBNr22RslzONSnL2BlcTf9z1ESMUQYgs9HqBT+l7isHKuQjgaq4KrufQVPkKDS9
F/wJq2xNQ0MWzevCjPZYCV4tbndE+UaT/FyCsCnIHMI88WbzXxfWGnxlxs3TFsyq
x844iJ0FsKcnQrYtKip8TqK+I8rUdh8gxMVg1LG2SbOJyKEk1Gd/ul1qI0Za6jWc
STgNvir1woRn1Not//g00UfIVPb6xoNPpDvMz5UTmkdPcb5lQ5T/MdGxgc5nDnUD
f5Brfx3iGt/jF9YJdWCZGIWkZGPHL4ci6yw8p87Y0Jv4zk4HP42qcIieowZlHojJ
tfcGqV/C449EHTSYcFouKT3bPzHK9Vrztz/BPSyM9j3OiCpSkZCQlWmNCkAH25+l
wqlDTl1qrVCCYxnahH3PdKZnnL/3N611aTSKyfKkMHpOrimzgXHWN+C32eOdXhQd
QYcecMMOHb+lSaeYMcmBVRHHwf3l8osXQOCFMoKZ3keOCT15sX5PCDgsyHoJno2J
eIk3jl1sK2qB6FAo000DhScJLMF/G6a/hf2UFPgisWm83RrCb9P7/Yd68SufL9hb
iNg7dtBCndUyJ5HuR8cNYi1df/Cf4xt1Am8YBd6SVeJx2+qwwO4uOid8K0F4bCuJ
Bu0GUOi3HdeyTFJY0lHfd26ug7max6MQ+LHM9290Z8b1svmkmIYZo3RwBM66L8W7
ljxJgk9Vzgfgrk/kDkQ3QH/r1WEOnJY/eHGZtwbZmUTwAkVu4Ap07SNHG38MIrmB
Gx84tPQsANMR+7Hq8cGq+DDUNM009xB9wYiFo3rhNlFpVo4DNNTlIJzeUBnwNeCO
yRN+iV/StUP38cCtFTUhtFkeIfotFWB7XwiEVrJptpQmX0gbHrVUk1q4pUhB4IBb
o8Rwp5Gl/NfCOQIuP/s3Nc4FVIL/5atPReoG+Jolv/oIu6u63PIj1J73AtITUCJ+
+CuUUO6DyZ9/yHXkFhXAaTrl0viNcN7nLZxH/z9zlawYgVuj2ovOKTTA9gQGfzHO
dYUgKbVlTC71i+zKz2A9Q/w87/YWQsWqtBuPrRysXmDDvIpSRkz9WpLZODMm6guv
hD1oQKOxxdEw16vRe/M7W/MXw2E4dVCAcrRvuXhpmQwA+qheNtdybOsBGdX9+zEx
JeRSI9OdzaEXWrvzgthWwMM+d+4gZfWxEip6oHrcXT2bQLra0IDfogzrtLLf8GGU
FpFeSktozTM7GAQXiBoa0uveqKGw9R1gR41LFIKoexbI957RbP2woGouY6QNVfLP
lFQE1NAMAz1Y3IhbXLddMXtbsSbMYHhzJL6bBjFkUpTFiTXkxQnuIFghMo5Iy5t4
uP0p4ArlLSp4OvaKdwoLxIq2VLMFLm6bXGu1xvAeGLdmGSs1EJhOyxvX2GV1xneq
FRDjF6k/6mXqnlXOl8CD9D5WBS9+tRjHjwmFy3A8sKWvwXsPvmuJkUYUPcOG97hv
KPUdLLOIeby5rWjBNPhuhhBgB2LefqBVdY/PrOWhur+Hb5nX158QdGqYq9/de89t
n4W0UGsEvEjoTc9oSWZT/Nhc4+UzqSM80Im2dDvg5ihEFfUFpOnyHBzEDY5VEFl1
vGPmsuSsjiI2OQs9xsM6ceQRk57iYIKPe5ry16pNDPE1eeUdMnO/hSIeS4iUjcCy
CaWQdZl0C34MpGPq/dj1tceWDVhFUFk+wBVHEzImKK1ON2vJ4dBOEqkv1FabN61F
+Wm92rEcOVrC2t21Z7jSZ+rhffKCHCgW5n6ZqxsUcVjw2Vl3Q0nZTkJER4LNA3c6
6x+BhXV7xgSDQCwHD1MP1sUIM+8OEt7lxiqYBy7rbz6yYZfABqE/Vk5jz9ujfoSL
IInVcZktPIEg+fSRqQ+DamDz1Sn/vb4s2dk5Dg3XaqznRH3dXQSTk/1sgSzbZWCA
`protect end_protected
