-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
RwkWBHbv1ELkvLemXWjCFrSwp48etfbPANNZ0CFmOwMIE9rDEYuyaED0qvpFNy1O
nez7hZ47BLuNhGomxl0ThZK7vVRly9UafwxnpEJFViJO5Y0OR31wpNN381/Evli8
C4geW7b/B2AbTewvvs6ZABVl7SWMMlLv4ThkEIHbZx4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 1661)

`protect DATA_BLOCK
mwchXOS3He6PgqynSKdxAp0yKv3kln7KjFasIGGpt/fI+hbusUkawP/YuklyYJ78
mAOqrANz/IqDz1Z1hjgwNqNgQLBdKo047G1viwYEq/aNLVHRB/5Z9ADKexr22e1W
WSBlJSsnPoSaVHMrwMcASU9H+9Ov2mVp51qgWVzoTLrzi4GJ6DvNdhRYm+AwO56E
9GKWINHHSltk8y7bJzSGwML9ztBhp/GakCMVVOJ6ODSmu49IsJjizwVQdqkZsd2j
2QWqjMW8u0gFvURdovqKoYanqrgifKSkT5iOe4r568Dl0Nar1LHqIhibkWgytr7R
YhlbTStU59HKFZfEDlOxjaja27w47JJyTf/qkSewirRB7A7UcpED7PHoU6JWsjcq
LFrQe0O0EVv37IwubRau0UaKoW9MsUixnERZGQPV0xAs8ER64JvXMjRMW8vf43u6
HV0qD/Bv31eOEsKNjmN/x1awir/GZxNihGE1ilVICHJr4fo6IsfrO2WgiuABv0Nl
g15UKEZXHYoacbaV/+G9VPgm9kEfyNveQvU2eQQC+05Tdrhi0W4pSMDjIA5g5x4R
YIvqxz2yhSVI+8IBq3XO5uHmMOvr+ThLOruEb4wcN8C1loa7cJt/F+3z8RIBrZMV
qIGADzJBkYn8/K1wZkonolnr0ss/BMjGRbk8rqVUHN5Q1yLMLZNCSh5lPQoFJNjU
IzYx+5mIvvHVIeN5yxcVE9REwitFdD3leH6cdAB+jrQYfwzebqLNNwUCMTGpEfX0
71B0xZ9d6uWPIWXnjU2qLlGiodgqZtUf5nS7dqCfEoCz4Kp+Q9fIteo3Prmhsk2p
wwjEpl6a8zH7SGJHiNuyBmKWCw3yVPxnanSfuqnzD/6nrDT7UKt+QZk1/YVkfEpc
n91cnCD2gQYsQc5aUDtY3w4B5+XNv2CN8ArSGsSFai1zn7E63uR3e18CjdcoJ/7E
p+rzgv9rDY+3CjWe5FHJ/WIppo3qM9lJ+3JAxQcoh7r6KGUzVyZMZhWDfZNY9LrS
T68+VlyZ9VM8OMx8XcMgZk7mFZ9chPa/8CGrSNcqUpZesgQSaZQ/HMpp+1Q2DULS
889Dni7XC2nOsrfSVByV0tz9W04KDlzBEkABszepYp+Ki7b3X2vEATJmazZzrpHC
inedquTdDc/AfPpVTTmlAJozfUVterBayeH4uaRIz/BjPiMrS68pn7xXbsmLG+Ki
GSbieQGtbQs4moPcPFlhs7sfcMBcenPen7dWTnQeu6+UQr/NFEvvMmSeLdequaoe
+1gTvwtVTg6X4z07S/UtFTHg55uLe4E4+mz1jfn8zsLdVCUdky/VrXZpI27BN3qI
V/MAjh2m95oGIH0ZMHlPjozzBQU0k4zkyiaLNeA8rXNOiRhQycGA4OmB6cx8nWf0
Q8wNqFhnWY8WlRC+4aT62uc3DRDg/OueZt1slak1ri/90XH+6GGnJw15V6cth07e
4YS2J35tgo5tjazb+d/Q4uPTCxCFQdCS8NBA2OcfB17byy68RarM2jKDUk64KQ4C
jtnGpuNh5sQQK+0JceLmit1If2/fJQc+ya4lXqsigNaRDOf0+iHlqZbFslxsrEdB
Hhen1zKlCsOTeDI3PKDH5x0eT25b9psPmw7qsov6avfOrEPV3K0B7zxmfgMO/17a
up9AFKBV/hQP0atfu1Hd+YweBNOxqyco+hdoZzdry7hBwIaek/R7/53SfI4X0LXC
XP1HV6LZj4GFIIDwXiTTC+49rG7P5exUzfcO1eUHiF++ZYXOE9eSfpLq6oaPY3oo
et/iQmNOmS1j1OA/MPGmGbdZNl34dJfkjtoI3lOxFAQQnMEF6Ri+qD7yqQl8IxhD
Fg9Vjk4fNg4qnEHp34FFg6voY1Xyc1KJEuYUHEjwifmOB0Jvt+T2jnKWM0OcKZBD
Wd38JiON2NjCOlJx4GVV6ip38MUBww+yBCfQC9rhtPI6GlW6REe12+XUcbw1BRVC
CbAeCta/0I5+6ZhujpBI5jRqSgGRCiUR0M5P7pP1wxd5hzsLWWKmsnJdCDtg3cwm
nIubClQLbLJbVi28dYH1X324A/bJE83LTSfUnPO74CoJTi00hlBRG7oujG5qyoLM
wEkltlzambRnEHOf/R5KhCk7VUIHRYPOpY/qArLKB7lE60lw4uSLb8grcTX3dJz9
D0/tsLUOBDsBrDeYhCOOLr3iG+lok/knyLTIvbpy3z6JQCHjgF8xA79dQ94/yytS
`protect END_PROTECTED