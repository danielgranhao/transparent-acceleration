-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
vK8FdkJLlEN9AW72VP2Q7sZdYob0qmDeEb6lIfW35kpgcJNfNTMPiLIHvZrenbd6
eOCMLfkF+DH3muxpuIw33r7/oML7ZJSQEizsxlSfcyzT+hQNQ1wKN3anLP8vEjS7
l3Zz7Em+VeUQ9yKzPCcf7yx4Gq9zvUMCW42rWPfoKV/h+2uJmTDL9g==
--pragma protect end_key_block
--pragma protect digest_block
HoDNmas/BAfKjp0yGxw9D2QXMiM=
--pragma protect end_digest_block
--pragma protect data_block
tFCiqvaU1XSuQNqavPQA2pT21s1bJmKb5/23Ue0aqIwbOdJzMV1hQMgH7dmChZF+
T3bWvU1ZdEwWFPgGu8OjYw+3SpTnF0zlEDTfFK1kLalCQMsCqRYeGdPnRZrQFDGO
UM3VANfJ2pVmSeOZwVhpPgYMcA8pa65r/qzbQv1RNVcC8qJOyYI40+3s/lw45HR5
KvMuNttMGBHzImGs4Wi4AebYbs+LOvz/hp+n8l8+IxSdf4bvKDbB3+jYkktyzvfe
eVX9BNNnd52JxhFnS45H+KK5Lfg7NPQIczQsY3qgZ5AKB/snP8ySek1ltosjqhfU
3qn7ENJWRyhFneHt4OzgIB7J7rSIWKMs42RPO7u1RgdiLh7bZ7IGwSqO5s18Ib2U
JqPYvRdkLwwxVI1ot4isn4TQvEneGH3HSsF3EcNbMHeqqP3B683aWgdwiG5wxqtc
60YURvmYbPwV99eDLY8RpUNMaVgDhbb4eJMngazPzyM/CSIV2UXBuuWjwfH2T9xg
cK25wAOz2FgbeHn7DesYvz43/2pkYI5TS+vZxuM+3Nr90Z2Ou33Wm5Yu0b8g7cFu
CZ5L093OlYI0qOdb8MmheiIO0sn67LToeYYuUjCWEmqQ3JS9M2NQJ6qDvb4JXpFR
Sk6I119wY6LjYZKsYFOZ7Op0FlYbqrOqxKaKE/Iox8SrwUKyF5+o6OlaJ7f6SB1C
eIz2DyxG/sorqyLFd69kFyGNCPbN9XQvQ8BwcIvr2vkdk2Ru9F4AzjFLUpu5hQCE
GoIzcP3ETJc3I27QglB7+IGKKXdlbdNrjet67wNv/iRIB+bigYRFyNg79mVj6YNZ
Ry+XTeXXRbdGjvzS5PdkjDDzmHqyJsNGgFNa44jFbN8XQzOR8mqWsGP/cXh7FIHm
X/UmdwiLtfJw39FMtE2EoFJwVMNyX0PTy0r1/EOzcv9jhqZ+oHZBWib3SlX3b1k5
YPTKtpaKJh9LF49dxHcCv21m8+mDKQaB8vGSzvfwjLnKLaQKl+1+KEdSh4kC2bwP
XBPGCmOlsK7p83b908u4fO6GrEQQ9+tE7uXG2vFR1idur4wtRBXCNW2/bi+Niet5
hFNBU/o6D5WtFx/9S18THrZQ76tEOt/etut6ViLWFmZMCMrH0NmUZ2+ZlQZ0hv3E
fWRE+3OvAm2SbvlEFzzx6S3pe6pCWAN2g8e3iAi3Dr3r/48uRa8RCRO0z9OM+//8
OlIBl4hIjPwTg5PMl9W22O7PvsFkYtX6RTQvchZkT+8qhtqAuxLftqCvk0nkwdaU
Tfnomv/UvbcyDWwdbHx6XE8PrIChH1Iuy6VjNOZm+6LeilifP2q3mX600T6cIg8w
wZttVv813adAEWx4Vn5/Z5tqIoTAZ2LHCfz+uYdwOLr41bNfdOJZljwKGJ2MrIR1
FDwaH3CXAtYIcQe5Weji80JNpJUtwGkQ5HtCbkisI4f6KuJxrXgxVsHbdBUvigil
XTkjlpneDLqSOcNIx3iQat7kpqF4h+c41OSH9bvlxe/PR92zkoQMkVfeYN9ghJYi
q+YsX56c2jRCqSq9LPY4Y6/Cq7iWxpCjZrYwNg/HE6F9hNx6Aqhh/+YLJq07/kmj
aDj02apHmXlaiopkqKmuVfEn/97wROCCq3K7SelWk+ykmhQ/JvNThTQjeQw2cEey
v47T1gbzwCPm3edkMKQBjvhlvc1JmDMwtnBuqM0Ilzl87Ih7L9tGQj8EZ/x4G1iv
vX9NExw0uqc7OZFq0V5C1YF9zZdP0+PXKtjdVofcMEx99CNOPaF6/2gPhGCfsBpz
C3oU1OU3BChD5h4s3qk8c1+naGXhcNtOqsJe2wFvRyBJXVLzyKplQinPeCixUhRt
oDVI68Z6vOCn5+C366kDfstsJcApKF2peH8ozAHN7319Fv9/bQ4duHP29e79Lqy4
UDIbKIDTnxjcJ86567mHG5if43e22/y7QMHlK7lQ78DQ2KtjaxmXZffmZMnOxsGL
zG8jCI9F0lGVPdBIiLhpfCaWYttqUHp0uUSgalLirTa6JIyyBi4R7tqc8bFLQsUY
OUgzRzIl4hda+fBkYbEKFfpMGjZ740DG+H8xpkwW50SgswWahe3o7b82b4fQnlt9
rIrt0VZQW22V8qLlswnxhYXm6oq2OA3qZPx3oTYH0S3vvsrlKqrwD1QZybZR/V4L
2Vswh5BTTYWB+G6D/l/Aqqt7hX8xHXGCOsn6vxvofXUtkHBCt9twaFQnWAYKt4hn
us7GdKXh23jis/1+240qWw8+3mFGE4Bdf0Powdr65VIYkaDiubTWhX8NXfqzKK0E
RuB9FOvPTaflf7Qm/CEJgZyX5RZ4BKmMY7eyN0CMOeD/GymdB75Hmvcox/lr8Kw6
Jn1LIyyWhRtBz6F2vWhSVO911qq6gT+zQvK00e9N7JqaUYQyCK9sraef6Pf7DApO
uz3/kglx1iWCD5jzOCcil8MJUqvKWnwKG9yANIbFvtRcv8A3Cir0rqigsQy9el+6
qFokTQ/DSiRGJawUYDC9PDSAt8zT/7pGFmG5VGU9SLV8LaJVF80yTRE7lxOCYQz4
6GmsC1DnzOsVu68OkbQpRbD9/KcDEVdGHDvjD68P7J5Zs58THsmBQp+Du8w4WjY6
05m/U097ZudqB8PRDaPB9gOSY6+ur4uYem4UABfVRhYLrNTBRRwYc4RTrk1CMSXy
31hjabrwtHFQyxaO2zaL5vuo66pQtTqj1F8OKpoAfXEpCZL4yyQjd7PH5IgVi7YR
0Il3RTLyJ/Fnou+FfSdWaxzyPorLpFtBkJEukBj9r2vdq0IxOUKwij5bsnn8P5ep
Tz6XezrG4d2cE++ty5RrgFjScp2J289uLCO+2kKYTXaxZdAEb0Rylh97ib/D8Sf8
Py0ARthDY6qhDzPFtjbyCyYAg8egsoNK2dXTRUOzU2ZtEW3rhrCmk7iDh0IE/ehN
ycCA46Ey6uSyLF+++jCrCmBzhaB6kO2lCY68kbyBYnoy+qyh4nM0XOkP2EW71wzi
mbcFvQ1b5hVT7aVkgOlYmQ4ogxp2ZYGcH8ZeuobZGgMcXweBn2/kpWRJs0JpJhuj
xJfk7fh99paBo2245m/ltdoIGM7rcw8lMYqF3rGuabg486Bl8vm9HLOBwKGMEEXB
R0orOGTYEJ04FwWREl5PKgMMH+F4x2ni6+c34D1AgwsRN0uOURIKORNIvvoPsrPI
zrYXpe5ClfYJ4Tjd+uFOgAF4uzHsbSdZMaaCFPjRmGAIPu7uLiHFrHWT2N/5I5nu
reT3Pc751JtPIE0Oe+Uj00AGOCY/9uHuZdGGtRHNBJoG6+m1U/nRJOTMXibe1Ftd
3w9GoWNVab1K+onsS91bX6RzWxRsITiF3a9Cp0yTWrAtRdtiKbb/1/G5VG9WEOUq
xTKl5LD8RXpRqvwVaYkgZaf3KH/4cEi5ICUZuAT9Yv6VPZQ0FDZ/annPf2zMo6Fc
ExnJGqeUlCJBGMGPJS+3wuoYbJzieUdfS5arEPD6rT6QZVTIIpIGb/+e0kGZAvQm
FgUgysrTpy+APgkxoEEccOf55raLKmvYKo9ll4hqBUs7n/ZnUuJNsgBWkEpABnKY
VYtV4VsQx6MeJBRJB9+FH64iI6q70oI82eKgZsdrb/H1tt588D7ladcgbtZg1DFC
ql2NVcSkUJg/ISHT0WZD8zGReZyqLSnMqgC5wRgp6+MGs2szKVCD6Zy/72RS2VNR
ZyJXvMhzVps///VMED2HENGK3zjb7lPsPNRE4aApOnjSLJknh96Cg48AeWTBxVFM
7Ei+u87RpKqVMip7l2FgJV6T4YR0onWwb4mTju5XE6I15pHtG8Ui+bUzin9yizg8
8lAg2DdKrtcpCSNvXyNzzm/XuVvhN8Q1/3Cq+VJZijnXUVQaw45MgaUpompzL+m1
gaXtO+brf8uTnZdg+e8SWGhDQ82qTkeEsDamzdb8HDWQWi3aVEnsZCP42NgB4Wkj
m6oNlc1YzhFfSfvIdvnks6DYGPLWWG8FacPl5s7lyc6m44Imjq8aC0GExz+ZlQgG
NtiDVFF8ma8h2YoYWiBxe/hMb7EmKs7SB8MHMsxkt/VQNSbcbRCRWVLYnrgiqPyM
aByAv8w1EVPAp05gpANdXcWcz/6h1032HCmnvqJijye+W7opWpASbLKmmUp508Y6
e/mMUlVrGbUUGt8dsd/SxsXV3ULT2Erwg0Sv9b6XokFvSGH48fYqIUEbAAXxHd97
5vfZnB6YaiCDUGkEQ2l5slATsBiwi0xCpuoRLqPX22dyrkLG/zKFb9hEx6iwl12u
2lv/WSn9uZ40NoLNf/XqhozPhGlxRfLyzXACCnvnVct5lEcZuEWf4lE4KYt6XOB6
KdR3HTzj8mOvy2qh0DIV4BwTfENk1/BvGwEqxvz1vlAwTWa0/B/NHGvBTmDUXydO
qbr0byqYnSsgt1dS+LjMJdq0Q+1L7WYDtplQ1fQVqa4cwLYbRuuJZHfavS2P9Y9P
7ZyVJsOyGeeO8JZ0l57d7J+45FIBuGm9gKhKzyabFCXaIAMPMe1ycAMGOpjSQKlo
Vt2X+IUEqWg0+1j2ppHk0fwDG2BsK5G0iugAJu0/c/m8BhfLFPq1JTzUF2d4Nf5P
9ViZSEN2itP8Nv63uUpNC1vObqVbcZ0BRbBnMjBrOZYJZsSW59Ypuc36sNYc8NO8
/OANaPQpXGEUvqEb7Ojwrr0RxMPu5S4xjrdPJ1yBP1a3GIu5DDYU15WJ6xhdD2br
7d8g+muou+cZxUCbGGrhpgZ+MrLN3ilwIxglZ6nuzZzmz7Q29bQmOZKGXk/sVlpN
xF6CWZAx/2GN8I3Z26SyejmBIGP0N8L1E5pGQpHBWT8bAxtVaCqYeciBPbfCq+0x
IjGzwH80IqWGA2WDfnGWuRLElMmIv7Ug9Jlu+d4lFLyKMJcgWnpALWikaaeLlS4U
iiLg2rixsBOnFUh4NCH+QTaWssaDtyDA8sbPMQtnNwZRlTwTwZI+y95DWzzEtIew
6iboHGJIsjwkvDbFXdC4uWf2WuFBRX81Z6FXawAPkNdAMNz1txgo50dPXu4DQXee
hg9mMdTnOh0NZrXYi0yPQYVaCCUSMu9JSCWfPxOBd5/IG69lYlewtazYJHNy4U6T
KkUgOMll2CZFSWsgpeCkBJJiHTt/EcultkZZCQA2hiD9EaD4Y370EOqvf8FUVKYT
BE+l6VGD+Rs+wnvA1robnnqIDS9kTFdetcJFzIzRMXm6mwbyQc/qeMPq4dlK6O4B
190ACTUaOwnU/kFIgw5XbDHUOsXMseh0FYZsgguAVvjPOWGdDSh6h6CDSvVb6NOv
L0V+mTti/9b6/EQjtCdYhjOqvxA1O/QSLTRL1LmWQ8cHJpNHZrHjBDZ4rT90LaaQ
2km/b006uwUEF/a+foyPIKbEekLwOlcdi1ZKpI0GKFKKoFtKmRQxj7Rhj80CPpY+
egOB/HuBvQdYCnwXTmrhH88mDvSCqh4gZIoOizLjFqQr1kkzp1WQNJXS4+mz6ei9
genlR/rt/0SWrcTl2I3pga+EO53fLl168ONxYZ55YwWBsb3VCcrSNpcrpKwCcjX8
mofuO9IG+w6Z++3OwHJ316VlbYcgpOuP6yhxbwbRh9yA/bzNuBRfwsEEYke6FKj0
crN3WCNxbvErykybmcLVZLf1wOqTObjHcTnSZXGVNFMC/iv01lZ3kwwmgnrWTf4f
bk9a+tnNhMUw6LusicuQAi83XiqmQJ38BDCSz8Ton50GsSnX88TLPDwApBXuh/OK
77Wt1Hbuo7k8zgGnS981ZcYIfVpvHJUqfy1vIjXFnn6SqbS188WL4bVN90hlQMdx
qzcYeOdH18I7IgmbOmh1JT8U/aACfpPSulFVi1vRG/azmMaWgM7umWmtPiAlfY6+
0laqzZxh9nzxBZOegdGbYLBg4Mwtvm07CNBM3BullCHIYh2jVwbOjDgOCjm2FIxo
v1IjUv8usp0CsLoFCGh5Da2EMRcOooaWmADs964gzts0JDxjYdp/NczRz5OcF0eT
t69LQMvy+CjzxKHvwpcn0y39COvXx4/UcSCKy1EQN80Y9Bq0q7No/+YHR5DWDtcG
c0VAL/1JO9cBRFKHMsAx4gKGV6jG9EEbcN7GnBjZsHMqofIjHPJMF9+yshKQavrc
iJUfSPWctCMtoADhECbh95NbSWKQlG/8BSWwilOa5mMwT5o/N4KH2zhf+jXkOQ23
2o8gzjNw/JFeMNCIqzB9KpbnSOXlRB0EQiUn7qbDSmNXt/+eOqS/JYxW90+rv7ZN
Y1Ouw3qj+S2kB/1bhc2At/fwwEMbVrfIJRuE+znaTIXF4tJO4KcjPu2WuANnRYzu
vgFfexJpKtvCjzbg+Uy0MUIhzY3O3RvreEA3HqzuxjUjAWcGaW6KR009Nadol2PH
dfG4e+YwBiXpczD/QuGJNT8jq14ObwbhFazEaz7wHbNzzXIrfdae32C9bS7BcpUI
wfdOEwwQ5nLku9qugVol/WlR8yNjJCtSk8SS9MVwlYZCIB311pO69ajfs77BdiWy
InuilxaHlZwZnNWPPKiW0dGgjzEODl6/vt5BQ8yaUQBAS9h/fnTSfaoA8qxoQLFo
UHc340hP9Jj+lilqlLQ6mrJX8CLsuAyHPA/L9j8mqwIkKLubDbg+Mzto7vOVM/wT
N3OPnft9uKr2J/23IC5hN+wxL48ShmvWJRRNZc+DUxCMy0Y48MXez75IESsCuhZQ
vd7YDdZMO9psEYQ05/haNdUqsiB8nkjxdO2gmGEJ+Iu7a3WrJzI37Z2zH3wac8XX
pLvZ8wD6xnqsa4r8wR0nSO8F4u4JJmOS4B5DOyiFiqSD3ghcB8c3MRZYuQ8V+wzi
ibMt/mZ6lwdCc0CmJUknI7hrqPNhRwCKEB11U/489WFg8hpbKpn9DKsW9C66qr0Q
U9t3foS83dirSRIHP7ARzSRYKy+NlzZHwRh82feoy2xl6+n9cFY0lnCUjW+XJmIx
DwjqvimlL7VeSE8b+2Rg3BN2THh1VmA5k+Opibxr6UzkXJ2ZvaVQ6ZWZVFU1uOCx
B8fICeP4BHIrCCkbgrBldrJJQlI/McYnI6/+0XgrK1/yAX+uR/OW3swPfStutlfy
Vx/qn+PXpEK3QMuhhdVm6b4dtS1bW2o7z8vYom1HBWtkR66dotUt3NjpwHvBwdBa
x0kH5sX/2SWNRMP1QOJ0EH0GdC555z4BetTGWtceDEbuJ7U6WaVqdo5DexLZNLNC
y9c0ipYNccCvcsGnBBSZLskEuVN/Kzl0/68A90h0TZ4NgFPkrheh3/l+7+mFzCg8
sP7P5k4cqF8XHiBjBkIigY4thY4a750yxllLD3Z7YmmE/DLU3OhpJSW3w9cLL2PT
iEOnQUJGWdowEkTRrAZ/aaGdeSJGjir0lYOGzS+k65f34vG82RwJF6q7J21HlhDL
X0KWvGbofA18qhVXwidYfZStuy04VdsxcI17O0J3+FLx5uG+AenrQ40C6cxUI5+k
B9AU1FHNq1CcSJB+D6rO/EiJ8fgC40CybCtbR+E5kfTlD7OTHfL5Kz6GVlZ48/BK
pwbwdp7F1/KXxzppwCu9en8QTfCOz/S0AhmjDF+XYlAgouzRKUcdi/05GVSXRo3g
Xm3h7RIy3KRhv+UaJYBjCGGgY7gstA5zFe4/ZGAhSlBEdrzAnXuxObbEb2GeLvdj
dk5zlBJQhMxZl82JWrVDGxAMpDUxGXbMlQEDTDA286FbaZDZPEG5OIu4WvOSiVzv
usIEoSLLsGXxfDuGjAzKuzzMrTxSs1GntQ+CYfQAftsKfYFMPfoVyOdD9sl4eRaw
t/Sc0WdhuqQdxqpVyq8jUCyEdPklKUfHNjfdubAOzp4cA6VSoh9t8ZY1jqnfNxbS
xI37WSnGUn5XYhr+kLP2uF8k0J4Nu4/sMppKYKI+vLhsU2V/3n6YTrWPQm1keMZc
7IjZWCR42BRnrIY71KTEiNy43MivrolUJ8cxFQ8HU6LFkdhW3Zny8O5yR2o2yyIj
ympll6X0Ihrog5kMpGGGbzm7QGcS7lxdoK5lzchrMe0a5BFN5IVxc8Godo6TsF0G
mup1sk7MfMQ0oGFHrUJfzQOF9JKgBixpeIw5krc4necba0QjSIMJK/6gYE5gGBZC
iUHJvDvFaeMnjiuL0in5duorlUJUBoSMtJ4NZQ0dIQCkh6fVucgDz7+3bGUrMMGf
MRCqvz3wb912j1/iEoyGMocHAPJASFrtDU3F6ZX/Me191MbQk9n5iC/aLJ8MsbzP
WsfHcAb7ukolXk54o7RwgscgDmDd1hzhIC5i6Bxkt25f6YypAXiF63RQ/A4Uh+Lm
TjlygLGL0B7cDNc14zsESnxmNXUGlRTJyODOc+lhqGKyycfj4ULab+XG1/NUT066
ozEMVMB30Sd3DJunwP+UzCUr+/9haUlAnP4PfhYssSEbcOYF19S4kgBisTp62Wk5
AqgRq6D3e2XjrJ7bU8QiddcmqKMmMTHpv/YEk6Hl9r62/RJsr2LFQMOFEjFX83qN
sRnJ8jvLyF1g0L0RadQ0ibnJ1wdBjPmIX0jEq298vkMTht14ao1zZuafk/qvpJ2L
NaqizuPQVCeQEXZox5JabJPBeS8mM0je5dMH2EFCYHecgyKxcTRLKW2yF3EeD8di
Y3uIBWDFcrCSqHyL6Jsgoc+vmagOB9vt9GOMiwF9ztVkj0eIZS3GQZTiA8iRJ1hz
BcJrBMCRvDbDlVUujik5zRFormcZ98EpETv7iIby6JBCDd9OL/uDhp1nrb6Yqstq
IlS7YXg+SxIhqj0g9PqS0y9gn2qjpMRjgaBwcLhnZC4DojG57n6OyHDgC34TLSR5
js9KLUhzXm8mjD6MV9g6ZvvpvqrjgeiL1H2Ra3fJ9K8tRl6eykCldlhjBSM/wcOZ
UeUKYME06+UhmzhgWX1+aNgrMbIvB1NZ6DMpF/4+DE4f2n8Mk5Jpjf3JZ7aguPhN
Wo0KeV3DSuV4quTDzXRSY0rMbnD7puq6eqZi9d/MxKk9QVRuF8MoQ1s3gOrrt+nY
9g9gg9X2Dr/5DsnDz9uXXYkCAHqiLpNscmGSJIG3zrkwNLawiR3j4gYJAtmtErA+
O8lKHjz/73SGLbqSvOzfaMZ5U8NwJsOJ2IOr176qZUG1xw5uASb/ZoH+aLOP62E4
/Ve0/oT6YIZ6KxZq+zeG/Dlnn14rGzibtEwDc5NuIGEl5QI38t0Mvr3QBHioTrdB
l7UFdaFFeLemmR3RLBqComEzCca0iAigEtxHRdVJtgu1ViIcGMYBxkWswxZA+flT
mS+1D6wCRUS90iZPf07SAUvzKv+YtAlnLQ8F77qYf39iNPTPU1sOh5Bb0+sRt6Zo
OkGuZKZZynkrDhpQrIK79k8EBqWnzVNDLSx31HzrNlpb1tYB/MG4Gfczq0D69hTx
Np+TjBUmznpBegqYt7gvuh9wEfKt3xx/jg0nYIFlA4yFlB6PAOEj5VxFsx4eJC42
nZT7OYJRLuBKd7urgc5lwL6Gw/EBan0szaEKgnf1S2TyKzIE8LGAQeMlwcrLWvyi
5aTQVUNXfqPlToQiXmo/WyHiyHLfojS8f0eLYppwMdoayLktqJ84x9KrJOx1TlCO
biLhK57CUc6s307uU+28xiy7pVuVdZcu/VxZhCBquGvTqRcDWdkJ2tHMB8dsfA/4
cGvq8eKWl5Y0j/4adTc3k2C5waQnKtPr4SqSsrqih6oDfrInm8IjaX//5H+RpkZa
JhOM+lmxYn6K3WxemcpiVl6J+sBaEwtF+vAABVgcmJX36xK4UFJBMQaZYOC3HIyh
kmIjwoz7FqZ0Gtwhdqy3I2hhhazu6N9oEP6pbFph+4GBI+wT7tbiDXnpNqcNthG5
fTB3SZBSddjF9WzWw/nTBbN0ge+UBZJpUlCqKxkMAZSyZ+Ors/wkD5EA/4gtytF4
Hj4V5lYWlH8rNnEKocbURggfI/GonMQXE9JnB+BIeU3BVICpbweyxUmFQEX1lpBw
4YJ8vr8IcIRlv1f9MKp36sCPAH9KU9lxg1z3JmYMGDsDl/IuCrh5Rz46PduZARb2
hRQMe24Xiqs3EfZIETshPA/B1bYdJe1GiQP3rchWuoY1FMRLaWRH4GRdWwSo/8sr
8B/w8Pqov24xyUE8Yd7qhjJ7Ds6ampbWSY1gjxGmK0NT5pOcvqG7I2XW2MZokz0A
uTAsir0NvLbPnnE3tUGbVEi8hTOKGXFEaPPqEXMkMjjH/MYmdwVlSPSavvH9eNQ2
qpUkk1VX5s2HwKZ/RtWSq3YqECsCcYGDjLlyyhTgzJgXcBXKxNBA1irNumRlHvs4
Gs8HCGYwDQ4yDNECyR79mf+BzTn/Y6h1NMX6S0oYlrFqU4BJIQ594gOCYf2+rbIU
MNp3+kYSE+6v/8HlrNxpJSr+sEB6PXizohYAmKfA3TRaQwUiVj0eTHfZZOJ6ETPr
+dbC0jVIX8BycTE90qRgv0a30+zBnHAwsKRMMAgKdCHHEJbqllTbyd5jME/vwmwW
jji6c/q3P5jY5qjyaCQWKerWNTpP/p8jFZ9l6LTiohQevjVorwIn6+YBGwK35DKl
sq4hT53KUjee1thFpCoQY6bKNFM9S/O/iSP9yRsUg8ducAnbIb4BaS+D2Ou1ywbM
bSvCu/d75ihSc1+472GL18QdVZTmUc19ZDL6eNORiqQSTyczBdCS2iaLZYOX9s9I
5BWt23MLN+FLhDAkQLiLEYuMEQ5sYbMI3dGZ3fCKhhfUcXB6V1uifJzJhtJbDF/J
yp62JchBXvFpY5YU3QYaBHenBwxaypMLX8JNDzikKoJV4cf4txchdG8QVATUslT2
UwzD+g0dOLDeSzftcXIJ+ulh2wtvgGXDuTkfQe0/6O1YxSWuDh0oU4YW8MOt8wRH
M6cZpGjK8MiEjmqU//7BVFuPJu40ZhYgXsd/z06lLusD4Ffwze60d2w/+s+TLhGP
fy1EMoiFD7i+MQ8iClvrSSFNBT9ljM5808igbrcwzHilD09cuiH6s9UgDsoP59/9
WybhvZDo2CGEmBDmmybjXkOnAMyNp7/1OJSOyfRiqynRGCR3d/O/c0l+Um1Q6lfm
X/itJh1wgRein1hmWnEv2o7lbgKBshm94FOiwLhGhECtEpAIZw982VDDbsvsNieN
PrVnK491IK4VHhCUlHOXNMllI7i5ZIluPOUGd8j1rpyMqihRF0kFMMpTzrY5Dx0T
EAat5iwNlm6+5AX/BzPkGKSS0Udjil3pGxC8G0x9rbRUzdRZUOZ6o3Y8rqr3CS5I
75jyxLIIjywQeLC0coLcD5Nch2c/fA8aVerdEjQrih4kETL8cDIN97w20mOSYEpC
mqDzUgKmxwhBOYFHd86drSNMgPOEzmrMP6M0r10TjhPNBgRbJJftXOrBBFgMuDfw
r4Liqr/vvCeDjp/+Jur7BENOeq/LBCp3uchnd/fV7WPPFOJUe/el2au+mE6P1Iz3
ZsH751cjrPDB7mDzk/Yj/pKvK8EA823DTg2ZDDANinzSdCgI82fLxAV07wcCf7E1
t1HzT0P3Et/XQyhDt0luF45QYot99UHN/PDrSgCsvhBz0mzUwLlEYwgNW2hUFTeZ
LPwdIjGQdnep2A96VD87KIe06zsouCHaMPuZvCGVydTnjW5Q9AtyN/GJLQjdwuqq
7RkYsvej8deiV3eCvcP8P+mf8nDjal5vByFrB4mF+Z+XeQhgbvmckljwifeaPfz+
Qnb4xDniTGQwnNENOgsBZA/MMMQcmKob0sTQ7GOb+nWvZegly3+LgEb9JzFNDIiW
LcLVjJ62UuMuHtgNyPtigjIXOmrfcK+mFCf5qn7sIM40f8btTdbDMH2hUR7mzNOo
tXY4BOg0Evc/34LdNRr4N+fobkvo/S/VjQ4ABB8dFip9M3FJiEMS3+MonhHKf5CR
SZnUTcoktUmgvYa2Z1r1C/Lon9LqYoOs1SnbbztN1nJyMMQdxfIP8wqTMnzVMLxB
v1KjHLz3M0JPpoTaYYoWod6KYckFvHxHlSCOda/fKovItij0g3p0eRHhDzzchTXm
MkIayGLnAxJ3vvX5gCSdFWs9ABs1kqLv95J7mUWj7NB2iXi53BjLTDOSgAzaC7ZI
JynNVa6SJ6SJYSaVBYwwvHbC8W/o6H4iM3BqHMeMqxnLXKMmuH35fTSKsm3N/Oez
LHK3JOeYhKs5FtAQdMIZt+i/gfoZayS3hdrYCuN47WwioWndB4UUVx+qh7WWSHLA
0Z+4iWbLXHJlQpO31Aic+3Q0FPUaFx+jeKKRBCKGj/umAiVBxkECtcqG5HpOK2aR
P78M16o8/DOcadyMMocPqR7E/Ebt2DVoXygOvy24twLJKSGYnnj8sxav2HnX4QLi
caBZnG8uSlxcV+gu+PBaY6UBRn1B/7SiiPpOALMBFMJZL+l8/I4IbrAdkPP23UIm
7ZvU+d0H9TTry+LTHB1x2XXYLB76+bafYwWoIbj7ONt6eDWbzJjge5ahjo0ERMcs
RQEfykyR1nCm0aS3k95/9o5ePjJ0WNQSQ/YtPFsB/E1Vy0d8pSZUAvKqkj6e5iip
XGZIc2Cl+kGXBF8ztlWfgZfLLTGni8+OWAmFr0NpQJ3HrcRoPEvV9sfWI4foum+Q
nsXuZ82Dkn4s7AndSriu293ktRVk2KNvrFtwNVwHFwK0oiuUATpwsIBQ47xcVms+
AzDZWt8y18hm6YYim1PkSMfWWYudBl/TRVcyxb0j9MHHm+exeOVcVRyxYhX5FNnt
q8MOHsrQBEZ+9drAMW0xJzOvIHUJHDmSGWFlpbRXZhbiX3SnG2waMA5j4++D9fEw
fIo5sosLfWOrGWDGXKnRBm8PtxKhUx/RIJo2AGPZ3pW9YPPNySPWcVC+CRg47Jj0
QqhSMozH7YBTfyDGWOdE0JnNlvooUiVsbh3Xx9+a2FnRWWiriSGb6BB1sTUGmrfy
ZjBjGgr3NpqIlkObSdOx0psoyDMU37lzs6kbUL5eiDWLIPutiza75KWksLqJelM7
dMMvHQocRMuva2qQcFmROkc1oRulaqZdePescFhGO0chDZJJnDBZ1fKxHxGO3ArB
4n57NO362v0q2hHbY6ZP+gv7l1+yzCXsbr7+v3fDrWur4UxLxNZuUSZjSBlM2xMi
01HEG3k5cCmDrW0y7Y/d1zWvhJZkwGvmJ++Kn5BtFYfCdc32AMNu/lggqSOg1Gzf
xkKNXoRjptmxxyGgy4VbgPLqAweZ0wZH4lMscC/f4bO+OMeTSQfxippWCX6a9sV3
8pwKbqE+Ahx9fvbzoaHs6Lc33eCVR5nBF7nRbLecGyHicZutxEwh7AXfkOhTnxtr
GGpjViFZJYg+WwDdcOvy8sPGf2cFBOPD6s4vzOeEESdq5jllutvTwozr8AsGG8U1
QVl7Zll87ZGHfarXckGjAG1z/yKNAyjZBkkZE0/Mbtrc7oBX8Pqa+oDljalJizkN
8s+fBsJt28hGDED9khTE+Cvmg5O98q6kGe+KTIIr2lPsa8CL9WOadlbRXZ6ba8YE
ig+Pcwpw7aKHpKF4RHiEMXYedPAmpn0BfaK8aglUnhTdbxJ/4UzQLiAmGeVe8RXA
RISLrH3LfhkG0Oyr6CmyX392hRNO1bU45XlUHmWhczfnBuYjKQJ97N4QFhotpwL8
3FtmcbNKenVKCsc+oQgl76wg8pMESLVSMPP/H3lmcFhRj66FPg8KCjpCRm29fHEU
mZUEI2p6XruVIOzhtj9jMaXfUNaeKvvVE0mEhZDDN+80+wgF2n7+m9nrL4X7j7Bv
FxTCjK+8xyt6l0nUAmH9leaooHvnw7qgBxeKbNHqcyJu8YMjGarhpWwffOCu+WRr
61qiT5tPBHrTvrSQE/xdSadnXEBtBtJhGGaL5qQkGfy8DBLqR8iXpqMmKVN2U13w
Y2xvZe/pIFDgqXZgFBanjc3BRvEe4fLteIId/1R6tf6WcmHajirsYqXmcBPVHIEj
fEFqbPOLS+HObpUgzOXCxihqiyttRucixt4BrVI8VP3CxxlpClN0E13olsahJt1K
9Rkp/Gp8+TbCCpzTeFz8eq8cRyQZkj0c7XmIhp40ojLsndLYefdK1FVPEfx3ZRHV
wNrCyuFGhKHn6OG394v+ZtWsJYrafejgvaUpQwfTHmg5Qpz9TdHhglOz2hK+hEJ1
b7K+Gb0a344OZDRyV6mH5xruCsMyOzfWgFeu7kp0XfIdTs1/o7/3sD49Y9otxVWL
yC40Hm9k6+ccwFHOtAj3LD8GUcpuwCAdZvvMdUyiYlH7KcBg5F2CYROcRyNwaA3/
XBmzoOVYwu+qaTA95O/XYcF/pjuziLFRSbGbIcQkx9mTVt4aB+Q6idF4gUzvGhaT
RlNo5h/+/sj5wUF4wzcGIAdP0psY5Y7cK+An39VJSFAqq+mZFa2zYqZ8yU+GRJ11
MNis7ewFQfM8k+UTX7SvetwSIfR/tLyFVy8aPGco958G1HLSI1egklCrlYFbsOa1
AhRct0Y9gmddFtBXlJkuDFIkSzMudqNTtw8S7oH8jczQaAsuj5CHPEnk7D54WFqW
/Glw5VS6O02Xx5cg/iyiROyTTwD7PZRBvX747TilToGm/bvinYT4ebSBvnYkOxjM
x23kKE38HzMnb6JD+XWnSmnP/GrSPOufU8eiFj6AwFTRXiXjHMGzf94KuW58trMG
OryWEYE29wWzPOLgWTKIZsbO9KCh9XgQ9IrV7jyCUE+b1czsYHsuQO9X+8UBDzGF
Vp0CjHonMIWt5jmFBaCUH9p4LAbo5H5kEkBzw/vtId4zeCPtnbiZ2gj7fzcmPkKF
7Wr7ULOwHxbZeBedJNnQxJITJptLIKnJ/eKTlIOLVt+taniRZirLodiK6gq7JJOg
6GRWPF4PMpNfRP7CZs2co5v7Ic1kpm2pYLHDuR7ZBlIkNuVXFxaPdL00aMDGqwMc
pATM81vdlcBI2HYvo3ugsw93kTmpZHjyzGaMrjxThnPl3vHDc4gmp5pGpSy8CIMl
wVUd71YWxHjI/OSWapf+ClztdDh37hQiczYl/SsGBvH0bYBL48WlXAaosmaSbFrC
8iTrAEviXBq1u738wa2JvaKKrBTcZACnJlBATGP98QpNItwvgigZnB3vZF9CooFN
L5bFDAYWVbjhZtfCB233x/Y+E0OUFay8KtZIVYHgzg9RpFAsQ8wlZZQaESh329i9
Po7rh9NHRvQYsirynd9wIR0eP4bOrDkVQ1Iovc+RPm6MfUTriTlgnEMFZ804AIq9
mmmFb+0lfgup6lA398ErnQqw48z2IJuHOPdHx3uCOVLk3U5vkdzfSh+GO6sMdEWv
vfHnpFsd6bagSxsPyOmb1NmX6InnfFsYTbL/tDdi31lsBlA6KAIASbHyPMw0adgb
ZbMgIERmjosVmEohpcSJ1y8sUjbVSuFq2gt/dQ3UZLHar0GZudc1ZlyR3EX6nk6W
mtJd/TIbd/alY33jNeiJeuTYG8QO3p7Vp1WyIJ+HrXRgIikw89/jniGxIBNavjoX
61R3Uyc7KdaRa0wYuoMs4hYrwlJnPvs5dxTCOSq1bnO9VP2gkTnTs+PAM0SH7HRZ
NwUBHY/sc6Wu566nNUTJlG75iijjx2AiRrCSzmEw1O9Tgv+gbj3ENl8fCfAwUfr8
tIQN3WHm7HwX4bLGYYn57jtYwUlWn84WeN7oQxsZyhYBXydxZfMoQnqR++auJDOn
SOU547PssefT6z0RwT6XvzPcXajQJpMRVOBEO85sMr207WwD5F7Z3Ymjj27hnVne
CEcHgihNeUrMx389/V5H+DS1i/ZOIIlSOvkypCdYy6eGNlO5dKgW/b+2NGkr2jXD
RCkt8EID8VAqX67DWclmhpzplH5J6yui5Cd1qFaKr9miJK35i0aF9uLlte7Khr8w
sKSM75GZpiaSkg6Xy1Wc9zr+afYzGcmpDexxzVfCYP9aWvx5/p0nrPTyXUgsYQFG
P8b9NEhogRW3weQPNa7x9HIHpkZK9DWvyHdqtt75OdKuo4zxGmwdAwVGEySpzgfM
17dK1e5LY+B85XrBfQ/iAWxQANWbXbv5lOyx6orp84X1ITtT3x3udFlfHxqum/kY
ETVTc+pxqHBumz52hz1GXElEGNejW2UzHZgGGFU7kwCTXeQIv6ts12clcGVMuzCA
4bo7SjrYcc+duHS3jd7iU2Qnm6OYb/8TKR6gksdoe4jwQDiUsarJLU03uA7bO4yD
5xpHG1//RGXWTl+s37iiQpAuj4sI6sBGiCWXbPLCOr0qH7eJO829pihvYHbmN5Ly
GwIljiaN6OMcJPIfiXxB7eDC3gm5F4IbAO8TCf6dXpy2K2ioK3PxmWpNtva3BWd7
ggi2Ka/yIlJuVFMUJjjUCuAHPCfpd/3/8N64iPEFLmm1l8uI/8c9poVCkNSqaN6f
UDETS1mT6UUfgKcNXZsHaCictsXhnB0caaSK8hGR+E/ALWnapkbSy03USJd8vdMO
QW+qTww+PjZGRNnNMGRweWEhos5gWlbhF+z+PQ2orWmURxQ+8xHNHZxs5IX0ICm3
pU5v6pg5+YmlN8ApQmpFXvqE9gLes4SjyShKvmEFPmFIRvJNDDvDUi062creaUw1
Oatq/m7h+t6j/oJL0MVGsnCNKPSGMlLFzoXINpBcDrpYr81AS7AviXosIdzE8mXM
bD8ijDoQvkWhMOVgJ0xSuSm2NbQMZwTLGrGZX2gG1ZbEdRj7tYarHeTa5va5EvWE
8JAJXXqMIwPx0lv8CoHUJs/jB1bptSC7WqyRnZH63nO5zsaxfido7UjJkk8UCU+D
IS8pdLPGHRy19TLfqkI62wbPczEY3W6yp0NcFG84N2PU+L0LuajptfsZYaZdBI8W
IbpmdkofR6cDFOZjlc9J+T3foT9yvV6AGRBSIFHpneJaV37vHbUZubCdeUFqbHAn
7bfZeYKJbGXu8CbBWMkaSxk7sOu/plYGIaO2ZPtvME+lhxvOEuJf+8BgyvwPvpUO
xFqIztyDbtPWwBMU+jsQTdRlDxBbR3e6uePW0clwG1hbZ5DBX3/YnvnhOIhQ1oIA
lKYyiGZAlbzQcqTJ+csShc6uAVVo8mVjA0FIXhyuMUiSPlfLXOYfWbCT7p7F6GVB
W6AA6PeVzrwjCsfHljOELJoVu/l+mPma6aDIktCuGOC4OR3yrUbMYbO2scS2vEFG
mJKo2kbMvH/1P7vKIW9PdRuxPLBFMPre8j8AflEOPnn+7B701XVSzjCmrDM3jH/n
vjWJ6SF4xEHP1rlVXFrfVxJ1ShgNV5AddDkUhE6dhrNo7o2mAHOlU60/caIJMKrA
73zOJNmBxGNn6VMLitMPKMifbgnpSQYHH4PlocFKKBMBiUVUR3R0acraKMNDeTmv
PIvt7SHjS0pXJG+guUJuY9xQMVwMZ69rbuoTseNVr5p0GEVlimiHCPPWOJg3+jQB
MpS7wpVEoiUS9LSxQPEoqc9I0Te4rSq+BPumOGD5Eu+2LLN7QU0t0EVbxz9ewg6T
YuXiyTEPj0ke8OwgmDu2cEOqp/MgaLxprMtobYSDcvuWs1U8+THbvlF7/fLMPH/r
FPSw9W6NJgwBIjp3hN9xahaL25mSLrRf7ZKes37GVrBjJv+R/gzsDcr5gu3Kdugz
1p1hBneKg921Nce4CjJNQSJjyX5jCN6AfoTHBt5v6kvB8pqk+7kB/HyrSnD2OvRz
IapTlj9KYDBXCvLmAVXl0sXL19oaupHN2kdluUdEX+lwM23AFV1yOO2D1B8ltfGX
LSqhL3mDYNWEm2cOQT5zaz4EKu6JOeehmeUBsDZCV6cneCGp+rJmkg0srBqlC2Ym
XrU22kWV7GueoNwy1PQSHd4MJ4UkHb0TsJ59f6DzB1P09UOkBNPm0DL3UNeyXtB3
w84BfADO6SOTuBBocQTcwheCCMAyKlaoDHN7D1+YknKVB+YVejY0UdB74SZhHtAm
yK9MbKoCu1hdZ64i1d0yANI3IhEnodQIzPShq1nSh+z7pMYT1McSRgcUn3PSDZQR
+NnkQli7XWmuDRq3xgM1UwDfWj5h4nNNJ+q4pmbi96oB1Jifd9NKd3LwY/Xfpdu5
DBU1KAhJ453Dvau3Gd3VrSRPYhjK/3tbET+xeJACoViGom0JWKSGDN8tj+D6lVnV
1fiu1Fy3vKFd7OBhzpN8cqIM9wv+48G8BjB5L/BLwe8yl5oHm2QtsbSYUootC3LY
Cprroo+kmuHL4kpLd8s9WLbVe8Bb7wddEBJqa+IlkLKY073QsXzDw7EzGn//77Ck
hOxaf5wk9uqZoJluSuLnUBOM952aMRtNCKBtsOc9XU2E/zRtVnzfZ4AN6GxV1960
xaYIf8Zgfg8c0O10gXbqjvg98+z8TPxsjcU2wbr2Z9L5byq80yDrK/eok/+CbwbD
jgSUCMcJirrpeo6NH+iohB51ct2EbBdWJLWn1JcW7HaNi9QmE+KtcxiaKrlNrtKm
TqDNC+PKWqQSjYIGLutaasD5CmbzRXu0jp5z4hTzjkdaiUHeVpihhr/K77wU2A0+
pg0BiG0hqclW9x7ZtRLgoe7JBPwfaCHV2VBhftzzJFsJLdCPE1gZBCvH61hQJpFt
eoXWKw12f6n5MEW/UqAhBbgTHar2JPjKGs7yEymBjJNIU2D2qoClhB09u2aefHeH
1swzULEuYtMGlp4ifmt85GIatnbXNLRQ3vL4nOEmZxJqnr7t6PkGq2xWM6lv8aWn
UlK5PCESEkXEbmP0NGaQv5BRgFvWpEOgZ/sIgYjKHx9NPTmKzAAS6d1gvkGtwIWs
j0Ei5QnnSx21DNWwpl01Xmu+gFWBpFWeEYbqOxvFLAzkpQYIYvMMj20AfmnYsWGb
WDfkVnPh6eD373Vn0rHEspH0zBuIBDhWVxYidSzD0B0x0RdhsPtt7mIMEJ0yY+Ns
H4o9IEkI0y3W9bugyGg2toeiVR9NVqLmMbZ7hk9QyIgzt/HcOQr5iQVV0Z73ATGH
GOnQv5Puo/fH5b0vhvqQrDydUoa7V3CGrTIcFzF94bNgIXfOre7IHcfM0nq7SJEl
GftMkbBMT5tedA0WUaSNSznIqKx5O2y3jKkCx9/V2tP3/ECy6tKd5ZeeQoSTDxE9
6nWNyvYNFTCRJAIoBXh1wcxOqzrk0YgDmRgUcCpGn+lBKuwqB7TV/h/OrqXciKQS
CDdEBMSakWuXEsTEB+NF5+GMufWIrxo3zASnX6DAy45KhnbYmeL+u2WQuzhV5dzj
tlLugl+1mG8GJKCc4N+1YychNaCBOr0DHfAPuJK6dhSyiUCIA8Ue5bg09xUf1S3M
cIAfbgcx7MTlMiJCHumSGYMSCR5vkXMpHmouhGPf5XOGXu5ySuJGD+H1ns3liHPq
boHMkSmyuArV0MBibekqoIsATdDweR1JNLYMwa8tn5Cu6GjzGuoCthVIiWcandZQ
2zDFXpyZyzFIwHJjTyXjwIJdCfY07CQKt7pK1ylxEzjvDU17etEyx+ZM+iKOtyPM
p99GTca/PWSOjce4NVOC/+FElkrtA2rjXyxEkStKTvpjNHTBGYTnMcbVzRFpREng
6J6aeZcuptzReKb/GE9AiqtDJrcX4LeJwLqK4XG4+wZ2mmxHZR78bqKxS4utsxSL
pB2sZ2x42GXvlZ2oBvhP4qhLne6chkgcBXF2WZErbdmXlZ+vE/lAD7SxlwL9PQJE
m/iG2MIwYlEjFPs84PqXHz0BMjFB4couBNSSKeu1DYI0myrKU8q5pHnOO5XhAuFx
bQNdyR2KMvyBKRyUXwvq9wYJJpRT0qsjPdBnMGw06dYHU7bOyBSo4ucVBwS6Symc
YvjUoWyXlJcosT2Y4MM4yd2I8CbPpq1tFt3H4Q/2V5HrJlHBCvNcaVN42hKKzQPo
HPl+RZjzE+XHQTpJfB23251W4xEgdlioV0ChPzgjoqJPI/jsu2bsOI7SPygi9+Lh
cEmsTrNN1wBiBCml65G9CCQWgmAIP/gw/zdE2m7Rk/UZWIAeYuiIF1xlcG8oi5PO
vmWDieSiF98CuA1+YxuFcsCi6yM+GEjZXeNWjucjPjMp0TTvLx3U8+rsG00Tj9Eg
H3Z6ujtZamjBvvGIHxVy+liMd2dEblDTRVjYShUPSBSB556Z5LlBhAUcnW7XkhV2
lnhPRki+viIdzGqO8NClI3XlekAlkIHxfPtLD5hmpXJZzDL55YiS22l2CSXjKOXc
OTsaIOBVnITXHOqNbZv4DVfmgvnRl5ulJmlDiDyYxk3aglk7mJigCPDV4vCzF9+g
c4UqyqHA83Akng2Zf23+tyHdLHMhjJheVM68MmDGNhi2tjZKD0BkyrZSqass2psI
4rUWk869Fw+ZkLCjyjLQvo2Qy4WcrIFQ39OzVY9u6hRexwZB3694bOdFg3cQ/ma6
WF/HjuIr1jpfw6nAuSY6vsh0Q5SvT5xlrCFkdloEoQQHXhddbM21YK4W67ciC9mH
HLX3iCGf4DgbL2XB3QnsVjzJl9cgjyzZ0dGNblH+j0nqoS9bS5eyX3T2qjVy+kbG
VJ9XlqMcwfr/KRUrQk/RIYataALPM8raYjU9GVOAg/1VBF+/CDBGHs7e8ytegjnS
bNiuv0L8dAEKHDir3tMLqn9JwzxS9F6Zy4VsgRBMwb7w12gR2bcoeCV1Xt+Obgkl
Xd4FOpuH6Nz3Tfqmmu7sjSgua6ynp2S+dDD7i+t5mYbiEygMKhykZ2XaSJxUm1O0
rKlEeVX4vGguZR7uiAxxu8pCriI9GU34eIByJKmh1sLECztfMwmzedi75pIEdXRM
ncD8a7EtIm0DNCdG9LNwDEP0y45nprGuOo3msj80nae0CvZnZX3eJw7fD2M3LzeM
pr3fMT9MPVDP4HWkZ+p3bZ5kbZIB8a2PBeMysXwxukK/3de8R9vHpn/CcPaXeJre
8+sHs4ujusOiu1HBRvnfGK0yK9VTYvIjuc+lw1FMxdxxRGLoC1TvR0FiIJK025dS
YVs24006iVq2nsYRz26tidVfwlBs0TC1Qfm6WEeK9pzF35my2JfqKLZl/q9IVdlT
pRe78Oy3dqYg4D7VDX+hfvAJDho0ZSMWKaC9jKgsAUpKxrgKFexyC7uIBlgnv8Vn
LIK4QOxZqU07WEa6S+uwomXD61fYew3zn2Sm2ZLY8VafiG+SXPGHEu882G+lYfob
fs9KW+M1EvGEgJa6bPYxzPPlQ8Fl54mYBQs/y21wxZX2Ju+Am2QT8s7ZzWMQPH87
2qlguHokMRp9BrnFnQUQG4300e6DzNS8ePimCf9ikboFguuz1YR4vds8dWCEW2cQ
ZWpQaxiyip0bLDCnMqv6/+Wyfj5Ao0Jh09qZ8652+uLjObsZyUYfSeh7RuO3akE8
bsmZ7ep62f+GME1ZX+xcjG+wqCfXigbZQToSSpZ4pJHxti/BiirW6sg8WBzvKsQK
MAardckifDU7BooVlL/ITF5i1uicBTkMZPDz6w9gwEreOn8HgLIjln59Nh4pX7EF
YQQjHcCYJtwNT6ryidRz4EatBt5M9KxPAN6HDuSSB2K5qT2u8vIqVnESBvtZCgv/
DLuBmGOFWnSElM+tgVWshcw70fJ83S3RxVtvTXQN80lkSl3R9h3ZnG4FVXCHHfIS
uzEkChHUhNwKFqxQieK6y330kKrOGCRvNHfstHM90TPz9kbRNx2RV3DOx5CqruTi
D75BHSK/ishQSCyGfndl30D2cx98pF8bIu9GaMV+2pNzrr29jwgG8dEesIRz1pKq
fv96FEbEv7NLX1PTUtbTd0cPY0rxPcCtdquoRqYYQQiZrjS1LKk+gHCS8qsj1iJy
SLRXgc4QNDzoUOKAFPhESJc+QP2MMoaClb1LL/4z25tCQgKZVRqU9GH4VDVlhZRM
YTHNP3CwC8zQ4LIf/iYXNid0U2SgLf42MEW4HY2vLa+B1rIyzT1C4vnpiu80Q9IX
MwDKg+jf+MQEDh9PE4UXgM4otikg5kIlF7SZKuFos0BJDIWHWenoH5nFeJTqYSJy
Tc64M/4s/dpDirTeu0ziWcRR+Numrkt3dBe6MklOZkRR6cqXrcdcgQo88KtTRihc
FvHS7CMhPd6ZdwlgFlD3Uo62nW/ueb/NF5to7mTD+2x5XXJLF1UGRY2GPe6HUqv7
bzKUB8hzWuNjEaAEY6NQBqj39ILER+MF7W9KUXvwuYAMQvI3TcQ9a+8j1QUS7J6Z
xqWFIadHQMPQoMHS5hN5LFPXLiBkbrnQko3IylxGuXMiX5wwMvrkHZd5HeWtzMik
9itdb7ym/M+Is95Wjf/dbetSF/5e0S8VdYk1seOYAXtlq58HqXuNiK9bQoG8EeLx
yZ7WMB5iNTKslmzCjPq381lzf5aS+cqYcXUqf6HpTWRGFqYypJemlRmA1CsERsWc
MejrDomW0+x1y9n47Okwbsx8VfbgAwnmxcgSdVSckHzz8MNlbOXxU4CGJQH8JsJ2
5vQv2ot+tkhGqLNxrG7mb/AdiAW/9iYviUh3DcYbVWdwfd5oDywQnlbt2DbGsQiZ
Kvx6fK0CSOPrEbujqUGii4EXQ/IAnINR5BWiA7XtOlwu/e5ym4cM5E/JZx6J93Oc
Yy8vkZVUKIpo2k4bpOBmYlZ6fWz1DLamSK36K0pq5R4Xcrn7ptTKdplkEgaw8IJw
7XtqcOPS6SKPGTxEBjjNxYslsVSPKGlI3foe0wnvtKVu/jw9n2sCTD3nlYHHMx2D
FxjoDhfGkzVGYv//2FtUPleRaVe+byffLbtYfc/e7Mko217+mmsuyVVdikdsREnz
ARiKgQHdp8Ukzgr2DgxMRqF63Ry53e1F57vrOUNW7CGgCgr9ApfSO6vi/qAX1ZOA
y6gIX1hJu52RmIPE7u82vd3FtT6mYwFJueAD/7Uvl0NgJpk8o4mtTH1/YYUdVIYk
8xT/SVcHqpRCvYBLlldrIZdPdrExWpre4MKj4aa2pP9sEnpjkIh4jA8l5oBQZjzn
Kxy8fSh84OoLWNtcfmghcF5Tv9D8qDLFt/pvLFkQuRJG9dDgZAbZSx06DkoTvyag
aOKwY9mDqWTPoarxJahX4kf2WewVP5sdbuiu6bsn+7ZYDfEuTKgWuudqoW4pVJaw
BjPUU220/iVYU6X1jMq7oilUV+tZo0aRaEYZHsUs9mkgCwc15BnWspzh7tQzWXjg
SynHIyg7pO09OW6xB0K4rWPuW5MCl9ZABdgC8zueF3ChoNJ++UBCbpYVnexf6XLa

--pragma protect end_data_block
--pragma protect digest_block
KVriV1re1HfgET0UJNOSRDqguNA=
--pragma protect end_digest_block
--pragma protect end_protected
