-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XIv5DhcW1osZ+oMSt9IbgRNj7udycQcD50USqFxn2gLscefbkpR4WKa12q+2iGo75yQDhLxpCzji
P+oP9hvOqo1rGVlwCHRSMPsURCMSyELFpx05an6OFscCdg8hUgMXJvUP0YckHXawvkJZOf4MWf7f
bjs8wQgr5zvvgF9S2DQBhSZB/9xGz6GrSPpZKuPXYM8ssnOifQ8/IdEcXW7MS8T19CJ3heQm7UKR
IfUCRzRuELde4GGKO2ywBPN/ZXcen4qyBejcMzVvwjZEIFYW6YaqmQnomR0KAMmf4jP7wONksMV6
LbJyiTWlXoLCUgWMWwY9gQb5D4ID+ZnWzKcn9g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20096)
`protect data_block
MbswHcdYfzjs48xWXF3GILwelcr+3BDd+h9FFk+MukYl1bYOt+Dojv1II8Hi/IaMp1JFUDx2GOgq
WidC8W8Hl2NPa1ETffIDXeWi0R6HOFe10Kfb/VAdw8HLDx+RDb/9PO/1ft+OWdFXTDW31E04qxw1
bJLSRboF0G+B6dNCia1L3nIi0T+VO7WaqsZ7F/wD8zhg+v13Hs6qSB2G7T3Jbvuez02o+Iypryxq
OBQw4p7/MNFW8p4CSjYnVNjnSGNi4mRZQlclLNg2jJrrkRXwi3Q8A6HcuMrnH/eTkviWw2+NEyuH
ifBTOo8rioODVD3anygAq/bSYFv2PugIYP6uOJQUyKokkbXyTzAcHv4he4zbhIjXXcKv0gODYFAh
XYL7fyE08+jrgbJRsD5sTPaJ98qpE18vO6w7gr3ZbXKHgINEt40qlucWoF32YHQDNT0Ppo/xQwdT
Nbu3wk+LdxzReAvMGDA6g9lTWMKA35j6ldS94qj1OThuLMBgQ3zJ4/lmy+Jxjl8VRnwep4xf+Kl3
cJpsmmMEiXAglZ8tsrS6kog3D8xXtmne++S+RW9kvsSwQptLhgqEk8sOsc93nmLzeIoq5IP+XjWA
RQRqjyvAdcCNEbemdPrd0DEGRoLDTt50RpCypLQf06K1dZZAUzaMunxQoSa/gqZ0zC9y0zYDxhYY
cYTaV7+mW5K36xAF7NiTmxGZKBYsEkOCi8F2fU/Q/TJgkqfIm2c6E+eR26lps14ZYZt4rxeDIuBB
IfcwRJ7fLcYj5fQ44xvjZUax/4QQKYHrWM0REXXrhEUr4wjb0q08UawKvqS3dqigHbmckPNAjkBJ
mMhCO+fzosmUXicwI6aHwX1A61F4Fhpcac+5FyetrdTi5/Eg2DbMtYKRJDC3MG1/gsV5rlKC/z0D
gEE3Rmc804aFQ1v4JTJ4Zk2IFYIJu5xbr89JZwzbvPgMXSvvG1vwXMg61P0B6Z7U6mfmf/Xayu+v
I/iFHNu98jt7HtGxdGDiVchBPG92Ky0em2cqSxEbYqUSO4zmVXQB60/YcQTqVdsw3Qv4PFlzLeNT
scRs9skpaWg/BStCprvPETX1+/XdLl/9s3oh1rdO+qL7KEcRJqhDa6KlIzQTzU6vpuA1Cp+IaJDP
GHKcOFW2oCFf0Vy/gzc+Zoiq9SWVBuNxnLwafbHsJ4rmW4n7ZT6gOZC/PvnwXTpHSfFgyh+EywNb
229OjDNlqb8YrQ8i4R/K6GKSNciHqm1XrgC/ZLfRbReSvZzksWQZeFxfsbGUJX6utre94U/G9T+a
6ApE6tU/lXEybu92FPd300tEP8pYLzRu7a6UH0ShDNgcLRYEMqN/BRCyPu7mSKonMI+qC6mTZop1
5CS6qzrZHMkww0hz7zBFwWjrgbXNu/LpBN1Yu+qezofVCkwHHQ0HiIv+JwMumakjIByZ8xdtuUFB
bm7gTuDEbKks2NasJ4mELKKguee1kJf0fD9D6JwB4lX0fXQjvHx73Ta5JnBuvo4r2IwB2NW/QNho
U51nqZfx2zF5N7dQXh9tgNTpB+/9Dlj4F11BFAE03HCQpe0Tvbrsi0aA+NhFfYVF1XtOqZ+hICpC
g1wqTTXTzW3l+qkiz1m2FDZjaA+GJoBhmXDgSsqov7+CtZjSurocgh2bMna0+mWSKiq0fVdajLtw
HZTIpOkedxD0e1uE7kOtrCh4m/rVveIT3wwKLvx/1L1HdDGok8oaWdn7qaRsQRJvplFJtiYIxu+2
3Be4ntkqWxlpKAeZL/27kO84xYj+9Gwei3/uZlQapdi4Z4XsjJ3M2FZBKlcnPmSsE/uFcPEAQ/R4
JHWulQ2q1VkJT9DPBq6Up2Sz3NIvc/xLTPqQygHmjXua6+sO4Eh9jsHGIuwWAG9R+CLaupYqsv2G
M+WOg3OIo0ocNE/BvsH/yaNKYpnqXa4m58wyOs62ZFz4SNi5JjpIeAcmRyDIP1tnpYFKHA8tTzzS
+sMZzNFS7RIe7bctPZ3hCHOQC4emKLggcF0nkI+kyzjyqWcjbyPp+s0m/abtOOcbTscUJpGNZJK+
/1TkrLVOkM5+8mtws4xB7cbmpDsmU8NpofwwfoNBrqn0rTYMga/hZKFJnHc+l/a2z85SDalyTxpA
t4kbjPlLCL6ZZTuzxnpXqxcmtti+fUz5EnrM07RgKegYIzqh8WGOylCmm2hZScdWg9YhmdzKpYaM
MVrb50J6PQq77ojMlHytIYe6A7aFrkMK1zEw4xgATtc5x8O8l6iM7LnO0KdV0X61cKYjuTVV0wjS
JGucwZ0FPuC6fI1pU2zPYrTxMrS8d4hCviP2+96SK7f0py0MBuZdE/7pngmbYnIk/cQk739iakW8
X0K8sd1IaORPvD+EDYluVoZtjxJxT6LmfExzCuaALyw5TajaJ0h2wRkHmvXvVZit0s0E/YR+Zr5y
J4MT6oHbhThk7IsUehFvQyFJE0FWy+wpR37WmjTVw4mSF5wfwKAf0Cv1E0KCPJf8iPokRnfi4lTJ
0ixeIyWTJBvvdSu9iJ4jWnVGrh/PzL9sxf+fl5GjxoM9CelC7Gg+I3yclH/SqqkZ2IL0sYG21k76
f9W6OiqAS6RsrvOPXlc3PWBShzd33nWxXgRaQf6WBqdu6i9QpgygILq5dXVMbfRP9YM9r+Qetv3b
kZ+NttaXtMD0v8Ay+9GMnM66yDgdylqdq2uPn+ahxVXQzNaSs00WW6NxrtpZUhDxKfQ5zNgxtatk
kl5ST5Ow+RgMatUXmkmr9u5efoJRU6ght9iA/25U2r5PRsObiZZdM2/z1llYW3+PhvfpUrIYptQ5
JXkCVT1OEXoDbzdnbowKG8VCXFrNUj7KGaisLatRXGFJRA8EZ577AMgbQaAmE+Iw6cBpnBZ2FpQO
QkLdjbsWEfm2RbBMl1YX+v+1GO4eK6r6eo7JA5vRn8G1sJ53zs7raB31KYo9O/dmFO4yD0DZXLUk
BDqpAbldE/XVEx90XTHSoO5kqNxU5YI6YnyQh2yWonzLNuqSPgtHN4DLKDuM7wozswAAOYvMpdzm
FBIsTG96vOo2tGoSOcUBYfw4LhY7FRcLFt8d9U1qMGex2uHmgW5nfABR/oHqPUXyrD35X2E4iJB6
nLvABHm3CU9je3HYJWk+sI8izfVtg4KlFMxxdWZX8Sp1sJl9ga5dkeVF1wpKgcoBIgSaRLt49UXu
su6kgErwmvrR533ueXGu8q4dDGXQiNTHPBNm4Utrx1XtJLDKrT+tk/RPmFUrJgBr4AHLO1zEHJ0f
yCg1OxGAIidcgiCTsRdffWPKffZd7ktCbZvUZC9Y+eKaoclBimy51xllZY7UBlc8yx93Jos49zkd
mS1jmzUIC5jjZsSVn46rhdhRrb7JQnEtBsNZ/DGYuR9oMXkhF/NHYXvQaGVUjxCHj2mq/EgbarwB
Z5PBUiFRroGVS2sJs6rze2/UopzWh7B2dcG6I+PW5MIyjNX/+YDxyt5CXj3BDCwdRSwP12D+wsKu
0vM6JH4AtA3O0o0jpYFhT8JM3y+8FphZqyU7jbbNUY7hv+bwLRT4aj4n5mpqvQTd2fmvGtyePc6J
lryZj1CmPgXyi/helpa2RQXokwQ+BfGYPnksR/1XKIvgLudPP/FXuKjaZSgMNPmb6tytq1trVidV
S1IcVegVf40kBO912L7zc/rkrZ+eX1MA2WF1+aahYaxKd/IoftSUTLMBwhC8Jdz8g4t+8plofzcD
v4XBT1xFo5cYNor7y7ZUVeB4OjvJslzcjXUqsVQHVPK8GFcx8pp3OT1C0YRBsw52LotLCNgOwMAr
J+yWE4/JnD8FY6xExgBYFzPiWzF57I2IGAdEUFae4igVVTHKKfrGWfZi0TReddBO1tA11eMkba8x
Fs69G0bWnMsd7FE4YfGEKfyB1z6RmaQYFKW+B7KJ1bHnDu7I95s6GA4/m9dLrdJ+rNO7WoNFPk/4
SqX/1QbIJtvGODj89iMUbeNtqN0tKPB7XoSLHVbkBBaQN9dpgWqooydtsJ4rqsj7xBKvK+Fh3RWA
d3amui0VWoMAL6J6ztPS4Ev50LX4hnK1VIKAvJbURLxmXJTV6vNWLOUqKhfQeV40qo9ZR/KAack4
mKdrKH5ovnOLlja274Sckg8cb56imNxzniSxD9DUrUYz8/diS87NgyA7xUaKsT7vQ3E8c8VSsGq5
/qAWxI6a+bsNeguxVFm1W8FlkZevGf0paLTC0bRQfYE+XpSFx3xxrFcI20uP7+xccjKTyFeXSyw5
7YxI/J+svxODgRB8camGfeXFWcCCl4Lf6yZ54TuH3hax60kavB9pkF7ITOWdTPGm8fhvDSKXTmUl
qffmVcBI0MdVXmOYQMSkBlYN0r8V17o0uw4gxM9sUeYWxMbZN4iGYtJjF9QWewznqweFgQIW6TN4
fpnxlAVEu1BvdFn0Hwboq+1f5vv9gtv4qTeuqDadbW7RGM3+IbWCsuCU4q073EVw7jJG2/xkyv/I
cJstnDmHC3bmjERW7fVuAmIKtOHD5DI8YvEMRTCRzoNTYnJvRQV/OuaKD9eJbsgelt27YQ4v4ZV/
xrfkNqdaBQ1FZKXgNUczBdRxManUHHUqEEEOgdELJFRoE7kARAmBpGCc+R3569YHH4c3H048177o
dx/PesoCbJaq2L3Y0+mv33eDvRZ3MBaw/hGKwfDWL1zR1SsUzBh3N1AmMiYbRYf2GsOmx7/IIHOe
cnbqmTi7KO7Dcl2UhC3aedUFdDg1rj0NDCEW33NUvWeoLceT0xAK9/KsnR1FXrqfb8ylak09DizS
ME4mjC7ue5lWy9LGBV+AwzzIO4YxSkIdxyLUSk4HrMo7NRpiQc61fCW4BZwn72fku5snfa1XS55+
jTtBKnluagvCtsLdrmX0R1ttQIuVJ71kkRmyFDr/J+D2EWXaBpE+7OeI8SFB0RLPNHtP23vYv+Qe
5IpbfXq6kyQjnp4n6n3yOlYWkZfhoxCz48ck6hP9LlbH0zisdGhydFFJFa79B8XWgsP6gh+rpJ5G
5qH1zVIGQwWDQxFwRL2MzbONe8+56UgV39CBEri0wRtrnp++FIXLKs2yvKKXMKBOkEh97OURgCFm
G+bWSbU1s4y67GPlgzz/NEDRNlNLjt/d/hRalrNyxKU2/oK48JM5ABFjAUMWU4rghqkHdHiivmeH
1SU0AUgzqy2sJ62OmZVEO/0OyoVvMFrtldI8IwI1mBbVjqE+V2mPm6WIwadStccygdTTXWVckp92
cr107vgagZa0bOlWz3Z2gO7VNueB9UdjMeSyQdgvSb4ZgoG0r/t+zHsU34rnO2zIiYwuOTBr426/
F2JudnugGaA10S54K8g4NIqnCUsS9M4qEF35SaxKE19uvtJF7t3Jr5BHADNKz1cnFaiHbT/WnFZc
F5DRrrmCnmW+jox1pEij1PM+UOgX4m/bLuSBrw2xhZyYQnefMaaNtfBBHhX+2cjwwpruTHCRNe47
l2oRoIpyNwqB+UD1j0qCkmb7Ami5QAcLhxVyDpqdXXnNVSa1u7hFHn/OVHGNZ6JgRqnUYi/ipR7H
2AsIES1uL45Rr8mWjLNuLEYsmHrtDxHwoh2AN46IDBW53LR9QnkY5NMN98l4ctNK/pDYbHA5Eayl
YkkM0hdP/LHYH0Fe4KqCxXBjJr5jR3V8t+tVKwhS/SwJvjDjyZwWnzzjrLE6PXYI/JQ+Ul4ynjwV
J3qXzLZ5fE3vrCC5lypkNuEl5iRCeZT243+C3DUWqX36dnGJpd7aNpXZas7HQjOyQwMhAxUeuOs+
esCjZihl0+asNb+thpA0HA0W+LIcXVPOxkztf2K9wJe1DeEj2rfX9GvQ9LVlU7RPJXg1+gBWeGxv
3+BJfR3Uei4rpRMmY2bjys+VDRN2EqeBeGF90h3J5NtnmyI57emYhJG8yDUw+UpOb0iPGqrm2Y/f
w5bzZKkrJnapY/c980NFRUJbmIudIiTRXbryOhvPqfb4O0jJsJMf0+lqzJIYW8/IcfGJpVjTuNZY
+pm39G5bTLouXzeWuJRNy7iopGxopLGQDzllraivQx7SojMuvYTHVEQG9/J/Q7rC0D9kZhY+SVyK
4BH/ZgkX1B+2vrtmKI4VCbiY/zvaZwd5zWSLJ86GDYUBYwv/SuXda9Ii+nqFOZFYCsiZ7lj9p5EN
8JzTpgpuLQw/xQM4m2LaaqMewXIH8GdR24v0Oxp36KsVvvyhoLQ9TKS5TmSNBFfRxelFJjkfbGvM
2ELjifZq9YqxQ+vGThWqiqak/ZgUbRmTUzJldjPoTHICrWEI0jwbYMu9mhPUMXKieWFIP6sgvpy2
Tl4C43i1d+Vssh7VhSEYxV28g1NkYnfEHtm8okI+WmD+/zPmrv4OQtzvyL8LFHLh4gpKSetUVH7P
bqv0Qz2LCNbpAJaDj508bH8sa3uEyJSQQPj4lXkf+oKlSmDKk2YbEFSZaEMK2oPUnUm+DfZwiX75
YhtYVvaG6TTDMiPTgj9MOe7cA/p2royuLlYEPa7BF6CcFtHQJ7HGTUMi38xZNLcsGiSgCIgcB/FB
8XbnWUhCD48+ZnRtWtv/adGztxzfZke4GlA0eHvnnsdoU2qa88ABfN/jX48i1akzPqTfcTGJKyNH
GFyttxSb3eiHT9cGbFraYAB91QnpOGBD5QKwubmt1VjaC7j18N7IUFsQBQZhfEQSEl8BFTtaT1Ns
hqubeO2XoZd7UMA6S/YmosOl/Y36bXeDh3SGiUvwbQdDUHzMA2PCRy82BNeqne06zWTjlvuKIQ1D
CweJUxqRs6gAnUjGOFEh1QiRlQ4urJvoXo6/QXxeogoLNJKYoUJbCXyBD49f/KV06pFMhLo2M3QW
DO/LcuIW4SZXSPHz5R1Ar7+RfDS1naXx3mm1uP8M/4neHLA2Kq1qF7qzBpjHaPtZFjMvGGFiIIW1
vOHv1X99CjzqQoHCamlc5/rsUpFM6LJ2W/GysQabHKNb4qPamvdSXj6bKvxg7Tej8eFMKzLk2Sab
u6LFJKakFoKU14Ffw933m10XFnvwFcns3+ASzVn49E5m//5tKgPa7WKm0wtkfQUT7g6jmZ+zMfs9
yHBumlXB97kY9GFqwAo42R+971DRqzIv2/w7xbGdDqDegNCKm8rF51Aliny0htsPZ6iZmsjAYxX2
94+0POv2BAOHLiOWGZVTxtOEyyoyPFfuv0ReQC4U7l0zLYwh4c19UVN8sW9OjI0zz4flmVRdzrE7
yIQFV/Zzfh9tzUjBFFaxdQarFfgeAkl+H39bSV6aFlsyON2LKk+ye6g8tCVO9nxGBJN92JdZDIEG
ZSdHb1IJSJoWIMiFNDNqnix96nyknLOa7CaR/Bty0BJm8jFA03q4QlmBs+ZnFiYa/JvFU8AZufg5
VsVahhVFOjLofzainpjFVkA6lpCKlYabqRdWVvsTrB+npc969fH12CBC5FnSDQJ2q2UnrDxf1TUV
Xjb0xI0WKODtXyR7dKA01LxDFxuXoF9R4KUNb6thCegTEElXcOKK/+rfxJBONX5Eivi1bumtI1j7
edfJ/uzasBvt1Ach7iIIGmQE/mRw9twkPd9Fj4/IbBRaWk94irD5RllCpodZJfxSxdH2f1kdWfnP
dpkYw4a5Hlk0KqPV/MkI+Cj7ckAaEKu2YhsArC8PGOdsi5T8ia4iBeM4zBAic2NPA31YG3uFmn2N
ZiioOs+UKq6VALrWEjV1DYM2F89f3FZ/ud25ZF97WYbDUCjK8POL+lcq/9l46wyqFqNCNGyUWNZI
XFvLirUOtLXTq4ccZBwY/hAV1IqmsVS0jv9SD6t7u+A8QZpwQe+/pFE0XbG9+HKGrSi/Cq/0imRp
g+LI88/+gyat0aJchXHrYK0hG7KQXWTMTnNAXyDo8carwyT7WliV1Po0ueembMgwzW9WYOwypD/V
MiNrt1KiBdPRn5cESgHCvIo6E2s4DWuyE/yb6+8fuJxt1MuzgtL5WsCD6O6DTDffXzofxkSlzR2l
NO9onQwcNy4AqUo7EV4V6KZ61C7ozgbv7KPa31+n23zgiy0sfAj8AhNVMrfMKrGgkDDaP1oDDUiU
a9IGuxyf0EmRVcTMvHgfck4awFNjM7+SH9vsZbQXobn1zku3Hz83Qlafe4hiizgtcYsgZB/Rjb6J
qw80F50nN/lJtNRWfB9TJQOWgQV22q8Vx/m8VwcEg3cVhvJFg2XpwdddvFYWucEU0wK473pBoLqz
ey1Pi220ekNq2FdFwzz5/UeprPEn6U5GjbCZhLOx/nnw60DtfAoVxAHrqF0jz5RaPOi2GyGkMOqy
LauhnpbeVq7xUHdAyeeg2z00/VfQRq55tPLfIiMwkFcqJ8Lq0eONraSrI0/SGBhDdokv1qIYlpyk
anTz/fcC86rQOrTjpwQEsHvUQP2QllUJj3hZgcyWyolKNx9eYeau2K0thRlaCukykcEL30rCXZbk
h/iQ+m+wSL6xGSIAWg2Q7emgT90rmPIfN7SfS9pMIxjsQJVmRAV/v7mSfPXp5Ei9e6/xXFrCUaSP
o/jt7+M4qymv0HzvW3hWJrcpSRgfYFHN2H+3mIK9D2Zqktow06zNlUTT4G+mqkswomi5qkZKShdV
XOBG95J6i9KG+6panefWEi4fsM8o32+G0RhyQdBq9qjLHl9IdBkc+IQ+E7vQGR4gCkeEaagOcPgd
gRYIAc+60s0DWjyHwKrFGQL42IVNKYa6KPLxSU9XwWnZb1nhVcidyE5g1lclDrj0i57eEDj5cgoO
o0WJSMrbcR/pWbuvuXnAyOK+bD9TJxjfy2zGfeh6+fbk7cqqjZtYqOtLB7iJCZXZV+YJdC8ZS0lI
ui3qi/1zx27/hdCJ2bCMkOcWXob7XroAlyWdWWGVoLVicVe8tE2GozLioDHfTl9xMqZiC/egTj4i
PIO72Yxv01IrE2fUiizO3F2DWaHRPgr8MW4LT7S6vVkNJD8XL/G0WtWVVvB/kUJz+NnL4iAw3lDY
UYVtpWlROzmH0Y9rFzdwzMvzPounFih2B+PeAjhM2vHxJFZ1RjlhmoylAR1BqzycPdfILb25P4Dj
rT/cznaDer3mvzmDmyxxk+HEUMov4GR4QqT2AdytfhD+3KYztczFjlm584IkkESrv8LESLgsd+VH
gk6tDlgUgIz3BWj1E+6zoSIT6M3wrMN9NrwVJ8SPsIPRU3z+sr35CSvIko5/NoowAOqkqvjsQ3Iu
xet8dg+YiXdxplnBXUNRvnLV2p/uaChT+l/TU/kymgLd5A219LHYEg3I6GNXqIZ650Vf8+EoPi9q
OWS8kweCQUeKA0NYkpJ+cAXm9t/3NtmGe85t9/xBdADG1I8QGBQqmPQyk6XRVDyC+teq2PDP+qnC
JNnJ7hQIdLLak89y6BiMV7xRC97TMc1Dw4lEjZi9lDMnEgVVhz/ae2NvGfsJ/vNoxwKFdgmK2AVT
UXxMPh41pF4UALVE9lnITqZ/fduUuyby8B/tj2SR3cjX6tcYS7VqA4bEeTomDg67jg+L+OCBraDI
kWkfxVhAEj4kq3nrgiW7E3D78l3VGrFKQAf1SZdGELQ+7WiPqLez+bnLrs9JDmn5cgEnjo9M9rqc
bUGXwuoQR1X7mKhL9GP2LEb3WDIhVLLFvrRXrX17qW0QyYAkLxRSDKeMeNeJeedOUzq13HrkhLMG
ZwifIWsqIyu/ds0SkuKqv5VbYVTzv74Ctr4MzbFf2BroGBtJC5k9DJpwZGl8XlDGCz6YOIUg9jEp
M9aWtGAjj4tLYW07NzqkMrn9D1HVroYQmriN37kD+shYr+VZCZgE/tmh0G6smjMDcrLzUXnTaZWn
2FmCWKkc8261Hn9VFcO57t4PZFT+FKJmS6zvqJFy37/uknH+yIK0kUH13vr8WgHmySqQ+k0EfImO
jXyu0ksHAQDak34TQoIrAIhyxr98Vr0HsSm7QJutW8EKKCszVMW+lOjRP7Fdr4SCuQZHPQNwGqBG
jaVBmlCDeRdN+kQjYHuCQAUkHj+LDzeISCrBmsSAzZXpbJLbOKqitxkkAFGp1/66jEDv4H84w1+f
VY/2NO/c2XC0JT9PH3/YaRyW0dZX4cAgAubLyRdqcNZIN1i769CYp+xCqHqF47jHASNFAUa4EK6d
YqLMpS4aLBpIed1sMVHYdNgzq7Bkc1FsKt00dHnFCIsaEwNCthyIOHvqVHjDWSFHMp7t2E1bCcem
rXh4F9S7dhIGr4fQqHdOWAeHhxQ6x9jbgX2tLVsDzy1Im431e4VeHzPwToT+41AhQ6j6ydhRWIxk
vIu8mcTk2n/S4xfoR0/o4uHryrsXDezr01FnVtjf5iPsx+rMOuJ9NkHlVin/EUROmEwQqKldfS1o
PdD4blokqEV+joepBaH8vm5/LO+kKq0M4Coyk9tmyzhQFJKA4fYdc1mw0jo4Fq4/QvAB8XVgoQN2
imUc54VgThI5WoFif3NUo9ObEa0WZZE+hGd2X1ssZ0eTmk0Cek+1emFIUh0a2TlIXnHiBK0lPi4r
4NKA0pyKjJ5o53yGgSuYpVjL8/7iMtOmKH5tmb5e+dBN19GY1foOJDQL5iCcAviPcPQwVg/bGQSX
QzKhZYol5Zns4KcqJ7Ui3k4yqC0XdjwMIRX8GDrvU5iRhLGo/06LtfJjIllWF2cOudwWGsyNt1wI
1aCkXCahXo7jeRXvTOkz66YREs80r/tuK5XvOkv7YlhMGdwHPT8SnWOkWhM7tVTnyXbxwXYxA4IP
3gkvHa3Vbn9SJeIhDe7FujwUP+UxkKWVjM0kyh/b1yyZxbenJyi75Idt7cOxHZwUpyMxZ3ueCukH
kQy4z5ChCMpaVf1reLcr00kdN78Q3TZvWxay94Sr/4CD8gYN3SpTJ1xTaiY3rXO94XsvibWfTsrO
ilQBx3rkB6rkeMCZLqPksJ2LB2u4fgVTpVSX52mK9R7hoLmLhIvthIxScbk0551l3lQk2vSqEu+z
X7Zn00nXF/BA7rmhaRwXqPDZeVf4kvlj5EIRIc3farVTB8fWXqS0CIgET+PQtzlD55w58F+Fj3Sy
HwfthQMd6qgALG53x3v/HJzkX87BBhZhA1IE51xqsBfzS7uTo+KlS1UFBOPXF0J4+fhu2Chu+otG
9/UVUiX+XgAOzT+aQcHC9TvmJReqCrwY8wbABueFnHpBANgR0OVkZjCwkBDKQiRVlnZCDEYYV3ko
xTw/xl2KkEIbz+P1zT+7r71qq3w+60i4M1PitdkKShJYSuwIFj47DnB6HQH06x5m2WCDot3UB8cJ
xTNzxQQOqwcpc61ut17pknN/0QjpkwOzASzQ4mSCm8JWyhx7cTSwgoFN+fmFJ+11aDz6rTU9BN8M
SgiWCjLOPfFvWfiQ0G2/WDdspmEV0dZa8drao+FthtZQqKuZHv/PbWVeQfOKBBk+uMnAeFJ70xQk
RSvTUx7ELOBjx+Zq+bv9FAm6dKokvAL9Sapobq1goVfhSe7P5qxW/OKDeMuHAX76w/JFxSjp4N6I
IwoisNzobdR5Qew/5pWt/KuqW0m86cdCm0zphZv2tPxKuHJ5k34FqadW76y/quptoO8q8pNaGHRc
0S/jsfIvY9amCE/ybRzLuDg1GLLly/onctrJU18yn8P0XIg2QbfPZ0CcFPQpkXwqSC4GxQROl8yc
SyKTYvx70Wp6vAYo4foBY0L+HPZMbDFwuzEz8clfd0UWz4OOrLZ/688QRoWJumQbleKG9f1Hrrgw
g3tvFDVjWRWH+TxE1P+5nsyUP0yRdTt68Ifer6MVq5AKVfHo7Oti3bAFGJ8IBHY+/xj/sv7R86Vf
LwLyw+r0W90bvBsdUTO3tsPxCXiuc/gupfXnZk2z8Lv7xYO15feso/rrNwYgCtd97iBCQeIplac7
rA2j0WQDtHHq35hLZHDVowpCc26TE0w+qqCqvpZ4uRfU/yn6Ac3RzKqtiVtPILnOeyy1NgBdaFMq
5zxtlhcJ/TVidGBz9zcBK686sWSwN+W7KoeI376tqELNDWFuv2WOKUgatkBIsrGU5t/F3eVAHz8O
mlEHBLQOvpFxaRqb+feLaJ4rf3p26FUVA1aFY7RIbp+Yb2f5eIwPvisLwrzAX7dqT/jTLYmmfdxA
M8/oitpar6qDNztpu04twjYd2KD1h0LafBG9A5XpqvElIbplapFc4RodOJnyONRcHFjL1kNzJn2Y
tUQEWdeYUIs6GSO+GDW/15hZNHRUmIHjKxMWbRRYiDb5Yx4Q52iqG79GW38uaRD1mHk0p0ykJNmb
p4ZGPc/KZ7ft6eVDXs44dDH7x/9jHWwDPGCVa0m1UlgmBkXFsdBGk/xdfc7s+kq65q3Bzko4GqF6
mhUAC+WKZtSrbeB6BJLFsgdBTWiBmw7suu63PYazJ81r6S9Ie2N6BkziBRVAY31duC0psDReYYDM
t3nVxSnCE+wKEixLgLKHS0TyxnKMFdXsGBam/esONIjjy0s8ci+kgwsCF05zvM5B6kRuKdPjTG0L
J83PbiWfGmVGuCbBL+5uwq4oLVlJCC7rKxDWXo+YqRqjudpu6jsRo0iYpCWPXdLYfk9qPKm4YUkN
nARmvwu2BCRDxiwI43Dugm8CLcMNpdzTLMHnL7DMxvtJajQXijIMXhheu+YbCXoDJScKG8ohp0yK
HwLLdwBiofLFR1htpqN4fTgLYXJY0lIOMJJZW2NdpchDTBOjBvWAPBS9nIGwQg81mluSSlLhw8Zs
irYEWOP7pQLcDJpbxh78rFVKrCEo/iDq9cspwiF6pyiTR5HnCGZeedtdwdIinceDjzWnKj9x7QEA
mb1RilutaYgs21cWYQhZ1EkOjXXyPZXJzT2aPgYZiOEBDHUv4ngIBb7dEBHvm7s7vC3Hptlj4Xrc
HicLqKl0/FVN+SNenPq8S5zNGOMZlWHDyKMimHMpCaYmmTWZa4ECVY6s6Cf/7cj3svmic452vRY9
4EZkylnYRHmNJAppi8rDLU7Ke2FF1ezybvAPV0OpTTiPIgUZW/IAxyyQyMkwmN3cQ5woTknxJ7r3
pHafdtltByj4JyTygzYHN7LxO0dtwbZuA/ad6MllX242clcq7J6n2B3kT9H4aJzZ6ep84cjGmehH
Q6UeN+xtz6EknqJdugv3vclt+iDOJoQqc79nqhFWqU4o8rc/N8wmDADJXGRlgdCZ1hK0n2tlTuT4
U9cVQD+T0Qew0VgstiJPP9D8SJJ20tsxt+gh+Wu01+hvLs+tgR/itl7PQWGUtJOSit8c69jvVcaN
OtPu7jeZ1xZIsbJ0tJvG0nu5301SXRjHg6oeIKh8rJnAZKFjkPYBPWNjiz/PDiIMu8ugk2ECsgYx
LhvoeI0V3jEBSBtxAEeBg/qZ1slFrEAqfOf0JJfAfn9FUQQtEdr3o3rwCZmwmCZ7QfU5l26rcsvN
6zwMK96/DTqC69h204QM0d+vobdX3Tt6JtBSFCYHkGWtF93l52nbGRINPzYhAHQ4SfNfMxa/8ezq
gayrHrgRa/qC3lANcdDAER1YIpcPWFATUMTH75HVCe/t1saXbW6If1ZEgdjIpTITVLjJ3ieKYoQm
nS/+jT6hCTMCf9+z8nEu9+BVP2ohoYs6n7jGXc6qMV1LLJEeWKvr2r/+wvTMLwtw+4Pbv9cH0RwC
0gqRpK7bqGkFURRBJ0A4kMmkeQrqMQL5asAJK1xPyUUKu9mHGhzDLqVHrVDdycPIW3v4WAWuXspR
Ar0nLEjvYTiTQsecv3hdEgNT3a3QaQG9MMILqUMsx1fBY84SM+gbAuMY9h6uX9qvRodWpe2xxIMb
EHMQUGzROjsLBJsWE+fEc62zgHrawBrziFP1snaZeBNBUp/f0L3kyD6HpfQ7PDTX+c8yTO7UgheP
d9BWcNgHhssvTavZ7qRVUfT+6hb7szi6XJhTuu4ZeSw3PADanwP70EkWR2sQ7JkH9cT98hx91Z+Q
Dz0TbvcKstaSiDWN2Te78d7jjh+/tPWqIGdNn9IXs6IqYZBpQwJBkSk26laQi2xv7WjugQAzpvU1
OrhoX3poMArVoYOBVsFrwX3OeZcESr0L9iUc1pZUSATrjpzw1GksBzFqU4KAH5EfOyM23dJg5F+s
PDgnx7W9oKyovwDDIVnCd4OQswtZSAB+wDgAY0kn5nR82GWpK8LAgF90e552OEYoZOHTDVKOkQCk
YeOt1dAAsFb+thvZTaGoC9RpnTQlByvqAdRZ50m+rnesuSqt2PTOMKUUkyrODpFU/Ggc38jPoiXF
iGc0cHb3J5GB2rWCxGGL584es96LsFV5tXEBhD/my0H5eyO7BYsoIypKW5QkShdMlNiVgCRjv++5
jXiEXSmZn+mgRkYGf4QI97eifZ4NRhnpPV4K/f25oUWMe+C93A5g5M0OYlQrp4UOjNLlA4NhNSjG
Vsc3PR46xwADZh7SkE6cdgzg84F6jK2K3CakoRbdGb0HEDFsFWsKDc91RCNIhmSxlQ1OyEn9zztU
HoCozBJurj1MCblBzOI1o0JR80L4ZHD2tymD2G2fFNm8FTHSWvMGcvfqaTZIqMw7FUAaHw9WxT28
WLVDPXFEksErR+dBCcPi5dNUssAnTX7PbELwE2sO79VOKU8+DvHyG22JN7ObhT1xuv/AfmShR02v
UoFVDnmbPsritV5aekvfUFyqvB7+8t/Vz/ZhmH21/t5CPSTN24kxXY35Aw9mdXDns/XfNhaJSLr+
uDb5HaBUYFXddLjkB9sTeGQmIBEoA4SyESyp0rrK81GzHHcyQuMsqXCSzBcrZ+J+pc93KvpnJUNR
S+Nd/JwbLebyhRpGXjoKVxBSJenKq/MKU9hNPpq2u5MIZv56duRVPM3Qxn6Re/fvXzRh92wB+ESM
Tdxd8XZe4ja/UE4ROZ51ggoYoEU8DsE3byo9XOL8iR0r26qsoVsAU95oqVLbOx1dVZyv2lGYNSaQ
pL83AfSTC5EcT7lmGYvSZ9unZxZDMwQpFJ3bflY1o7DTSGbT7pdmCjP0HLL54F0NeaJ3nSvnk9kd
AiozqUWfFgTYZxuE64dJk/foDCRnz3AovY7x1UA5GqjE5V6c3EiPR8gMXBRCso2WGpxNa8c3mft5
o9IlmSwds7GCmxGlupIjDpdWDZQABnEF8hQgOOm/EFpUBLsF6qfYfdFiWv52BTTNxCIWaUnKtcp3
12hiVrNr2LPM5v/7j2n+INnIPi8XdoaSatbyyRrG8Ejzg/S8amIt43SHqUKWosWbP0hWr7Nzsxu/
w6aZwYZqcnyM70gZ+LaBKxfo63evY8o+Juhnv1Rv4GjaP6CobtlYHp4Z+vwd08Fo/B503aJ/wKci
BFF7ysLFoGhtklKHHjIYY5JjNhomceAmScIQRz430W7k3nLPpRMPTgiPUoIAa9I4GReZAYqGGpSp
pXtCdSn6MahQnSuoZEC2cHId1slei32vwHGCGved/3hAB9B0aXtvmQ238bqDiHOjiEY4elRJdlmN
E5aFZ8Y/+MxYuCiVithJi6p/nEwkUo/Gn9SFPXpY7GIn21+Z7cBL98ZBFhGcB2Yx5M4NpD0liwDN
qE99QD4+tu8a59+rlyWdykKfd/QrBnNe4b9aNpNnkxJIk9R9daMPWlQQYlqqy1OAS0B8prMQMZOE
T9a/D1az/QjIT1Aofe6e7eALFjHeCXI6h8DYz2uOHLAdHk/eu/FkiP0zpY4gfGZnH5iksxucluCU
OEYH29UPp7XyOPbbSoUXwOdeF5HeErLpJ6JeAsKsRnZs7hnGD6gjEU678V1O7Fqo+2GBoq3Ih0qo
FTq+XPFLmfAqvsxuhsSSf4L0BscVQIfKEMBxu66nrPW+pfzQ8I8EtsZG4NPtvZn4JN7IuF13uesv
szryoo2PqxGOoUu2C1Dr6EP3wx/lP8L4pC9xC2+7hI+6YmcKaqDv2ZEO49Xekvm6Y8Ec70603eSZ
ctFAvgR9bLeM4HxkrtkmiieUfdPZD9uXqwcdw+MINwcNYlmYN76ULlEuK9YVy95z6CIlFMMwqHMz
0z8ENWjAnadWnArPyTtKZFz+OKUpaD4Sz3wwn3R2YxpFf3Osw+JvkiTjh1QjUu23n+d519iin/lc
pyeH/tytBWxtd5QjFCTr+fizbAMuQ4pxBLs1sssEAO8G5KWPXj+lQ3tz3+nAi+sUlt5DLjKBW3t1
q5u3djw+uaiGQKO4ejYhux0mCFsCfQCxmv3NFQd/h92+etYcQsTSDePBiMBoHy83bmlLPKvtR0YQ
xMNk1DEzluNi4Bh7jC1TZb5etD/rv/LaQFroaTc1n50npiU0JWDiOrReUkjfoLAip1pX47eVgWih
PFb1jLyQs89nDegWchzNZTTD40oWykCHPFWP4JKOfMrDOVjwavygWf5cvZ7N9NgOvKQ5cwa3yo7h
liXEmBbaGuwejIthTIKKYQUasDQm2jsuN34xfJbmTBWFjmck5IhhFozPcM+QbRa2NiqY3SYsoq6S
hkyi9TSf7jbjGxSRdSbCUZ1Ok7Q/y0LekK68JvNpGIgVivBnXcDuhaEW8uSjq65C1vJD5ndPY9Ro
yvS8ejEYNU0aoC+EfxiHJOynJZ//oEC3MBFxV6UNoelj9U80Ju6Zn4PQlr0Tei/pbZxidJJAq+Q9
ZjohudlYdojxC2NJBGQIXWLS8njFlTK9V5ANBpiq+AFklb6pwViDO1PPuCnNVMNSN3hz3Jx5PtPk
1YtMACxzMjOP4Mw4MBOSVEYJdvYKiCN+QpdyjIZVJD/CTGvyNgR3V5nlQ3uZDO96mazB+GZMLQIY
3GikxVX4d3nJ17o/4FYrv/ZGrtoQGUoS8PvMXKDKh5luOumPuvQTTgkAisa1Qn7hlyF/lWHjfHKC
Ypyg1huZMq0vOu3rURuvMEbm6aE38Pz5Fe+5JzraqCjPoUeyDmqJxUHVR8Gekaa0hFQm7An3IZoN
bCRoIBe2K6kartT3ZGHD1UXT69UleIgcRZqDxqWs2aVZaeifbCNxIFQAvkLMdbSUCbTUQU2dfPQx
mVZY6NtQYnlNBF+SXrAoPK4PdyauocdavHbYV5Kr+M5mCkDe/FGKxxWounHfa0PDrHnnmrW/vdec
0V9mKDGa364cxkPuCKeh0QJJZgdU2SiUutrUvznbcSVpR+fMm58kVrjPyJZ6wgPnQI/G0Q/kevGU
fWJZN+4lZpozGDm1NCQCA2826L77+TYM5y38QB8UEny3geatDtxMYyNSZ3CRA19F2Qt6RIfjA1Ej
NYMr/dZVivXbSqM7IB5hqFgCXE358NvsSsoD92q/yah/aHVUHEF4Ibb4O9c9j2tKG+o5d6toW1ZG
Tnc0jyKw9RsDw9KWXhe8mpociEb0jg5rdnpkPsw7sPwBvfzIKn4Va0c/wwk3lYtxKgZirD6SR5Iz
iPOK8CGVHDpoSBbk2zkImgdkS1B7vpnn8A55Y6amBnwnbNesOuJn8AzSEqm0Dt7E+EbbPCF+Y4x+
PfHroePLhzVVqJrWwu3kD60l/c3hHqdD0Zo8Dln4apXFGV5MpRvzgVIfWeRbCXqKpe7NzU6Xo1Mx
o8QFYruOiVeoMVUpbqOmTCGirNGI3tHQ9ks+xoVpgndbr6LwRCmlBaPEwidTn57pjVNewtr8EIqm
07IaNPdxz3PWlqQn51D3ariVFnOdn0vO2s74t9QE1K6+oYLMfDLDNa1VRC1tueYuzCJ+nQWTrXnw
V53nf/i35uh/mNxDr0A1q5Yebn2tX9aajfg8d6Cu8P+XZ0QtNtNB6AuLwzvq4lsedWAf5n4aaJH8
Wci+KxDIMsQgM+24exNz+5S+ybQ91etSOw7xEqoFSUvwffCRHSpLaHpRcj+kD40CkEgtJTvQLixo
Z2vACwM5rWhOV2WNgE22Kqt/LPAtqRcTsHIi1JXsR6UTpG42pAGg5oL2xUlKAKli5G5cxD2mJH8W
KrhbWG9jjlUDJi54Q1qf3eWLmDLHs4BSoCuctzgMhqDZ49dxYrsBYF3Lqo+M2UjTv6uuS8veftXh
T8w3tXbFGsOx1ro8m7HiaWaMEFdxsmWCAzqehqs+i/r3NmhhdfDgeuF1LQkylMKWFsQqIiEC4g0a
7cvroqaBTXPmS8o6QfKR6jfAupVxLCk0Voo6FfjZnNu+6rs1Yh29TS3Iwn+rBvpFFMNYQIBCALC1
HPOBtN31708LuwWIO7/SEirX3zeGHXwAxLAou1HPku3KYTTb5wACd9OE+1I6kakHKPKTYCX0LrXB
D2GBia/8VcNSw8BgWhNRwt5qGJMjwwMvFiZ6iixIt64sWklbJyiCt6V0zHCp5bqq6MidZAWG93CE
zyQ7j2mZV8d8JERYEp4XpLqNIVnoPPCRwbti2mlpWy/aB0WJf4eEbNZsh9gpZdnk+VSFTw83J6D4
pybXStp5dC4zR1v3oXId9lnQ3nWHso3NJvaXdRsyFwZ+V39cPw/C+45HZD4viytx2rHtvP7Bug4O
y8Gsv0UYaE857Eg1jCyqO+eh908x91jK1jclsPq8E9oalxJYCBoINMmNI2JBoCeGJRbYFBhPkzdH
WTKm9JSl0fyxSIOLKud+FlG9hYQ5xMoZgj3Cc4dR+vcmE0Mocoo4kWxpuGzozhmG6X9xY+fZ/NF7
BvNObLFquZRlbinifZwoxCYUKFYz38vV+TJCxpRcSlPG+xGvY1hweGPsiq9Y8A3uL+PurnDgQLdu
NIm7k6XgANhNCTc06pgg/B9yzQwQ5XE7gcFqPBv128NMwM+MwDdfyhNTART59LamE4H92YNDn8SL
l24iGJThWu5VHawHeEkYSre97T4AYVRG/5vRCPSKsOOnpLi0a7XiwFOX+173LktKqEdJcudbJlCg
pqPWI+9MH3WYysw5I+DXHGzQWfkVJVQ8q4jxwhr1HGSgqGx288y5WPnS9C/uVtnzAkzHtW5ExPBH
sirs8J8DRvKPWOPIloEGzCQfAbToIruCD5tSrA9CC/L2jCAymB4c16suPryyD3M6AHzG0OlAytLf
urXj9qutMbV5lL2r4PCwQThIl8grOtpGyqu7oXqBSylD3p407KCa4JHpjraw0oHr1npJr5xkRYQN
8HKDEaD5YvNadql1CBEdtmImxGmIuG4903pIA2lWJq/KV2dLn7dBMzSdCymlT4bFbG0XnPq6bC5s
oL5igvPNbFn95vfz+K9cEFbT7C5fqbRSKROR536rSKS2kZkqgwT7wPuc+IZ8op5omKO1XaR02Sbm
LYNPax7mGI6rOveJTwu3F8YIOtZAYBTsfk2rlcd2OFy1cki1Aiy4Ijlm/AhEL6V6XY7979fBk2hI
rqgDRBmaaRrb0jTJzwvyqdwaSPcBZPyGKCuBwBTujfol6b1n6XnZG1eKwb23yofULlp5+Z1iy/Yl
SmM0FtqCqLsi8wgHxSbkCZ7n645P0AU2GgiSpLaKysl+nRboERg94AqdaF/xp7w/sF/5Z+zzMsJB
fS6jg5NytC4ZIg27eTBT8Y6pJfCYtzqGGMEFUa0U3B7x+6PdFpNg6m91gBZA6LMnK5oatKFw/YiI
5dGKN9ouygfHaNc03XKCTGoGaC9GDakTWLybFwLxTSgmA4QOd+QK/Wh+Jlg/SGlMWqr0H1ESXQb4
V9ODQFAc/olVRt4ohso5Y8ftNsGFjTON6kSQXs0MFGBd9ffZafXsmj+o61/sFPOU9GoV1N4bxonX
WPVEg/TG93lO3PAFKjqsg3bu6TYbFCSXL9dKel+VN4ru2ETEEKLmSBNyAJMdihPExACZoIr2nuDC
3Xu8vssGmXDXG+QWIFVfaUM7aUXDv0s1O6WK5ad0aCr6m1I2bclwCyMj3jJKwJhv9xE8BpF3GO2T
9WYaNln9KFELbJey2UUlCFHOAmEGfvxAVf+5nzauUNyvOBj8JvBYIuk7qaf2daIaH2+A+Uo80KRV
AyFyqebHReNDBFdWq7S+gHGe0hN8PzqsaX0ThbHl0Of+TCN3EaqnoyfXht6OawdNeZXWvISOGn4x
3ZiW0Ujz2vjSg33mJ+OAh9RKk0fEgoY65d6tFnbaZ7BcaCs9b0mulfOnDOZK/e4N8j+UgkJoyMND
2iI4EB/eXDEe8rAwVpMDAZxa1wKRJbRCaSf1ud4UczXrgF2J6IlyEcNuKtWEJppfZIxn6+Zvdk/q
rP1UC63HLpBjvWg7118TfjUUg5RwupsFvOtsaPxtKyqsKqYOPuRZAvV5lC0i1RYOKHr1hbvEkDgl
FuaXBoNp9l9UIU3UVMr+oH0OsxImuEXZgE9s7aOu1Zl9LMejKUv1xjw+HJ9GCQ1zfp5XLTyyUfVJ
jvaJOvFGnjpNqzET7b+xUuu9/RT56J2XYbJh31wUh3EwTVqyXpUZEsozN5gNWN16Pq1qLREPs0aS
FSPh/FyxHL4bVjRe/MFIfEYCE0WEknuMBzJMNeh7ZdQHTVYzAMOMw0wqSCdWz0eQmq5RFTy57FZl
YOirrhaXYH49ADo6rQ1NFg2NDpu6zI24cAv8dE8RaIHnJHLlGcvkWRT7xu3IObqKC9p1jo4KMP9W
MZEEF25aqw1Tju4VWmMwxdLD2Ga4GWEKl6Xdc0zQTxkKANMLaRFup8QTn+jx9vbSFGHD+uIcyVKW
04RmP2nTSw07Gnuk9UVJm3BoAiIiNMnijGIHSAp/Res34VOeoOTqy/cs/xOqMjFzx0NWzL0RjXkR
DCAMVRdMUovMIaFe6bVCBfA26k91Yxskb4R1g0F/IpVM6RtQnfZGqPnfGPeTRW9rI8ITRKOHtsFm
28istk7RbaaWf0/JKAGs+as5OkjnHe3mHxa2n9ksDfRVhNBsoDmnxUXXRYowhlIJ+Fn5Mx/gDPkN
HPcVzvq23cZT82WSluLArQlSMVgxfgX+ns9e5rBCrzWp1/39szK3DuMf+Lohr8ic7kTXmh5iVbYP
aoRs5PHvIIhHt1O7VOdVBWlkZcx331az8WElXMDnsVrDd99H3/JAAeJwui37F+z3O4X7RE50UdHa
ri4qn6AhzIpvTAnFfTcxFnd/DfZClcD6g4W+hSu5bw7ZbhAbZSDNFSCRvSh7IPqsJyMc8TML75jU
b8ZW94lOkCnFprx0Y9aeViATbtp5RCj85oC67xlbH5J+iBCSMEVI6bT2siWzBNEjHV415u9q7VzV
DEIZYUylatLImIyDE6hv+lwPFPADmfDuNNveU2Hsfe3PWND2gkdS4ltEigCoxnEY7VCPOGzWqben
r/jEIR5rNReFjDuZAy1DEJUM/zhcrc2+KKRICwi7IoolrA7qFx8vgjoX0erxafsqxTziqr7Fm9LW
zSofJEqzPM3nZqhOppJKAe2jWyDGzhpS5WHObNRH0vcIYUR7VUX7HrV3XQkCGmP/tJqHuVO3Qfo/
DEQIL0FaKdPEsUkWirZyNQjJsYaADFWBoiIK21FRDXRE7NkUNZYqnpgvqq0IAFONG2tE1tPag5sR
52nfLrC/HYUJxw8Pq9z35JXLLVVNqLBIGSTMXdtZZFjcIn4A+Lbh85zjXs5u0KTWDADNUufB3iKx
s4Yc1mUhabyqLod8JmI3ZdgEktXPfBJ+qVyzCTww+4Hhz4OEEIdpXvys69UfAXkYocqSsEF4KXsp
xqIBZH2LU2BSIRZU193NV5xuaCifmDyuwWDC6c+xttbFaepGFnO3eC5S7RSv8a2sI2blHrfDNIrT
C0DadkSrmY57qM7KyvmhUxcIvd3yGXI/bIXn30XleNd2OsgYPEsGepowcg+SN8FTC+vWRAO3PyFF
j5vAemXR5GRupJvUuMKLakkkrUGiJU/dyPHNifCM6PUaHwGHh+VuytrUype4a7aTtPLPjDAUZUo1
TjG1Ysgif4jlMECEUzcS5QMioBr66IekH9x3eBh4ofaB4/5BnLgMnDD/gQJIzdaAKZsTFIyF/4fd
m+hDxi3YOQzXYktJJmnyyeUv/MwdilMrIK7FAl934zX9bW3rW5fyYddXloa+jRsb5Fpl/8gMi/AI
QUqXPLg0/41E6/hMciHd+tfg7R3up+SzxNCIonMoQ1yCGInZPBNUtJ8sPd/VwqIA4OPM1MPQvL5w
cMtzoLDT9IDlwbCW1RYdmDqzQAzhounMSDvFOCmS55Na3Oj8rPFQefn5EwOsd8TqEYAJ5gAed1ls
NKtfj6I5QEbFJ1qgPLtozlvyh7PFceoA7/O19ZTasPLkaHBz8Hpu65uV5/qMYScZAE4z3KwF7/WR
MIme8duMYUDrLYizDg7l68cO/pcYtpLMNlkvG/qXhd227kjRifwg4YBuh6/1SYHq6RxXtsFQyHnp
am1eeUQnX86pn/pgg5V6kbE3Q5AgXmI9/7BptG0PTLLUQ83u2H2ZxHpLctwWvPHPLm1+L+cl+MgQ
76nTsaQJBQcnj6l9AnWruHtpvL3+hBgtVnuxtDE7VxhZxO9+cIfPjNWrY7GcNtaB9dSV/rcPtW5f
F538to8UKubw7OB+0tsu0ygcYxCJkRkKAHVcd43N56R4up5Z32N0zco1ataMkFoqhZ3xDDdLkoWE
UGpfEcXoiQILZx7vXsSwbRyqaolz9TiEcR0mUtXvNMEW6/MEOOQ+ZgNewc/oZjbb0EnV3oLAAJjP
eYc6Zfo1Qxxj8RNUN+a5eyzizsQ1BMLCIacs8q/s6KKyKsD+msquk0KuKwqbiGyze6USfT0MtLUJ
XIejpEziSg5R/MNFrb4ttRPkOsNCbrcmsqvwKzxZ9w4KX+tP4K+oq7i7SAVWXCXAxnMhLhOCAP0p
fLCSvI37bkUXxnP+iGxPPCA7+KbWsty90yVRKI2yWwX1v7XpzzgPGjPk0Kwv0nkvDoDu/bYv1MaO
fHTPNzKOic8i/d1rOBMZJH6hjQ6QllSnUR7BsibvkU0KOZC9gsi9wsDj4l/tqJ+i6wagI5h/2DV8
hOfWVw/ZPduO6PkYH6T2Se8z7A+kBjq1j1TVKLTh6d5QmmWlxxSYwIDnqSh/+dHWHL7NyQ9MxYod
eTApA5/iniH5BCS7m+5B/j+JslHWAC4CWn8yLkBkKJgfDq8DpFsOwM26AzWYbRDdAbDvBFZZCs4N
+O70CTXe+hqxm52Ls1o5RkZmf17tYAiXgHrbsbw5X4x8lGbMcAMpLDgSzLYMv3roVuLOfiya1nww
eI2oHNu33HOviuUjttTThlJ2PWJ5BUTo5MJDnGVxBXWPT045AlFxCdyBAlKxJ/slDODsiaL8qiW0
hTrnxi/qLYh/g91iDKjUHlv5U2JYIyaq13c4JST+W0KccmjTugeKMhkQjRTU50Omi9urFzAjZod2
/YYUS8l29BMQpRyU5tRAdfNLYwHUsS6JvczbFuuSfwnWm6JlldY/9d380jBmWSFxe6yzzE02rCLv
Q/F9X7Nkiwfc6RcH5aa6lQCLWriBbdnernaAPPGxArPInCmMi9QXPdarVJrz3CB8xtOWa2/Uikym
zY/VnmiXDzpcUweSiuUyayeZ8fuki/u7uVJ+StoY9w3DR0NQUf3DSyIFsdwZbrfheekbMcDhJkKm
9CQwEJ6TphmnID/Mo4te6MMkVVr2LOHIh1cnHSL6SJIXTjbtKlcsBJoxWLu+gSKdLDclt1qe2urp
rYmP4ylhf2dOHVsWCZJZr+4MNYo3R4LUy1shlhrmcMdEmeiZwLKQ11Jm5HPqu8hdnSCDppM8P5EU
IeD7sbeLWKR/p2ojdIhQtXkbp4dmHBFvov+yxVjW7NfZ5NY2hvozExmqowNRBVc8kaPXNJRYDITX
N6EZ91sqHd7X8fS9mN19r6gizaI84CBMz5LYi4X8IQSogQG4VmHcUoj6tXsMAn+s+6f+51L7eTTF
ddreCQUQoPAt6ZrFiE4OOQ/M3iBhO1nsRnRab0dkhFsLSJOVjqV4cUfoxi0M4eM2wYJhsM5QfVot
b6+qujKjPdNeNZN4QloHR8jPNfzxN8oC5TZGh68Tcy1vD5sAwIOUF4Cb8HQfFLIQCv2r2pyZ6sWE
0hvaYfzgYoiNNBxoIqZn5oAzI0Hfg1kj5SzDQNa2bJl8wCnCXVUupJGSUZCBaTumAaArJ+d5XqXc
ANRpsz4DSqmWcCSiQCwzSLDxoNRYyKmV54TG5tl6tq2Gd9HT9JUTdk9qyLmmQDFFq2QWskGGMYMN
wO4DgoOOukb2l1ftzcofnrFNgIpwxBD3loreeP008cY3tJkqicFWytAuO0ISsCc95UVkxKdZzV3b
lHdEBEemzcjpCYubY3Lk9CoKZJEZhxX24E834iD4GAqT8FdyVd9qERjEEZVYpkwo/gaaco85SaS7
v213ENt0fasfLg9jmAEkSBDgi1MKqoohJ6bFUWVJAGv3E8fGh6qCb5Co2vaXTGNPwl0SxsSGz64h
BQWqvoWamgmzs6FAziMFl96PZ2ZcQ+SeE4GuaHcwtXZ46vjibO4dhHyp80pBQoFg2Ow8zs3zb97x
LIKggzTE8T3AJaXYshkvypelJoKV9psfJ+DKc63/EUHLq3AZJdlbVeT8WECjrY4e99zmH8KAxR8p
kG2dqp+E9LAN62A7V5GpCpyCg36Hf1yGuamSRNBvvIDkLqjXryt9cbE3gCjEzLMPXXTHeiren/Fk
WmKg2qYFPgaqUUtWUGGYud0kN/VeSWIbH7Kw3NQQg0cywqpkncpyCNDhbIFk2gZQQurkSMbtaciu
RLweLeT5ETsOKRkJkdboB5hmG1O68jMtG0WnBH2qMwZYo+29hlgIyX0XtKdC73BbCmKKOgt8wszj
eBgBxCQ/FE+rUPhVGANEJArQN9g2rdWnGTd7eOxc0DW5zUwtagxlYnR/7GEvJHNZJ2414b4fgLqj
V1kKJrk6VkTTR5r2zCXLVr4nsLYL4FswmkMdVsaKpAeWFqWy7jHB7isjAfaU/Jx1Ta5TkCWQtQzI
yDxx8y9dQJj30n3U/VIzJQjEnzazH976AFRHvmXt+5C53hJ8OrlLjNhJx84kxWXU4ud02FwQusIU
v3grsci+QiRAObgccpw8SAwJO6evOPcyoAN+YhoumLlO/fxUBxa9Wzc+nHWoFGIFiwj0kh7UieUe
XsNxDCvIwCNui/zpiGEsopiBQAwqTd8uL8xGfR6hPYA9fDOkdlt7RnAUWmRZYU+rQdRvo51u8NhL
IyNENI2sF/slSAENvM7WSJQGNF0IU+Mrr8n5TxciaB0lLf3sf8sdVVgba8youeb/J1Vlrfx5kjtL
0UEt0LHB3xw3JKNs+dGraGvxjO33+AZ2RRpOot/otDi4s0Eqzem52+AxN3UF2B5Bik3ISQ9uP8bf
YY6uLhPrRfOhTl5JXFIQtnk3OhqEQp4nDaMyfpb3OGj5J9T2uEcZRoTktkK2oEvONsg5nGn3R2kR
Mp1HLrSiF/nqTSzpo4NWhGpvGqFSPYeLe/cBSrIFVaDX92zr5sIFjzUk9/fZtG/7Dh4i6WzZTTZN
lB3sxfEBha8TYczTUtZ9fexw292Q3nv+J0nJe3oUAjxtF+/wG301ngint2nL8qVdHcnwPnFosj0B
mjGbTgIiBcc33yBhWMCB3fiYuSyctz7VPrbJMVRc2pe4jFtUo2baUTjTVL3K3gzQqgiXRfzy5s7g
UMq17G3hFSSyR75j79CZCDwmwCFK5LNckJr8UgJ3NmGyMuoNSgHXUzBJAGD5+8m4wyfglr3NQGsj
DA5hoslb6qqZ2pyiGZnSUc0/vdXos/xzbNdJcDa2rI0AHabunPjKlpplka1k1qbnj27cSKjMAZyp
jEMUaSUXPjoITbKbEJy+tHnIn7YDms8wnXMKoYE2tT5bycEqe+KBGVbumsI3C93iawurTympkFm7
/C0uRVmvBXh0yLRZHlWl8pXZa+3QEKDiFOzwxxE2nm8RSyg+FCUDNGIk9O63w36WlRLAy22GV8gn
4IVKxDc+AYdLUNAelOrRxgjU9eLHHtfRgMUrMNkujQzSPS9Pr0aW9hGF6tEenDceFe2BVPxslsG4
LQATBUKD0dVal4DI5AjI+oxA9PoW0iHC+VrngO/pnfo/RqE2DL6+ErBNrKllHoVVIhWJhZ4JMPYq
nx8YNu5IwACNVRRYLSAdiNSEeQvSmAS67MwjQycgXwI0yQ1wPJhrd1S3YpMafN3v3GnViKfyaCml
waX1UQ7oUNGxSsM1RBoBg5D4W45DaJIqR6JUnZ3+Mp6Uo8T2H1O8wIho3uoHk9Cp5QBbu7niYZn2
Amjsqotpvvqf8XkfM/7hcR+NEcnP3mQr0bXrkvy9sNeyyL6PqcVVYovM5N35JohklTyIbGFQce/T
g6Ljo57uYc9L6lfxKHS3bjzIjWJN0ideIbjtOj/l1CgpfUzAgsqrp8pkG9bGtv/5jdeJ0MY/DZAu
i+AV8wUBRJSnFJq3bwiHtVC0Foy9v4clh6O5+EFk/Z44LdK74UM+Nt1S8a7wng28BMoXyJmRI3bG
dO1Ju2maPJJgFCcM70CxhPwecgM02meLzjsR0bqKOUKBdo1HHhzv1Wg+swluJpvV8Hoda4e29Lb+
GUXYkSvNeAmmU90Ogv/GAxdirSDjPY951Yk5MYUI5XRytCd/ZVhD25YFUGmqyL9EPhLjkoR/dU82
0Yikjt3Ac/MJ9EMKWiOr6X8YCjnVzYzdz7BRN5k6Fj0mpvWVQSX0h7v1zaiiTY/EG1NnjOr9auaX
m6vkg7mwfJ0sRZiKbUegVf424MRr11pYw5IJDCWui9+brNFvoGbqaOn+0/h+nWAJi+V67zV30dMu
90ZurVcjmNKEOMlhq9GNEZJHhZcqBRxl9/3Kgau4/dovaGqr2Ub/kxXYuV5Eafidv73Ld8GAFfzd
Xvu9g9TVFVJNayuBAOWDMCB0WKxc8Qlavn7ULoqvbjoI8Ep5rURNEq0jn37oiEreITQcs/RunpuA
i2B4a+4tRjJOMnHfO1htkIbAu1tlQDHFqEMcMkOE/Kw=
`protect end_protected
