-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
X+YgT19WawHhZKqrqXuAP8FmJQCmo5BFPQ6lPhbNksPGMYa69D7xjpbk1tgNstds
vtnW7Bb+uUYquvaP1eP+17QLhNrXY/ueJYDd+JIzYYhm4ww25q3ZSvSPosBoKU0N
IyAiVhMkrDQ8JNy1ZZybyKtl/UjGY6f7ldAMwFd/3k8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 7584)
`protect data_block
NBwY+ZbUGhv6jYitKSh4Ps7rjnqbpnen/okxp4fLn6CkjkdxI091YnyNfjT9JGWQ
h0AGqkMV2E8nLiRCR+aHQLAL7iqvFlKQE2ySPOUbPmDj0m9plK7APXT7NaIsPzuG
eXm0ygck7UKnLJ2D+b7k5Cw2flTwNraLRxYIKWD8MNP/1fYKgEYVjHoecq1Oh3IE
/QKEipAEbfTD7hcTLk6lQeb0MKObVCuqZPvD9wckE8K5p/YnViJIOB9jOjb2yPoh
U8TrVuzJ61d17lJSnD6ZJPGAGZgb5R9GZwS4N7jZ8C4CEPRPvfkB7ZTiNtBB8wG6
SxVnOKZiU6t3wFPF+KCpcPIgyUmE8simg0pUFIwmBXzWAqiSG6jJsQMXwmzEZtvF
7PJ0iIMj30u1NZMTD0+sMaMsTmB15d//nkyPjqG0pDRNAuy9VGB7Zz1xj3+vaASO
in+MKwmjfYRQ/Bt8udWLGejnWuxpfjaNr30Rx3jzj4/2z7koA6qBrlmmTnOm3DTi
xqwKK3ydoK1lwc/ULQ7y6wdjoRZHGoi123SiSCvYVUMlUsc5T6OJ5jafseqNcyBf
JTEsokEY+VPrM5GRFJ5irEQXmXvelxfqlXdiNrujf1x8mrAnWZrmLImjA8l0l65x
W+aULdHip3K6L75kvPHsIapowXfn+MTFNG9VzCmNDjoMNyiLQTaHv0lT/NfLETQc
f+kavnuYdquxhDCbbZJP1DcbDjmk1Vey9zfn8YO6paPZtDqWYRL0Bwo36tNqo/Sh
nvhU52kk5kj9I2bo5At7AlQLrMHEyNYP8yThpUkFfLO0PSQE1XPYKYM6/0oPHCv4
6QFzmS/dAgfazzV41RaOmfgCCX5vUH78+BAZUwZCrQngSdV3iZFLBM+0zRSSznpw
GhhUhHCkEavK2QhvqK7DbUKzP3/afJr479jOxaeH4tNTIBYsbTpkSJL1VYx3Y58z
DFPeWu1LSHeuE9UXQCqoOorhIJYe0/laGeNWm1RY0gQ99GgqvMsWDSkCiJHB3+4I
H/Vo0b3eLdy1dR4sj8Acqn6keMDAQisVQ7lAcMVO8JeJKEmeusmm1Ro7UlMPA+F+
RHiAS7sjAUd2AZZd7KMTVNdyhCm8iaXefbGK2d9o8lTMSPA1vmiI9rcbHMIc3sQE
v/ONZYH9Tdohd+ZBk0bX71/gqCH/lus4zoEgwcqaCbaMirvvaR7UPr6/Wnss88xf
lVKxGhk/PcbVdI9J5HCV8OrcyYgfLfk3FxxoFu4ohsh7YuduPBSGQzUAvCFOWqwA
Qy/WlehOeOxxO+REa/drqeZLTFM0lPD20N4HW7dYVt+5XbrICWmJD285L6JUXut7
RTkbZZQdWRxqUcQO3JLXEsZDMt31EJys/10qe9cIImSSxNRhX07u9dJ6AnkgAoZh
9xMXghZoIF+bs5ls/zs+IR4Xgr2pJ9mxRqDfFID/fl+Te8E1fcIuHixLo9TlibY8
LioPrtsfd65lGX4qIbxLa09HTqBwl8don8cMOeIJi7hcw+SrbQ8UsTXNkECukfwS
Y2A0RymuJJBafB9LFNNCo6nvyfTJOH+5KcerH4drkc+TfzBfFJPTrSV99a60Tf6l
nLI0z3mo29l3seQZm9KgllxBu4J88DiBB9LrHpn2JOCEXJVtp3Vr1JWeLNSNIsxD
gdfKD26h+wmCasF7GBWbaineyvW+c6HUJwT1Do2zIxHVqEzkxaoWy8DbpEtXbWlU
DcRp1fgbtTvbbOZuL4vzi7GvnayU+MaBvyDSU2u2mENrjJW0I2by64Ls5PDV38qG
nIdru/wEK88k3Feg6TCQB0Kmszbl+13mu8T7h3EZcwmFxgAUIqKoeBk6l646Y+My
232Lo89S72jEKVhA1ALqYLx+Ibo1zrCFf9a3QkjmFcCzQmZHACSljWXKUilguJgi
bpUD9CgSdA144G7ajGxYdrssNuwOYF6oK8IWJLhTjXf7rUvIDuFsnyu11NuAPvsF
yI6dsUGAYuf5scb25EIaeM88Q+VX/5yms6LuS5xFSkk4w4V3bXn+Y6iArz2E5VSC
UTNB+rBkVmQC1w7VnHtWqgo9sy4l8BANfJa8wg7Q4NZBdBWGrHodQVM+hpUK60K2
rK2jsmdW3y35hznLf2n5nk/BJ6swYJgamIutDi0lkK3ObndOItaORLmGoPzDR+QB
9BXH0GO/O3Gj/og5MKK7wX/dAZHwFkTZB5gMHLUgrchiz3NNyuye4Ro4dsKVbtaS
80HE7CyJzw16mk9Gl8vIlrPPZRdWHBhRtZpBsK9XTJhiTdSMG4uD0p+X0sUyzDS2
KxdCzBVJN8BIx52LwJsT42jG5rBA5inkdgL1RdVj/PtL+82soHHlO9OI7SCTBqAf
bmcpM5jp6prIZwXgOgkmvVHoT6Z4rZeimty57Co2FJl7N0bH0tnlIb068fUa0Uy7
+VKLLpvGp7nHsVPATulEI2M0HcUEUI7JcQaHx16or8IWUEkW0PFo/xexYP6Jp/xj
DPnzGVNvPZgOzUZ7MAXo5zpBdW0VR05/C5wOVcGlwIOovuej+dkXoqy9a+IZwkXr
F5LB6PYHpIjpBK8YZjdmROLgIQkMv0fGpf7mXN3+pcibf0QPDBwL70TPkcCEXaGm
OlsdHL2Bk6LVe2ECkqPDLdhv+zYxvHRsBrWEYckz2GkdxDYf2dS+QdofwZKaQLNE
VgqIDhynMCsYUAptuIyfH9cZkedzl6tU+nxgCRKKZjD0UKW+9AF57E0GqdQ2Ws24
751rrlodHNR7/tAbWeqnVd/8w/djt/TUaSRO6EuwGF4G0zfamIbsXOQ5Ks7o7xMN
4EfNK2CJZxeH23Nz5jHv+FFkAGtaoT2a8tmCzC4fCDmAkD6udRWeDV2/ENmkR9f9
osT1QDRDppF6VOFYlMVHKYUXYdrgQcvfqmAEX1WhrX711ZKWNrjuGFyA+pmNnVEH
edpH/NTfjWyAzteZwQ8Roo1E+mBHO813l35GjwKLKQvNkd/m4q5s+MptDPx03YHt
yBjXU0zXDAlgGK1V7DV1C1cmred3NvU842+klhHygc2H0PfbhmH4P9LZ8ueF6qkY
cFS/oIW3d/jXQhMcZzhrW+yVYqmXcXavifB9aRK618+tQUeYYUbo5KeyBciN4Z8Y
9T0X9o8PeK17HdWZRATmCqi0EeUtSLu7wj1WtwSN4brc81UbzyBTXnasWYkKtMpS
k1CX3xi8pIWYtlVmdhXcxGliBUp5zh/p/GLXYm3aIcHU4aZ4Z3VS0xWYVHLeJsvr
W322ixo1+29YEFzP7PmQ/Gt0sHnftbeemeprcvdaiqhhc+VkMRFpXRZhF2vaHn4u
/NKHqj7RPhJlDR8tvUC+eSYLRM0yiAOZ98IeIlGsUG1w1ii7R/0oTsIYinyairnb
mddzxSw2cQHWLZ0q/fmAZooEFnE9Fs8DvTUeHJELEjJ6LD4WSemKhTOdKT2q8W8h
0sbcLkDsTK7SmL0ko4/j3idzlUun5MhfAqpWE+sxktJ8iVuD8jOx4QkQfSGP6/SB
rR0PJDwe1qauKyQnfbOHl9BwEOb0i0/ff/fPNEr2KK5K1yrxG5HCkPBid9Q+a+vU
uIFedsEZPpxRf7LwdpId5NRy8Gj7pLG8+ijiBOD8pEpE4AhePPyAE/Wp2kNU7LxM
vqL+AnqANzE0Bkwha8E9mzQhmMUhqwsHiCwWL+YeepBYuq2Tzppqdlq87mjIXqNY
IJb7cBTFjTPylmMbHpEd1M+YwCAqBo1vvjRTMS8YZzgiq/yYpcjNygrTCXhkEJj2
dJVUk2lI/UvwFWOcOZ/fH2sGq/XzMcTmyo6C3ZNJMOTlnOJMpfxCl7EaCf1bqihc
oF0uQRed/xcw4Z9cw2Rs1ffuhI7Yr48vTG/ZpGOx/kGhRXWYzgozB/QjYyPmQwor
uCfgtRJRsbD6SNeLKPsyVNFcf1qrtJMRVmrC26VXZtFh6s+/n+FqC76yqHAa19fk
RGLvk9/Q+IQ/D3pOiPtoOxnaDrpRK06EifwmWC/cMnOhPfSUF3PiX7uSI032jeNS
spEcM7udENpCOTgjNn9nNncIfrYSqnfzf1iMATn/1Amx9U9943Rd4oNsjxM6Eect
wE6VmOolPtY0dyTKtJ/PmMxJ61MjR/H4TlPRQQkedS05IKmgWIhHzeFnn1l9QUWH
41RgqAe7jLmx8GcJJmsiBlYl0jglz5xqdDyByk6FEIznO+Nk181Rsce+3fN7QeG9
6ST5C5QTWgXG1/v34Th5BCcWcTuPZZewJN5RN59FsS4CYmPpzwOQmLuqjH1hlvFc
ngrbXpJEr0ZtdIlEU6Jl9Y8c632bZjEaKeHkQ0+5l5VnRPngOQx401uB01ITGNc+
oT7DIEyOLpS3wc/7B4jhSF66ZzfwPDkbmG6qdbwI75lRDiPNkVZ2zYzbAI/+LHsO
dwZSVizU8i7DA6Mj9ZIj7lBBk0WNJA6WTJJvbsP/ZT7w86SB4v/KN9/Z4yQPpNsU
6PVaVpjJbKZF8oHB5xRiz+bMn5lpX6Oy/SB+Jx8T//kACmDfdVrw6siQme3mqDQY
gmgsALmez687DQjYtDpkNyJwExkM7SCWv72knSRrBh74ZH9TZMBHE3af20jUUI4m
7/24axlHSQ0fIcU5M59UoKpDiLrNYP1hAqT54cBEg8jyoPuY4xOGdCddS4vlRS3B
yqyX1kBKOCN3h1KnGCWMlaG3wDJ6G7yYbII3u7dYQsd9G1B55/YKNWQgnegrmq/d
aMVS4uK5o9q2NMsPFzKe4hBP74NGT6tpjEnI8n2xRknNf2BcOOhyyEv9cp60sWVb
wBdn9VXxSxFg/Sgf+Fdytw+Gq9fFNftbiiOcJCUqfS0Pqro/SkZNWZN8zGfsLbvB
JtWR5flE9qdYPvYGhogqrHzTPiQmyT4JPaueEBYuNzh4nZG/do3pO+HNgC0BKllK
Ps9QZcUiEiaHdpf7viI7NvFMs6zNdvhVwJilF00vT4LHf/ntHto6Y1lH+FpMx9dU
b9DLzIz4zaCKqk/qG711emUG5PqRMoC6F3Cs0iaFFN+i/EozjXnuOwKhuFCohFT4
qVi+0AMLqgQ025zm2C6RjwiEWWom9fwbKklz7ieBvMyWI8MTkhJomKPEG8rTNcPv
rcOylPSJv1UJUN//Wd18dDbsDdUSVZhJDz97VKXnHQJ2s+QOKL7DTCya07DMh/bD
ZEoo9x/D234Qi6C/ffVwxxjbcTWX3DQZ+LfQ+tBSV+91R5uExk52dmWN12hthxBB
82pViuP7BuXw+h9rpQr56wcBvAVGoQYm2OA1SRMQSkqUjv0S2tm170BrGPjjbNST
z1s6Gm44th2Hz7bJ5LAsHMaVFkNwd8Nb7r2PeTBu46ebTY8dH/zmK1D4F7XrA26c
LRjw/eh28JhCQdOh3aiLOXBGwhwyNraDVi74XoV/1oJmwYADyUFsC0qFX2TxERJ1
aeQ/eReWO+lWQqYGmHWnSZ0wbusgS9LSwTfbGj7QB1NNGwNsO/dX286xmGQpjyD8
pC4gO3Y11Jj/f1bkxX7u6RM5lbow86JkzeHd9GTUwJ//gwmlPEZhDNBeLKFXtFur
kDIr1gnWc+NQjxQGfhlGKO+Qpocx7NN9sCxC+dSTVayOGj2fsjtAy54aY6FGNctq
QvHSkJe0lq+O5gfDp6y59cizqpJ3+xAf44VD1nxkLzZRXyocRG3Wc932R95NrZzJ
3UpSeZ0xs16pAu2S7hfhQsq5Zqb8cziUVp4O2RPJhxZ4SR9yFmDgMY7SaVCUTbzb
aJSOcy2jsfsyW4QsfnCZtWtd8tddmPS9xn4f8m2qM72NX4A/k7du/xsdlyo5BrQY
AWXuCKGFYuzelHKHSGZ7B1h4Dc0CWtTwCVIp0PYod16j1+/K4Mp9oSu6ex2CrE2d
B7M0lUrMKt+MT0eJwZqh6L4KmvFlVjSp9zPlrMJp1sh42y8QdVJY3KYNAR/9u5Rn
BbmQI2m8vZ7WikT1znViMD+KyKdp8FJtTvGYPk07s6OADKeF/TVf7jM5q/LoJIfn
E0DTzIPYQRN6ud8JQCjse4DAAY9GAYRLgCthUeobZht42Fu2hKQsUfuY+rkbY+qA
nu4huCIK69AYDVYlTBjK6r9DNZh/C6GCov1/VomOfzk4AjPN7j9I8FrtluJKWq5E
JC6rsLVRwsAmxw96GRiMtvtHCKWmL7IVPzJgeD7VcAVVgeZYSwb2d+sZf2Y/u6xP
XBGYKoAMCY00zeYhov1MafxKP6qCEF9UgTEiBCchV7V7y+0MlOJHVek7c9syY8on
qr2ZQjLB57LWdrmxM9V5yQ8DvOIPRP9ZlPq3NlkIOaH1Z4IUZlUBVheS5h8hmXMu
z8EFNlCrFojm3STCCHHwb0vP1km3sL8tY+H4qeBMuFw10wICTtuwhfRLYr56cfdk
raBli8Nk1V6ierYGXIat1FlN/hFQXajSxYJ3z07bxX0QlSGIs/rzxXdsd/dFaiBp
EQjlG9CrqroR0MPAkD9Ny+evoDMD62rDHSab67FPdI4JXdQ8SebETVSfBlyUKvOE
QZXDdhEehpcuOBaX+EhhFSDmdIvRM9VIhT10c9cZmG2HkQCLZPnGEdEAu3LYRnjv
4zNxXUmjbWmYy/wUYxCS9IA6nu0UJTQ6RKqIZ2m+/nNJhZ+xSu7mibwyt+8vR526
l16s3TyntGKAYzT0BHq9C9/gXSiUX2LNj0WZKj+mPJPmqgZP0Y8fRBQc0c4NJ3cH
p3kx9qzvIeJNimWw7raj76L0XJoTjJrv3/n3pw17CZQFgA8Ad5Pnwt9MOFt9anuC
gfTA+Mzav6d2JTzXcRlBw8JpTtIdAAOMoKSqV/PbEL98itm23ppMdOHaEyIxIkrl
bu4Y2ueCZntZaDZiE6A59mmnVSJNdWKScbm3JzCAsck5AVXj67RTBkdtWmvbh7XC
ZlgHF9r0YgSkmpocMc7aiNkJmcSBuYIFRQAclcO1ndOXoT5KaGyPuhJOPgyh06av
nqmx248Wz6XhyiviLnTttn3ZH1LoIDaJP6fF4CJSpta7b4VVaYq5Vlu/T6T2XQSe
uJOCMm5LeMiIrR0DzY8kIttKWp1tnOabG7lH2pqk/XCVmUVUneB8ItfRDa2bAAHU
D63swkFTMEtD36NkZ2gtLsHGLt4vz5StkpNvPNmRJFUHL9cHoNu9p7sVxheLMq9I
nZJtPN7pgdVLj2HiSvmVOYKiYm5jH4oviCZt1MPaDdYcg66OUIupLw+Ifw7lKI1b
Y9vvFvPbK5Q/0VSkfV7PCc+Nuac8rX8cqREAga4dZGbQM0T3g9NU9OHwRmsxWLsv
h0wnMtfQyIczDqItdZmqLb/VaZi7rygs7SwajFLHECPYEe4yoKor5RF1TQH5h84N
t/o+Nm5uoUG75xvE3bxvGOHSS4U6Aa+ugXyykWkqiHSSz7u+Dkn9HPR+e6eRALad
9JuRSoQVYKtvIc0I0bxZ0qEn4rY9fuegQOVIGyCv4cpmxTL7/zNX1s4rPTAwki6H
S0CDeOZer/s9Yd1vOfcEvvJRSHYdZEBL36Aw3bUIa7hSoJmfDwZK7Z2PEBQut0Zs
lqbH/+im+QboBaxyj+nCixlCgDL8HhTb9PEr2xsEVJdtbvQ9DUNBecGdR+eEMc5k
AtX5gMKzrO7CKsGW/uneWquy4+kW5H1A60F/HobfZIfukkm//Ax/ZC69TMWGlVet
wqp9fUt00MDxoSgLXvkF6qpIKXyLfoIKThYx4CbCO36SXNTSiCS+2v2kFkJjiPR8
xuOnrWJx90jhQltV1vw9C4oAckZu1JYxJ2VF/tr0vpZms0CraG4q/Gbd/205rwTn
cJ4C8qjigPKwDHFjmQx6vEz+JgxPLhH4HGhGTBphOT+TNQcQ52YzzOTCj/wm0Knr
DfdQFBUPxuJrktlAKDfUvArucqzDe6nAs8c1baM/r7bligjPu+tsQSeQui8KNS+P
iN1J/DfslzFwEN4s1r1gvk/e9WJRFPbA5QyhgZJNZrjWYslSNvF6QBmEyB4VgqP6
DRqBz+NNLQwsv44ycpjFFHlVwDE3K6O7adHBqJsBe77qb+mdLtpNyv8nwsL3QrQJ
XrOCDjcceC+PX4ibcP0ghBxx2iZHEG6m3h8wJCZ8ZXrYp+ih2g4ZhuBSqqeHc22e
TCzb2dtXUxW3x/AJQ81emu4Ca2LC2XDtJbJDthvMTHbi5FFNeKVgBIf9+W551n46
S44ja2iVhPtJdtlit+ZdqZpkzL24EavTs9VlYOzSDPSwHqtoGI13lvlsEIyN62V8
xMHAa4afwPkAhahOo2Y2mkJgLuQVal4xZMQnoVONZSuT+2bgyQvQcDVEbmJfVEJ/
43W5U/XmGqJgyGHEyeokM/eUEXczM0HPgUG45tirfGsPCgAo/Dx3bO15mktDT3MF
5zo/hqmHvwBsHlQ4NK22yj/0nGP6DAi5VSb7q3dVr65iNoiwp441g1s1vqAOBKW5
/mTzIU4sp9yst6Kq3wv3vaYBjM+KYfE0agf5G661HSjgi1FtuP+C3J6i3aUUplv0
m1l/+1PvM/VpC2TkjweoK5CjejQRIHaMJ7sjRmqllLYgHKf4G60CQYwCSIJyuDpL
u/YHiXYE+IsLw/O5ownYMuVdMs34LdiQfIKoStiSTJ75ZUNBUnuxzUOXIAOSWFQU
442+ebIV11GGI7aKtHjbhK2UQuyLeuaXEelbILGKIXhtQQs4bwLbt4kRE60Ue9ou
AwNf11aK9JHb8ipn8+a4yOLQYgATMgwIY2Ws91bm7NmuAJCaS8oDPC68trg3V2Nz
tfmVZVxeA+BSwUi4CEEZlUg0nhH4EF4b41cz3BU/sa6MGgl2Tk9Gu6NgNmt/q1EQ
c1APVacTQ8YGOPbnaO/0O7luuDpudyZV4oARCELsE+CeuPP0YlYVD9p53SwF8rZB
lUaqCNREIGLAny8A9Y+DS2lE4nyYNktB1LNymJFgLa3tCSJKVAyoifmFRpLeVPPS
rYpI2XDUOu7RhACWN1iJRuKKF1g0pRaxJ65sIb4MnUUBe1qYf1+V01C8Tj6sDHTg
R1pXAREefXqKJwp4I09ARh3zPwEiE74mh3fDMoRk/MiSfbUb3V51l7KrM7A9NlTY
wCZIC9kNomsFIxWQ31m1VYsnNXkjR7DeGrtDquVRwIgxnoDe2+Yphv7/wUAGcYxu
/PYi+DG8ql6ms557BLavh8F5puN3ZxtxMOffiL8q1cSyPFsDecHwRFWUWgVVdBm/
iD7zgNZ2lW2dhbZAgCdVssPQYPO0N0U7uP+KhXwQfO4wm/O5B0Muhui1OxSd9ggz
0eyyfKtYW4MSG0/AvjzzsSkNSiBZcGEAS7uXtXdk/3VgSis/NhCRM2xfo/MS/mu5
cOi8Kly+79Idkm40UCoWOBPkdWbZu5MH3rleFiDCTrRIOi2MWPabJ6IexE2U2bfr
lJztNvHalasn6jmnsCQ7GkFLN1VpegnAUYyq+fmYtUMj9vJkg6sH/XqRzC7uW02N
KkZfar3Sah5al2tgYlGHPoLwxzwWIhuF9yf2CEAnEAADPlfpjHXYG5mPWetLVRLE
1OQbZoW2OS8Uw6BXaE3Gdb02HAkV70IIKZGPao3e9U+Xa2mM2VstEv6SfujsHECw
hXgaERcGMtFCxEMDhe348hlZrv5fw0/HACFJmBATzVsUtTh9v1S8c0vRaWKYi4dd
0KmNfmWwpR3YUqIPNi3zwvFZOt2thxPQ+JS+oRH367aSBb14Dl+qCnkEhESXv/qy
wkiFvB/E7SXlq0fr09B3ZBYxX2XP0lFPLIxl5M421jqxd3MwktqpsmRLzvzX0tKi
chd5O5tkJXNkyfFIm6LAzM69wd8wW7cWLsEohVOoHjC+MDDe/WYvHG2ZitWfPtfc
gCiA0u1w34FG/HEhlPQbHs39dUr8P5LquOKuXibq7gQkO0lAfCFkMxoa5oaYtYms
9NIdtO+kUD6Dx2qCWskNa2CDI1qBQtwpxbVw5Z9X81z604nfuuWF32Yydi2wDNS3
UOxd3gpnUKVkbCb1ekR87qfuSXnJjZxSG+vBLkWVUJlShbRTxN3tkEPER+Pbt84A
iV8x8f0DZ5WmlbYoz551Uwox0ZVkq1qyeQpK4LVBcAavs1FBbgZ8YzebFUcidrbd
`protect end_protected
