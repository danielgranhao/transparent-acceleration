-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
VS+C0U2D1yy1cNvxmh+QTOxbfwwFTK/bijNTzH7eHSCepbaIax0IMK35qnAx/yJA
Mm2LhiqEJZnyMWt2DkbsIcMLHsjWC1/7WzVL3GJS+HSmVgSwepCJMiq08RT297aJ
RcsLO6IUrlst9BQuQbR73mKAyrOHhc2QNsAXSWtFAOE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 12624)
`protect data_block
dPuHa7BH7H38vyY5y20SefJbnrqrLs47mDn2ZSSB5ZzU/H07p+lI26k/0AkzHGIl
W1cjMVEt8tQMQMECbB9Q8UYXIbSfYYugIHGIOm/wmeKoiEWtfPD7AAb5oxo3DXZE
ARhla4DB0VFWnJfwDKWlXXEw3rIbX94mDp9qMhYW1WeA0W9qyRNsqU5UYS8R6vCd
QDZ8McueGhRb/5CiQx4ClEd9EU6WY9OrJGbAD7qrXHCg46K7lSH1OX9vjDcpgz+P
lFRCwAmdVrpmF93bmy9cZZq2B3Lgrs/x+ivdWZvx15t2XOhL1NAcpoksmv375ciV
FlSH/7Ua0IbmMpFv3ze29w6YCUSDJl19c1Gik4Mc8zsumZM6QzBATaggOx2kpYec
baHRXWWj0FTkBkwkYfY8hr7Q9gDGRCLj3zQnsNJJMaxfKGmMJJTkm2+h7P42z8ja
XnXQuRNxigMxzVJK8grY6q6dsF4srPz3AOQLkFWsGaRQhvQoCyyNvvNyYuYw91qK
8O6wuHc3HALQdZIetuNIQMtBtY4Hx/BiA/5T51bsejDBT2PDzCLjcNqsmtk8CXUn
B2nSDaLikIn5XU3DgEo8Ga0XzfxvjGteKSlYSFPAdkbd8WRWGLyr7RHobJ0nl8ha
LaBN4nd7JBc08BHxr5PAxfN/B6yimcmLRqMPNYPR7S/7xVYKQTbrLutMKoz5SZ9i
n+/Bu08Qzo6GHIN5CaBIUWPckkvklfYyOuGUZQH54vFVKorgm28Vq9aeRn5SsEVj
x174IHH1qDlZ3l6SVHPniZsd1o9Rdp+jglzbe9uOxFkd2XZi2OhFsXE6Dtw3/O91
agCSeANybf4zGlpLcVRHlCMgkvi5KG2EnqkKkINbNgjwuEVrrBvh1N6FnlwLsh9+
mVRspINwQ0nYczZNMhOfad6dO5VMu1UAE3bPU7ge4J4dNU8BS/PKezTuBOjzTgrd
LsZ9VC2jA+dx01z84u8btPgGANTVr7FXai6Ch5itEO4fMzzKVKnR4lpG0nD0gdW6
se5GmJjxdBD25yF1QcTcZVx4blaIxMc2b5BXReY5u23OWE2ogF5AoK7wpCeeRdFB
wpQFIvGm2yTh/reTSemg9MeeW/aDJtNWi0POjS9FzyCMpraZ4j4YBLdJNr0pxrSw
/7guzkMc1v8BBaBM1WwMQuY9BbP+oteUqtMoNQJQZM39sHgqww/Zd89tSo3v0t6O
qN9oEvAY4HQFO59O2HIf8mf28GUhhI75nc1D34oFnjHy9KSGm3HuCDAQ4DNXHnk5
9xz3naogXazh1VjIORlgzKJRa/rVN+deuZcUmPP9SIiS3EmItzgSbpL9o3kUV4bO
8pKyQ/dvsN9b3oG8GQ+1GdZBzkk3YA+lSxghDfIh3KGya+Cs18lVM3SU5J49qi+g
C7QQALd8Ai+Bywa6heKfnwKAsj4RH9IyDogOybSDkAGHde/W5hShe09V/9LJbWdx
BXh9Vqwv0FDe7kNxeWssCUbJERN+hFoQuUeb4qoEyLokf+PO3anq6wz2EfWWpdGM
VtLzHlxNekpnAd1OazK9B6q/MKohXRFy0vG5mn830QBhl1pC5mPutg6D8LKH5tqd
LqOh+6INmmfCdM9nZA15gR/cVFEGgBwL2IpWT9lmzLxgL2CI0a9yzE8e4YP9PTIg
CTK7TSFXf8K/VXOPyzywRGX1aIdGDJdP+tqhaa/V2dAv3z9XAzbaMxcLfAMOQWYt
8eISNQL6U4dZfaTbAkbkg+84eyF329IVD/BbggNJ5mD+6Gvo7kcEl+LtCpSw9dYu
jHyDM1P/Yew2XEdhZW7f/xOX+pR0lnOBNO6Uoew6FcMr4FA0SD1P0Qnb+N/iz1li
m8UevpQUPnrjDPp4nHPWkEeIA10ttN6S8tNgdvogEatTAP0Xpun60zxLjwsjP5Wx
kn5OvOY814anuGeyEBV4FWKLkJQLDnw9NpeUaOuA1pEufzBUM+8OCBxIIhsc3QKs
o7PevaInosp7Avn+DX5h03/T3mT/KuwbE5B+7mAt5ehyalMn1tEkdTh02ptyEJcI
VCsGgE9kAViyt0hmByXyGXHW5OTim1zriT+xv5qvNekKUsZRqjzu3i6u6726WPiK
9kllxAvJ2EOG+JJs+xSf/x7ubNSfpgWulSaEn8nxiPRpC+fqurvV8rO0ATboQWt2
vCbGSyQ4hzlSJ2pi0BbGxnCpld3eI4mMq6iRjOXHLINTSors+/smxLzrvJkOw+yQ
xRNRgZEun/1DCD7eGVZkFnQBkKbtsCIF46448ueKelkd1f8pX703Ds+nOx7r+7NX
QUT77n6n9J4eXLBH6Koj5GINdqTVe5pXpUrSwLBi7iVEnDWcXB5Kj+K8c0vypVGE
VOdE4L3QlyIoffe5Wul3x3mmIRgHIeF6M/7TD2DjvkUrmSL0c4zPu+X1n1x2FMYe
rWlwa3Rib9eWhnOdoCNHsZVysm2Rsu68AxgclnAa2J7BLtK41+Uxf1fX08ZZoA8K
E3neyvQHCZOW9j4Tikj2Ut/OOpIOPtmQOYzqVbxoYfQGQMVooyN8dM6gLUKPJezy
ZmJb/nwLovB81kFckHWXzzwOUA3S9u7EoZsmLE8z5n0yqG1m6BOgGIZuGYoFNGUr
x/a0Rx3ebc+nUQMhtcsADhB2XV/y+HFImJZR+cGyXG65gh50s/2AsMto8k07X2hf
eM2JFsN5zvCj7ZcNtDHUL/yxfV2g/9cxV+b5FES/0+bTA8rCV34QkifClgLRo7b3
V5VEYV0DJdU9fUg3foGqTcMlLDPNe3/Zzlvh118YMVC6YSTZlJaWJmWiX2RWq7Yj
s7Uq7UQPT+oAPrlwIU/YI2ub5m3yok8/kl+6BfqI47SaXE60PEB3FE8W5I8+B0JI
rH9BNKGbkZ4xvLZViZ87G9KkoYlyoQSLl4pypn0acx7JWUVASwfssb85Qdiqcc+C
7MM166Cr+Lg9LIxFFF4NgvvfsbnQypnwOTRRc2lTjmcWAuEd9pjkSvEgFElbUU4G
wrw+0b6WAQ9luM1lLzfg23rKdEQlccvR8Q0R1jfeiGBbW/ltcdcqJh6lBEf1UXUt
u7f404amFfJyhkLPlD0TdFdQsRVBgwv4Kc9plSNcdLanUhrsi0S1CwKF/z4QJkGh
3PSCsGnmZdwJFs565FtRJXPVsMCERBSHlWu8GSxw2fERVwmgm/k5qiN0ACvJAbIW
cpL6zB6dArWLZuXLpSeGRAi+zjEz5Hdo6z5sySiUz3yIAbUyBFKbW+l/DdHgMwbH
TOGE6HWVz4hyXeyeNd2FSrbsNlqlMVb3IZ4gdh8Y8MbF6e/UiljyUa40IKqnH/fO
x+u5fPzQOgjgGwBoD0RE46j0/0PJLw9xwVF9AroBT06gYfRQypKdMo8BKPaYx4S9
lllKzN/mi4bBsrcGmY4Sjl6bX6AdieW+JGakYN5VIj62DV0nj2ZgwXn3j9IyvnF2
ULsCc9TfhjKaooa5gy1VsdQoD1kFqXcUM6LvCTEi9tMxJvpY7wpfRjTYzyhOvNRw
s1qROR0k+WsVuuS8uK9HZjBi33S5Y/SmCMSHO8gwLS4M87IoHCWF8TqBo9jSA6iW
hNsw5pi4x8/VdhloJEJKjtnBJAEx/zM4sqNYBDzGA08cppRfL7QfGO+6/EVGPxGR
PAH8LKwdqtillp47JI6cKeryLYCSTLXV8PLe+Otk0ia+UXh3BaUTk//T3b4EmeI0
+aR4rdNoP/u0AlIpAHi5gxBrGuyJw7nGhuRu4LNttT/5LgWo1rOv6HZUT5ghdv0F
Ul3YD7O01P0VBpkvwxU6I49AZINfcVnPD5Ph36mXwthDU+0tXFoG3scVlHEKhI8L
TNwfsUld2GPBy4ZPyQe9SNhvW7Thgvu7Gm2l/XwTEPQZRi5qg3b1PfH1Rf4L8m8G
y3ndrLawAly8jZIO3OaVPPpfDiq42Y2KaBz3OCIXBbqyoKAs1gXNVWxbURx7IY1Q
2KV/z+5CUy2JAF66NghC6eQj54bhqrvm4QXfjGzP5xVOkGHWAGQiyBSQeHDk3CFL
DBC3HC2S9I5XIwOzoGf9sNitXAjrqu65cBaoWNGIJm7UbqxjwgPEjMeCwETPAOW7
o0sVb/SBJKJ9VMgWjxCHv+pgi/kzZ22iO9n17FxWo4RaxnP0iMT7Q2cCIAJfnvA+
oEKfpdVlyMbA4oJP5fso0sg+QtWETt4RjoqUVGTV3xIodv6k8FSIQrLF8Q/jNHAR
9BLIOpzo3M0eOGue8yc+A/O/xC9r9a3m55YNszQC/7VQ8NkRX+Pw7PKj2TR4uvyl
GHANxsZEt9AG5EpGM8q+hX6oMdAGbcJO8BwZD4BITnTNj0kWCttnuAjqutwShIVv
QAiODYlcXXmBYSBdkJp9Xi6EAjp2QPL7ms55iVB+t83lsm/pq3w08urnB9s+DigH
rrTt+/rm4xDj2veOb4Rl0SDtTs+gt98DWujlLRS0Zs/9SqdbFAV6vLz/UAvHWv4P
iKenRBGuHq9iqpUgv46ksUN32vJEXrddxMDjHgtvP3bjFEH1dK26NmJy4a4J45v7
gmmLK1teJ6aCxOMKslaAqjTuKhVPdoW2LlIZHjmTLbVDPAHMyAya15c91A/OXyeA
7zcasfTTARzPvPYkTTCT9axv46dT5mIi1x0PJOG8KfQN+WQvVYz6vPWA2+TtB56g
JDF1jrtOpQnCc6HLsDnXmwqxxBsguXdwHBfnCylEQPTrf64QSF5P1c+iIOjhP7dp
yjIuO2HdY3Xf0nuHEVBbgvKaJ40qr2ElNN/+vmNrNhDmu0csWGhCk9DLW/4TFC+/
lQWoemET6Y/+HVWYJ/3QGbQlEa6mkLqUO5mwYfAYDSstoaPytDLuMy3NI8u1INDd
4+QS+uGE0Mt04CLF1aigxzoSy70LVw7v+V6LjPwDTDZceTHMlsJg505le8KFFK0J
HhB3BH6aoW3VHO4Vc9IHKGP2nk1n1I7NXKRLytWPggDrbeU7VZzfefKgJLma2/5S
gWhJz5rpeGhesXuOkCCQYRmJNoXIlWOla5NfoLK/K9OK8G5PSmXrJHrbR5QvhX2d
8knc42Fgf23AP95D4llR9uWlUsyd7rIjmxPHX1JnezswP91+XAFf0Oyr7/4fsjJt
m8PDfg3n71+g6ah8IM5xGhi5kTOknrql7KKDtVM3MHXAIuhm06XvQPzuzPS0xzjr
QnTH1Bal4f3/C2Vbt1VP07WodjHARGU8UEKsdczdGGUwCLuw7xSLvD9Z1gjJgxYi
uoeov//KOJwHK8LNYPDrDMUnc1C4WTKLdxVikTVuyCEO9F2kCaZcb1NVG4B1/jPn
GXvDGU5jDzU8XV0gr9XU6swNBSurIDo+GSlSkxZMo3RqUDJcW3v1PXKZ0c4FZ6ap
miftM+WLVCi5WxieApN2NpZBbdP5O/BEQpUSMYw7FwBAF+OvBzjOHg/SBzdcBG5c
7vcUD5H67PF/qe5McfjI0L93NqTqn+YP51JTxJvTCFxMBoLRlTJc9TEOG+lMs77P
LTYloii1f/JKCGDts/zXwHPmgCC+gIUAh0QW1eyabWTDWdtOepWYFue29zF3oe5C
sx5rYNTouzwPItEL//xO4ZYV8PygBFBZnrY/W2P6EML8np8DC7EzvIwChudSiAIV
mbkawYIuMwefVHQAr8NlHeujRbeHQTETzv7IZLPAPAGIZcT0cO9ZWcwf/5Lcdvwu
hC2hdPy5qbdNNKBJ1KA+6nB2OVYe2oMI8CDkQ2BKQOcpglOSfD6fd3uxazRRdGFf
R+ATNhhdjZ94kjoOYIhgHq9SFdMZB2yhGZYrO/4uvJrrcrBl3QpX/W/RPWz6ZMW7
oJ0PBNJnZoLh3wpxa1cu+UszTA1JDRuHnuE5sJHBNEMu2tVZ5gjm7OOkTXkaAf3b
gZmiuy/cczVhS5kmJHzArD4rSQrBZ8bAerm3D8lgwm6xd+l+8ubH9ChGLti+M+qL
L1zYuQ4WBKWKMAnPMuS6coJ9Arm1cXvQ9n8i2Y2eXJATCCh+SrvfDsdSw1a5yBG1
+xP5YfBHCT021S66kCoaluq8xg01dRDNavgjj3R/+toiOGrueFPDawa9hrr4woJZ
yZvmGUfzsU4ZbI2zrZwEXnwgQxIhyL3GPewnkQlkDFNLsByJDHUz1yBkybBiJndd
2rkYGgH6CIbRZ5DEvm4wgLdy5jqYZEpI+wIYUYm5uZJjxR2tjr3PUUc5Qd7iA84J
vdjTvvLcEGDEA159gcMnVoNkfljGJnCOvcaguv2qBnpkBVbmfnauLvbVZs+7poaL
k4mMdVO+6MfzJ1UDeTudISJOWjebZ9FoOltiPhBXRDLor9j7XSyweQFXjK12xX1K
iZFH9LDfsfnr41lHFS/o6yJ+hbbgJtrTLRTnOgAIU2G2IP+gw71V87XiSihPZfly
s522XiTVYxPDhiDEviQZCKfBHuh8exe4Jy/aHetbNCZNhStTKPOSJTPEPK5FE8AQ
vr6QiE4DW5bK00AgjJYoqmQ3NI6N9m0qDA8gSDvSZhVKRQCE4zkb2kd7uDixE4MY
MMQhBUeCkesvqHBBoOqmOWkLBrgMpf8QMZxk/r+dIU2M0WTpxT7YoA5cR0ruCxC7
kQolDaZES+3ownw+274s6SzaRpDOHzALwEzMj2MQ9TcTiqtHw6EYsRn5f3vZjUJG
QjIXDRHhZ8bqeo69dxmRKpYUEDy5j6fEgggJcrfxqywG0tvX5H19uvd3Xu/XitW0
8mAMPprC3xTvZmlbwdvZy7JpUYnvOSCdtppjfca/LwQVIoWAr536uHUMp9K6CJYU
tOPjNCRfGNS9DHwrJhdqj1tAJYmS9qXwjPxP+T4FIGu7DJBIqygoYCXyC+zMB/tQ
MG0hs/tsnJR2FjPT5SoWjatOEtfap2U7TzxKNwJGhJxCwRxYmmeWPs9HPk9Z0VEW
y7dOcYck1bS/k1b0JlEVBMaSNDNBLXgbt/Fx7mnVrm262DLWS/5Bm+JwtX6treXC
S+n9+QN2E6ka5wmVmEGCMcYxovaq3r/tcLfOFXAikMx9xpz7h3TCViHMQhJUUvMF
6MYs+rUOqRATT1GRcwwwifhvDl6oJaOlVzpUlauRGfV2GG2MBpoCtJMl5nyO75ZH
aWFtciDl3oO9f6dCyHhqHoqKYcmwKiFVGMNV32oyPmQfsBZnagSxnKzZ9yZAmAnd
4+QUH/QCbYwVDlJD7dDre10wdYN8dobVYiF9UHBjSB4hpAc/djpz3OKRffGcLadS
eekyzi6uCnH6jiHD5DXxCGCKe1q/Z2v0hk0RLcSA0RByrTcd4mBBoOsTyzsUYmM0
zYpIaT3RP8pJ9qvRaAuV8sMCr/hVDmU01h9sZxIuxIbPdr6WfW/cI68DjwSnLCQ3
F/sgmMq20CpPHtI/0Y2HLPVDEuwsbate5FbGvvll4o+gjkZQSwCEixS6sTU7vHAa
FOfTFsrDYGP+Nvxxay64gQm1JmtK/1BIWCRCVq5XwTiEujrEt6Ur3ZARjD/xZOID
zU9cu+XXPduRc09Rmtev+ot2bLWzgXeM8D90svWdFTK4jhmo+mXyS003m2yXYSxM
vBQ3kAZnTxDj71Zc/fvMwsLwEH8ezIV8oYvmiij8ZpE+TgWY+4rpNW4/kQfGBqSw
lekrbsMXf+YA1jqtPz5YAFmohp1fE0ZDqMDwKQgHkh0Jycy9tWfw5MwCbxRNxB67
D+aj+o1sQ45PlwZoFMomO6iQS71+nhgWEYhLMXxl5ztGEjFjD648H2yu/Svz7ZeK
07AxlvpsjaGUWYNVGl3SITcH9uU23QZhR5HH1MZ5IEzM5ubaf2bs7V4PHNoB8JJS
yB+osTmqpMlXeeXjGG/0wGYmD/J8tQYa13IeC5hVGM6YIbmOJG1z5k3LzJUxVgNc
bW/U25cz3kJe/LpaYrJyibNYpEUtYV+78HtydjmFmDwYsioQ1S681xDRjucjuhi/
lHSO5V6W6XmLOVOFHqMw9asdWXqWKwwLGlaZ4LRhIatwJ2WnbAjqaMpMD2nf3wMy
7hJhzpQiTqBiv8yWWzJFYnhS4EIn7bDjRSOhlU9+0WwoOjCR/61Y/oe5mZqLRjDC
4VYBoiFc/HNY6vxl3ZMr8vFPg2TEP5+xoBaT80e4XKUa9gUZEfXpTYZF61qTTieZ
K02DhyCXaDftsMC9M494oySuh6iAYZiK5YmJxJ7uW09OgIDzouq1pDLhMuSfFshy
+2DO6tHijiggbeo2Bn9cQT5osG37kM5BDEy5+b4cYURbsF05aXvV/1NNBwGccED0
E88N/3XwlPjsTTSaSXCRy/KGyWC1CfscLOTFgg8Asi4FeHyUJSRwxsWNHg9bevzE
PnvaL4VNshPjREyEXcSJ+RP9zyD5x1VfOXpKn3dSDqSwmOv+IWUgj45Wq3zPOQXr
h7HabUbFdkulUF/LFbKBgPbeELq7CSSdOgwJA6TbDw9913Gwm5QkQdQCeF1l+KLM
qOnXihDA4RdW9XdD3Q0YCUxoqUJQDnLnO9R933LBFzR2EuLaY3h/sNDme1YgLCxH
LPaR+1SfZPYt4ZymNufMt5d3H1mdu5O1WhIlrAGgVYHZpcG2w3kfST/jyylLaLGT
b1MKVNOWLLH9PPCJDuxqneizerRiBQAUM1ktl/B68u37wY9fJi7PBVdHQgrQm6YO
EH0E5+ux+X6cG06AkLb8DpFkUtAoL+NwmBHwmOuTQR/sMw2ru0EvqinciqAmoOzN
2sPOSwn/QkXZGtVPbYKHUCSzFSqfD+OIIHhoghMweuBwptYRvFN16mTYi1/vmAy3
GZizQoWvKjt4vvUKjAY+pByPCw1nD4FSWT3xWWQHkjhgi73oK/Oh6MC0HClH85uY
XHF8oOln0lCAN3FoU8EgMPX9xYVxHvKuW485Jj6pYQ9NazE4DHCyImNnfWt9Fzuf
SVUkl0gr6Jml6AHeaByF88P9PUWg7BgTZ97mqGz8jDucGILhPoPh/Rs2eLYN2JoG
MoU6TgqmLZHQaFcqb+BBcUi0ofQavZqpC9TwklmC6thOZ/wDu1Rl0UVEv/jyqTGW
OO40q7trZHDEc18OEFO+gAoQUz4KVyIkg3atvhzWrqRgKOs9tA8H8SSW/rdXTcMX
W9Ue91vDcTC/MS+gfuQ4J8WDEVs2+cfkOcS5K5EQP/pJq4mXFnN8z3JCQEH4ad7T
ncM/slmFKzdwChMVJkkilWXrE3PLuyWEBjErhvCmZ3yGjTY2m5L5TiJp1CJuSvEH
lrUJAUzKZ1goS0WoPAKVZttngsT8zakOW9RZfv8tiawbPPMGkOfz+6XXvxmrYeyW
i4P57nJAQ5HPXhnUOi4zPG+sXGir+MAvtwt2HWXYk3E97/nNHTthH9OM9RtIK4xx
OCBHyK8Dz85za+1hvvN3ZMlNrAAKVJe6QFIJvSzWOQ+qUWebdcVERPshyIkuUqv5
ojCPYLrHl1aA4tpZ/tW8mru9wWDHYzsmkE1vHCqd3rLJKBvt2ElTkTbAKrVtek65
FXJATOP9SMsQRv8CdXGhC5AjNrzREpAA2cX1iXjZzaGDa0KeFv1l8rYhqwEwRyO+
Ef18E6QJ1YwzV311UrUTZBtsBN6oLAAUhnDLvZCRmaSYeCvlbSZGkLu36NHMlSFc
2bPv0t2ZN5TqWDiFLLvSufoz8XZThxqrbWqhPrQXnlBGTckuC8Fnk/1pOJhrlVTg
JHTz1IOF8QRemQNaDtcvViW1HEdduNRIO1p6i2TsieiCCPxU4hey+XHk2AI0SLM/
mc5JKtueJh6kW3GvcaQfj8LT77SmXjzK5aRstikJ7AY6B0krZam7xlN5KVVafNMw
+2tGhjyoiLBq6dejpY/NHuUEfBrkfTUaHNahivMUzYREqNa8/4nSaXN5DdAi99Kd
LFZdEY01OD7G+qinebz1Mr2IkX8m0ZdLVP8VCWCmjzQXhG61nGKUAEtSJBYu7hUW
Na7Y5K2V8NNcUkfCD5eIw62gQiTTQRxpxvLfQUyxbXEA0RPNdm1ft60S3QgBEUy8
DsIJ0ir5y09ja2xoxoLKNOHfejI/8SynmnBWNGWjW9IfH+DabwWfyj1fi7nNYY0v
kEcgQxpb69kR+HuM7vPh3vjZFEnB/WROfNWlpZ35HYmY/Z00qi+R6CP8en2jQKS3
gtZys9PFVbNUQTxVktx/Xfne3gkrK5LXTbVryXasDV1uD0lfpGl1DXX7KPrgPAJb
lROQV6cWruwydH123meO/xC/1zs1CCbe15qM/Cp82XLoPeO99JCPWumX0OHjq7wZ
s63FYfuoQ8r2dW4ho2jvR6DXRdq11K+1skybc2fWd4/lu4fiQ/hdUHgASMKD/+bT
+U6Sv/5DAx3lJ5XmgRaFIn+enJ8wwi7+4ceoBpznlaNyBHOxdlp8zbiQTfbEgI9u
D+ssfI+HQxQB8VCP1PxAcwnfuPmTSpTxUS0pfCzV+xMCSXgjMWHzT6xF7gUAtr3k
g3eru659lcRCRAMmMJBZ821dtwR8+UaSFWR0+V/TeolneROE3+GgOxJ8Vc3YktEC
I2sRRiD0DZmLB+9GSf/AJ37uDDOIFi+llfz4c1l2KzTAac36tXV3sdERpU3BWQaP
pAZF9M+q6AwxNhy86vgQ5vIgBuA8lQFK6EYivTjYKOC+KyhzNHrhLPe8G4Qm/G+4
9e+Z86BnSwv/Zla01TeKP9ZZQGqsIQX92DPxltpvpCkePuJnxwIvHyuNQWYhk4/1
n+GxGFj+3TwqLU6AgcF//hIbwlMxGl5ctiBXOpGYqqQUmTKykXRdZxyVu+7Sefnu
grRYMmm1+BV4j6DSDi4z58+jfbCglKNhHGqUpYLhrGK8lze3ZqXgzEwt/436gNhL
wWmIXWb7LSd7+I3+NBUGmr90SlM+53FkzYDkRzqbnZKoqzCcLNb45wnXxggUiAo5
uF1ba/o6Kn1aNLLy3JKjDbswfocmP76N9yPTb8b4FWjNyP3lNV+LE3GJxwzS01yi
U6J5v7UcoFgEXhHGIRaepcfChhLbVLs4nV8hqgXmlXSnVSI+VFiFk/5on01viRKn
4COTCUkkJJeZ+a0VA0eGsRpRiDCmnhHZLU3i8SkQ528hEBeylFMAOysz/GtGgTZh
U5H9Emj9Es9x45/Wt/vAJzNnur9SZboBsL+96oYsftteV4+G3AfHfuy6O03L1wCf
/68kF6A6MH7llRBKWhnIou50MKIeMLj62yrh63vcTEELlKthIpmjuLyqPNXxrnTV
L9eomCwQx598BiT6ESigCiq/U4JKGOTdd8nwXH+MiEWLC+M50sla+3hpBhdNOnTU
xpWb6mNuIZu0orhVl1TsgPFI1AL+VdFjj9HZQwFlUZDHX58GyzQR0ingI0QVOhad
DSi2HZvnLzgC6YI1XqqyU9tOfCM4hhljfIUldzYSko6OCV6gWmAPXw9M6XaV6BHy
Ai825vrrKGkyII01y0TaO9qZq7G71iAtCSmPb6V5/0ow8xnbCJ+ntnaA4L5Xx7Lm
/lxws2R9c2JZ8/2j1MbWNCL0tlQlHf3WSytbPQhg7Fu3LGczgdcPo9Le8+dAKDcu
1ak/NfSqXvHj2am7EVqTg4wpMFSZEIMNbQraQe2q4mzEBiTUgdZynJtXcwoDADQw
CJ8n/f8DHRvdaUVxDkfT3LsciZgHtHSCBXHTfVweXHSgTrBZ/SAhVjPRXq9XTDjL
Cs6Qx9iTwLbo4vz8svtNU6DXOCAOg9pUwEqTkq5f2jG+nUfUsCVPbV+ImHQoKBLS
cltNyZHVTdDUNSaOdtvCqwXxeQYvDFjm5i1+mZfkR4jeXHKjW02ngdYtUquwYcbc
gWXfngbAGOdyS5ZopH8D2flNy67IxIkOVIefKunfb8MjVJAqnfiw4+TF2uWnBXTr
sf49LDvqofmY8bascLCg7S8b6Dn2rwGPxRqHFdWHA2Oves1Lqu3HGWJ+qQJRiEkU
MNNMtvhwzISLcIDDhDul0zc8TZxqGGSKObkb7o+0HvqKAaEMBrtApGEjOI31fK6X
MPINrBNtFpeXdgAiN0xGidU+7WgKxmWT82z8SGasKvcDW2McIzNChkyeggRlcyNP
4vPny4Hiu1w/gaPFB+scOdHHjYfItFGIT2y+zBZg2yqpDTF5tBi4ll0rnNBNDvCz
LskQny6h8LTEYbLL2ZoM5bhPH7raJj89COSIRWSDe/FDHXDp8IRAVB4inEp7q6RD
Kj2ujEdUI68a5HDP+58q1aGWvKesbUcbUERAkKfJytyLKcJzokwdYUCj2CG6+0tp
+flY20XxBjlHW6lNRY4vJpHfZjJcw8cfT/IgDckKKWH6RNaxnZ6sanOO5o0+Cogm
AS4szkOBUKewQCkWhYI8f0e+guOjCCZIa0GzWiubPXuZWMpoLipZIj/Mwm/zir/v
udLsGKT53/qTR+IKzOlmV19BlQeN1H1Xzaa/FOnQ4r3WzCp+AtgAqwFkMXSo0tK5
8OWzVs1NAVWBe/WqS64WkdQHPzw4upRhBqY6pDSfFnGpiJFGBEEHpB7nBmRnbcBZ
DOYYlUvVE8RyfRYsUXXtKNokihqpZ7/1YQwuzjC+gABkiYguX6uXxHUw2ScutoO+
FhfseUbu3Tfbq5EzcrRdNRvq4OJWwwu/G0cggJ64bL2BQtoRZSAGNAOiePgXFFcX
Sn7nqQw3HJAZtsX6nBODxOouv2dCpNAK4ovro9lVEUVdY3tMz4hato4u/p/Bb2dw
j/TicQ8Vg1bTFfHjjuDfF2ouLZY3JPn/eTZw+uebNixBSRUBm2u273Vs7CMAPx1O
JiSeueOG7Rh+P1dC0t2eSFpG19knqjh4SkFeGMqbIKwXyAt49oH3W9gv3TAaY/XX
qJS/TP2BgnmUvwU9oKmUlBVbo1dGmdwIEiUh5or02pf2XX6w3OnGAU1yAbUqE1AA
PKQ8/ZSiHF8y6UQkvNhm8UZ0UGMojqQrNJ/fU/WWSjL3+c9BH/wyJZrV267LKekW
hDny5biDBSSdSUipO6NaWRyI789br89GsciNShQReVvYNNjIRgMReDxJ+Dw0zVBl
jnSvKvciioJmgGNbNE34DPzS8FUU2TFYwQE63Fc4ANFDrCkRZggTz/NvOiZoLVrS
x7Az51lQlpxPbUSuYJt69BkVICg+bLYkQePZG5OtJ+ezdq4Iy/vX7vYYmKokLR+/
45X9c41sa673Aqprn18kJvq0yv/jFp2vvYas6YVIJ2zeemM+X8pNx9qerrZ4NUaq
nuKPCW3NGuHljIwfqOHwFOIdYvQo0foIuTPc/TSQAS/uRdOQe1Y93ZxMlvu7v0lV
2ctboj3zQeMtMGuQPHk4/MuUZOpDGUxc+jlNf3SpUmhDcLdOJn8jkbkc96jyLh6s
/uHwjxSd3qjx++jsLBDkkve/PHo5SQNeGGX0LstqMWyC/naOo4XmPULNJIl2fPy6
eKgfwDhoeJGOPFMFrbV0VjcpYtmZHyE5rRmeKMGRrr0Y0m4P332bFhEe9ozdSIZc
zp/skM3XEzNV2hWKag0dbUNlNcviAJED0QjpxcGzcXly23NqVWmXsMFCHSiWc2Rv
ISm2n+QgDqqfRc/kBpeWVZATJTcuSIqU5UNmaWPEfdwPisZ85hTghq8M+XsQhnSy
xXmzTwTEABiyoq2Q5Fc1NTnrWBzJZa7oBN2BR/XPLBlfudzPzx1DdPFGkfB66xa5
io+SKwhbITk69aRqZlbLNuZ8yvec4XRP0Z06jk//sz69cuY5q/yKEzO6+cp7pLAJ
vn/4vr/LLoreropbnkZi8CJ1Jtoi925YOskkVFgTZV0CoJwFsAjfkwmIwvBjKPzP
OkNn2y06oOMcDVAtkzrxis8ONuIWMAnWVKofeDXQSSSRk3ENCcA3ddYVSeW/SIB0
nW/NJ2jYa7cOf/qJSqclJ/Olduy69Qhrzc2rXZjOlYeV0C7s4B1uMyRwWejaAMKx
2tajGVRXNc7WDijSTZLHb/YQzm4K7p3SzrMP97qnIjMKA6PHyr+/i0aBz82RVT/4
+xa5lmOq7ci2EpN5Iov2DRzDCHwq63Bwhb70s92SfIrNFMx5VdTl7QAnV4IQuZ1X
YfJdHyVdYD+NO7hS0BAkUy3EPf5Fw0F8eVA7VeOJ6s0m/dqYfG8qfROwJhQLaCl3
tQJQKHVfaIyYWeJa5so7p4ALaY/JPhL+9N59Txjh2nhpzLfJNdlLzu5P+JjPQKIE
UsvBjcodpUI2/bLY3DBWaNqv+8+NIM7uictk1vDE1rNJr6FpLwW9k9lsJW9iMCjJ
fsdGcQLWVo/3T++q+hWf7dmz1I6D/VR2P0UXfrvdeeKLrFYS/O9t5A189jkJcCMt
4DVpjMI79F1GkiWUV6gQPIJAJA1VUNKBWyaD5+K/Zp4vuAMm5OKA3osOwL1r/wt6
ClzNi/dwJ6yDAq6pFH67gAW8GFnx+HRgp076ftPXesOWpbxIWJntpLnzIaQzFa17
JPSAWy71uqWX0Cgznbwqc61B44ZanMp9cbi+C+p+rNVLnlGxeQ0clG3HUNDjA7uz
2Fa/142cVo8rCp9PdNpbWRQyTStv3w4k3jq/LW1ytvGKv832zw+ec4OoTqp0PhWn
yZuijfP2fGqIrrV9COCkCQvGtPawjwbi3LMDGp3N42AbUgrYJv/WjQphwxuvY/e1
nc4kEo3lJrphcya6IT4gQb84y412FbqIrfafPsvLjL9BZAoZpvujQLyASThaPqZa
PUqnGZ5okL80Vt4yaDn1MwB26cn5qFfX3+HdfOWml0Z86LDA2no+ZG23XNpV7dEr
fDpDsT7mXml5iLBkJ+u/wrg8Im6ns7pa5LwoZjZUPIIVrKzJarNEe0YiEBmFD2aU
/phQ0nN0jNDeEczGfp5qUp/tOejLkiUa99ZP1s50VVdoUy9o3oPMy+LwQYYOqvvZ
n5VqeVyQS6R78fmEP7G0wasqx+ynouBjVxdr/iWSiMDzOkQPB/qkt9n7zzv/D6w5
UjZ9U8ScAQJSD2OXJZRWN5y3CRnKsBeHrEphtTN42ZQ75KOjBjtIzpJBBzDxFA4F
4fEFzItFTRi7qfB9xmnYCpvNkbgYW2WHVO4bIzZ+t/2cDjNWeFdT5Y4Co7c+qDQr
33DuvN+IaUQ6FW39WmEPSyQUmqM5xqh8Z8zXOXRrJ+LY72LliIf37Ati9D3UJMgc
aPecnozvqhbKnJO0xZa/Re0JYmd1KLeszFPjDcdfSXSmQzyqLSOB+7EJzpjUpmkt
uTbrjC++Md4JYzGwNDKlHTm/onRbzHuezFyCO76TTwqmnb0k2NDE4HjMFUp9XC3W
f85wXclEAPdL+TzUrE6d96v6quO0OZNskVuZnfWHEpcxrH0+Z022OPUubk18atmy
Oigv09+moBw9sxd3Hd5AvF7k1l5bjOUPxMaLyaBIu9Q3XEsIkA0nIYbRW/dUQhm2
YE9u+7Wn6FCMbFpy5Dg/vJuz0z3jBasGy1FdVbGsulf3IKcjzCqBEvJB745wkRdE
IqgUVUsAC1KyFwlxn9BWME28DT9r+dyj2py+m4iqXR63p8T36oLPBx+f6v/G1GxI
oCSBrDNueVRMXpfacCzQyTzMQjLBcmVyr0k2gkZGnCFlu6YawUY0UGZWoNBdnDay
oQaNEKzvMgdPNHbo7tnDUBF4TdkfGFgG8k8s6LD+Abzq4gM53MwLpAgd2asbpx15
yN+vnEgXltlM6Mtlh3ahqzlNGs1KcpXJDyk73fU6GOAHUrvDSezq1KlxdApczp2+
MJLZz4jWNbXLtaFRQrwfCAvSzIoEllKo9nTII0Yt0vjsGMDShs6U+VC/9kl4UVDf
wqgZpweUTijUjNQMTotNWJ+r/BV0OKzXMpdKA5QP0/kD/90ZcQC0cRDVkzeed7C0
1QCqNslQXhqT1pz0qNrE0y1HpHbrrhuDlF7HZTIcneqJbMFph/+IHs3xhJRXUwZb
HPZzytKbH9CkXjBtmHBid5BQoe1twhsY4pncIp/vM16dfpcfsSszzPAfNtN2gn7t
K+YP6e1BpuNGqwn9+68l/iBDY9YMup5/LjqMfA/JRcx6hRLUXLVI/HYfpR+ECt3u
EzdxDQWQlBy6TOamxs6VFYTspK1kN24+QK7as7TUVkYIbt13eN04J7hOZH4w2pTw
u6l2WQZYAPuaxBOzm4uyc4BDdi9uH3/jz+HQz0E0j+JUkZFKrGPF0hyLc7iK+0uE
2b/lb4Ta/2r5nZq8rhe8FPrwN8/5hzR6ovhifCjCMXw11KqfOuT+2ijT/D0lQ7dY
PdkxBMY1ERTlPdyChDBqncxNjDSppWE1K9DXXZLEJPDVA3dYQjic82tl9eOkKm62
jllc0pesO/TlnQcql3/sGTV19JHCwvQafKodDJnKZZcPAwPd47Epiq34xONjqKKK
Hr1xYZfHMmR/BtzeVdAiRHMLLWUMpIGvnhMpVePwEikObbtG9nt5pvflnhhYb2n0
85/wClvijsGRKZnZWI9lJHgNcS6e1unb7EXhNQhF9KDm8eIozkwYMZRvRdTSns/d
Rxa16NLpopQJI9zxT16ZMuihr/39B/ofDWmIs/DibpsDwcegkHSrM17f1B67ysXR
CHoKZ+AQX/FLe3eEV8gbH5kESEvS7IyjhROBHxzuBUJkk4xnRN5FdAwRxa3s1NET
kSGufqV42mHB9sW0zWgKoTyE/ynD43WX4ybtZ+6Ceizk1lthWyHxlRifK5xvFZWG
1MJwNhweG9BZyKPuf/iBMgICMzxfx1Z/1bWlgnOfAUxN3d5qtCs2sAad4qvcSzfD
1dI1pghfkO4zfxFclJAO9n8sAaLBc+6SQHR7w8yj7dv3ZFBRCSD73qphEKNVvVyD
gFjKoVU+fa5xE6epYnCJOBnvgrIAs4r/qUROVKJG0y9kwgR1KQc4s80w+qSnsxGA
`protect end_protected
