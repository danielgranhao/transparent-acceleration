-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
KaDdpEq/NN9pJ9+jhYqr0TOYtu9lcN4KVcZu+P4RchLghhotJ0bhPNBRWjAruZQY
y6uPrj+AxW3UkGT89HfykCnD7RR2rrTNdTD1zbfS2pBUPYtdWSv+PFKsmLplHbIR
pBHuq0HMCBtkaMMULrN7vB7uqpsWy6CEFx+LW/akk0ydtj85OXdd+g==
--pragma protect end_key_block
--pragma protect digest_block
lonhXs36OTEBfTlQFSx4bjfjPEc=
--pragma protect end_digest_block
--pragma protect data_block
RWNWE0v6glUQbI7rLy51SUVe+QEmC9VPfsHZcb/DoHnzl8lHQfqIWGZffGRZrYf3
XYrbqDg3atVDpxnEmqL1g3lYR8nr10YIVur+yQtARxk6Wjo5K2f5xVVghk6JeyjU
ytvmtBrUTy2FL8RNdqUNI+Q/s/NoBPT8GkGd83HkrcSTqngL460TsyVowF8laROG
Hto1qwiMzGjyxv1WPwrbUUljKX1EwXdQHQGmnOy/8cPJ6nMqCV6EE3VkHvo9f6U3
kThT1a9JrFHX9v9iAaCUPftxuGD3xOLQ3cUM7EKi/tQUP4fr5CXzX/TgA+i0vV69
F/dHQS5CM2QZ2zN1HrdB9iz7zNtyJqjDc4jRLpI1W+mFHeW8VRB8qVL/qkmRwHBL
k4AlXJn7e14jXkN2sBuunG3eFWrZ0AeI3hTNrwkb8J9sco9mrpzmkZitNvW1C0zB
tXUIptgWLczc6USzMD16W5hUNR7Lymo1URorEMO6RdZG/K4sIfHfu63ONE4RcD9n
AVqr/jnmJBcd2wqM2FxUNm3Y3gT3pr0vjyIGxO2DFtTQlB6SVRwO971xOEAsfelQ
NHXOKCVEWTwqRACpMceH+x5RybHkf52+miEkduFxoUCOcQiRsDH3x4Zv1B4e9oN3
5bVlezuimAbd1qpFlTJDcG2n2Q8jz6eZcDOO6a7KQYLPZsKDVOmUjYZsjXv4lzCr
X6EiymiL6N9F7hFKGoEETWP7VgO/EilppBlnWI9uW8X0OLZed8Q9zQ8wkbUgGA2+
Q4ebkQ4yOckcZUJMFiOucj/7lV7SaeiUnq9m3EPsXQ3xEQYErxJp/dr0ndQ3InVn
2NZ8QyyDiTmTQ48NCmS8spkzFX0LX7NVN8/SkX8f5W9kdmK/GpGSACxQRkfMQAEG
k3tb1UkgAKDgK68qdTYFCoSgv9hw1ATlr1dUP2e0feFmfbuXII4/imgg6OCq26HR
7WKp2zC4VF7wuvecaqGJNZ+/fkjnhj8vXyCZK4HNMwNUIQKTHTxI5wUUH3u/Kp0g
2mmbpA97XsInb8Q+E1HMbcWlEbyCxZU8nt2NBcEem0fy0kmn/CE4wcNo3VLBA3VE
xIzgkHC8NeCZP5o7qYAZgR40ZB1weye8mMxd0dLN9MkwlUqredCasnVGOa53g2Yw
0HV2btkzI/z2HNCB+C1mWTgbjbUtcp0a0q4r/1S3q8hv5XK6434WHJrAfBZqc9Qn
OgEj38CFM6vy7HoWS2CZLAehtverW7JsFhaLKQp4zKnMmA4KjP7FJDAF/ckYA/uo
n7rZaLrlF6cldlMQOXiPKVMDYIMFC+YIit9or6osIckS5Tds6mjeKpV6fb5zsD90
+leEL/u00+OKOlvtp3cL6hq8RlOb3mS9BdYl2I8XmOiu7O65LmvTPOgK/powp7r0
fTvO9NaPL5zXYH1Ybr3j+xAxOz9sFpxJjaaNyE+oDL78vBPWPYVhfZv4YvhczIKB
BVrUnHcTOjmPV5DLsFeLNDqi6lJRTh7ipMBkfTJjaO2yM4ec4/QwXYL+7bQKORAN
kt8mEDBO2am8rUWaVXvskxnRsXHGfNP/MRIeER7guOmMybbLN74SFGICvinraLOC
tJr/EMYiEAIO5cxJ/qBs60uw3VJ+5V20T3YH6kJswG/4rmq4V/4IDuuiSQMWwUq1
JxaFTRyR8FPdzx+jbo47iKPi/t+1Yfk8zgMG2brpJhhKgAikEIsJc0axwA8n8J6P
DWuvHTL30dJff+xS1gFDIMbNcG0MQVzJh4TSWpiuhh85GiBP6/zyOWUOwl1Trh+P
IqBqTrN4jtzz4lVfdLNNP8PTF6ztM9KfAMGy/KTbtKvIv/NwjeE5601qqdeNOG6W
deMwYe+FZljNzTKsY9Ztam56kxAmC2J0MHQDdXZTl2PuhnIhrkV1DJItn7/ZXoRb
obdZTw+2iud3XMT1lVMOpapGd5cKaTmqZ7IoFVtzWlzohWVnzD2R69PTGtpA9cFs
2G/ZfLF+N6YK8W8jfrPZl/m/S11oBjC59Gq1BkLBj/9/Y9NGMPvGjRd+g21rgD4+
ip3tazInbhDFuhSmbHXNiO/+k7fXDWW5I0r7NUaORBWWkCXLu+NR1hB+y/gySoms
JxyNqqh22KSEmSNUc0ox0SaPpMGDRk8NDLSSTjzclNAQoTZN9db7eJ7cMXAp/t0p
95pmIXzYvTVNeY58bvgxa24B3cLJZLmW4TzC8s7X/HLh5WzIK74icwpZL2GVRB/I
Oz//6NNZhtwbk+SuYz2sh0GDlzT3xCMLDSd+b2xgZzTqmugqfJ5hv4PnoXZiEfEx
DIbjJizrkH79fFrXKcEg6xvjX0C03pEeaacKOHWwkt/zofMMrHWygZ6xR7gPnCDd
sAhnnXzLA2FrVvjr37ZLiwXhC0mknwNv+aB+ZmxpO3x3A6O4GZO8CK9lEDw06Hvc
pzrNOI1O/cFZ/tnlczOH3Sr8FAlw+6UcVMcmd44QMvVFTAbW2GLRpf61DMvulzIC
gg8wlXxqrlSglzeqD/fQnrp4Dw21t2wC/oPNALZ/ChhJw6Epsscm2ahHY3dTjOF7
KGDvLnKnuvz1ZGGlY6I+mHqaXLdL/y3HL15C2WrHUMKnp0ANvjhe5pcpcqxlCqv6
b5RAQis6TMtJeM9LKzSshZbD6IP8N7eCf2TrQOSsovGvZTqqxNGcoLRfsqTQR9Sa
4MmUSZr1hhKQSW+/pJaSnKA0GkTp1rY6uuuC3lwTTlLP+oVh1OR5UudxnLogsuYH
fIAZPtf0VUHgExYmsxu3Y6OQDdyQdzxaE7t+9ETTqiTbDnPRTf8cy/9h7dwSxg0I
5utCdcxr0BSSvp4TGpLoI8+FFAXNeDYpBRdkTbHwCN5fXU0Y4g24l6RmsOetuGns
V1H2r2Cce3XWGvKTmXMO0Iz3SH0Ui42aSWu7FzWa4Nf/OT0Y97/dw0DDO86Oaq/X
88R96IO0EeLr53gex9jBKa8CGKGp8dHzRR1ccpf15dB2biL20D2sqLcOYgjtDSSu
E+zkWRKx3dyw9o4/IbA1U08BcSZdpbB//N/l0LqMO1mCycJegykeE/b31Xddubzx
aDiHydIRate3HRk3HzUHY7yoVvPxQhfHXZUP3e9Opprzpb1U4aEVkfzrdTEFbn87
ONREmCYWuR472Qi42vUOlrJE/BTQXp/4Y2DPUnT3IqUUSlILlZazdWM7kFAbegOO
n5jigroyoJg0AVv4YKBY1vF4OZKoopZ05UXjQLPyCcHAbMm+/3QDkDD92ypce+pL
WpxgiLYohXcqkTGDIC4NgLBhkgkhgU0xaaIYXE1GoEDYdl4lxU3vjm/+FHIrmKJ7
bg7SwwEeZSNtCEGulKxJsE6zSufouwbFkC+d9D8Txnq0vPn3WvMRryi2YFIrgymd
ICubRSBH5V6eM1ezIEwPdsUryxuz2pUvmAI3pqVZlvH7WNdagKVJncwvXfYo2VhO
MzWL0Q+teMneTltfQiYAv0e4rSAM0aJXXi+wBabaKyo0sxNNspyqRr726euvV/28
FI7Mdn9qkwmKVvpPcjWesjAnRCy0gHodtvfVnI/n4iUpTGpj/BEbUmpormJkAejs
pGUH3Vw4gSC+NGo7wkweN4bi6bVC+GEWsqPoK5N2yLF/xmXaf+Z7iiDdxwRpTcFJ
SIH7VLBXDJEnoAXn/GGXTiQv0nme11O67yNMsUcN6cSlcRecoxXRA5RVZ7u6Hg0g
O10sk3RlRzHY8HR66GZ8NijJlyxIILwwBNLZm13dehMwut0tnYqgNk+rWUcYzpF+
oeyFIfp6cJGnXxN4MjYgiPA0lbw0Cbu7xxrnzth60BdpHiBSyJgl9/JXU35QHJRP
V1WdRp2n9xglSwg8jdjToLPpRPdRryuYyLY+uVFT0NZ5mC+KIQAyb3JCjthJlwWr
ZEyobWM3DPW/GVFhw5Dv8AT1xs0P69o0Z7rf3ZPZuciZ8BrxVbCzrzLHzdF96GI+
8raGp0ren7dm+mTNUdTDqoyji+7/NSJfQQVvYzE3eTa76Y85Wo6yyLFjTkIZRtE1
ngHZ/INYFs7gb951hsmpHEesKfBO3vKqpn9guWXMJt7SHkQafR+okjats0MmtRNj
k9XZhUhCWZFYMvjPktJt4qqNqImvWzhGQSpr6zWVGAAjGsAwOktS2UYW6qHXTcrQ
Mgk4NpfLn3HR5ZQXNGUpStpnU5iiybd1WrvljB19B7Gou/ph8gWQE9lUDsz/IByE
HWAKws8RzAfCQq0b90+FO0+d4nm7zjXzYjfxh6C4b5lysf7XgzlkWFU29Gy6Lmkd
2o2ElbtT4zXfDIccpjpr7Hn5tFzwosPT3A04zhGCmpJ88bQEyLwbU7kHEKnc3uY8
wkt2/xaeY4n5wR3s7izCJej2QDZqtnMpY9J36Cwb4EineF832WBKoZ5Sz3Qz7MAm
+2s9itWbvmjxELnE83MmzXcgUyuaYgM2mbxhtcuE2t101cmhP8kGmljD8Y6DSm2z
WCvYfaIm2zBnjbOxm/B3x0/7BaWZ+V34dlFick8aVxZ/xnePBmvgc6jvXYZQTgmy
RU5u8CY20qUn/CE2O/0jRPUVPkSNjPe800S8rJ1ohDOD5SeiXlRGtxBt9cmGux6t
80TH2mm7hEBRGE16sgo/krBrtSJsr/vkQDG8DSjWP4UqgVb3ITxFJg9tFfiHkrfx
paNlX52BO3Mmm2Ic9DtW5I0oduXunsgB/kNIAqrejxUvCNtYg+HDcjVlNvJD4Ngb
f954ftxxnK5n2m7yzWqaETxgGvFG9T2a3FrDjj5S+tPQOcAjuSV5w/3tttTOG+EC
R8ZJoiTMsDR+bok5CZifRGfUf3vuCCVU07fP6+ZoLiMqO7HPc4zeQmA7RGmi7asX
zxudwPKJeDddkcDHmEWXhk9rWXDQLDiP2+uQJllivD/t430m0eItsaM5hp7MlEWn
5+QHRswx+/iJd1T5NIJg94Q57MKWwDwEfwaL1TKLlPN91kzrU96DxdWyeqd03CrW
jTWXPb9e1p5fSSPGEjwNOOcQygEh+E2Tqu2xeOzAEv6m0jrQ3zY37Vrn5rw/5uLN
mzVipoosHK1TAHF7Ss0fkD/04BKjL+nCpFGgSJ2o4mhfXyxxbjn3jpBh++Ltx9yy
sNTxAYmQ/hKRFvOeqDjfcJbmyuh9ZNREL9cNQGUGIzxnz/3ZviSrIRQOpBWuswx2
EjoA8YEfaa9LpOYZuvFHdfVCvOwFwmYMJMmSzDOY2B8UeqFH9JFJHwYh4eJPbwU2
3PKOt6v5lJ+E67+0W19CIdZ90ie6nn2KJFTdd2kVE5Wf/HhmElsI6H5U91xDfPsP
3mzawaEJH7ANco5Nc9W6lMynddBQ2KwWAu7KqgPAcrZp+jJAGjT/jhtBRDYCt4m1
euHMqZUIw2E2zvxfhFGDiIHXBCefy1nrJYxb1JwDo8avC0UulEr9H/OP0+QmTPhT
oPc31nE5/HaUUHW9x5DAQzduriiXPATPWLvEcSHWzNLVW0nNFZvgKqi0YPDKPuOu
8Nd8On7Jj1sEki5SgtswZB6HL8PQ/MW6AqylY+gT5HMSX0/H9bFO4bgP2uVGdNDZ
4sFu8FgZCg8E6TWkzlLAT6Xe+7J1wlRKmvEKd8h5PWvdkrdWfdI1c+ydSzrREaaT
phStiEBX66qHSRUnDn8eZGdpBJz/Rx892wd2DrCXE1TiFRpUR23ar/VNwGwzA0jN
VH/f/+TPMJJyP5txqtCsNCqQfTYYxXqn/GwFgCVqGTa9yLCFYRANFejNOExZjWC4
iXbHXS44eF6hIyS3h8gu1IoS9YkPcdi1jUtGGBRDmhsulTvfzho6faEJTBAnEnid
NOb6RLyWHVqNxxr3A8UlT9PQbKxM0XJ9e8GgoqnF/wLrhDJxMltLg/TQo62GmNly
WuoAE4LKD3iHdmarruP9RiDCX653rLnwY5I7HcNL4CBqh1vaWoYLJ7fwP5LvVzi+
wrxUCvAiFVVnBArofT+A4qF5dJCdKGttSsjqYvhrbrc00GlgnUzD2DcGHCtY6LeM
gHEqohVsHuCGI2vYRNwkvFuBBCTa22KN0lmnEOjDFozAGjL+XwOGcDIf4Ky6H7iW
Y1/B+7wXCBGM3j4PUxBm9VxzDFLt6g92Vp6CEJasXl4UnLiu9mIIkbsj9S0+eHYc
OUIHUGMBT/3H4ov2R3JUn/PboKnoOvkOGZdgv55TdPzW9hqPiSbiPRZ1Nl57ASIB
Tckl8pO6FNNXg8ifJvdKfP73jWKjPwUaGM4gVAzFMcU5A/vGouwp3rZ+mZx79qRt
lLdhTpkMxKm33vSQe41zL1XAjCNrEHw7i0IspPJR1Z8tdqDBXdYb6gqNrPo46mij
vV1mP4OT3woJn8IMzTmC06qOgE++c94Zy8aSRbNPPjh3tkL5WD3HecKh7JuapIbt
75sB7XvBbb9GeUIK+P1G+IdjfekcPWhhptOavEqV6PXWqp3WQCb/HZuYwrI4grsg
n6zK/w21wqG++Wy4C8NoYoZ/TRxKeoQ75L2L3xc4rIZac5UjeVYnpXVVD3RfCvI0
M3CnuBbNuJSiIkkWTz4CWLREMpO7o925LyluGothqWO6J85iRw+ImZ4Jjwk6cx8E
6IJPXd8INr3KA+LKwMOJeRlPB3KN4M7W9AnNz1S+bm80HMJa0BbqKGG+mZvTwUSo
rjVqDX/Fpj8fCT86B3zabMVo0xb9ZpX2y6nwKRvoWdlODpObUA3UQJlCyJDjYO7I
BV0XrIKiZ/xRC5KWxlcL9NHhHlBTrNrpVCpA8QNwKL6i9NDz5KCxe1RtKGmYDboE
2HrEPBG/l3e8UJm08rqheZp95hbE69M1d4bgZ4N4XzEeaT+f3+AtvE+3/1YkXe5v
VUtMZRYFTXhWYdmm7G+vzLEGRUJ6IkrxV3QvVeW9wGxdN9V1AMWHclqmm+S5yPUE
xA1GQP42TUwxgY0a4y9IkRXhcp8E3/tTOvLO5P+m9/5MHWbY2lkHJChK1pnlprfF
H/kB0RW9QQRZoueallFZoveHIos3Rd07+JTpcfSDleqqcxpWOoPRoXS9PSbj//ZS
h6N5ei7xM6Lk4AoJ4wDcrdKXkxg9YNs1y/XYGAlRsuiYbwOHSEKTBsRdUR2jtNow
HpzwUcKmJ+fp5VCp2+myhm8cpnygBvM3iSyk1NOFC1Qa+/tGZvy4MCLxRt0GKeKL
6B1NcWZ0vK9VSyhKnPUvu6zAamx2fvl8GkHWJ+o0noQiXRUfgDZqqMtcDxMcsjmu
A1ZrxduRHDlMA20ij7fALUkHZB5oJhHIdf+M5VjcG7jgsBr01nQARapU5Q1QE/Yo
NcvZVa7I9ECOoz/0YOJeAU14pYMjWu0edkNJ8q3/vGSY+13UfEG7xm+miSVm2Tkk
e/Chg9L3bTy7BCJEMibNCFv+3aGcFSWtAFSksjosmwaGscrtMAO0R3vxrojmu3h+
bs3yEAWuPgbPJ6NT86cQeVytYWe19DyLy1gNNH5ZA3HEIYdlMFl/rP5IQl1JI0cC
0VrZgGW6Vu2KVHlEZKxBkwM4ptCv9vBYnSBR5/6+qfQ+exW819tdQ68do2gSYY0I
FrEvGD6AHjDAHzMI0GaFTW6aYjkhhyQ3E5n61EzZh6JXvldUbIEN4zGmPWQTdWHh
ESa1Yj+utHKi2Gke8cAddOyywkIlmHAchXp2s/xk/Uw3yvRbpBtEi4STMYjygrPG
iFmU/hdOHgCVa8GFxim2U1xR5BCt3gMBCYzEpQsV0NRbPb0CQ3HZCECYVmRlEZI2
Cv+xyxbPgzPMILCStM4wI3+iwHYb+pifi0975Kt0W/q4W4e6uM1r+fNt9DTPb1Mb
xoSNc/eOlBKFkl1bAb1QwLP9u8+gRQF+ZkkOunPGka8DZ96BhCTomvggOc9yDMxx
EcBZz6ZclnsLx+VhGKdfYZ6n6dNNPShquzEiH99BiF1pMwTUqFFciVqRcCC3DerQ
iCvpTvKLqOqeR0JKulmbveontaLMzPHxohuUA6I73PeqwEAE4nEfEnea9ayMA0KI
DTRDcOkHeqHq9KdDoVwEWzO6Xkd3SCRM51TKKWCaar6Y05otKbNGqFVeoqTKaaia
Ccyt1Yl6NzLVkfncasgF3O4cvURGA57z0ks0iROEVMSd9I3Ztj791rjPgcU6u2RP
vJFbINiqhJnzuL9APKVg5QCJzJsJl1++SWAoEyoLJvUoLXpvVaKa+pZi8E1LXbMB
w8RHwPphbYNL197SLtCv8AadTjjFz5uYA79Djaa7FO9OTFRB9oBz1qNDmr5A8GFX
HafGn0qU7gUppzhKtVM7WzfEROXjiGlgJc3uHuT6bz2DqH3b58Sa5XE8+J1Fcoax
RzRccQElpfV/jN/g8sQtN8T46EPY+3GDgwiZWeJLB+re5kCxztsdZ6ecp7EhAGg5
x9ix7nS2xQPIkxZwms+pR7DOerkc7pJ6lGXdn6kZF2z5qTzwCZZOf14/jMaJc68t
50ctcUy+keHgIxMW9gCQtQ8xOEFkfx0Z4FJs6x3eiTNIjlEh33KCTbyn0p5TQEFU
8Hde1+mpSFpoHY3kZ5p6zYODbkoHeYOzT3xRafjUoEhMh+DDqoNQVRJYv/xP/aDd
rKi3/JoAifIEGvnwP6kVjf+y7q93c2RLkdH5LjQeHhPQM0Ea3RuYlgheFbFQuV/X
/AVrCwGQ+sC3vTfP6qtkoyPmI9tGFbSVTSdQ4mrKLS3mjVW8rLjEg+tLTPsgfOds
T9YYxjRrBKYV8tiAknm2yPjN7XY1naN6lrvXlO3TEGXtHj8uA/h7umoYeklEfKuC
oyFdxDqoMoSnCxBZyRdAg0qpeiSfcDiKOaDQFL0pvmgguOQly3W1sLnnXwk5Xa3x
QwNa8CFGoanUbM1p9FtWzbGUN58RSLs+aMvWNWTwh/MPfU8bLRAsISNT/Y+cotsw
VTkrK6kM4iuc2kjOK9ga/9DFhqiFRhyDVBalauBlu90JfYeWfNj4WkN052PRTWXA
hF/I+0o2opcRSyh/eyywE1Mp7x/4e+cNcMqQwR3nKx+6y0652Di9I8ZA6VsrVFx7
6dYhJu0K7DK2Ef+mr61Cn0KwJEEExPSHMs2vbZVdqcaxLB1CC0boOOQLqQryiTcl
VFtd/PTSRUoV/eftsQazqpdVt/9UL7Y3K4uYEAUOTBt8vpJPQBr6dWtvDy/HYLeY
X2WvN4yZY8ALlHd9u0kJrP0LJl64ty+YOjWqNRJGZAMM+dySj3ZdHQrBi1xoKUF+
hgHO6TlcW7JfwJAvIksL4tsOQi/iN6F9Y2ysEQ9KDQOnEKl9KZdMl03wAz4UH60z
BIu0ura1jHF34HoD+BuEzSc/QRNteWQghiptgXoY4CCIJx5xYEhUiEZMSCfYa5WN
gUH0wLmviLQBeYU7wH0C23sK8gLn0Yfy7zaCmoHixbMREKCPJb5crbqUKfixJPb5
2KWnWJUBVtWsmLoh6LXE4fWfM9t270TdXVyneUyaQQM8lS8aW0OkF7VUXY4aEmiQ
IbysLboFvCN7Iau62heRefIi01Zjy/0UJMNSkb0JVHp1FO7oLT2JEwyTeZRcE52S
WULnbgKG0/j2Ks2B0nk/ZNSvCzigh9PLuRsPC9LALCTnf+O7bGVKKf8LvSUsOKjk
c0PnFhvH3Yq26dYc6PTc7tVwNbjLi7cwWFCEVCwiKzaevHS6+U5cKpk9Yfv3uK75
JSK7p7/PN4PlASP9EacxtEJp3hQirehb6MbmubqZp28n4YS5AdYYgSXrMMjWX7Hv
nS+C2AEVkm7FrjTJon0Q/s8bE53/N0vNV9jA1OlNLWtRI4PUohUXsdZRmrKPWmf9
JsZR/6NSsEWUzcSLpNbJNU8XNLI5jqN690He0Z97JNr0vGqaBivFfIuMe751pip/
fCyBkuzFQNcfvgCuxcX29JB2WRHcad0kuTJEMmh1Ljs2b3BY9uDigFrmF/wuJ0AO
2Un18NkRd04aLazH15vff7LZ66WsrpHkfWk1IYDzDAg5NgLxxtp/QlKf4xLQJmEg
kjyFts4K/LQ697/zDezTAwFShBn9FuvQ+u7Dvl0hPeAacr7BnUp8zBEfPzZaML5B
v1U5QCOMmJ7zTXrXUC/2NxaIsedAzHukW6MteT0OfT12g/MkNOKe3eJ9/Sy1CQhl
V8n7bnEBQeTQvxc5V98BaRZj89XARy22L3EpWiMkvGTMMt7kYdwCZqrr1C2IsuN6
AzjRtyVSg6/a+DQQtPaemvgWE/LTr9nJivSnzIzrQSWrsc9caXb+HlztQ+ZlTN2G
Utr6UxN6ODGKxTRZOtg5PDV8f3RMzj1qgPPCv1HsCM4A7lqUeVhd8/JipMeT67fj
3aWVuGuWNmUjhJoy3kGZ/ntlqjr74Ep9AnRQ7P3hnLc/KpRLaG01eWshbpatkuQ5
uwykG9UU/XRvvnqLdWbBgX5gE1IoMy+X4d90n0PlUN9ayq+WYMOLcdegzFqhOt3V
VgeROr1Sb2qpK2NTL3qsJ4kX1l3j91WHay7vsgBv46xmo8qEp+61okZ1uLC0qvZF
m6lz/Lrez7l7mUdRCzUm155XCCYsHYWuyQvumFq6kTE7QS0QPLb5JmEqz3ycpjnr
+7jpSvKz/3NvfP5b4EToTAUfAdpHp34ydk+vkkxia4huR0uu5frt7YHYCA9YNVKx
DQiRWkNMydaq9hU6kNv7qhUo2O8ElEaXXHx1K65Pl0WprLFcB5tJYqKYkwFgMCse
R7nBrpBT4SRNaeQKOzAaaF5mspNccntcEKvdtcfopfocGUnFaGcr2eUvMwjQqugh
iQDvw+blFuz1dAOsT2htVx8nBktMMRYShzo2Ypl9HMsD3BovLU42pH3D5DLMgzlU
BErGrtmWluvDjsQoNQXAKZ7PgqLjme3enKceyifGbHBxpmKlUMGeWHaQlNSnM1ul
S3znT8y5qlLlUVeBSpIiidESX/KJ4EOMVucyVw75XmOfLSsqcSodzkJQ6IW6OFPh
ULVqqEX7jZUh+8VWkk3CN8KN2RV4DUvP2yHsW1MLRG7plxhjdiTsYyYoF6DQV6y9
cK5rK52tzI3HjwqiOWuuDxq6TOuXy5gkUfJ90gcdPspUK0R4ylNJFo4gHH19pn8b
/1np9E6eBeYUpu8lbAuXSrntvcppBd0X+lLLPDhjLORc2jay2lqIC89qWAs9VmJa
Hr0MicdYQ2wNM2+E3rZBw2yWrVHvRKN/yz/FuI2HT/yA5s3gnpAa8ndyjKiMOMdr
mSf22wfkuEGq/xjtwygfsUMQFwG0iMtS/+w7Wignp0q7qTmg/ojB0r8lFNOIJV8f
WwXPkejg9XwhQYsUEKOsYBKfCdR7nDX0YM/CV1DCVGcJ9Yp5CYFqKEhVmooPf+/d
1k0R0Gzi38NO53S76B9v4RQ1KxH/YramnyFRy3vRy77JDsDJ4aauMRWCMzu/nXfW
39+TzzIKz1ggrF28e8tpLyWQRKl5r+nVOdNQVN06JXa7n4deGThLBZXXzLm/IoIG
S/jeh9sLjqIc3hnlzk1EZ0SNESJZwhVYzbRTUBS9GsiyNF5xVibHpWm0xYoBcp09
b/6PjV8dr4Phma+k8E2/dTuGsNUL2dzgnKMBURUAzbWx5D+RAGuFumtwfAwwGSEw
jNobG92kGgg8ZAja93H0sP59Cr5vOgf/VZJLtmWb/NiAghCEbuVJJOm2KJuNPOiP
elcGHe3cx7Ti0YAXPtszhGksMfpxAqXLbkZ+9VT+no7eJEcH3Tmwo459506BzudG
wGzTmm/D01w0dz2gKa7TcghmGnaUuzWlOQBzMLOuXhyf0oJLFCe4VAR3joolWdMI
zzU9m9MEh/KuhHZYhjSqXWZPfoxXbugrSbXhfIpkVFOxphs38uEAX0tmLLFN7yxI
CR9QVbLH6u9l9w37f9elckwogdexT7/hkutKv3dMCGlMxCtR3dW3lBJG7Yl7T+05
Nn+MxQtczuu8gAVFbn0kJXe1QBhobOLoru0Ql0t0JBb2QWLvWYyOM6WTFQXhmUk7
HTnhLfms7qfpOg1xATUz5SUqT3Nj5+M4eTHnCKmG8dv4AHt2+tlPfKLfJq+KGaJ6
d4/lFgPCxCt1RVYEkG7mhziYb5j5OgjTtJLP4GcnTtkY1eCR1HJCjakZwf/yiV9h
SJSNCQJlMVkRoojBPzlC6Q2w6DW90shgL+mdr5NZTnx3xRgCSE3XyzlFFuT12ybu
mejfJXbzsIEb6vRwqdjkRIz8FqUvDusDT64F0e/JDtQNZO4hw8CBQZ3ClpDKCpbu
P3VJqBqCCKylFeYgM/flOVp1Rruq414hAL6yg7FI5JxER6DLQOcIGn9S3T0VABq7
hyf9HRRddmtL1+TFBtpISJxC3ZjfEaQnqeHG8m/fo9VpiwyocMSGtc0JlP2mGnmN
jf2zz8P98ttsKhUw6nHuPZU02wIlxoE5TWpLLqLBebnDnTGeZrpWfmGCTBZ7BVeD
yhFd8Zt6V0npvkG0uXyI2LdmUBW+7dVY7r776N8Z4BeJc7MsjSDIglcEXr8UJZK7
LXKafr3uw1EyzA2H/UX0dwS2D9omfn7ao4+HlXcG5suoBpb46ASHPBKvfvnTyIgt
jqjzTO+afsbnVhXr7n3tq5tqQatif2ZZYBaQVPclc5VcZl7H3bzIOq5hHicFIcYX
eDZfT4bqFQeeaKdpKoQfe02wWd5L6ARGq20PlRyL6XeLfAeAD86p2j7GtdJYFm5C
iwjZowRYGiulaIwMsSBtfAodHwJM+nBezG4Bc+b9blqWV+Po6VlanHXOt9YeLGee
W6ia4EKtvXXoxNCzHsNH0vuxDHltTnrHBiHYlPUpVPhzP1BpKnK/0EXMDaB2MbYu
kzFHkNgJikOSMom/BDa65dk16ROT2rgpSeVBkozqmNCuUXbzzX7Kdh1RFLhBRcLF
aPYr+6SKE4A3Q9OBqMWBOPgD8CveIqtMXZE6r6XLXk3G5NwgUvPpKeSMakxp7VBI
o/wljyR/qb5GFO9qMkjHgWGrHVds/CmYl2Ny8I8nv54gKp2aUQ1ONd3kVNDV20MW
D9M3eI5WFsJqKbEnuvwMouchjy5f3pFRlXDtbAOUC6RdbJk2ohwIFA5yucy0f5MW
zxnQhxRxp4olt8MZaNN6FRNcwzH1XoabCAD9tyJWyUNliH6Z1eR6/NyzDkqVeBsG
J9Sbj4SJlPWDMA76Qjb4vC01SV6FozfvKNCx8XGYPbBsZo11fmdKGtfipLDckJCN
uGn7SO6ZOfVtMIuzTIj0CktzHQBsa4nWDgljIpitI6JAtb2WZuhpszeKxOMhEhPX
hT6JZtzd6gi1iIQxnnHihLwkDJ8l2BLOwps0rewXVnYHj6GGrTN+uF0GeaapBzPk
8XPD0ZLw7mJIx7i5wVLyVafKsTzhbe0N5gooK9T3rg9jRlo70Cy5Zkn4WP0DqMlM
FoPTYyXzLG8m8cpKCqtvMd/cI6vSw4Qr8u9Oll4f+XnCAYrCJXvX2Qy6G6Us0RaH
CkrVpCiJsN4toPAV1zRTOw8QdP4jEnIxqhQxGblIjfI5nOetMpWS83PKo8fULaan
BAyO/mWD/mbVG8hZHUUMH4bHpHG2rIBE5Wb7s2nQE+kirS7PDH75uy47AfwEQKTU
xyYR4DbyOl88Q/njJpZESX6G7wMGXf3McN/RVcY5pdATUvUzSPtEoA2RdxUPQnlS
M9E5iUiQadGi384G5hxnJ35VO2Odawj0iGVkbwyWlHPMvLJqCqIoQMYwtnH0REk5
SDS9lj1gcF8qtmRkRgwtdVKGf4LEt0S+0iXXazo7nRxeArJPg2KxnqDIxR7imXsk
L9pxblhcSmODmCoQuZR04IQ/p38QNXJxQiaqy2lzninBFIG7rEQguAhwRX5AjKZ2
iqOS4RrtwK1CAzfAEUitnpcFmpzYLIaY9gXC/oaS3JvWvdhHYnj/JiVSQgEpI4nw
3PUkOSTm0DsfojV8vwPSeXyK2esjPmSuOnEAcESPc1slXnH/a1HA+8OTdLwliKgG
AOHTZKQ+yfQsV9BvY04tt7/Lf0n1uV6iObqG6YwW6s+608TRTTKW3StgkNucJRpg
nJeuWSWdKQvmP6qUktQWdKxb6Pl3Gq2VvXFZ8n0cplvg/rlr5cYNS9vXplbTjOAj
ixmKv+wGFJtatRgTVaIU24i6B5c1W78lTBX76zPOxT67ijWjvX0zT2yvgvxrSBJR
9fyKabfKcsowLNN+7xFEdbsFMmcCr90JuQdQr2+uIpdXalltE+3AT5KmdvcmBskS
5GJMCFoxebzbMkBZJ6uG5/sqX1tffJ8slrKvkj3oezQSUzjKRE33ItSaToVIQetj
OwjITOC8tevCqcSHqraftFDaEgr0aWehBOvm3Tx9bmkq1ScpspMkjrK+yLARFOPM
/0d/vLDBUPtcDtU5x3Emr/UywZaOelE7qNoTRs+e2ZtVtXK+MnAP6QPJHV5R3mJ1
wivpJZUmB8QwKUMS7/tUCGVFcvdz6bMmpKzd/SMuzSCnB5OjYfMPRPdEWWokDkTO
3n1kdvYqcI9cs/XYzHo/eGxs4yRWs5tp8oLeCfDju6Z61A6+lgm7L7UXjpJMVtMo
0Z56qMlGOtW3vzRYtGbL/SqI3KHJkgj1WeQWwsbSe9yHR2CyIkOsKHqxbDD57Y/b
RScpUjJYUjy8CWcd9iQMfLp9jjceqaTva6S+OY5OE9veYlpX+e58gKyaNJjqwGuY
+C1eRLCu2CjtfXrKCHInFIySoqGDGmC8ONg6bXlqniD1f8mzwvOg8GK+mmfOKAKA
iw6pk8oNhznHdNBXc3Zk2mMYaLLea7TZw7THx5cSsN4YVdws99ICDcLadP2qK+8E
mAs3bVKGB0+GH2pG+Fz2lYJUiqG6ou+6dWOIBpBTlGywQHW0AjD14XU2wKn9Vm7+
V1FQxB0A7ezu1eCsIKdGF4NwMwCkDLNRCabyrkEqgW8Ds8OORHu+2d/ppYX3hAUX
4ONr1S+DMMEnb2xqS6UFXDjVu+dixvT/7SocY4UFbknFzmUaEUzIgTxbEDQnHcG2
F5BrB+tLK/896u4eereiFXpOBAshotNvcIDzzGmdVl9byVdMwGljRUu1FfI2BrAu
4AI7CQ2eh4UH+2DYH3RcwU0gTCVoHPZQEROMftzqPXXENbfOP3fDCCruirxjUV4o
HOhR79HMMxche3E4wOn51OYnyM3JJc6phXKYZRvwTD4yy9HzMMOrj/1Ccpc8pVPO
m2nyzY3ZoZpM9k/jtdI+QRGl244/O3BdUH4SSeZdXiwWxM87JO2BX/pAzGty8nhK
S0DL+Hdpi0Rxoa17QHmNGMQV33rtSjAKLyTmLmimY8G8IGhDMzNPmV3qnpf5gYEI
wvrMsgqvITfmVK5oX0ohqSWnb99Ed6QlEAP6BIBmp7oguRabPYa4tCMN9ExDj/S6
fILFUjvxcB8ie1dMonNa6XQ1eGE2p4o3DtQzTGYusAB4rA+VNG9mRup3Gk2isyzY
8/XOuPfyyGux9DBBlhHEoTTZbmK+j1EHHQ7xHV7stuG0Vw+hRFxWhpU4K7LEasOk
uk3ydWTvqIKJ5Ex2QyvqfjK2y8p5rc4G49aPvHfnUIr5H6POHOgYfxInx++oHzUo
q069eyzbEYZnQ0/G6zQNgI7+NC078lvx17/BkGYP4iwI7JBsPnVx79z5/NycKjmc
DcW66ZdDuAFpkt7QzG8r9f7bi5FP0U1VVftco0qHpGX6Gb+4kVphx1ZCBHUYCOak
BMECi+nQJ9O/+JkXsVCfb11dQm3FEwhMboGNx7rYQtCAtoEFMSfQBTgjF7UhiCjD
f50peA2+sXTQEEF8a8lb4NpRAdghx2aAkT2n7XKQZROiluEH/F7lSLC0JcNyb4dC
0AG+0q1wQlvnT0NjaRSbskvhhVDUOScYm8IqHFg16/929rtRCixwpLbIONz5a/5R
vjUmFO+ZyA0IWeC9VCM6tNG+1l7C4eBQ/yMhby9HWT07ninWnLj6aqtwbLYi4h+3
3KgxcBknu4nrBoEwBv8xUMfayf4MlFajMOuZX4hFbFQC6ly0UKQHJ/+bEmREiHBz
lHyQNDDJHxqaq9psjG8NHmk1V2nYdCKCHU1TLxWcHbc9rbcwEbsU8GpKKDbi9DBy
N0kd5k1asasIJAW5xzFBFCbBpyWAYMlyYnYS7R6P6NN5CP2Nwd4ozM/DstthYPG1
iiQf6z/UsRA8RZUQ/fwJL8Ge75gem2cByH0Ua+Q8N2fpABZUkzxW7Tzwa8i0CBx2
d3ppeqOK2GMtNVKGMWWRG16IbXqXxNHQIrjET8pXMW55oqMn3TFYR0lkQXJhs6TR
Zf+ppmcu+8sOZLGSFXAGqbMVeSAo2PxCJlTyus4uobAI20unO9Tiawdl/KPuilkr
Y4hqdh6t8a0um4SQ8na6MFKNxkNfnKU442gCkPKYqkpPKk49Ifn9z3GRgu4PT1iG
s3S7RG2t+Yvb8BN3eKey/oFS44yZnyARQYi1xByrU+Vc8pm64NPAEUc3drwgbmmA
GK6cDOaQXCHNWOk8nHUVP6GHvmLwdnEue3CMEBQYeztO6XZqQVc/8dI1+Lv/6rKd
enN8C2IUuAUrm+0+q2q7T34uSSA4nMwdoU2FV3PO9Q568yX4mSH385QXWwkTFGRO
cTsctCGiX8mwQ1E+VtQbkE3eR1oPEcCJSrawyggqVJvOreDqlaw0vm1E3YUJVFUZ
wTAIbNsnVFcUm3c2lpUZRWFulN/33cPgEwwg2bTqxuuJzDw3UmdH08J55NWONdRo
rXUM38UTpoJlnFn86vSWTK+UyXmPFXLlOagHShdiXyHsGI2IKVWUdgfV9mjJwGce
jKClCJRqWBJAt0HxL58mwl4jzJCMKpIvgpBAwsUaS6wEx+qh61GPF0lnnlWlMEfK
bmSTCB5w8gidx4ORCAW0CPs2XU2iayeh+X5IpghHztkbzulbrlA2Icvf/CVuP0sm
UyGq12/o8CNsPQ10kzQGTuff6h7kaRHv1MQNhbdFsfFe/QYdS4Xnw21ADpT7pA05
7xo/yXzAi+wab/e9lYj0qT9+sE7flT3u2vvMZu66M85re/RLfTHDm35NqCYxE/uh
jduDHyxqs9Fva0/Gke7VRRbGCLGsMqtyBwnqG2aSaaYsd08riPumDrzmqH07Zxrk
ql65ZM6y0fKv4hJznYWdeMDLkNxpeFYTslQljZJEG+Fr7E0K4lsmCG285Qjk3DU3
BoznDYLHVny9bkbVnUy7HiP408MCmsK5ayG54taQdBR9A5ReRKVYoWoenjYwzytl
Vn2g9IM78fOwpgFb4UZGvW6q5BMjFwAYaG6dqMdPXDT+B34OKTj5c0WRThlobF4l
I3KAbf9f+SCYgZO4tWyJD3Fqk+9UXQmNUYPGzK0PucpSn3zhvz85c2JCNzn3Yk/v
lFMMF/3TgoYeH+v9aVIj5WGrerkHX28zuMHVMTV0du0fOzzHyEDafKpOZa4kYFWf
A3AAeic3CN9YidB7qOQcFF5/lFYBMhmiaAae480l3ly3ASbckZIifH20Wmt+sJVm
cq9YM7vYFWn7P0hvG2rDEU/KdG9k697k/TWKIXwHUMcarfVQbBE2rJJQsDRdDdNx
QRuiZfL3xadAwXw1xETNihAdHngAhOBYxmXBJbxCEn00p6yJ1j7PywdVE7q3du7R
u3VCs77kRKTt21DKOh8Cl6Hy/mfxQaZVbZWFG2UYR89Ofptd5+ddv/yP/JOVyMF6
/mFov3Wn2PA3je+HVV1/6YuyB2Rm6wxPPMvSnxFzVlu31sUp/QHgidq41g5MZ4uG
wsUcofl3O8s197Bqu99DRugF3L441TGph1qAs9kd4qqk6soXa2xqNuT1W5zAMP/v
dIXSbeMV5EprS7Js5fKjFg7xUw11uN4NDJnCw6SLVmQ0sCX+186AtfhTIyuA1Bis
Ol+rmBQ/0b/DxEz633WWJ8Rl4P0Ma/9P3NdVNCPCvt4enO9q6kmZl4DpTFlff4Nt
1B6xI5YhQlcfgnt0U0Lrm1TaULJqNyapdksy3Lc0/D7aTi8mA6IVdI1bH8cTyZqD
trhmz3ehfwWvXnUaH6xck5c5dlnLfdhN8iqW4O5WWNIrEz60KxJRAF+0bD2okvAU
hx+Z/0aVMle6tLTalcgS7HdJrMCA87HwYQG9+SpGfQTkPA1MMi/8sZhcJB+2oFxO
pdpoImK2+94HZ7pIVdFGZ4/pOKYkTe3Q65zAHIUjWaYad9z34qU159lqXDf1P7dc
hG5LHfbqNiMz2JiTG9KtKix767DF+DjmSVjNv3WWoEs61Kx05JFZVFV6fvzjW0eU
9a/XWeDmVAwsDAIzOAEH6ZZB/5CANx1DCXfnhAQoW5Yycc616h4VGBBJc3eTAEBz
BahziNvQAfOrlzVitdVt3d81L+QtPfppvH5t5L+9VgBMLVLawJJI2SmKuhvSP9Ht
AwFb98baoFep/mR3US+Vy17ktWVCw/3A5OuApXe9few=
--pragma protect end_data_block
--pragma protect digest_block
5GBnD9DLRnnWqWQBnFfnxb8xTTg=
--pragma protect end_digest_block
--pragma protect end_protected
