-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
jSGoPabGAcvAYSGTL80U9JSfsNNNbuno/CzDpOgNuy+Rhh72upqSXgjFFdyXjn68
7Ir1PlWf+3oKTCAS1/fDV+3dGNpjnhK8i2TNblPkozIs1+DkYSnnISpLIIKqePwo
IpIwyab3dEiXmEOBIeDwK3oGQgPOf48hIT68W7HmIYo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 23298)

`protect DATA_BLOCK
+o1ENJMMkgjV7p+aq1sW64jYcfn09waJhYcsbNxgnpXIcTHbHlEeucrp3Hfy+7ci
IPVaoerQ19DEVNdDNpFCP2iMZhBFatLSzKxQIiUbh7C6Gqg2Sf7l25yNA/gZAqRd
JVdPmms8GhY2fMP7aJVGDb6HQ6XCHlKa7q3WQvruZ08uZzcQ2BfkuAUCAUIslfwd
dO74402+OM+aW9g6W9hANIW4SQaCeEnUiR5zOqcSKl4ohezGGI59LK0SAUAlZR9Q
eZG9xSBWC4qxwmjCui6aSsJ4NtgirOzRzgqqnD8xXodVJ3EpbAfwVTQpy7RuZCM+
i25M6Zx+YG3nBTmEgTlCoHgPBVGFTk9qytnbb7eC6vbiRpOm+qXbg/RzQVlQdybQ
VQmWgFE5654//i/0PYgEYJ/Q89d7sJ0CSM/GpYNmJgfPWdfq5zPWRHz1LuzfQDPZ
tq/WhwtQd9GlFOfvzf9PhdnImU6WK17TU1BL21oAgedufPO/1CEuEcN+8sAT6m/Y
dBipAwpJBaC7CFZbcMwQ0j2XJc4ayyZp8DMl5MX8vhZjiU/Bv1B/wqDX/WeH8q3S
HPf7a7UcId34UA1YceOM04Mq7+71Ej4ft5NHJ7IN57UgTVbLTp3iiy1nHheXCVVe
xzHkSCkCGJF9EeZGnzB4WIo9uwA/nRDWNc0bN3WAYUCjUQ9GvM2eGUBAr4ZiV5NB
NHr542DzBPmf4eCtUDtrIOEc9fjdN0gC+RJPHsBsgXzMbz3Xb5UGl/pD8/ZdKSm5
U3FcTgcFzE7ED54778njw3nPkkOSNJ/NFFFHynOPtsA6Lt+98aTMIyXwjW/es6xR
sfekKIoBYtxzPt6kY7tmt1/jPH/XEAepUclpTbhuGiDQk4vFDEc/1e3AKSnyzDZ2
r9dBME5c2HzPCsELHqVO8Qk515cGYhpkbCBOIm9cdPdWScdOuKYUnadKxexR7njv
pP3wTGt0xpcB559L+AbtN3XBPkb4XzScXay0wiWE2GhZpCQq9ealoz4Kbm45VSjA
swB6l5rKjZx/Fb06oL11UdDXjju2+Ql05AoRvi8NvdpIKyHXOzLrl/ULAK75H69E
9fB12BPYTDOt7BHaxnfHdtWMwD2gj2mQO/x/gSJYpTEPc1IzZ0hQsOcii7DEiEXR
jJtpyCEJZZpZ3slnteFaIQ8a3Jf20iMGRPLtVAHypI36pgsaSynmH2LpcQW7nkp1
KXKorP9IkhwESgSj8ov4CfCmEmN0PbvzA3rQ93jurIdujU+ivMrwENQsxCjgPrRJ
Fh7Vu9BMKIFQK9bblcrlyxmPgEuqT7JbX15NVxXwR0dbBkSm2oKBARIoRXc7/NBk
uqY+HPhVLp7nh95scLrcGGNAsFVg8BRyaH55uGDz3ulRzqZb+8Y2po6YPbO5Gz4G
4sCZPKY9KKPjJ8WtGvHfKn2cSGRWJYnYJnxHfkbSy/XH1v+lOUkXtZ/VMQt3kwfp
CbfIndDEApeLUi3TBzMelOlfijHK9AJi51JnxY+xtBlZGUE4lfFuy2+kbFRe3hek
EkABIIRG5875Uo7falu3PubmHKXfSaSsn/jUabWJzaB/2wwSYbPlzD1bP3ivmE6N
6ZepvJus8xHMWuyQUKx92RBn5hvr1O4Z9WhMYmtQ6m3tNu/En3z7P9TatwY2UBa0
e47Y4zxReBMl6PSy+ac9XrJhcARuriDzDOLllrZ1+ccw9SJY/s1hKUnVLukgrhJu
vJyw1HW8W/23JEXPcR8Mn8ysN6Mxooq8HT5e23NLfZcqvgsDisgOQsWmMWS3AuIv
om5WLg98wxm/Rpp0d0UZ6LBB6yWKFPVCHToLX3gdUnhd1U8Gh19J3TTcGsefbbio
EiqZTOAztBB3dDRDc40c9f4iGs9DhpcmoBJs+g4JszANL0jgd8OEVcCK+DreNkBM
3aheMJOHRBw/cW3HTzFtkJahrC686IoZqWntAXNtC9LKEXxUdULbqvcWSRM6x2sE
35eN9DWKV3ifV5ZQGU4DTgbcQiAr/TCTG2Bc0RJcuCsS9k2ehji/Bd9NQu/WgVLD
hG4C/ZMSmCm3h+MWhvf6h58tM3Jmf/B171oOwILrhMne4/P85OEKY2HA6CskFdO8
OkWUfXAXka91D+1axJvrfGiXeQz1cUNkunwj4/U9S4UFi72qP54Fc0WPzphhsLks
TLSRC1Ht1fGLw2Z26MtZd+LQUZ6lHkFEBXs3oVk7ekbZvW6j6U1aPcy2Mp2KWkxV
9Tvf3ajroJ18x3vDAUz5+zT/sSqKJaODzl1fofCLNhcCTX8c9mxvqxbjpkyDBxcS
PdnIuA5aPfh3jNYXvsU2MOC0KnuLXIVaBLHbXaCLF+Hq2BMVPDbs2AqXu40412MK
M4v0wwBaEfEhjIHoZoshu+VUkMeTMryHQa3MMGhXCj7BTDceVDceidk6sbBwSDjj
tr9JHt5dE8yVtQ+yziPrW/CqY3BJzXXzKXxJtbzdP7MYh9uS20CrSTUrt9u+wXpO
FzCPmEF6XVgk4FHNhTEwT7qsPwNtJ4NaqJnK3TrtMFM4JYWcvwiaEosR1qMTrvwD
EzKSAOJSM8l9zaQp2e6QDR96mck9IPZlyhxmzsS79jHdU+rfFSVs/cqwY4WXts38
HVG+BrJApqC3Hrv9yiGRFDqqMPFOJDzmejeRwpfgHnKcySMhgaYMTen1AXkElFJL
yBHSHpodKNbH3bGcP7MnCyzUg/Nrz5vN9Hoy0RrSsDsFNodPmPFZ40ke4l83QCj1
ie3BWzpcSWUtde76QdJ1Zcd+5877NpTyHSvOM40eddo3mbT+v8tPL0zyfS0TdQ8L
HWsFKWVt7lTRUaeBxjo9hJHxIotfA/eWhml/hunxeJdqNAOw7LOCI4TgzmyaeR2C
GG9HYNHPo3LayB7eidTWxKIf4Po/oSDLCwUXKRBmj0ZJuLFNQo4JaJ9wv9uyOqTh
9xTFDiC/sRo/K10jqZeqMLVjEofeK1KGQCtdIFiAaZiSZCK9aV66uaFiB+mbYJr+
qSIZmHrXLNyi3VSVmrjn6DXeXSesfd5sB09JTG8iCYGCUSzmE0y9y6cKuE8S8Mxm
OtxJlvqfSujshMGs20P3GkvC97umnhHGKrSmGXy3ijEJZERiDzJyrlhiNzxlcGhm
zwrFAzjVqS9onn1v/eaZ9MZc7JbNjytwIN7hcWkAm1D5vU6zlcQF5x1/WTY41PXj
xjROIXvS50Cbe0ro5SQbnkU6tm3DZV8Qgg1aKl8LdCFU3YjxUjknWX2m0ZFdO2Oq
c/UWp723Ji4eO8xsz/4fV9YTYvJwlGYFCn1N81g7id8jkyphIbdsaHOCvRXp1r1B
0mB0YCEXlYBeJ9orEpKsSMR/9ss95kebu/phV2KoBjmJE2VrfkHBpuyltV7ToRMV
H73AROG+8b7dBxURGgwn2S8BskRn7WNGBTFjdihf3YYw9fxjnn5D+10/MV0OkMHb
98ROxSYwA8vzlSLBzv6T98cIOvmbLlQZjVkFwqXypFDzaJ65n9BxdqTNOIuLIwg5
PCWUn00xf7e2D1IoZLDnB+8LqzAS5grsuEjN8q2+FA4zhRD2CE2OE80Bt70IdC3M
gKxQn5opHCnNDi/TpJYBRJ+Y6sgCSt8B7z+Ip7WF1MeZXmejfoiwXj2stsQFD8z1
xQDtEAnKVaOZ1XcPbQA8UQgQI+np7+6v53RyBOnSdYv9S1GnNwd0IV2mpTFz0sRQ
QCEOWOLOVAJSKGvHg1zX7qHojaqKTRQwXIFCEpHdOElQR1MhxKgL7G6VyG4YOv9o
upvli+2tR8TfrMDIs0h8BQOSE4lhfvlOs0jiRXtAJZcBprolmkzV3rquTHfHDhUN
K1sXGRTLA51nHQ1gUgPoW2E7y3y1QHGPoQvniMTojacQZQr63q5bKfFYR98yVoWs
XxyMizSJNc5HtdpkrFgOcMkhoyweWzNlXcWQga0YNmb/87A2CIxPZpOTG0DicuA7
gYzV3eQK2y8sIqEvn6Ml9YPNcYM3EU0nC0DuREaucly9Whqb7FfpLT4duMtVsUSy
YBjijBb5v8lLgKBuYahOVh4AkoBWnWp854tmZqjKl3zKl8aLK/PbuzKznJ+gkvYQ
kzEKTUx1YBeqSZeQt3wx4WmPxSJRBdv92AYl44g2MPQ2S/I4Ubt/+50fedItv/A7
5tA7t5W6m2nv7PfHHKIAY0TLRyej5Ew4xNNO3xO47QfqiVpBx7Vv564TpPWNDFf5
xOQYVslRqOOY/tUqP5bno48g5ShEdlkwYMuyP839nXMFqXOxlUBdpInPhB2y/zyh
08+oAnfPQYOyut+jwgqjfHIn8ttSch/rL7uuo9O5T/C9wqPLl59Qi3UNmPWqSdug
E1+pszgnxVim41JbVZ/dzw2uvkGoooVf+S0BV/7HzhTpqmkG2b1/yhdLL+G2qCp0
IOL32fEMs+8eGIEJtE5MLfwzrwBWvPv/RBt9UFWgUh3+nAoWlSeK813EhRKW7+y0
P+neJiah0wIJRPOPRxKXAchbQL/RvO+GjK3Zmto+EQky58RA5ssGAKKjDHNIjpko
Y7A84PiJt2IGjG2aqtV9t6td2t21xJ/tamC0BtAZUJo7RokLhNPh/yFh5oj7zHlp
LjvKyrW60dkDlRX9VHoqb4QDs0xcjfSuI/1cTu+aemzq7avVO8KzFti4mVABuRjM
Wpmyr87K7HenG2Xt8LcbEVx8tsnU7cUinDJhzm0cd1PCoLJiYed6TwNbgoNNWn2i
cSym54915XMNe52HeN/mG3MKBjUNmZyZuH8mxae+pSqE30UYZSl81CdB0q/6YWJ0
Ui+AL/sH607QvxqG7QkF473tG8oECzGY44i8UCSCR1jGoPBUiDajd/Lle1NQbjY5
FVXClYkNits8lR+NroRccDHfcXJ4nXklMI+4wqPGqTRp418z7jaGQKad1z82SevH
c0oIyXsExjiANgHNh8y6OofY2Bz/K3AcI+aWu5Wjd3hUuSPT1qHfV0b+T/i87JCy
03HA6WRZE4g583apU7m6lGDYWC9W/xX9mWcZfE/sbpPD3TdTjASD0VRoJ1lF7bDS
adRA4mTwH8uXC33F1Rt/WccdjdqeTRmN9xYB+PHemGTJeIiYlldi5bBGb1Z+XCn9
dLU3h1CcEDi6vHmOuoCY4y1LHFoGNHEWaaOaL8uHk36AdxlNg0RYeZGjW9C7gSdo
GTD56TsvHq7ProuuzgzGnijqR7jeVddJbbhTF9z4I/N1MquyneeXr0K8C2u8DpOZ
YpGEkU94BmGSMUrwSZtzpeIoS9lqZb7DaTi5STsC3c3Iobelrj5VDgDDL+rwBCon
HajWmleh2Jt8UiKu774SwONOtROxSG8VnSz6KpY5RgMBKlrFCoTG60Arhf2aO60I
t89uBucW8auAtCrvjBAo3/PPq9cHP+BXwNZhSTKx/k/2swcGuQhz5QkSAsQo8KAz
UPtkBTrMT+IILkLToUXKspCUFirZs6jEzehCQZTdOIUhVhxqvdcVmIvU2/rVDptu
r5kCywiQFyh8pg/xYQRABeeYArB8IrSsIcTbBQvoHRso1tVL0C0B0WycNrsK0dQj
shPoqYp2yV/c3/3sHqXS9jJZ1nWU9uG1kifd2WedPI9Purp6HgjCIFlYUg1qaqlw
GIRQ8EgNgl9rIUF6NAEguhTjNd5FIv9hDIjgubvWrFDgZeuSAyWMn+4E0XtVOGJj
N8TB+0pRfRz56sooRJcWNwm71mVumc1VtM4ETYA32eujO99NBv/TUMsHfmrbUCVG
WwqGvP2gaUuTV1VWPPZ+P7BxGxl2tAY6gILTN2DTqBwrx4WX+MaljUTMv/adVBYK
LyX1wBchu643L38sj8LC6NbBPdKIJu4TqcugTli61k6bKQCAJAOzaOVLtRaeStdT
WxhzoDUkQeAzOQPABqBwQfw9aiyOyLcQ6ZiOU6cMjEPx6PihcVQhVKF8kR7LSeh9
7WAOrp8wOwDTWKZisY+KxbWXKOAa2viGAQG2+/DmeIDSdoMq6igWBxeCClJFI9NF
RLLL5FZRZXloOM32C2S9S1n8MKd/tNFJcy8uv0AOq1IRzXaEfp3dl6q5oj2qvHMZ
eG/IlTS1o0xdxSnSRAQmjiyPaCTBeyeXVsAXttWX/lAZAwABoCrtzYe3NqssVNm8
2V6XNbLZYbzEufkpYbjcA5l1DV9SgFoIx77QCD+LGBPsuaIAGyHlOuurKoP4jGaL
JfxKWrYMWO7PsQnGSDX5zbW6QwW/H6IceAcBZLozUHvqlgKvir+1WEYAoTRSe65S
dFcwefY3xUFNyW5UbPLY9vCxMRP6JTjaeA3yORZqlG6YYxSA6KFguuX9MPmIowKc
8yUwj+9NNs1txWyf7J6hEWLRG6CPb/fmUtRZ6/GlSnaR9BKM7PqKKY7mh5GxOrpS
ifmy3CmlOcKegdITteH5T1jNta6MJABvJgieU48I2GEVwhm8pfPXDFvtLjcNUw0t
npbsFsJGEEQdtQPYDmKk5jUehEQmGKtWqYIrWM+q/tRyEhFz9++4A2g8XytEkuPK
nauvzaKDmCpqKEp2qFjPK29z6VhVY9WaPklYnYofCtamFig0LZDFNEGGxQdO0037
WCMKlSZlxxUAaQJGRvUXp1C3Fla0tqLnKcSs7QE5GuvONQkzoaE8k4Snrt/zcLSV
1rZvMn1GLOsNSKCDhwjx2HE/ocHRP6gLaIPQhkHS+zYWLdZnmbCRgf4BDIKSsaac
Ie4rKgOhEXnL6xzqeQgA3P3gvfvUd3zPkr5slRUEjs9F8+BOrpqNSs/B6XyFSEEl
1muDcMtCsItHYdYH258CW+508jy4FD3Qe+Bgv1fc4MiGldygZWO8wEDMyPTsRDph
XEqalMv8XktY9akf0XA2MeHZKp6ooqvxNgmApOS6FSHqUIZ7Bq4O5D3qiO3Bh8D0
ctlDM+rY1F2UKxFc+RrTWe7J8gHCuhpQ3ZgJHz4HU0y7SIfHa27ELDMrqGzh/YSq
VKsJa34XYuvTjoBEiUrB3SfY6p324NGsTEsbkSXs8nnhFhJx3uHfRgOSzeg3yqw6
hqvGsXUuuj8FyAQH1uWfzYg1p9CELytuKs53YsaesBQwGzSMgZCWKwyBApVUVTp7
G7SjiFMdRlhQG11e9URBWLVZ31BKp+qbyM7h8SdhbIW1VcBetYI8MZnWPuVEwLZI
PFBb5kWhg3hAen0l8YqXyaG+IYQBEuOAoL6moftqfMYkIm4mCVf7mOSv1WBNr+UJ
UEbOASaP9d6L0qZAX6OBknioUJ0a/fSX2rX+F4dzSerI2BT1xzovs8C3FNI+4KUJ
qapC5jc68AqNkcW338kigB02F3VMLxY/F+Efvtxei6/PxUNT1MHuFBTCcj/Nnzy4
hAdtko1f84DFisvsKGztuJSc5yT2NM8SiQ6wY7tIjHQqMWpqIP6XyR2rGafXbRqP
Kut0a70vlSsvFvhplit4C6DyAGYj+yMIrwQQymBTfSKXWb45P3gH076nS4Cp7y3t
rvTmG1r8zCx0YplYIth1jX8yQBKZbgtQMgzXEv6mY7hPnkTgH1ehyAMzX/navgEQ
pqpZGGlf2YDcm3arI5Y0RfBR7kxjO0Pe23sOj3DV/9pAL2E9sLTRyDTbxeFs0etz
otVUleoAq730RGspwv1TbYZ/N5VfWu9DQTWYxMqpQUfviKCHfz6UwzdDSjjyMwd8
/2I5QAFmGhnMR09gFUoqhhOD5LVMGzZPlv9wGAinFPX+uAgBRm4x4VeN8TgaMWjk
uEyJzuXqwjGZAmBSkckqdAcSxTo/JegKcx/qgN0xY4D//jbJD1EoYoG5Md9yqv9r
w/zSTdI6mBq1mYdq70QRN3cQc33DBC2zXdfJQvbI0leJ+cB29BgD4fF0u3RItd4f
qSgAi84Ow2/koINi/P+jFT865OSRICjcNQcqMEV2o2mBoXLEeESAQBRh4njoM9nh
yYdC6eZlKkucXRFaV6w5yI8AcyxeBUUNFMxX9smIsP9fKmhw0v/NbxAi+gttJIza
2Dorz4UuzHvGqgKL5CLtwvJ57B9iFpCalYbTcOIGJCDD8wkbQ7mWk9YQKbSuhMsj
vchVSjO2ERS3WbsemgvGCTPZMWoBufWXDq+2EOluoJ+4TnzZObHuf0uWNdv3DXUH
PDTqWAL/CJYM+vwfrRs5RGxVcC3G1o+YZ1jEzBgC8tSJCOZqIrnWa1DeIyyPBpN/
ZAyQwRjvmII/byQ82wlGd1mWxU+2AOksQBcHoAxbRmF8mWwrYbC/eF/Pdhp8sHkw
XRTSut8J+3v6sMW5rpxLwsDjE47s9z4CBe5+ldXhjtZIioZxl+qQqJUYJiP9sPY4
jKosZGVeB1ieYhYKfanTYjqzg/vTy+ccPMuXesi+VozA2r2B3HHv+dP/mkj57ief
bKbpFDuDOVCLWfyEpS1CxFS/EvZk89+tpiubJ3AbcISx26fAtkPFnKRLaIzNozMK
fJ4Ys1ZqVtSYFXOoFQu2fucAHav2NB3udUptoFmThGS8cMi3c7eUYzmZ0IiwOK2i
URLzXKZJdAYsKIarJc1/T5j+4jIsL56CMaI2lazcP3JH2JoqIXZSf3MpvP+bBHHf
HYlleHdR0qxmOiHoHPAdBLQe20KV6kNSyZaYAqVEnfdrD4E/9yWRnHcXoaGTrPJA
lqzmzUYa1P7Lmf9eVKNzs+iVf3gfiSWVS5/+paFWwG9aJX+PWWq/gEGGGnDA6Y1G
q/cgEIOTiWM/8mKhMWzr6NNWDY3kdcIXIUC8PjD4RGx62eSsZwO61How+Az9PXfN
cwaXPoKknBpE+mJdtE0NCnZj1pZrxNcGTxgj8wsBdKwHRVpLiqJ3p2UciSvncGte
hKB+w+iS5nF3iQ9PVIRYFwhd14lF87zwiQxwhWZA5UAi6mfPiox57UTZhty4mj6w
adWQTd/Olv0QLgOU/WYYTcsHyX16NCyXA3l4C03jpY7fH+l/uQc8vI0mKBhgWJY6
kCmHPQpquO7+CgTQQT/7FiL6uWz7b9Tb9+EXRdtS3JB4V0yowBnDN9zfymLnO0lz
Tdpu10llnPJpD1U/2FMayPYfXOqm+pPsFnUpoXtJpcvZ3haJlPuRyZ35KZ9PtgoM
Cp2/5iD8kwItgaRN/AIngo+oZhmlydmLVaV7O33cQKVgI7aGzgYVX6xi7cU6MhGj
UEfs29U+tPHAqqlCr78pNrhXaOvBOLe5mOVl8HCqApTfVbv/T9xuwD2KBGCKFB/A
J72NSaTTD0l7nqh3TIEeFn5ZIX0DbQg4Rq72+yg5TXoH1GPpARekKGrpQNejtUrE
4NJzbZi7j/uCgfSMbc8e3O7CbsZe1Q1VsaxmYSFwlBgc6sMSbagKbXgSBWaf9MCC
razxboOqW21KnASWtmGtHmp2rMhdJpheMyRidRUBgOL85EhLDWngZjoaxuaLaVdQ
ektoT2Qzm+8doov52IyxoWeVrzBKiT69+3Ka8AA/hx3KTZF2QFMO+KzksmkgCN4x
iNyY6pG04hrmm5BRazX433BUJlE75tfMTNdVPcAVVwSsmgF8xVZn1lszHym1w2D2
1lKm65d3i5bs3Gba+uj0rO3R7F5cDoGFxADlWC5EebsCHctT2KeBChjQciFUpaN5
TTfp0FwB5/IzJ52CgYsjjJvmw0EByrRMPQng3WHtX/V8kRLF0CEP0Pk8EwCsxf+5
FQ0e/stf0BHEdDv0GEDR4D93iswCNUKjfNCvLShVmzhHoH3xn8mOnA3Zc6+MNSv/
L++N7ItYn2NuatT6qX/MArjWm2+k9Z9Q5Cjg8HRjyhUgwPpRxHKxO0QNeEHY88n3
6gxLMoLT7QMxFC8Sv+PvRSdEyOZkoVczhtZriUFkNsj1AELd7fUu14tOihmY5h5k
RG+155Rv88SmbQUVzfPZ7aRvwOzq18KkhLgjHtQ2VSukgJ7bUSwqLsdgKuCAo9h+
Oe6kHXEWWpUhcIxLJvtjAg9LVoGsscT67kMzw/6q8KX2Ce3trInDCiwI8bkQkQ8u
/P//pwR/R9M4/z6D9k2LzM+4w5lnu2KOEKEeIb7q+jcgf0iIkTfxTlj9gfxBYXqX
ydKLFg9Ny2esyYImhVfui1nuRIpXju4Y19KiII5/dBN/RMA8nF4DPWSktp33T0xI
x3DQsyFezNSfVUJaIzYhcTAA/NLZKx1gncQC6g6AMpXnoJiZhkA/0WHZbd5MmefV
mTrSAJJItSXITYaYIgLSDiQBxAIyRHF9n/rGUgYvXqZ53CLc7mfplRJBeFfN50lD
6J2SsMr5h/c95nLluJVqMxihhyS+YQNmndsvUeRJBr9cvsslPHO0becW2aiN23Yb
Wz0DLAQCEiaPrniBsb1F4HQDqKH8sLadqFPCUJa+gHQJCoySOpFJpY/RV5vn5a3d
dPJVfo/B/dAvnPWrT1yTZJDOVD4vhUX6SEkx22xLrDTKpA58cO3xs5Ikz6iJwcgE
Xc5WSlKkoXH9fOiM7nlhlUk1cLid3l+mnIUtq9SRm5uukJJDxkc5wQJG3IX+2KEq
8aN6iGC1rVfGhjMXM0MhcV55djWQ4WwD+Cwnu3otG3Qq+IKlV0RohFFdLMP3Ka+8
O2jsoUWKYusMIr+DMpUTKFEkJfylQiYR5iULcjAV4f88yScEcTR7KTWleRL6YxPD
Qo/GWiaNJDuGInLshzlHE49l9OYJ3TQ6yj0AKjqm9SySaUh/DUWug/aL8Cngo+qk
AQBiE1y3mNqnUfvqJs+t4TmKHxsUDECFTpuQaKHvQbSkMx1THDmNKYui7BscgekZ
8hm3eQe+rEGj6jQsvdBEg+e3m9imSi/dBE/hpbCuyosukcw+vvSsFcA87tzuF9mO
PFEMcJba+DzqAAqYr6EJmb9lhsPgwLnZyLpZRC6xsPl72MRGAyFIGcKl8zMhKlfZ
jQamuw6pP13I+9y1+KIf+3DW+eIw9ouIjkuQKKcZhrrkZlU3bqQzUqLo9D3B/7qe
UEN93NZQh3mSzAs84hHX+4Fb0oDndjoo+/LuHiFzYy5pvbgz995GtVwwil809XxG
afnjbWwoG4a1etsUzgwsFWGNu4aXVI2f/Tr3Yr04iEYSH58vwT/hUiVoGgDG/jCg
betDB1FDSCmxtM7ORBWInzY4lX2mYUbf0OEpYfoXQP+ATCOlg3mTA5f70dBLw56E
pr5GRgr9xblB30WHmlAHHoykL7ZxjyVyevi3gUNqEPPrgjo9mLuWG9HWBcvjKtyP
IZj2mBa2zId6hfh4xJWJqQf4l8xkaL5TwbPhT2R9EfLtVDHghK3oMEGL8tmyv9BJ
JIpN26lw8Y3jCKlnabd3WZyLcxXq8BoCw949ieswAUVM6QkqteVvVEtnxF6hZJo/
MraEHI2eiTP4AgRTHEGBNLu8zyKtiHOvrajNW0WrkSFM11nODmLcY9YCDeES1i6x
27kDdUiOardBi+UF2J5knaT1cx4qMApseYACSTAC0R6kS9SgTSv0oOzxLIdiDPfF
zWcC7Oe3S21gxR4vjeFg2AEYRX7hMACMTUEcUe1pdzQ8gmekOTbfMvoqbaYH7WkJ
Yfv2HU7+y/ZFg9VmWtoKE1MI2AXleo0uJCOAi+6aVvfGtzLVidHwlYWwfEdqy84Z
E8QXE0HcGDT6TzpS4fKUVpLkjSW+oE3jpHl6g0XF/c4CVZX6fNBYoSi1puPO4foY
AvnScFi9JQfHhz6j0VP1UiKlrbSiw9GtIm5CPS8mYgLGDQ4WEPSN6fO6YdxhmWpk
mwSTej6xnW/gB4F2tk2jfH6mxEVlqHG8uH5t/GsPI16sfEypwYXvUPaqC5GsxiZu
fZmkBnorJRaQciF8BF9305Fi0BagwBd3VHvvT4DeRIG7HtGSHI2ckpy6eYv5c/9d
NCuHGa0Cat3VAgBmbqbzpKvpr5SkAGN1bytL2+zxG5IKnzoTPxztWQgrpjCcET/Y
h1UaPCEkKQtFPesG4UZbpaF07fDR8U7dibakLcP4Hrh7gBaR2JARC+mKhkM4oVt+
i7Ijl3ztDepuYF3Wr1dWfVu6P3gwrHbUDYJznAdrdwDyNPmWRAED8MjvRY0CKwj6
PmmlZ+cnSxmTx5Gi24epLVZraBI8LkNrf1tkNFbHqvwNra7xl5/fuspsJKxC1je+
qh44dGJOUGFlpsnVNvWKHhdOTavPV/9RB/hnoKy3sIRQqrUgzROKciNmYBKif+fl
V1moi6iY2q8qrGdmNGfSqMZRyYaSdZg1uCA6x+0WUTLHXsCVtg4YhdEy/SfKmMBR
CaUEC6Pj1Nq4d3rRdyJtI5/Tkat2U23VgEsTmcktMrRIi4z/khbqacElw7G8V5uv
9MWvdsMXq7iSQRefKDbYGFrqL5/NQcEVDsVGnp9SIY+uKTfOeiPosM4zk8AqM4Nl
/aM7tnxuFNKv32mfAxEca11c+7mUygOWlLNEFY+cLUVDSx0KmGlPd53MlzR66Ef4
BW/QUXI7j56St1GxGnjeArPgOdOSNRQpwRGoiJbaVP1pnDsa1To65+BHi6CQnAM+
aQtff8i0eiXI67HZEcSJ/p9zOt7JB4Ln6hZAQa4Cq8JHI+zXe8xzIB4ZoMlQjUhs
GpRhD3T7xU52pI8IpNECRh2HyZk0OSd716ka/5LwW8bJTWwtps69tyahnuO7l7sh
sJL/ucXMeMzfa/P6DJtr2w7p223JwXsAaY+brcEIhXOpoo7tB+8y1lilhqDZupti
euxv93oZPmLHVj9iApMXT8YPR3RAhaz+9tZ80/uR6d2wP+o8wAC/YbPuM9FvXrSd
D9J5g5TZgfnMUPZBQ1f4j/bX1HOTbQM7ug+gO3VAuydzAeRf8mEo20z6SCLq39eL
Z5Z/OGj+4qh25HzUuwIfHkS1wA9eIXRi69POVivEcLMDu9mKRpjKFwFjbyk9U0rd
QjXPjmVXxGRCA6M1/3posk8ucfVm7xRUeDjZ/Y9oF0v8vi/KkifPD8px87xQq47w
/VHWnjrswfHB63flAilSTduEWP+msMO1/ki1sPNg+onT2xdHO8NpWOhuONx5knMy
jp/hM2w2sr/es8KjStnRHb92rkYTHo0HQ+MjlyHGxyCP3YGYd35jqJPqGY5oxyJv
9JuBY37Mq2i9wj16dvz3dexXzk4psUazyUbfvj+uU3g54KS0qnyBd4xf3My+pW0N
knk2YCZ3bTzbeT0UuK+QNqVTYA7/repWbXE9JcXIa2/V7l/UduS7UqyetAB7CuNy
ciu34iphsB5T6Go6bBs3RLvUCorE5RhykRRe8SIhLh0qGM72iOycodqNt+qktomj
iU1FiECahZYRHST8eawlIy9ZF57wUeBAxgBHfc4T0VYmGkB7bk94Z6HDQdgb5wsW
ur/ClULrduiNcXRDivE18gozFMVNmYFn+qNtx/nxHRDdfsc9AGJF7VpLlgbhNH8Y
0B1LSSWVJNPCGKVooJYwF6Usvn2BVDLxrUMghYTyfL/irPMBIMWWMvVcl+tyQ4sU
1OohwITCpYDcJOMgnrBfBdMmbGff2oNQZYs4o+FUsUjAsTZ6hmuIqEkNsx5rlDlY
fRHwBtljWwlBhGMifduXeN9qWelBslm45fbZf5sgulrHs080TSRXa68z/CZwNrpD
eQTGo8L8aBlGjJ8G8S2mRiZ48BTwxE6HwAdDJEpj4yQ8KBJ5GuerKseYHzuVcK2S
uqbjyrKQ1xS+udpW4uUAvRWD0Y8NgpjabQvp269O2jJPFAj6V94ioZZ3qRV5zZT3
0aEy3rIdFh348BsaHzpWzAJHPVV4vF0TygFv+/2Z/77EVJbVOvgGNKtEtJX4O4+4
lwpru0AXIqdGVjNeUQC2wpsac3dpO/eK5VC3SR8qQ/uDMUnvgvG6wXH3Du9Scm+P
6LJ/d0pZioj66vEVOATi5BaWmwmH3KUARUd+lK/sse+xmAdduZqO6Fh2MqD34ys0
KsvmxQEZmLbMClImp2bEqmjnEl2R4mrNK7s4R5YBnQiWvQ3cElM3cRPLMzPntfdu
L6EN0NcxX2NFBkgRCxDwUmtkKuSQqRm2ckD7gTuRF3V/navo62y+QBLA+YERXTdJ
m+QRlcliTVFTBbKZ3bdAsNzGTszIZCHD2FL2hW7wM1GsNCjjXM25kg7SDbI0HpO+
TPO785S5CRfIzua/IkBuVu7XxKLLeXYtRBe6J2EYJs1Sxxjj0s8h4BL6KMCYKH7v
7GSGkUS3/w/7EnaePSXiymkI70zdqGMiK2R5KwAULzq7it+zdCRYWV4qq8sPh6mt
chYNc6clb0rBcobqO3vWWrrPO3dy/f6DddvfOnvwdGUbQsaxk9Hv4NQP18TH2xdc
7vfvyOR4TtIHnjDdB/jeTFxBMAjPA7qk4MBQWJi2ryWewMByf0ZIx04BAWBv09OE
40JGLpqkFDNNMlP1nY+RFr60nD/KERfBEx3ijAnzS1dASCL/8N4XPRxlX3yM81bG
msBHc/QkIAYIyl7qN3qn5pp3la2dpOXoLyKkSVZaaUbkhV/asmSq0Zfqto6GmwsI
TQiDkyXLHevIYYknRYy1hJ75zU3++68FSr5A0sJt/HwZKcIytGSN6zuE9xKrB1Z5
fCJB8aB+qUxiK4RURSKoXJkiBfRtKXwMx3xR/6duGQRQtfXbV7qWgU8ILlm9Xk5x
thmxXflh6+loSOdqubA/30RpoemvYWgnZGYJtnzFo8Yu9VMklMC3znzVLkUJAyt8
zWUZVLy5NKeJ+Bh3jQQ6QPCdWMVKx2mRn2uLYj5VD7evG45m4JoulEniwoyZV7zD
hZTnfZ4J1YERFIAQHqFE76VNYwjOC20a5RLo5u8/CA+Pf2FxN/inswV81hpVReFN
gACcIiYWLxDVgEW4mwgeP7Tmy52BbjZCBwDlvszF4xOAXcqO7yq9lGpNLoeIEfoZ
2FZ9u1e3QKf9rfYliUWZADV4vFNkWfbfiXEDfRAxSTB1QdpjlqaTlSTyekEIZ/xR
unRVlJhrV7vdVCrIlilNR85DyNA+DWGI3SLgxcauCVFpOmD7dypKJYk+7JRbJ0dL
cWvh+FTjpew8Pp1oBOpNpEtYnTV3bt9HZYAC44B09eA5U4QSx14sYd8jPW9Z63a3
qh0hL5aafXey54AZ+Bff95pgO+AIdtCJs8lcPAo6CEKuTPUQFqn1Nc4sBYtIN1ot
Hj+pN7w02A+d6a6RtvyGnS+lQCB6WYcOov/FSVbQzo+6xoLPibdQEEZBiyFd9jZ6
jgcWOFlZF1Pa2D6vNoFq8UtT4tXxmjqs39b1GsBqflmPHweQlnNn15jFRNtM860/
nf3hoHOSunf02DpbO2xJ61RymunBRSKZfeLzI9p5Q3ljQVO0iwNw9zfBdi4ay411
0PHlPxD/ohCQd3qZ5JKB8bGbVJJRhDLzDWshmvOIMKUAj6GHKxNMldCO1EjBG3Sa
QhXqvHfPpV4MkAa2BPnbnSQP2CsgBxGlLU4BL7Luvza4Vydm/t0pSi4h5oOPVisr
ug5Ip5NgOvxDcfo1/mi0Wvg4XkHQ1ZkyHymIdB+AzhJegGFRvamNZtLNI2dc6gqR
gHQBkX0+RZaEFydJ91nhXEuoVF/fi4KuGJhZL4Rufe2J13P3LbchZbOB0JQGr1VM
UwxL5yqN5FE3DWfGvxGo94lxSly+7Czz0AwtgnCdhx9X1jIJXio8SKizFXDWJsTK
32hAPAs4NFF8Nv/Jmvz1n6c1MqrMpNQrYO4I80zQqxiaYGiCBI9xLJh++Di4xTHR
HL7y8E+Lhk+3H7mDlCwtKbOT1Ru+XQMY/gpu1+okS0ZfC1np9KF21ZrhwhswLerT
QutDn++l8WRNg3l5AtzRv3ndeAcu1EoMdY1WwswSWPq1UyE6xNuzOoTmw7J971zg
ObVw0VKX9CNfOn2r17XIBiGOOjzno+nMznIhHa3gj1aOIR3nmf8JE4JfXsWGhQ7D
xWRNJG6QAG4odEGxCoKVYq0Nv8VccsYHeAl8QbEqTsB05PVc2vAZkL2AI4T8IF9z
kWU4nggVHiJe0bGs/0COicD8K6yKKIYEbfcy3Uvm6wEK1sNuYKPorGlbyM7pZ3g/
Ji/pIHXY5vum2aYK8V7RbaiSDdXWxhplI6M5zZA/lOLfkCi4av00dUX1aOzNBkza
kVxwnGOIO+VN07TBmpSdrRxSmklU23tsHlvW9TMIR3JDj5V9J2KWZgqq1TUoZcU0
pckoU3bVvSzuOIihzOc1j4U06Bqj9AY5170M7fKq9q2wYy8NrOqe3eW6B6f6WNAx
VBdIv8pZ2tjuD0vc/CxnFf/90WT9WVTrs/e/AUNs4IP3Hss2EhyL+rD8VCctK4vg
hOBzFHkYdlIIEZgijnw0DRa3P8JhI6HoPJEK3WtioW7kfFsk5xVyjmEdUqVWXQio
WUAKhe9ASyQHBrlQFivPDeR+Fg2pv7Worc6NhjVp2hftOTRK99jk0ul1T0vXKZmt
igTYWYeMy3DurPkCuLCQSYNUfX8N4ayV5gzPOPj+I9xm+cSRLLiJEbFu91E9baUR
Qi/K5P/BRdO1d+HpWpAwQUxj0N9q50ZjngSvApPqP54t+9MpRKDQp8Ga84L7pzmZ
93C0QXykeuVB4WXAwd+WyrAmXiJD080tcttyVlmCIzSkbFFl5skCacizCQ1cF1cf
iy4/RSistJdWl/0LcdebGzz2t8Agub1jbZRx6aN0RQiX9izwSchqMAHN6VvICSMR
eXvLcgo+vm+RW2MBPIhNf96yzk0909h1B2Ynm3J/kdmSdF1gLuWWBm8t4n6WmtJU
3BZNLFEw8SUAmmZtkeNXJ6zct5Rimz2M2/lNawuX6AaOiHlMrJO11GLFtpkIyYhl
ihaU3Yu0drbECrBRDv8aomMMFy3ccrk2+aY1MNNkaDvBGIsUVMfbTGzYd//jB7v/
HNcxdwvFK7Xb8Z87yzq+p1WV4IhuBcFODGTa5teUBd9Y4cEAyUVwWwj1hQgAAMMZ
NaGru8Plv5L2BBQxiFlYdoS0Kv/iPuBfR5bYAq6L3ezaVJ7hEG/0zpNUr7sA2/5F
wVHhcGTetfQnPUWFMtm3Et0HlZTcW+PhlUbXP196YyF5oE0V4FAJN3Nm3P1I0jWL
4waNXwDRKxjoMQ6bH8hqH48PjDevg0F9mqjDm7mZ8wfSlsg1P470+nmYaLy/1y+y
pDRlU/s/PiuaeJW4w+bypTMPGT1uDZvGvljbr9iYmDtTqwe83Wm11znbAD59tzv/
dCvMlp45uKQrNL0y3ORtStmuH6RfhAtmNrEw7XtQl01crnmxo1AqSaA1X3JvsKZK
ZKYPH3uRmeGdz4otzdNqaNZSxAbTFQVMdah8D1aefntG2FdeR6dGihkPdSWdmWJB
i0PscKyMtwZvr87Jr+50mpvWWBZz4ujuTpBZENqp8Ly6d+CZV8pFv4eayvjfOWWo
KrtxUw5dsVDIWjNDWOtJMsHEItC1vUXZVdY+TuayNOwVidT9IhbDQD7iNf4JLx2i
9vq3cEepGEM5zDA93AJrjCfnK6SLHXEgmpUt1rhVVnqMks1ZdkDzp6OHdm/iSKil
Fs15suF1JzbWfhHUofmORcDdvQJclPfy7D0JsZ/erwWv1vD30iESC44PRY/Gc0KD
URJs1Ml1x354piZ7oSSuUyOt5K6OvsBEHLF6SbLdz5HT98XSJHv1Ck/lppspv3vK
Utmw5V9soRFKQzPoyJ6WAZBAIEG9vHP9qsz3Ts0pGmJ89IcslfAtppg/exHk623H
jxsbVS9u7dOpVNEzSHGBy6TO2hEeubcOpuilWOtcXGF/glnvSK8ub6rWgnLtNAzz
09DA9s0qT0VXBDLx9xGp/Sg71H4xobZExylBtUfu09MDQaeBqYzOhVcaAjmcStCg
mVB5Lv0rsOWcjz0mfHZh6FEZlJ+QvMj6JVRmZRLhG9wK0EZXPicXB6g12c9ocrq5
M8ZDUb1eKzpvaotf3JE8Bo26kHzlnU9rnrn09uaX8NPf/ZhozXbaI5P3kRglo0UL
yXPRkyySjNJsE32v1D+SQ0A4A5bBHMPqF0JdeusZaM5z3TUHpFmMq/22ZtnzNmd5
lFLEvwgTxQflg1m9OBpDjGvXsPlWmXnqAm6hnesQsSe0KEmEpGOfRd5EWKzuHfni
nytWLxdnmWtkDjjQkc2vzgvxxqyBh0Qb0aH2ArIM/tY1Jb96qGx4fd1KwwSSt3cV
iJRux/kXNlxiEMCUFt1CrRd0PLfUjNLFJr2Wc7XjBJr4OGwApjm+HJydi189KHf8
uzJna3w37xPf8UkQjznTYuGe49tkPITCygC5OYlBuziRV6ERpm+JpSX9lMnM5Ki7
7yaDGfEramhnVz20foK5mBXMGs1w4BOHo5WgMiRx1N7VQL2Yyqk8WWTqqJScxt/h
p7TaONeTKDwWjG1Qw4d7aUAgC+XMFO6FIMJQQsA1QWOTP2vALsRT0rI8fwFfn1NV
OibtJ8NA6ax7hZrMLr+JUJQDJNtybLkZTFLv+bWU1ZaQjJ9msQN1UeDYOzmU4Ouh
RxttnyJnni4ykBlG+YikJdE8XJSrAoBDdHP+BYzVgaDGhneDBbYUj52rgCKPNzWc
pocwoQM0iPuLTJb4tyjnlb5plOplJBMfcclZHOsZTBJA0I1E+a+yiHPOy7g0pECZ
71oNZp5Y17/pOLlG+367m6I/JArEufRdBsZhOTFaO4YlW1ZKe4zW6o9vCcwJm2ZI
CEOhWOU7nh/Nj9PRUF7l9Di/GvuWT5rVsE0NssE/KEKnZmcF7cbi1IWATB5jhGLV
GWMp1iIjjSOy2BKooDRoOMNINqq48p78lzUHVEFJTdIHSsGeoIiO8DFr2F+AUf0y
6ciJPXmbxgzZcr+LY7rHOu7cc+3dsu0Q7p4ILfShAHQRbpAJdbpIl6UsnkLpOg34
GXiPFrRMwQhWDVxlRfHQ56fxJx8yCbAsCzJgRZaLY6tK6VHPgHLI5/ZNjSxsDD8c
+zVOR8F91zqSd1Oigkcmuto7v8APUm4v5E/Vv7qKtKPxUFEWk3B6ynBdrdbt4Q1X
iWF3QNc0/ZpQ48ABkI3UVf64MZwqqENnW1dNkcyMZmRf2apa+iYn7Pkek7fllsN4
zJw6y9XaT0bEC6h02B93GpdWHhodMXOOGNq39IO+7RsV+4tlaxAqGn6z9531FQNl
O/DMAtxYJ+8jgfIf1OAelXPRVqWobB2Q0utQxkf/r67NW9RMYdghoejRrAH5CJIo
V0mH9kakvRdxR/Nf8yGmfcF7VSpJVWkJm66FVUrdpOJ3MuLMXE3PHR6mA8ereO4N
l8wtN+uLj6OtaAi2f1IwMUsuYZdhwm8wwrLZUD+ov1ZZOy6G0mY2P3hgDI4/OKgq
xqTt03yomjfOY5eYhdZU4LOZ3YlEq+eYpfCedemWBpHziABeudsB1drrpljBuKI6
d5NmRrcQopcJU73SnQp6Sfk/W4/H29/J7miWIusF1pcdyntWI/cnhgtuDcv/Tk0q
35Tps0S07IokYmYhCiDgImaOo+dVvkacBnQ7bkRGU+fMsgfCn/cX/JkAR74tlOEl
sVGBhkbAQ4d2Ubs9WQaOdHSiKTnTLlMXwPqFt3iUj55mUHf1kDxsZ/HnybMA9SjL
cPSvzHA6UllkSPDkzj0Mh72kQtTNajwAST9R80C6wMmzro6La5VINhS+FU/38H+j
S4oYcPmiEWUSPGRU9AGllqKHLYo+fql0k1Zfst1Jqku6D3e5jfu+G+vnKTkjlIGK
+ZKTlLDK+9/oLlVovACI7LYtvwi57IcX+CQm8y6fZ4WyjMA3YYjcmGWYCtKtsGNP
x7cRXPtBljp65b0oJPvbdLYxTFV63Re74HHZK+rwrMabD07S7lugL/BtJp3QcCp6
yipuNn9kVWHpnJqnp+J6DLWbE2uZnyO7ObuwGMt5PHQpRemzG41tzX3zNpxCLYTY
BL53ihGrFNtnFGE11m1sT59f4fyhup+f6NwTZWyAtzTJURKpOF7GbP/M787QoJPK
SYbHb2WDjPjRkev9PwYDV+qj/8qVZ/rz9bUcCDhcfwPAOA2SM6zq8jr7GRIYf7XI
+sAzqAEbPG2WEXr+B3I23wMh300jdshH4bP89rw8YY6SpThNeB8gO1vLR2Ei76zv
VZjklDU7CsJpmxDoXzvyqKIBTjHTzXhKSM0xH1UdT7uRfBO1JTon317zVkoOybRE
Kx3jG+OQ4u7cq7lJUDAhqKM9fC3KSVjEqSPkWj3Xu7LGYLpvluatU9vi5a7R4G9I
C/IIWc31Vh/l5RDoFq7SauyU7KGW2bkGI2TBNbjOtBUoYPgzXN4HpQytH9WllHRe
3LLkvRYMQMZS2Yeeffu61Ip6Nc6cQDqJ9+ejJevZefDoghA2vB/zn+Z+qj7kvcfP
aCVtjYcf6LbBNVfXu9PH4pqpJ3IbN7NKWjn5m2nQXGnWjSmhEaslTADbzfEce1+Z
vyiN9+XutI8J+n1xUT3tlD9VfiHPkgvGBKlyJEyYdDsgdfgKFeGsMlBtszpyqpCe
uKPD8W+HPLQ9ckNcuSXKYQtCPeuoXRWX40V6lBZvvu8TY5W0np/YeL9r4ro+zoAo
PtppM2qcSVV4KbETXUrUl5P5tDYquQGWjNVxnWDBGHJgUX29Ta4sGC6f6pdkAMGk
ruaBzZ6UOxwEcEFiBzPHd9cfXx4eMs27PmPpEGMfAmHOW1lavTEWgme7fPi/zkQx
yY48BAylDBB+oXTFCzzSrFf0Skg4eFk3tH2n3J2f83sxszt2n9W4WYLJIlGSFOUT
LHmP5XEK5P5aR0Y4HYc/78gNRN3JbcyVxalueoiNcShSkdvy5BOlQRRT32urtA4o
oqXUynFZH/6VqEcQHHl+kzIuXdUAcLhjvKzeQOM+KosYKzSEtEuBmwngW0gGG8E1
XyMVPoO9T4K3S32rUsE9LZuadH6/7crKur81IF2uQ1LTNEg4AKF5NmcXpMXB/4Ui
8GQNTTQDUVKSdZxEp/rClHQamdl0HfcR1BfU+HGsk8xDUfhTY1bd5bCtIeJHxUkH
QyS6cg5fdGdHipJvxTcnW/yzOqIq3X9KAdHt1gHoZku1IukavyG4Bs156nsl2wF1
lLeUL+ITRd3cFh2YoEMDLp81VRBt1YIg9tRAlQYR7eNTM2g9iAZP8epxTGfCx6hr
EeViPiL0nnqCr/5oo3R/FMntIMdfXroYCD9PsY2NfcJcdixtlmjQus/5UDV/YP9K
cJ+7XchXjv5jI1b/dYInNlZcPJjIKAvYXzowHHPL0XmndXCcRPojyMC26zu0T/Kn
CDmYEzpBLLnNhX8Rq7tPm3YsIxOMCKvMNeFJvrVTsy6hRXRibbITOKKUg2xJrrP3
rKjTWZx9rz0+4fRJ8WT5YN5Votmkngq+Fzw0/UIibmuyIvDD9f0nVOpQKBGtmVI7
KHeWPswdmyFKKRPQik4C6zhwU7Ce92r+QemVbd3c/i/BajEqUKdBSqCozC1XNaxr
pc3Qxmk+sLJzBeEXxpL2TiTnYdA8opQFIEA885NGH8KShHyDbVybNfXi/aAh1Q40
kE0T5sY6+9DeWm2wtM/ccdTe8lTE03t2Hpgta7D/wYimcgxg6OYdeQggHVC9Acw5
d6uXb6uCDCgqqP8etEzM/QlKJMYjVFskOQWzTqvE1EGcHz7KZ1FyyQiCkUtif/nG
mlzRVtmcY5QLTxlgaG0EWypm0SOYrsq9OBgYG1jMuE5tTExKswJAglHy/Yf6OXts
bgNqgPwc/6fVzCgIkhYhu4l4IymLqbboVq6Dy89vACS5gtKMKJG36kh13ELn9xBd
ns3Qa0kgUoosM94BD3D/S9jNS25wTaBky4EG9pEAJsoG1qxpXimJH9J5JkkfbtxQ
nlMivZjM55CL4amocg8e1fsPxyCKhHDe6udRJ+c8KoSFtRgl/9Y19GqGAzAGqCY2
hwR1x6cScInnAmFz47Ja0+KKamsAAFZQcQ/ObJWYhzBKVTCg9LxFrz9MTSIFpZ8p
n2Jm4nDQ8u/Pxs9PgQEcJ4fWf4ga6s6isuLcep+bZCJEJJuZV1kTUn4cGhNeYB9r
Ra+07j8vW6lu/ROl00HM7BaJkDt6pCHVTWCo/3wYExL978cTpIyvVIqbfU1sVBzO
PDo3b7GN67nlniNQZe5G2G3w8VBnkNA/VB5cVPclB3CXuxsmjryD83C7gNsB50Wr
NJQdGvom4h5fday3SnUOfhwyYA47vELriFJ6mzelg78cBKATybn8ozgc5F/+F8gH
64SKyiiL7lEkhO2sGnJ38UBPITVp4EwZ9PZ6IJlxR1iO/8SLpvgJ08Dh89bY8yJh
8z7wvSf5KYS6bQURiviMc+t0MVCS9ssJT2b9cBSxPVDOHRF8TgnYHCwiQ1QgQgZy
MznY0Uy72BdKK55zPKBU5afFCXKekQaObvRaxarQQrSXIbKARxASiJzmLKqNwTlx
9oSouewq/H9yN44W69oYvaOHSItHwvMXJgSwxqtaUybEEkVWW3hkumeA6xQi3w+n
yt3iTsjAEMHmjkwxCmm82XN6/OkAxAHzz7e+ldZoTDK6gPeMQ4YFnjL20gi3ke+s
RiDgia6ulTGclCfJeXLncdX8DxS6FiAO7ThxH0vFUCqLw/EKjViElOWg0ybBuLSa
NAOXVt78k6EKMA+wILXrEJ5IDj4cz+pu/hrRrf87/Ipym3XftY7KCum7qQP5oSas
1cu/hDHahhEcSGLac9/AIj1uJGYPFzfyx7oMnWToNVmA2hhOJP29tuGkuDm52r2O
1XphPQeHKbXSyfmHBObsSTIs4jBTz7dPyZOuKC9LMoNc+TqWMiiuC0G6Jm4d/WVK
N66+W7yDLHYNFSIHTTwuahgOgPTeYRr+eSBvKrOG6sqjEHOHK7t676HZ+jCVUwcl
13irvYmb9lUejANxxdh6/tLdbdIAozX09ak7nsKBX1H6tMkw1orxol1z9ah/qeCy
hYsB/I681Jp7BEY6AdWHVWcg6qv6RJk6PPF5wFaEUGlofIVuk2JhNvLKDz9fMFvy
0aZF/ArHSxl5HAdVEuujUlA61Fr4v4YmMypJtg4R0bgrp2PRpe+MfYTsL4EgcXbl
CeISz1fsxFlODpL7lJOVz/KR9IlYpJAuN/FEb4R8fqDSx6aYdjxKhkGJdvVM/I+N
tlByoP8eLnM1lpiQoApNo/K7bULjslIO3atFu4/RBnF2sljf8XtbSrnP8dwWh90J
Qj2TgxAmLq7VWD7BdujNe0vveX4ZX1Br2MVT+/9TR3r9lmr6mn6vBTpWHfhdLMLt
rTvb0bO97Rylt1FUwtqALwUVLjzs2UYqrQWJhgYpjekjT87pzHVLu6Lj/C3hLo/u
K7KUHyR5+uuRDHknS3hNYaNhzieYfhls32v3KiloQIgzVFR6QBc3AcKUnUJnAY3C
TTNe2ea/z9ljTd/kqYvhIJmLNBxAjk5+bnswiaL+jKkgiEIAybr5nHDbe4h/iBlV
2QbPwBmS4XH/wuVpup+u9qO6nDSNHtItCWAMxiahJ4goj+T0FCiBT3ZYIcf9IKkx
JGQ/WLEcB+WNhdzfd7dbX/fWfU97+AK0ClLur+wxKoSmmgDMHSO6WadUbBcNiH8s
BICoJ/wPzo83hSvzI6Ddmw/3/DDm51alVycFW2RTYDcvPZjqgEyCWlBUbyEIoud5
tgq+bUBy0fjgq001OtojdXEvTfHTvT7KGl6wjS6bYRYPNEqjksJGj3u0bQi34p56
1Vgtj+Rl6zaFeysUP/FQyTuZ8MOtS1oMxi/flZ8tqY7UJi8qYuC9p/uRU4LX56CE
ZAJd3PxO4E49jode6aARO4X77NDhJJad6Vte0J2GQlfPDb3OecLwi55VtziZutMd
H9QbXV+O3IIjJNlTqNzvIVz+1cX1MN/uiz7oEjsmGyALwYwi8ELUFRo2rjxYvDy1
DbCan8AMl6z+eIS+y66GDN/KTvWshJ5i99F6S6/KVhAguLLkL8SfzkmxZFjKfK8X
hHj8a8KzJKqH9ua2/7aDTzz4dnvMhwFuDKqBPv6RrbdAMVMYQWf1ZlAMc6asHKNu
SGS0aVvwe9Uen/Rq6ZsgxNJh+Nbe0J26ryaImY6unYEj7jTR5Su1PcHXM50Gxih7
T/1Qv25nZDIxj0hGKzOMvFTKA3N0Wz1yKP/sb3aIeihyJ8I/+5mBvfI8HzaQTvls
BKKgf8eTQUAGO3KMoyEFIPhaWRF9us+cVtUkLve3TxcPs4DR5DM7HeUEjrfxvaJA
+dUop8cIgxXkaNuurHTHUcmSZmlSztg+GElH2dTd+zoX25hgbvGddBOe5EipJAxn
tLBXQoq8vlLaAwF0Fw7iU4PNL7dOiVfy4AEK5e/e2eXwvCU+X1fQyzA6JXp2obc6
9GcSNSbvnHRHzAP6Jixnsy71Y8vgDLdSkFKuFkErkEJV18KB0hWDjgVcieTniJH9
AKv6SGpBu2sYIOncs1z0pDillIbOHA13Kj9LTxm9YyipW5PxyK0QRGCq6lx/Ygy9
b4f/wrS/kWR1Clh8blHCEdbQaaFCdBESjHzfUnZjxrIckCiMZ5M4mDDxbDD1XGy9
8fpv/RZDnVjdZoZTwXcxw+x1MavVK5sngiUY+An/aqpx0rN6x7AKg8bXKA7KyXTI
4hv9eXbxTL00/RXsDnAiSlT/3SzrMgAHRbSSmeBKFSmUwaBS5oiHhVC0NlFQINcH
hHdg4fjemlfXPbV1Jckjoc/GDTqg3pVAhq3i5bMAdeUorfdi0uiO/P114wM4XeAf
W40C7P9qqvoPx566QhACcziSONUzoSPpzW4TbRPvHU8swMHnilVp/SCXoVakQGUs
jUo5b7Jm9VNBTyXl37VYv1k6G/OkfhKzJwucF8zHWz0pL937fQisoL+mifOEuSia
u4wnoeittQNxx3R4BgjBDx+Z6jCaWIbDZ+Jp0ROtz7mFEwLLsmhSZ+W9qc+p9v1C
8judnke50ibRg1k4U+ogLz8xJpP2rtVX0HHqoSAuMDYkVvQsXmlpqMf8sdo4UMOp
WZ0yY2zPxB9RXS4T9Weh63l4bJaYEMXnLMkGMxYeLnb0wuWPJL7rlJlDCZEy9mFW
GsZfg+DdBZkqU+GpjQW4TvQDuEYgKqrTxyP8KXQnu6xmdMg2iZt7uS6MiJHY9kIb
+0sjowOypjcti0QvCZIq/rtOtaEK7a3Lr+ZkWVRb4zM11mZlKMcp+wA29ow8lDUN
qTLPM0q3iM91wiMAhgvLPeFLp0vDkZk9gHXKBiqmdJRqi3ri3PTZgdxjZHAqNJM7
YFrP8e8FTayvxh/+fFYZlSt3f0V8WYiFJ3GwRZYTh92AJmh935FaG9nIt5Vp3lbn
xVBk5hDTtX2j4za8ItVxW+rCgF2FDizRG0oiHQM878xDS4Jdd53RDV1QJwm+2i1T
crArlKIBz1RkjYPRJyDgoswGmyoEuBpYzL6NpVKajVelj9np8jYWJyd1T023T8dg
BxOy3IIplvYSEbxVrkdcV4m446zjX+NMOa2FtvTYwuYmvAmzfTHS3xzupnzx/c5Z
XhpSz3VJwfjwCtMXT1FTPcLVEtCsA5LW2j8EbjxryolY++daMsJ/OHN9zRFcuUJT
H6CWzWha2qUkpK17ihBVThzb3zLN28Gc24sqijR/EpfgFsDHNmbsfSeZDGTehPUy
ZkRSZ/D1Y4g4QOkpF+Rc+MyI0DKIrfgyMTvqny9yKColbE5JJzqZioVHZiTcnxeO
jD+yVZlpppRj2X9E3biYIcHIyPB1u1jS79+47HZc+0n/TzF8MNoRbuks1Wn0DcjI
0DDufxhjENgZr+xt8M3i21gwfp5VmJi7affbp2xjn14t1HN9rZlvAXHGKvKID9eb
sOdkC99A1NJLOussq+BGoe3Zd8Tp3RoIA0f51jwfBwoJH9WKcvNzQ4cliXSOj8BG
5l9jPiZ8dsFAt3GDBlMOa+RDwHrDEgP+dcBTx4DSuHV9bB2EQLA/+3hU+fT4Rkk+
lh4q+KPSDWXbOG4NE228JGLYFQoK3VUrLidPSLFYlI627tXsSkmHWmOUh2Tgzwt3
6mw9nO1/3JQQhxHL0vcMvkc+ZoTtQEJdMCcsnGPgOCjgoiOH/jE7E+JcnWyTT6D5
8WWtYyXLOk/xGfPeQNwjXqvCJFquQi4h6pnFdq1REbo2HhcBBjMsBt068gBogyCu
xd8CwSC3I/+aEcNHShKG8H97N34X1XTnDGdjRjODxoRuIR/JPWtqqZ71mwWa/Lgo
HBNRH8pcJhBJ1Sz6bvmL2aYpsgORSdZW3qgqPH8l7Lgsn/KamZpZHBlxyMFvC53A
8brg4V+dP7LtaTeZb9po23ClHnKAOrwYIGBv+uYF355bSuTa480XkBQb8eHXLRkK
mcelINrYpxISC9VM8XhJ+26QxQ00kVZa3h2rOHpLcjJX//OCs8H4WQfA0pk4nfEZ
yxojr+2c8+HlMHkC8YZHr2JqV3JK4UOPqg986ScYJKo66mnzk0nlTIteSTZWtJlf
hRO1QBMoKExOs1rvetDKH7Mf3VZHIQ1PjQB9hPD/834/B0lEYZhKbK9NHu+nsmDc
Lz/0WBSztJAtBbqmPFK3T3vBK47SY4mqOI+pYNPrJ0DkHMFmdHvmWrpKYm+k3rO5
Q24kw4X5E0zm0k8Nk+BkT9Hnph/zEKu9vbta8Td8f6mo51UdDqXU+Pt4Y7XNNvr/
dszsJWF77MYAlZ+mvC47IzNw9aF6tegKfAeFd+DgZbRm1asPuk11hPb3vNT2Gia2
qprVwherthmmGX+CG4q1Xr/mZwoTC93tR3dkvE6N9G6oTmuJF/hBMbUZxOqNxkdz
p9B/pW4dFDvyYDgjc6rAZSc6xyrHuliC2ZNg5BtDTOOQWsLcbl3mOPge+UrG+VCF
NKFL186QsBk+Gq6qzQoWwNRGxJkvLFu+xn6YcqjcZ3U7xEzn1j/4UXA4IMceBFFL
xKhvKePUY/VN21HWGQlhX3cRU7eMf0gRjoH/X7mMnDCYvdJW0aXFQZ0CB5JH39Jp
uU2eKFvs546PrgR/iOyV3s76xD6RL/b/md9sVjq357nAfkYpCjDlAr8pjlfVBKf1
9Mh99Vp8eSn1381pJxNcR8zCtNSmB9XTdVLTWHZuZqgPYCDAzYl2s7G/E4xUa4Pq
wV0/RtHOIN8bXPcDXqZlEih/sQVdy5HGwGF/CIVTtHCHxRnVrJymisnVDTly5TdJ
VqOM8UDNdziotfSupD3iWoGm/XZuUmCAIjltZG8sDBqneF+5vxxtGk7KnNXvKxcv
1ZAD0A4IUlieyp2KBt2UiL7Ft1AUkDzKzg5WfqUYrjlBFxzltw8RxF/GZPkuy6mx
apcyQ5nXDRU9BGBxB+Zwf/qdcQnj/EqX9ID6BkjB/4nEdCnnpeoPFl4z2lgHdwfn
5HauTZn0F/yZXPhVc8rAflYpBxUthwSqzz/Ub8xiyUDEq19/FIz4jkKuydc1X4XT
dSTwdyEU3KBG8hjzQkEiNNveqgiQddnljUWGGmwup53KYInCzMOccGOS7wncQYBA
1d87Cvh8MnPMhNxewtQAx41Ynt6yg4ZS6ft3XozVdXOtRfp3CZxeXM1F8MK2eGOm
/laf2M8lLUzqGSKTzQOuMMVEL+pylrZvYR038HIY/Zk9IFrMlqC4cH3Kb6Vpxtv7
/wokrt0Hw3t+IWDjzvl/kq1CBfjk8we9/GL3liYpET7FeI0feQevaO+wJmp7my14
I+UU1R2JdA0pfYOM7perE9VmECST4j5kcah+yH4Rk6INodyvErncK8/07xaIY3Gl
LIoWe2A1w/yxGoQWLLqhKh3Dio2y8cLucl2g5XlC0Xs1s5wZBhNSBvKXUXlqQZtf
6KV3zJF5H2l8GNf0ryLmydoAZJffUnYT6BEp3awiCBL668DYKIRGgLw0tUbx6A1q
5x2Py17XKKtSMI+yVlRMAVxaH6ebXQGkH4ygggM24CZ8H/1bim9lKuLMml/OA8aB
H9MQfFpUee0JoWJ01CZu0KBWVEgEC7bKRzhJkKfvsxrSTKesxo9qhP6tIf+AmaNN
tGHfmMJv19GegAhXuLu7TA8mOLdAtsOjUvtAM6ixdWzetayGcUeI0gABKlDJjmWA
TLMlNcb4MhwPHtaZ7J0GcYGZZJvlgujwslRpWY0DCnhzn8Ta3YAi7p62F5PKdshf
sqKMhv1KsWKWiLccoeRxmcHkbXL9oocjfl0aCvervr91TFe/I3DCKfeuh0UiNMek
eJQ3X9LKMopd5qMeKmJ2ISklb4MfSCVvkg3qg8HDmulTzm57UlToR63EvAKLi8S5
URrurCc3NAYf031DSUhbYPj49m9RdyCxrgMYwV5osiI7akAZRMrQtyTjtV/nvrUk
pwGYZRnMjAw7RxY33Wv8mmcQTRsLM67AMzygIuL1MXtn46WJ4cdcFZgz/TiaedGR
Xwp631EVoOxEg3a3Vreuu5x19EiYnbXBEGwvVzhWCWWKMYmXMiJdqnuwSfoyG4Gu
PlH+E9DRER/j00f1TzMzgu3UsNXSDId9rzu+b8ARSZnS0T4BeA8QShXriYH+AICK
FGRxBy0cKXyinLmd4CLdvZpBxFrTUHkW42zEiBjU9N31pJEIILty3eDqwxIMlR5k
gnzIAoeVoK8dt+0kr/RQ3iO13bserwUx2jiFvSD4nM59eWZNfjcGDbf40IrGJVaG
ul25x5hLJKDGi+32o1f0j2B+EvMU810MMq4jEXxO8b7NQdQTp8uG6S4bjyGFiNL3
EWoKx0qdjwG5zWXb/SKLBDx/R3dnljUYLftMPAP+Rmq7dxwayS68U1NMf9ZLuWNS
vkneoxPzns8fwauSx2nIQSxfdFRNL/Z6gSPSMU3GFczE5B6XaFgurLGrxcSo3esC
oqVCUXsIlfEQ9Pz5aAUEbO7KZ2EvSZCFzr1HLC0P9MukrfpQHEGCLOrn7NmTpBaw
nOvicOlxoWIh2m0Wn7vzVXJ64eDde6m8jowlDaeVOsAg0uF9eK8Td5h26K2lyIGM
TQhTQAIxUhDTuyU9kBF6WAjOwXwNaoJ9f/oLQVHX9vWX8dYznXffu4/T6+aGu6vD
99bCvdRFRNVzwObglSkS/x2RYnui6wQqa+2xgW64TiwPTeNdSScdyiKv1qtwoWJ4
SQQkcr7MvTLwWnwrDI07AVUToWNpF2tJrjbKmRCEWDEbCXzccs0EprW7OFI3tHy0
/goS/3hewKgncSGZg/RQ9aZ6bJGNO6nAjyCPaA8w/9zp5ByOoxBPiBkFCk8i/N/I
9OEfa1xmk14suiULGteOZtMAWugV/QCB/QW4BOrLCVGedsJ5A2UgdbpNwm0o6y7o
meE+9oIVBsqGHDUsYf8h9uWJRUesy4ber+EZR3GNb10+C9EbUStHnmNqU2GLaEyy
fJLguOlhNGZTKe/pdKNslZMOArBz/xie/9TKCRTQOb26lgub27F+Tw+XTZzG0Mtp
+sJU/9vL9l4B4q1nGy9ySaXAXZGkI2IAPS7IMIIH8jwVek/UAspv3zQFeQbzCzS4
qtiUtie5CYYnWNsbN8OFzuHLkHcFsHShDupn2TSIlbzphDxlI1J5U2ysG+e45whi
Obx3nR1hMMbcM8qNfzAQZFFkEx2K/OG4FaX4yvVJli+EuJ4U2Z3nTZAqHZ0l3ZZF
HUZn370RA5f8CoNj+x08t3xw3CZ8LuolCah4Hhom8t6n5hauCbG79a7UQvZIu+Aq
3B/sUsJhSk+P8oKK7XypU2sujC6wKYjnuAGLiP/10vyFSa7XKUPQ8/1BeGVxYnOa
T2IvZzESw8VXBSApdJhqKmLt6mcTFaqBT/u4wZfOCEHPCVZzQkzuNwLEn0qTxm4B
J4SZymZDPxqB4n/TlVEwdRe48qmbDUBvWFCtuFr7I3dX9YJa4q+Pqh2BHwqIJyRY
JMrHRH+Iy4MirLWzcEb5dDN2fBpKw38QNE19WDZ83mplcar2F6dR4awEPGXGFWHc
/Tt3aXqGWNG+zyhCjo33UwvXzdVsO3yxSWdT0GCBJz5yBwWeXjJK8UNReghOAwon
reUgHJ/+bBG7YaoJioa410zB4DjCGjTk04bFTlx2PYwthLPibQelUbTuL9FhgR+D
j35yjIfXyrp2uIymrk5P7ByxOjQXG+3izhRLTP04Xi5dEshknf/egYvVcVKELy3O
InDiNkQtU9RLx7Nl2duogzwejn785SnDMAV2/SosLHkyyjVL/wXincN3JYyKmG8v
jFBZlVBXpH3YfYg04wxsR0NqKLau/+PIvFvrITtpUObahMRvd/ppy9WxtfCXE0DF
B58flbf/nkB4uYX7Shj5HZ9+TphYEyvV9iS0M18pHUyun3W1MK+F1AJjMFjsJuQ2
OxZSrVwtYCf3nRDOJOvfPrDRDNpPz82XhNaYNOZa4cToDLU1Cuox7IXr8Meig7k/
POEXH9WyGTu9yFB6bg/Dq/R5+hft9WsAY9Ysg4TZwJ1l0Wpf+TERikDJM23adf3W
3FTtrbfWuRX5DeDgMpb8wVgPH5lm6VGytmKkuaoulUggSCgf7BjyaIR3y/tD4EyD
99mmNXvw1CoVDDfZ91QNs0m+71ZmFoH/PZ7F3SZqyJ2dXuv3jLCwEmoBb2Pm5ytM
9M9ZJP0LPNxkgB5KiMNwh4U9O7RAJ36XsURpSbvrbdXtq7Kp6/Y4avUoQu7Sfik0
d2YmxIoWTMMKZ87HYvuh3uH4UwQnvHSoKIztJ+3yVkTpz9KpbZUa6Mj/XWzdHcKJ
gRVET5UETqKyY8EgSJPus+JTZq8VJwyTUV5eAST5WaDmi2rXZmPuq7ssAB8SOIUr
SmX6t8a0hMVesMK8pvYHagwEVTp4MoO2OBkWqdT1FyaKufsPIYUsoEUgGxxumXrb
1FTuzcE/Hyj8ZC7TRFYG3rQjO7mb7ILxJtA+/V/Vhr8V3Va6FgYk76gpJJUIiz4p
OX/EY8SIwXvIAwZM3abROF3goAYmlUb/XX2gt75v8M5eIqkpkzjIlk+09PwkE4UL
qQ9mrMQVIpFKA+ii5k/Gcmsu9SmHYQ4CZPJ1rZRdA2Ow72uaGDRlMiugZKcW0DRz
sMuY/2wWYh8zqvP7w8XjpGlzXULNRBHdZxheB432Vm2wDphKuIEaewzTCEzCpmmN
8UHaTuXQzjZovs5L70Jk/IQ4rKyoEqfuxjbKQz0MJnv5lUlPE7FJHfHrD+uPpK2Z
E55esLlljwAmjmKzFwTeVg3U+kIrtA/2u2/Ks7HTuCv75YA6kfjcf60N25qfDMFy
`protect END_PROTECTED