-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
oCT8VTbxTSXbTACMVyOuixBFxDOdCq4rvNxWb52dr6gCg+tsbwEZIjivShgsNip6
5YdGI2De2b6MlzBtJ25qzBIxA9n98qlm8QAon82lnvd/zFQzXMEeAOXT0JZnB/CG
AEJxGQfvFyyB2ScGF1E5x6ItTH4Z5AclSi7TSZDPve5fPdSCeN8a3Q==
--pragma protect end_key_block
--pragma protect digest_block
XiePkFSFGMjb6U8JTaAzgY5G33Y=
--pragma protect end_digest_block
--pragma protect data_block
JTHtFHh721t8Jo2mO32NZOytaWcN5msNddbyAEZmm4JnIWKGWneNJQED6jgsrTMC
fKUd3C306FueE352DG/XI6QodJ4JY6PeBQ9tI84YyYf3upOcfjQo4YKF37bxN6rb
FN6bPhskVJYEBfinhFMVf8sKnbsYTS6ZQMtPLj+EOnaJcpe6laldjrldj+LlWc/A
U2ffweNnFAZdh3yue57qiumGh4zCgva3XKmCj8V2mBSewG2+QbqtFR6b3ODHoPsF
VVFmbNMN6p/mrkaK1FXfgXwLAdrb1CV9fo442fTOdDAwXPgx0mV8t9OkRdD/84GT
THc5C5FUyvPMZ0/qckBtpkqOuXCVt4d3yddNcwl71rox8yfzT4AgbdtI/4ym8VSu
ej77Ew5kOLjC1YvZ2qaZC3ET1tD57yXqOLGebpP0tUu1b4sYu1w5OAaZifAO70RC
wa/7Awqr8U9nm6o6qOxT6LQ2cMvD/RLbrCGeed5R0hC5xo8KGd82osq1mrgyjMJA
5p8k/RMI+F/fxohIhEFqXyijxgcmPEaaSY66mHxgsXGLag+Ku2ULierRMh963Fxe
/iGcducAwQR7e6ZJQ0+xdUFiaCNbq3jZnfMR3eGWluM4wPGirMnRjgaZNXaHlQAt
LeiD9Nu1bPus4tSN3KAdnFYMoh5or7NHP1x6oUVGWkAz+IPRBSujQoy1XmFrmnaA
us3dIwSVRNFQaqSJQSX+ER7v6LX4/LWiFMy3hBV1qHqGgkdpnBffryCQUww2e4U/
foAJhzj71f3SATOVQBs54rez1KENrtErat4xEbf+CISD+l5+DPrptoaZmxO+15+0
yqqoSZPrn6wwvErFwTMFD4otuc1nDcPleVHtce/wLWMHyAoEomb+XLgNOvfwuiR0
Gut3Bj20I7VSwGtnBiv+8cXWzhPnz1DiEmptUsVG3GYB6olcuDmHttW7DaolZ5u5
l5M0QIbjF7Q5p13uFk3u5qJTbke749jl/F6LXexgZMaiNsZK5IiYnaXNrSsgvj/P
PWNfzrSrDyu2CSY+5gj4YIa+oQEdykS2kvAa/na5VFnNUn1b6AiDkwslQm69098u
vkoiTxlzl2voVIvCHD8+aqGExgUZaYWypBeBjocnWC2206psF3z+VFCEJZugtmwp
umPa166z7bWw9RkkUsREl/M1xIqNKq68NvMPnKLUokebU3zwEGFx1e3QtJk2S8mv
6GAMmrkFjDsyHhEd3PZs3dM5Y+ER6Y8YEcpJT6QWG2fj0w6bGKN2/GKWaiMbv8G6
AscDO9666TWimVjmAPy/RIq0exhZ9UmSg1xwV8X/Vvm+mfgUGigd2iU7dWL0wsMC
YLu2aWLQ7UMQ9oc7JcDel/RRO4p4T7cBMf+zvsW0rn9OWi9PtSfgCjbvt8IyJtjg
WXceAO7yeu9OPv7gtSI+z8uZ5gTLifbV0gUO9+uCQKc2NH598k7rTVPZFRgoSawN
Ch7r4FzRvgWKOVi5pjA4la6CGCcElATBnuzQxRL8Lb0tj3lntmDV7gEJYPpw03ex
6GW1p4Krv4Mp6cOGgtwwR02S+zebUoE+m00ju5YQh/278FnvElnGb+3J6e00RLVw
e1ywIq/mH5bmjQbBogF8EpAg67dd7kpjmZK9L2nw4ZRIWKjJjp+pzopv+7tf3ZbI
qFgj1T1u2U5VGa1X+4P9xI1oCEErx/tjGwVOY0kjhegsHeljXCTeMFmVdhJxznEg
CY9vci2eGpcuPEl6jyLCTTdEm3vFGpAQcCsqzkZ5ldxCC1CzjWdxqUaEXzCOmmXt
mkKfz5I+YN0/DBviy0CcMVz+5hC8gA2Gd1Dk75G72bY9/x1pH9ItAPUjSEC+66+U
+T8QpQGa4sp9svbAf6NG9bIiqslnmy4PybbMQa/GECLRdJ96UMi2ZXXnxEKaEZgz
bVuWlGWeLNY5h5mjOuGr9ti3BtDvcLMdyvXOVtV+zgirmGuqm0DiU+tDxC403+si
w0iGobRnF/BYir07FHUzLAzuOKqqh66oERS6Qk85NyOnE9trwLoljOv58DgFIwCm
JTxHjHm3avZcHbCQRWkJPMJiBdeHhCC0qNcI3OJET2htuOHeyqtI70H1XoEHI0M2
yYg9vtBdTRB5+T3O1rnoCo5YmRnteIELHo+BarS0nmvpZtajJcbB5MHHc5oTbZrq
/tHVB8msUghXRwv/jTrZt3KBuS9Hyly2q8QgQNPKzsvAtgUgSBL0wdzSc5N7HcgR
Uhx/5zWQypkcxP6pLB+VEtZHbNwgto6r/gwDvcHd1PVt1BY9oiJdzd24vAlIAU1Q
cYM2IY+ILbIdJS1oBqweFTaVyj/+RczFRYZzT3uw5mdtGboYLUPgdvlTJHDabUed
adhJLIrBrzS2E442PfGmepzWXizmq/miZhLKER6SYZ69mTAktXsQwn7m6kTZPfvX
P9t5dVvhhfost37CSGKJ1S/H95fddi1PnoDdef8ZGyUF3u3Oz0TMgic+MyWd7hXm
yumGpL/M/hGjhMyEEnP2DGyPwX+dOhkKInDGWaxmNv8omES8q3apc+QUqnB9ObKf
QAtViFg1yRSmuayg5IT8hlbFyPyuNYlFsdTMhajqVN3KvnEuO+7fgLQuO4YmsSYk
/qjN9/XlbrbO6r3ZHfHRKgVLrT7+ti2f3Oss3zhwaCzJN/uhKxrMuu0sqVOGygDY
EJerh/nn5u+/AH8TWzMzz+1A7Xep3eOqVBzoGgA5noGEdTCcg5TJaJApBnwq865p
szm/WviqvY7X78AX/TX5sUtECrdmuvYFJqhrUDBqYyaoqQG/JTsRO1NgX6eRjhnR
uOG6ctB+VgJvxP+L3dVMZJoDmX6n+H6mAQTbu5v0vxT422b7DnfTJycy80pzhT2/
ONn6NqA8GVFMUWZ4iV6hB0tZ4BY45HHCBK12dkp2kBZhksOutnXtnNuybaQj135s
1VLyXzfmupMeJJ6cBedCzK00zmNdCWy3ezGmQUx/1Uhrf6dlNAEifKciFJd0wHhM
TGzYwN0VU5ort2j7fKVXwdzZZaVmaKos33/IjBLos3o87mK/Ik9sjnK7IfviXIcU
ga15AoC4dpvDRIT7+xcGxUHIusdi7zoxo9U2ZEVRGCVCkXOrhs7aEja6SOT2n6qt
Y+1ugt3NCs9ruBKAjGRgVCObsVdn1ERUBdfh+TQBJ/gESzWT981azsUP9dPgUbz+
DkwSLIIMaegFuUHQ5TkDx5qzfLw8JceSTP3Mwv66QybnkjhZFYThrhJREvjEgppL
J4fdn1Kpc8SxY62SxjZd64L9CEWgY0Jq67Uq6mZ/wHSWxtrPFqXlHEFd1mkUfT/2
jNoJ/IjYUo/ESMC8M25ZxapIwaVeDHKRavevV1/UrceTSJ6hcwW/Iw9NjDR7HKyl
btlKTDL2Qk1u2lXhsVNjuMMQ3hTFhLYEI5wck7MEAy3i9pHrQqRSi3IqBnG+YFO7
2WmVeM9/GrwVILeokgkuLGFGHsKxwWzdSbJAGgti4OXJkEjTObqHpf8WYNX2c/Br
nY1qGtdvEY+XiB1guhdswaFvK8E4GvCwBva4HvBj5+giqhKz+RQfZviKs3v3xZAC
VVDWiKMgj02Av+EC3bQ2MYlBkFKqZPswcyxdjD2/JszqiiXYF0u5LUJRXXLfaO+q
20A42KLQIaKtBAC9aAi40cz6AkeFOeVEJhB1NOQx2eaYaVlzEe52BjtZFQWzmu5K
nxl5DU7I6TW2ZP280hRqx8s+g2mRErOOsRNro525ohR9/YE4Y+/HMU00OjHmLQT2
pJ1/dXESDLQ1PYG3xlcxvZutW2ueC+CBd6PaN73hW7R9MejDnwNFfITkHqli3yxJ
jVcRiri3CdSCQn1rw5u49MVLklRyMdTBpFE7ir6BZWKTRNWezUA1LdzB5h21fNhc
A2bMfaK5Eim3PYYB3xXC3liHuRSc8yYsAUU0Xav49/xQTz+/mUfjISNE+XiKHZNu
yx6LVuuuXXnWtYYIOJ1IWsQ+4f7CCB7DxK3L/W+tNbXz/eKBiNySLAqJDH2vNHag
X5lSVYjJgYwJltbujQiphPWQ/DMQWPExkRklr4tj7XzyVWnvyhqgSlRj4xE4NxBY
va5jQhaj+tEggiFny6Az12+fPpeWS0fkC/qybIyXeWAXxPT5touU+nFE0+1HvNCO
56g3On0luWqzPBvEotz1TdCqoCLpjJx3hDSFt1A4jUFssy7rrpbiKx5+OHxSsQT5
IeUuJ512GN5ftV7Ml+0IwO9NEL71BZmU5Gc6wThhXDqtRe1UqiSKnj0mLiWYqUEv
PeYdHQdZQLOUVP9og0Rlk3tZ+yNr0lcXG3Kg9U8oGRJ906zB7eNBelpJKj1vDNpp
+P8/ZOBnVeRWDTPJbuSvZXd7hcWDfogIkIc5saofUb8oGQ0e53lNyFl2jWLKqIwf
0IjZgggK87qtWl9IXyD8tmi4qzt72tO4f6ComsrZCXbQOVUj9ctcufUGqAhHzmtC
5X8LllmUrkXiUth9SYmCana3ZWKs9+VcpeMAwqxS74UfwB3cRGLhjo+ktDad7lv4
PRfKVNhD3qicjp+LO2ungVOGhUPBfuRTppm7u8MRzLsm3xAAbHZQ7kASVp2V14rs
l5NlXHQqbrug7bnobTlgzr3wQX/L7sypKm4PK70jQCaLIT88v1usTCxNPFpv33nv
/LfqRrk7C5UL0uf4624PRiVcNgvSvsGAPenP7fzqw3T1v/B67ojWUmWK6XQeziEM
YbLl+QXleG27BpGaGZZU4NrvHWFpmcsS0jfUupc1pvZrPz0oh03v2m1te/ing8HN
xBCFy+Lo1sgXElnpTM4tKEAuWK2poSIbDyHWVWSGs8nM45jn4RWXUq45v2dXB7dv
SmTtIursP/GCydD+CDPRkScar4URXyYmznPYlBshhV7iMvaxpzXpzH1/gZf3yZhu
s5jsu0jheqc4U4FCUlUE/J/Ro8PudiHOw+XeeGVVmB2wADBtKIEaE7w6I/QXOrmm
50iIViJvtBMlVwHm2qch8SkLXEX79lznz/AIBv8pSkKrCAhey4zE1m9iMjkM/KC+
xCAaz6LICR/fm+k2FRFFiDNfSznxaC5dP98QieakLVQXuLzD44ncikhupqL9i7WN
CUsa/3vLd1R7jX3DRXGPamqGpkcRS8kM9HscJ0QB3sxJKX71Kf2kukdLadzQxKZv
TpvayV1VIYY8esEFdMfS5vljs9iTbIYUU9guDsfmCqufWS1m5ovTSy7EJP3PRLiv
1+vS6qoCq63YvqU7tnRDHs60BC88N4vhOIQExHy5fCz6i8JqiJ5jCwlWqbAmzOZr
4Kpg6c+7Q0F4twbe0D4ISiwxtLJ1EK6zeSCI6Bexm1QE7bcQlRFFlVMsOn1xtLeV
iRSzpMy1qMlXJzTjSKf59ERHGuzyhCBoNgJbw1ctGDUEuylD0FYX/q18zuZKDwm4
btitAz0TlTYrOx5t+0iBPweRbl/cBgV28KyUMItcohi+0OZm9ch7k3hIcMgY9vfh
VN9GeOoZJWrKq1IIRJ+oXwQ+vZ8SosaJMdWt7S6+9Rgkh/PLAhbekagnach0JXss
Hxqncshg8jphjehFwcbVtN1qobQiCMEdvIEtdGor50m2bXUvt7gMvcnvn4ngZAtU
MBQpwXzVvxH8JKpt6TpSLdM9SEtnLcNAveezJJNimqqjB+QHgGsF0/ou7SvIyMw9
dr4u8a9GFqcT9BiqgfSg8kRTgw+ZuNbTJkoBoqRZRqIbuTOZWQ0DeVpHuB24856z
s3U4ydZjDrQDvFKyS2PWGkRaU5zNDkY5wzyCFYCSmt4CSSC1LhfN9NNi7CFy9jkS
tCMm4wRCnVVDPB5I9/1MSmg0dsec/JoowumzVbgSyPeFdW4iOMKADBK+AyjHzfNm
73EKn4MgkNtpp/RkMrV6lxXx4RQFhC4FV2cqmMOMNkZSzg7oCbDesrJt+mTj2FdW
3Kf7yvUsIokFlc0OhmduPy7+DenCmxwI7NAE/mhGmxJX1fDriXfyCs9FetSG/hxv
9SyQM0nG1FBXRCGNFFwkDtW1EaFMekkWtwx7OqFfNuvhxLcZ/jFz74Wq1ScAAWQI
rO5liLAYgNf7D8Cws5qVHwjrmFN05GbFnk463J7DW74E0T5JvFS3hekm9KKO0c6W
PT//vZw0bb+ABpTgoYt1IEXOBUSj2bc/CJhEc8jL39MC5LprRURYr366DjrwbhWj
cTO2BMs0oQFb/byHKnBTk09rClF02SGS3AxuFZ91lucXWdqSuUNLTncetEW18FYL
8Nu3ih+WUlT0Mzxh0wQmCtZ5WVI4Hd00J/YBA/NJmLKKmII7dSTfyolbIyICJA1y
QoA4+bFC7TVN8zB5DYJZpEe/pCHcDiPrRfWkHpb4eC0F4C5s03OOcoaCM5JJZ7+V
dzCAXvqNSMZs1+DJ/DItLRiGgXdM1q0G92PF+v+BTgc0KxxWsg27XLs5CydMoF43
6Twwq+yhBVN7duM6RdjLbto9J3cf22GlgT99sWWlrqv2maGOXTy+8noMlI4HijyH
IVyTxToaB7fVpdaBgBi1E5ywyrhhdld43a7nv373nd8C++nyc6eGQux+IONpVmok
3O71FKJNyUzpyt5QiDyy8haLwxgsfd6LNXAoJjpMvEMoOaF9LYGnTqlAXWYWvbv4
eya+93liSv5E2/6Z4giVTDaxc6PaTdSXtM+j1EbxdWeqDZqR+ufWFfGqEOxUbHDN
TwdVaNGM9ApslRhKnRfWxoRkW7+j72EA90FxWgChr6ewuEMf8G2Z4apytSSrZ8hq
jhvE69p+i0rIx+rQW+1Bf9a5ZOS3H6KTHTVAPwlh7rNYwIKDp8uf+UFmw1t8Z+Di
86Uxm9mk3SZneHm9/YaPQ58chXTMDG6qhKVxCyTGr/r44uRTh3Pzio1kwnhikFBr
b/hyeocb08C0h3+zk3VCQk+BjF9yzbSVkvwJu5PrQNTq3xwVOkOlD9VAo+2zFZZa
tiimYsHAp3/MblFwBWzIRgfGioXjD3YZOT2P+gzWfV+uKQjidRP5Z5BapswH4Axs
kZOWg9DRUqpyS82BDujNqtGMEIxe6thheJWHraoLAy6yTp+iS3n2ZWdchJUYhuZK
30yY+DSX2TS/Dr2MRQ2JAITQZ2Wn3adyLg/4qT/FAFh94tvIm92JE4oMbMGkBOKb
inAImQCKCwA9rQnZ87df6BTwbTcBfcHPESnSZBpbjUTSSQB+PQE4l/4sjt6yDdg/
fsqpm+GH8KO29VHYlHbeJUNF07Y5AOm25KdrUGx6bdtsi1sJ+kFJt3uywd23xA0P
fd85AniNKGXtisYnQK96npVHW65ImJxn+OzhgZsPMo8ThBvTQNTP3t/OUYX3Mj5y
uL1lGS4H5cpDTUwhlPqgq1xldE4KwuMyTBYA1oFL9Et1716x9fLShrPoB72BZtLz
yJnIA1gOjkS+KGP4o2BR+DRzTadlPpZjiA3bcqoP7ka8uW573TOG2pFGQ82szjXN
P4v4WS24DIRrWZutNY2dAw7Edx8g9S9r9lBU4+IvTx/tCIdxFcdTgaJ2MlU/cEBG
wEA1Zo6M7GZ8+OmxzsTv5pbdhMXXqxL96+JeV+GJkOWOU8fkcq9U46aDNxNwrfnp

--pragma protect end_data_block
--pragma protect digest_block
+P7/Nh7IgC/gKigeYeD9SgUfRdU=
--pragma protect end_digest_block
--pragma protect end_protected
