-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
YB7Lun/5fClC5cNvyMXd9pmOYPYKQhlWgD/fZD5v5LsXfEsAiX9IDmipElVMaOeZ
xviWU/FbP3zDhh7jlD/HsW8/va7PXFZ0M1zKFiPHyZvOWKeslVW3BIBL0hh+/46I
xwLIcNotNqdSM9hvs2sPsCIWQJuXrK1Fydn3EwvyQUs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13569)

`protect DATA_BLOCK
hj7yZXrZ4D3g4jmtYNSTFBb+usW/XdiKQEU2kl8Zo97gE+ZS6Wr/8MfhciSWgrhU
hB5eV8AOxvKM7zFF5pgjU0xIny2iopOxGOi37lzjO/mWys/VOsv4x4pQtIqlE/3H
sJ8rMu9ZmsPgew0N3PFPMBMSFluiknizDAwvT0zHV2G/OixPLGCvxFvFJItf2u/v
LqUK/kvtjRWLLPSXpyoCU8J5jkQwz2beAXeT6hpesriE0/muFNusrEoyNjsxaOhu
FQmOcm9jfMSRAFc5fag7NsSkHmiPqO4FfEV/Pd0+HFfV9t/Bw117BwPYbJ1iEQHc
jmWZCpj0od7iopI0g7uq7OGo7B8TA1cKk8ZLucSa+zxoy2mHpSpV0IHWU//c2/tP
G0/yTBIuZLjn6YgxBtnqP4sjCz54CulBT4vAdDGLbKD459XxESlmWvdles+8duFV
F/qjsGu54qbRWetZ6K4nIP7dbJwpQz/2EAXJaRPs40fRkPA6/0NxwOUVk5ODIbRN
ZGVY37UHNgrTP8OHyb29D7UPS5eilSQCvDw4qrpFvk1IpusLKgscYE0fUoS1TcQJ
7SVjWBLr0v0cJq2uRDRl9hWkESFpDURiLVVLAFHN11zTxUlgohHJsfuGYRGh1ieK
vWHksDT0k27WZbLbpjX6lY3aPckTopUhhyaW3gR2bLktP30v1thFXgRFDYYw5NoB
p7rIUFS47zKAAwHlmgn6TEi6N7mDVlNZoCKu/v5LVOmwnJSeX1kmDbpoQxAJhCUS
lc+q81fWhKT9DtXwaGHT8V0CLnuKSTExpvNFeoq7PELuyzrUrxi3Sih0MqclHiXi
gtftMBvfB4WrMS52rq1GQVawrGySHHID+mvbcANZwYDsarwHXCIu+Scs6HaRs0fm
Lu0qm8jq6VJmd+yDSmOb0CUfmrhFSxH+QRUwnEunSLMBh3jfbnOzNdMIhdJcDz2J
YgD/HJCY0B7pjJ+qP+/ASe9mmhZpwM+OmNC60tKVcpDaj54gtUfOKXmXUS9xTymc
4CQfyBNb0bZDjYiYKMwJDxyl2H9BFxyBMzTkvm/fSlzTeUOEZl91gUj9pPhsv+Fm
Izbnjj8HDeUTaGPYaxrm5o1iG4wxF1nmKyYkYQP0flAqDS1Dn5blJI/eWfaL6UDq
NH60fSW4fvsjexwV4CEhG+j1Hk7Jgqdtn5TVbuiL9H+l7uedfKWNFIkIfwP8mxRe
/OVNCCbwLmBDDuzw/trgYMCio3wNekhzaTJtvpWmurSppYxc2Qb5CrzU7JTCsMFi
UilFGEb4XhXJDgAdTbh0sAG6mrt25U7t4tQdrzFjrO0ONasPyCLFOcsKN6Ep/XWN
VFLhVwiF+m3PV3PX43bxcpc/+o+nbjeyXe85OefcHY+yYlXW78RwYLtx72THuQp/
xFVQ3xdQ0KopQcP71xp5IEL8wAW27tyOl6ovOt7EqYlBr7XMxKlgsS4XfZeSN1zy
7JPAkAFvlWL4niF5cV5uEC24F+eHWQw5pY6dRPPE1Zw7E3LRqqgk+g+Si9c5Spta
rdSbJbIWPPXEYHo/Q4bhR7oBPyMbMmRSOyyUzIeqxa4QMezZ6kzmWBjzcyzbBrp8
Btri8xy8CCIlTHTEzgT1Yp6aeJiqpSNUCIXMscFi6SJuhwc5RZnYPuYBXb1oSIbI
BwoTm72/tLvB9pHLkkIJVG1ghc4+R7tL6NAmGak9LXmQ3mnqHgiRo1SDitn4/BTm
Wk7QivN9PinBAPIgW6DD4TTY6JJzIjSPPSVL4t7g/ObqV2+nmixMZBa6SIdP5fHJ
FT6VMdhcRv10XxlL6BX0t4+Jd1jO5OY87S62DTu5I54V794bH9rkm90nh+WnCg0c
T2c9PDg2yKqIDNcC3pTFec8Dx/z0XWOjcmBd6XxrvZVlTONEbcwvIB7LQnW0tIks
eicN6KekP7z+1fkt0lnhOTEBTQOSJ0falHbYGGl7CcnxB7cWTqCL75ReogQJ96Xo
7pFWBaYqPNi4Ru8TLyPleW2Uo2TE+0poAeXO4OUOPyLSzZR0DXQmxx6fbpYZnhK+
xEcKkuXMH06QYgSuwH5qu504ETT3it1L845qdTe/CnWLu47bJh5jaBPShc5gq4ft
6CDuARVjKNX8qFOGdksxnYripYAzd/23HOC777sK88Y9nKe9XTbAs1odIkLqGT6y
p40XGJ/wF7ctwQNmoqI+R4ZqMk0PmOSAI75QtmlYxGonNWa/BpuT4AE+nh7/cR6L
19BWnYtzzP+VBCOn5HKZv1pp43VfAfXdB1fjZ5nWbw44ovoX9/AmO1XubrSRvY/R
JsNoKw2pwCFkhPTwNlqdfiyPToT7bKmflRge0jE9HSVrGkJrTA5Q42DlLDFRmYne
pel3kZCeuJKVpV+jSr5PGirQXSgg0ozN1cnsQMQPxmcmYd8DguhZW1mflxvLYuxT
r38lv6Ef+r0AgGWeWnOIDD65T9CqN4dw+VTTZhfmDU/x01jMwZ1rIg3k5D/kRi9p
OStlLeS0FHPdhM0AL2LUFMP3uaptR07A5yo5u2cFpLmtjHWQCu9aAOOEzaqgElgi
vUThg20+uThEXi8ycI3dXCT/hgOp9XadvZdtQl1EcvSNbQf4KCx1qiiD3o7o9np/
5Q30zqJewZX06nh/O3HaLHv9CV4nfB9mPnrl5bztiV39kWHpkgWML02mO7pKpbGp
IuME7bfEp0zvETa26Oxp41wiaY+IutRtX9lAcqZ5hSyz5euS4U0WFdlz7kR5X59c
8PbiseKlEC3bT6ZB7EGLeA1+1MTgjdBq/nlcsNP/xqVMk9y1LgX4vHeqd8+128jv
4jM8+nPRibiQvp7eGZATNclDFM1bBBKAB+yAZic8/p88/fMqmTjB22f1lHPleCL/
qODdpV7CiAvPkQsuVkt1Buj6s+ynJXWKi/kpn/v6d4zGcFb7uIa9jQL8tA4oVwPY
0/I2dy/Bd8PgmYLm6TNwcV9jKMNDbAKr8fh7iBDQr2WlyN1q9ffFcqwJdW7DVGRp
FbmdQKB9rLST19Oo9zxsfxoA3P0UnayNNTbyHhh+fw12fS/btZ6dFVIRbRDrIqRv
Z19YjrcsW7iX6h3tKxSV35caBtKEB05Ei5OL/wCPp6384uuiYzVRu0k6PABY0Xjw
xQBamLSzlQRTJ3qEKpGR7VOpbqNY7ithx+5qKnoZvV00gQmB4h6mHhEaiKQJN85e
lnIzBYBymqw5LIS/gXhT9XxAS0wJHeogdGGnorvLXgumtCgP+mse+oKqBYHDxeb1
ouUc/GBgrRbNGQ4xamzYkwgC+MLFUog8RmILeCTbMuqByK4cVWUdxehUMgaIkvp9
dN/WQ9T/AmzkAKdN3ku37muTkvvX+FCu72ZltAHL2YJdjwBlvUV6eTy7GQ0lmqQr
obGkoX80vdLRPXMD3hgGgjKgq9xOKJ2ByMZ7gnl1uwvqYfFVu9j2rNZ5gEbl53z3
OouwIkVVQba+OmHREe2mnRw29umDtNYOLZ/+4Ex2hFgSmh1OCzSTjo8GWoG0gWBw
Ep7evszOJ/7PyGfL/bbmJhYuS9GVHr99FC4uKyTH5PvAU5wNUEsu9J8GnADvLp13
6huCSDQp1wWEJxebGdt58E1HzIjRdej29LM/W4gjxD2FJ3NzmuL1d7pMNO65UsI5
flbA1cnK1bYHS2Y31Jn3FZJrlcPvuMfMTQcilN/0Bg+ejtQu1nJW3R42EBLuL/zN
TGHlBpYv/brte8czCe+4NqfcEaMpI81KEzfUDclJHUKLdWR/5lokOVD45/M+91E6
SHOU2FOq2weuGX98UPDoTCa6L3XK/7wTN3t379VgCAfeMO3jHoMsXsZIgHDJk5zY
wn9l6gxgNf8sjX0yhLdw7K736+uP0mAQMmfv7WSidEjPonEiK+27JL4U51XZ61yS
mfLGhZ/PQEHF8K296J7LcuPT1oznnCsepckeWxvMXW0TY8Bpd4HpieGQ6vqzxt8F
wKrB7rNe5JY8OswHI+FI8Jim+9wIWEIk/2OqFEr3ZADzQLRyOFs3N2zdIlfQ21y5
3FVeBAoL1wcC7QuXPxExV4mEI059mDYcMBLlLv8a0xNmfuyFk8sG+5QJ82Dvenb5
GzU79vNog7/nKFYJJtG86C6pRjHw1dT4HFVk8fPBq8slCV9QV30amqBCoROUqs2X
+5xkqNvQJVNMwNTcarvp9EK2kjymXznIuJlz8B3JSZxGD0TCynmwtG1QmP+KR42G
srHAUi66e/UH8CKHwRtSzWDnNonyE1pUeM35Vg8koFc2DfkfodF+krqjSEdR6VHf
z5zuBfSvQmF4FHRUcfV8IwOCUDuyJyLIOQd+FxIrnFkdbiRUOcRHLAcZv+56BvMG
3jckZkXOc6B0BSfmJNLBY4IYtkOGkNZHNf993Ya7w5fmjkgW/tF0dM7xzfwYmDpn
jVDDfNbi57Xpcux2ueOLmz3inbQVOhO5yA7V2KZ9cYfi6SDv3t0J45uUgJHIAm2f
HU8RBLCfFFOEn2ayf2sYhWu0wBedngoelbp8AZjcduLxOX0dHcQ6KOAneeb+QbHi
z2PCJACuAVsQrVkVR90l8tiLijTmR/VSZaSUyBx9NguZST1NUaEb1GuI5g/8tZpx
UCRRh/9FX2z9mVUaXemIkQpyalKdAYKgVQo4MBYuwVzwmgdJw88pMwUE0E/BSzKz
xS2Bp1VTIhDeY2BreXwS1egviXQdd/9oqu96H0HHSOYwZbFQcBy5CNGj23A7KAnX
7CjXCpVCbZ7Bm4jr0rL2GkLlDlQuSVSjpozDrAKQgTXoik4gERtK0hqqn9LtM2sF
aOTIuJxDQPDcc77G9OCNI5NLyyw/UJSK4ZxJCYYxy0I1QgM5gQf88tlyEKuSqbde
XJM35bju3umIhPwbZebKMvVsAkcDfy8AJaoExB6glpvjjDB0pVVuk17tZCEooshE
JNG7pCuYQxIIWTaBHCCdmFvAWsHtvReSPkWwLPxfx6uxskjyFiMQF3rYzmihJ3BO
vwb1aGiotL9TXRGEqR8yd0gFwTr5A0rESmyu0tX8JIsbynWnrHYoC+6qw1BcWXgc
3/zeu6yEdopIhC7OqqdFKusXch98REBF0lxVa9LLGKCfdIdQN/uqi0T7Ec/hPlfJ
bYpUhSVxqIAhX7IBdWDP+ZqsBtZ+KjLybAifMkOwin8kZMHLrGaC1hNAGuZWXCcO
ob3Ty2mkP9TIGaMAfMmuzdckYFRoYzuX46jxx0djRW+BN6+ghrhDxulsDWVnUyy9
gQOfnCthfkS6DuL1ya9sfKAy54sVjX3qR24toEe+QIFt4udO9W27vAhgTxzdIHxF
GEAwdqnhFi+bKW409eYBgyrE03WjBAedYjn04v/t1hgIqOn5iC6qfjP3EH7JO0DS
WSjFITOsaqtcQSc0JajCQbMMzFIOOFb58UoDeClbQG5urMnukMYFER+F1IXRxk3Z
/9UFAAUnZKauhVFp0NGfH70nzAXCSDhBB/6HS2zK99Xg4bpc+Cvasog0oyZtJCZU
3eybdfBo6h5jaOwe4cbY1IE/mdTsfKA0hAI2HhbC2NbqK1r9tCopUdzwmTAXhouE
0LHu6ttwuhnsgCWk0MUTwU5PMXWfHOT8nW5RG7qTZglBlS/ZUlgulP19gypXm0mI
lyUSnVGxL996zcp6KgCi2vCTszjRvpPuD7cHgL9oE1k3h7oz0+6Yfz7AS+qHIwyn
zZxB2/zzIG+EuKRop6sF8y+HMOLwCAuU1W2WZWfc3kegfeoMBZs7FVNTqaBLrOs9
1d0jHTWHrwLZmTTAzTpegmXHZIks+uuALfoCfezIomSimC5IH/9pOhrJEpsSF4Gj
Av0mXoOQtDcjHmjSBCzntckHuWGY0iyIXQTl19jH2AtFC3F95R7dhdrcGQgsr1qY
2avxt+spyljlJ9qcfjUPSgzDUaA4B+zdWJHmkJla6Pymmd5a/NwaVYNMg6c2r/dE
CGLLgbVkBQ3m4awEcbiy3l6GFtN4prEwHleGNo+oAR+V1qGk427RlGeCcSzUjt+w
BnpkqPW7u/5dg2t8Zn88YUatVp8D9TGPFciMdH/6iZWxN43x+LmzME+QuLfSmB+Y
z3pyU54Q4TzOIsftUqFQos6tD/7PKQHjirfVVMyDRdVbhH0NBwSIo6IP7as8OSs+
3SIZY7Py3Pa4pcW21UnrFE7qFyXnIIM6BQoZjx8gC3ZGcxSY2inpKe59l9vJSvBX
i0rKIsTtCFx/hRrhhqLlIrAaHigtPuEE31/a3gwHQwm99V70XWW/WZXFqzxd13Sm
Nr8MJudaW5U8hYqsFIThPZ+ZRrhzU07sIcuRgumFzSUgZp695RPBA5NUqW2hm8bw
7VWu2fsMIJY+vK8mNsU9QhZLD8x5urIx5glaTxOr64j4+uSxh6RgEzG2eOs0x8Hk
Co37y7W416iTF/VIwsdcRbZPgMHzsGUof7oT7SpZEzQFKWXFc4Wy19oAhfPIG1cX
BB+SbyAw49mn+W8adXv2uTpHs9xKdlQABIb4NWFoI9mIXHHk1NAFWwcCqVJT/SEL
RCBbEMAvdP1oWAI+sZnmZLanAreLbIYo9BLpHlRI0VjnuJC6nI3j1jaf1E5HKXdg
Tlh1xLMJBp73qRiaZczSBU/CWSOk59Kooy8H6aKmQJoOnoGrzS1W5ytl8Vtd4qSS
nw3b7sKOKgAPK+XiGiFOm97GExLdKZ8LG00vax4YHueYkgtXPaXpN4LDxcBbEWNS
tMiHn0MAX6GM4mrhcG6nJpQim0XknIpgHWsj4DCtG8iuvNMyYxC8pEQTE/bW/P1n
lOFCZfgE5eggZsvnOb84exDPNrs3kk4QXG6xR6zustWdIUtSY0dMugNmHXNYQhEH
05KE+EjvHQYERM15djiBw6RqwQ1J+iUSyVd4O2q8xuwatlR8c/OSZ6NbhhyIGcuZ
05bwg7EDN9athzyv/C14zCR7dgEo+UH/FWuO5ImtOIoIJvMNO0daDM42OGhOocqB
TTQOKldXf1zYCnHN+t2iawvsuryfN6YdSxTiJnaEbGU7j6rcsNmp7ehcjfZy1JjK
Lx0JYNAKPTJJdlwa/OsXyQ1Jsh+QpwZfYB/lTwD8El41coul5BSDqAUUJdLLgcSZ
DbbgBejWGzQ2f20qGFXsMurVFJ8bINCXRF+T8r0VUAGDWSkza93rG7nlTvI/ih7G
7qIfhZ3MJ+UUfYka0NL+1Yu1FyccGerRFMg9b209L4Pb/x/SX8yzzJJ5MOmvlA/4
co7mmQx1mHaj93tCzHMj5Xwjad7EGBapIYwfjrP5NrKevzmrPNxkqeCJUlUPDvn+
ZjaislB0a0SiORKr1m9wRhVWqxslSmxdt1RKCs9fNOMKPZFTbuKU0Bc1JYu2Gd+7
6jJmcxFBl3JnKmqVfAnm4V1YCLKY5ZhVVcCXeuCvMa8L+1/lF0hs0y+wl2pxF1ak
hHwyczEjobXAJO4TAi5N0WpMlvIeVwR+HuA8HeVQ5ZC6f/FyATA4tZP8VXgJB9Gv
3EvS2P3cxjS3zgsFitIf1I6YBBmCXdg2QBjGj4SwsAoPJ2nGLiPYFFDupioVd57s
vRXni8ryYErSak5FL4cOaNKZnUQUChXdHfIj6rQOrfPYTGR5HpgZdFcKpB9xNCA+
qu7b/I9fXJkbEHfd9oRIU1X0nyZv7Z61mUq+eIdgZPjv3Ez2m2VNJK+QHqXzTUzA
GWUZkF1A1uAz9+d7NQwy4bz240DjcbY7/59btOmk6LfSKwOk9D9MwKU2mYWrqbfo
440vW6AtLjDsC2sgMthVyVvlYVOy8cAIlM126FP6ek7k98hFU57knlvGzeEhk13N
1EI72B0gghKa1omL7+O4SOkwCNRw5DWfRLM1vRwouFdBcrfIykaXnNaiLBk4UjgV
ggnsmf5jWYrMn5JIr/DsmODiBM3beQuqssdEjDFCMO9CwiX2mkR35VxaoWXE2xCs
eB9c+5xayza0HPC180wqkW2QrDLTi2EKoAMoyJSxulhX2N4u0V9yJ4/+t87cPGSr
ndbe4kLQ0czk9WV9h6YmC0YWc7zMrl31D8Pgj5PplfE7eiW9BLAFL7AQOMqlCwp+
8nvFX6KKPdR/cbuUCC8QyIUE5MV5Dt0uN7w+HAD5OBXWnDtBfJc/d6Ud8bxLb9v2
NoDZC0+sp6NY9R+ZiZ3iOLF7kLSWPp+7zW89/kT6NQfknl6ya+UrV5YOXFuwruHQ
8TN1b23PU8OPa5vJbXpS1XtspbqNmaG0i9U1RtWGmuC10Vwd+mOqYYbBlC7vwtJ7
AZVPiuZHphG5qK74sVsWEwt0Ip0xQkrAaLGnaRS8NPCacfAy5zoJ96xIdbMmfGQl
wb++MoebVteq8TNdRj5me1iHbXaG2ZRaS0+150etoSyOasfG1jKYslv97t3UtAkr
emABrWh/XVRkiUYqfBJel0NHEzu6o5P2py7UIjYzPG+OGJMkpqQdwHivjQFJvLlD
rNAZdE342dWpNhfIFnE8niYrNyR1RarI3nTKf+Trfj4apTLMfsQ/nlqByI+bVsiH
EzNiSYR0sZ8oSsBP7ULzOWCRnrO9uECPWtw3HeF5xT3/aGku6Za6mOycy65wATvg
nhK9Z12dog6T4N988/3V1qJBFWrAIMtRIii59Q/AMk+6MRac87H5KxzkZeDqvLvl
ClEQgEvf9hGv/15+KRgZnls5DIxzStWr8/twXOeqf4ijRdtYAVPlSmBBj0T10GnD
2WJDZVVzo4Yw7ChbN5EUfSOSNBCuGsKHbb5l348+mfZENZSylKs3wNORyjiC4jhY
2pxEcPEDsnZ6z0Teh7gqc7HoiMnnIU3/fwV8T8A0GIQwtGtGO3IW4tFQAnSPyS4U
s0AcCWlV3lLnuPMovKQgYwXl681IWkOYl3zHNu3VR9/l1mOSOZuw6GgWwiWSFZsB
3k3BhKQtKRFwflcaRstr4HQ0Kx+gqIrY7pKDOtU2zmSrYiBXyDDy4imPSWbMTeFy
2J8VmhqpnS8o3PABK8Hl0dqaN6/MY+V9MUdJxpOA6bvhFmx9cfujbu9JH0zLL0pK
k+AEfQlFuEFGKwyNtThcTKLG3rr/w7sCfzYni+GCbxBmnKwjnfVAIVm45km58Esh
jPV5nKaQa1MpjkoJzDVtGFJkGwIja6gX7vXzecK61KVvLkmJNbSIdk7+8kMq26Hy
sXIeFwRVcT+Wg23qoLRBO6eUDo56mZp26/3In9/I5n+Mk8xQbYXX8XoZnNa6PqSR
xuaoNpxgacKAMDntZWBlDF7nsJlM+gAnG3/8B48YHfPjc94lASlGez7OmIiIfrKG
KMgLnwl0XlhXTH6CO1ZeT4gEn/gRmfQY00KVplC9L27iLaRM03q4Uijzh1RUuYio
TGuS9O6ff7qcx8y0w2A2fhQZjZzTrAStpRmBz4X2cFjTs2fAv0SwlX23djvL/eqF
hQn8u3lG3/6mxZ6N7bguz52yIH3zGHEE0cgI+0WB+IaPq5/M5D4PTk7i3iLOu6rk
iHzyviykb1k+GXXUSaHS80XWoixDEn3dh/oGE5D6tc3pLQyjYcbwcnU+OyEN8bMI
9yrlxWA861GBfbGnrBs+AiwQbDN6mYcgx43FrPT4IY1cd7Gkx3X7mO5qibtphG2F
iTxnVUs6vm/SCuxammkhe9s7siaLUbGR7JK78Nqk4X+MWVQdJZpjZI1mM+oqvKJN
zRGFZmnxiwE3A56UPd+0ou7kTELr5GisYuXfLitKMGB6wV+fg9r3MnN1XANc6RxR
IA89iUbz/DBwb0JjUrmtAo//MA1oczfE+uxZJFjGD16FGaLjHz1mugzSb/w0WrMq
2W1yMV2yoVpO682ghgagFzsiO6PxiLpcxoLfO58qzcXDL83URrRg75s29Cw8u8lF
GWEP5xdMs2jRL8qjRhpT7pqmW3tx2vBp+v9hXqHKxPLehTsFcSUw9098M3UcKnrM
TiyrwR/+0XQdTMbAOTOmvK28usFhqOQfnDoD0OkvMSBPzGcM7vQG96C/0dHL80II
rxFaBDxmbQ5HfkBqTShABXj4eC4bLQOkskvAlseuilFlJnMGxEhIYcCVyKhj0FpK
hCyT1Iwo3ycB6OPeLeohs/3Bk1skUHaQAKpA/wEv2oCAVIgXY2ymGwpUWBkof+G2
9Ach4Rzlo/9WjnLu+sEbG1cc2vuTDvbDiu4MiLK1vuq7scJLb3Yyb+2iAvJbPApD
cPTGUu8GMomCVGWkYdD2/JjtYCVdquJLL7VKEnIHutgfaq65J1XPdkEQDFPKsjH8
88lasQmu5g177H10TI3dd5RHx0w7eKtKTBNNRGYoK1M/84Iif4PeSZRTpHeoJXXa
iMRXk1IrkbkuCRGrsg4/qcDaddMv4buAvIRo1D90emH8q31elQGgAkwBMT0WFGmS
nyixQoSJqTvXavDMHFqy0hoIAgvmP/7Ej+Jh0cogllHVd4q9ueRpSvWAKzVW1npj
t9O6Ac2oXdA6V7KkinaL9BWtpzr8bVwaZK1G2PQ1xxK91BUd/+KdBLX+7mi8a3WO
CXCnNqs0DQBNcTo7MCLoOIKyneQivjXH5oR9K6VKzYKhdd+qrg5MVP49NcT9jmJc
kJaxmnx/OkPJSC9FZdE4T23KPUl0Sp+R4fA/auVxmOnQ5+buPV9zHTGSGnALvvO5
5FNjc1mIGBLDXsQw0xuJgYuzrRxfxspz+kd1T8SxJ/2SC4ofI+jvFv1prPDpivx3
/onQaOFmxYlVGsY9prtzjeUJpTD32evBdm24pwU6gz8ywGbR2iSzqXJ80Pbgu7V/
Sjc/Kbne32whxBK+lI1YEqBTN4vhlfAFqBE5stWXNKb+nbXjEiYVu9bHw+r8cwEO
ZYUZ3LeF9ckDzEJe9J1xKj1xMhXeTaF4t7G+XzkPggn+arzpg/rElOJZe4pJ+2cu
2Bl5e26Rbz75Po1jMi3KfDYuI88gHbBshhlXjMRHVoBi15CybHNFW0grnLPinmuY
1RkZnuy0roATQiXZfO0Jn2ZM0mP9MIgdb+IbrAzh/CP9lVw/UERu5w+i2oK9lTxv
cZbrch4vkZpgvaU8gW6I62b3p8KXz0q00KJo4R+u0c8JaM4pu9hvXpzxjvcJmEit
R8+pTJ4n/ThCv0qjxj0XsG4opd8NgZ/2qAOb3laUbLMfIsp2C4hHhqLSoLr2i6Q4
tftBO6RiEuvPHjcSoUMlxQTWWsBsZHmNR55MaYj4ScXxD0GmJBGm594Bo7gBTqIb
8cHJfaZtTys9Rwq0hSSr6r6tABVgWco+sbzAPYtZuKjsfxZ2fuTVfEifyu7AE1Rx
KTrYCTgpwjx49GdOo9AYGeobGmrQmGBwsZNDFD+VT7jW0LyHEmejup5m3c48pbWZ
ji1NIkiFrUWPpj1QJPOC6gkGIgCvlpbB24BOWOYGfiqLSGSRd96UmipTml4l79wz
muTInYac3UThBmjJmpKUb+8ECFQKqAAtAX/JjgZXSihjAYU/x0t3ANs+4zxmz3dO
AgMlGC0k8harhMXSWc7ok9AvoGW5eLN0n/y7CC4l1UYgdke3kaYx9RyAD7xM77Wc
/zK+4gT9FmoUtoCeDBUZlPBYwpz1e7Qfd8g2rAziAH6YSCsM/JCjTxV7Do5ITcbb
TW/A3DM9zNlUEpe25+es4Gp7qTBqnJIZXaVRCOWP7zXcxW8oQO+YZgNEVi8urI71
m3QTm7FVqEL0pmcJs5ao+zSiLbcerUE2P3RakjfvBL8NVYJpMpQr+d5Bk2tpbGYN
jd20vU888s0Xy/RD4FyaIVI/O+6lBmy3FVJsIMztmYRgQBP/K24hCX0fbJnruwOK
mmw7lkKzM1NfbCKn1bs7qhWTe8Bck+g+4CDhonnWH66z+wwTrnQFpm4dESsFA4L/
nVBJCJK6vhLdPPyD+DiqntBgG8UlAuWml2uhOuaQPOiw8s1c1UBIaFZvFWzJKAvJ
u6Gg3b4gtCNKI3+NHW5jZ2b50ARS6v/djlPA3ql/gtZfrrb/jF++UhJIgwJvZGzl
RfX+KTT4VsErHMuGopz7fAYhnbn8a/wbPW8qCpcFGM1kFEkRuA62+Pc52fjbz8P/
qYkCrDN88qxLHjpq2QmSsMvaREicxCGnX3uG8WY4v+RVJuvo25QiriVE+o8HuIyR
r91WvE60knemgFRkN2+gtFrR2kJU+BWuNI62fOlSWDGs8r1OdhqNlQVOdGct/vhc
P5/giaNdEOOemqcDgjtfERAgYLwaGVGoC3xbyaZwXcgWwittcB1wBApkHJBhInEs
IfCZH27gyLYqJwNoV046rqL/42tIuxqyVVETuLcmiexy/EEG5CAiV+tPuVMtTLWX
KeDqLz+6MGS4mWTfY8kDCo+cxSbCE25iYmxwDX68bWmfklqoifRm6VFydvxf699G
XayOzCNKHEkPnmkNalKTXjdBc/qbFA3b1sy5bKMJPgERghMhZwLLRyUhTVcnhYH7
1b/0CpbFPFaze2sKtJY5JSpKzk6t5aRbXOgy0NAF3ypKK03bQ79Gpb+MYbHT7/4m
BMKFnNAPV1T9p1JLDxYwfuQ3zkOKqRig/38z36TTfoN1szF8H2CbQbYLp6wWleMz
RBSGqP+UbT7pkjU4neyIvtwXP5xCSNtS3YReD/peBf6s91MGrgPwxPMRUGEOGUea
YgpF4jmxNwdbGv0qRWnJGjkFhtv9drayv4pDFelgiGcKdMDGTHPdpEKer+R6+p7M
AAGIDi2dPKNPzIouZXDVKagrQ0w7pgM4n9DNFghzY1vipfa0s1eFkoO0uupRvpu6
ef0fcKfZ1YJTgCL5PQffhbv86A/HhvdTM1pKNFNk0UF6o4+4ihjAuAJ4sSyfE8nh
vkDnnkoQWV495bdad4hzMZUrqSPXLDvQg9jf65TkyRJq7bPeLwCCTft4WHu8BWyY
O3i1v15HNprV4k1cokRgFjSwPoBSX9bpLzzMoPIg7ZfwKTB6yGDAl9GExu+jZCjx
1uM0yqQEH/8C+YmV088I3tVohhQ2z+rXW5tRuuQQst2XrF2jcZj5gchXzNMTFVs/
Ey/vZU3/6AU5ppqiPABiRQ1heeZpQQZUtYIFqoSPKugvS4F0/o18Kp+E2sOypilE
6oPq1RoQqdVqKQ68b0A3tvA7TSfFlWanyOWttZpOsyyC/C0H6PZx8bPyEqCNV7Pa
n5qAiF+mrs9mYQzZ+NVg3b3oFgufRH8seZivpejTKhSg71NojvswYRjyRx3UTmNW
PvVEFl5sQJGNgZJoWUP5B/M6u6ixM/pooqrRfIisCSTCbDx2J1rxP1+If5r+T7+J
gxsDhF58mnoiXHjr8qa6s6ROrNSINi0U9zNHYwRXuuGsnts7SljGY6i7RkIU0pl/
aJLNjRXGXirbdlKvmLo1OeIFnWRP85sJDHc6w2igcpoTc5VVLECs4+xv0BbtkpSO
cj1Ak+87uoV325UU79awKCKDiEnAf47E3EdREGSm1TvEnrkj5a9aVlKBE7nnKgOk
1qLAE13hIfj5gsNwxhTVCdFu/2aQws22GQGFerF6pBlWX59nd/NrXk/UO5xvfsWR
/I9GL9IykyazicMhHykZ5ff8xqHkETGAn+HcpFOWtZN0ywR1iUW7lNTHlgFS7Da4
w44u4vvRuEefYfJ9sjy2UU82DKAY/9DlzCB37cm8vzbvZOA8e0HurzXD6cNMXBYo
I7xUaTeCXB9G+EUb0uHIgZeSRoDJbwvxshdCdfk+jokk0MYW4TQeNZRDbVjTZkBl
yYZpTOUzrXDMHzol4EWARpy6wdj0RM6mrnTnx2sIwIxfVzzooxjSJye7mbK8nj9h
RSk8yUrrlsS5x1LHJRaE8rx+iHcdjMcrTfcJae7qG1RZbsOI99u/XYbq8ClYeOfO
vYZCchHr6jKxJCxhdhNZ++RgaWpdqWhg/6ZGrQgx6TcN39gKz6KM3oEZc5HNCmqx
DtXqL5ahrIeD6QIkJDUMj4/opBP6sVrIf3ZGeVwV8RF6XhnuQy8Y+PPT4vaTUWue
5r4UvdSh7ZxPQjHxiJWai77ECwNOrSlWYsOg2xNzd+N6VC9qwWzpcaGe7jyHE/H/
zQimID8azwoyzQ0EPq/dAleWDA5rFPU0pMFHA4Zte/Ym2uSdlPrykfz7ZfMdf3t4
MYnymiySyCb4HdsiabmlSiJ6cblSxjGKqlLhiZKCt3Tx66h5+hDXUt3c+gmqdqWp
ZQd6DMDBrCq3beQf+rgX2zfgxioBxj2TzVUp5X8pWy721fcL3bW8kXwqkmB6CmkS
APv9YbgsRtXtI3DjDDy7xgAhbfw2E2C5mRfo6iuxm0wYueYUnb8T4cZ/ZmfY687G
wG8LGh5jwrkgnKZQm+ZGQ95Zft5qgvTuTu4L560kjdSHIICUcGFiRzM+Y3bsJomU
DNoJOTQDQl2RdbZbneyix4dhI7OpgEBLRC45EJHtFdS63d0gFGLKpIWWLxKFwPCf
sN2vgBX+BNct1IIFHF+QZpOiBKVLGPHw4pLV5o7aZTZVg8tTOSXco11mKmrJ/dMl
pdEmQwnnzXHztik0v01dDo6pXtF3cS1BAbC1eCTAO+Pgo2Pef0SAiP7ewbdCnWuQ
eP7Q2hct8Zv0Vbl25MbA8POOtTIA8b1E3zfOp+PgSGNDL/erBFUyOJvnS1oCPyuk
n+lV1UR7beiL9hZwnL4ASvD8cBUpRAIDgcHxXgqE1orBc0xUHQn9zne+K5TNk3TP
Po93AZWdKcbvo3zyVzUmC09xS7TUxaq8oqqrClNeT7MWvoeu68fj7kOExkG6poPR
0EK6IAqyOAYWdY/ia/EB5vIUmGUztxwgiqtdhZLV7olS8VY75UIAsOulN1v2D4ux
3vySzx2WpfUk+5hcq4tNaII09GjsRQuZ3CfPoDAnaZ4taIH59vB0oPphCnPm/tz+
VTItAuR2aa7zvj5D5axCAM2i110ifzKXxUsH7nTkImIT1nSyLzk0srQooPf+FQYF
8NCJFf+WaCroDTEbGPfB/fjmiWA//AwfwxKFOV3kdG84LCH31e0JJ7uwa80iOHRy
pjb20uyerX8LaDclPoQ7h1lKCT4dNoFoEEbC0fXtFtShWBFWld2LVZ/ktTRyU5K/
5DBGYV2BvAD9W0ZrbI8STy5DY2hM/pBUBpoj2+IN33IDN0xSG56FKd4/cKDWpPTS
JWAChr7IFQw6oH0naUfud5qYezjBtsCjTrxMwYlyS+xy3YU9TEllzbTKU6lTi3Hq
ZrvXjnBplCYsbMYUXojdAVQALxpqw24E3Uo4xdX0xXaUObeQ8t+fC9OJ2qjbptI3
XCEFd1ka1bXtvgMw3mLFqFWI//iqE1IMN0UYmN5lROA1Amk5JFInTVvpGiyhcqXN
CEda9SdAxc4Rz49sFw0bhf/yWbfm4mX90jHVXzOTKnHhN2t3eI5vY22tYhonBztZ
roXtzR5SIl6ungwhjknGavXNVZjjLPUrgJJmawfPWpWGQrU57tRiS7YAREMiuPKP
SrtzsfT8wCxOj6theemsLakJrefv2mZHMfyDjRXB4txMso4d6jhlZcOxX2x2PcHj
Jr+Vu2FhCLhL531RTczdbQbLDgVw6kTQ0FhLe40eKTKsS5l58elkC/1K638Apqi1
+ua1/09WZ22X85I8tKmI3Vee/bOVbMMEuKOo7DvUNzZhSpYRNQOgQ6rFmUlGylv2
WBJ3EfnwrOR1iMfzqBY1tkkaDv83w69yNKSn7orOzXpzK0ht4/BKbsACxtbC0a5G
JQg+xmw8BdXlvQ0NXHqvqXdw2BFWyNCm72A3Oh4GlpoeG+R7tWNGrWGhGm7V5N+d
JRsfF9qWTaf0XxVD0e2zdsrhsrGgp00LmOx1g29cVjj8/ukGQv+Zyogp+tozg/Ji
g8i1PU2TszCgHTFTlVEDMMdxBIZOeGdihOgrfnnX9Dz0/rBriTIGt+bcXHcpbdt7
TEjriXaBZcYYqAV3xpNBlUDiurFIfHXOtwjSqAEIU4ETkkr3qST1CDjEYpjBGyEs
psRgO9kH5quWgmbpTRZ0G11JiUP6G9un6wqORzIpNTBbt84lFT+e6CwJPbS9ijlg
yDlEC4VuMWBct6QdRqxnvOTAJT+l1YeMzYefbonfl+ddJKDNGilGou19AzcKB6/t
vAWftd5H9QjxUKrrpXQSmhhSS/ojtIEOGjtMxlTDaaRp8IOkcdVGCh2l3dOGZVaw
fU27kcHcs/j0G9xFfxTzsiIc55MPP1/jgqwjSDMi5qzZKdcr1Mms60VbknQnPjH6
5JEnoevTLQwwoKaywCU9mtJvLFq6GxxlKmYnw1dxAP/5NYLflZYMWGkO1Cg2Gxkm
dChVoCoEsWS2Qecyygl7CWsoN5AauzLaw6AA57RmFgJiK2ZRolHsk2+32H4oyWSX
YnMqA+ydCaD9fRtctvlfxKOYsig7uLf+xKFK+bRVuHazhWfdVqJFCCGfpWj0o4wl
Lti4ORr1EwhP8WESpF1a54qqrxlYE2Q9xiF+0upfTtWQ4CXQuq3qlRrrS7FDZhT7
e3pBPqVQRxmSe58CI3SuPM00zVECj7tqP0LG2FyBihsogXi4NIAASuou8EETaV3W
MNTcvc7NjxrIvfRWd5UwrA3gIGRUixayXCAseZZ5q0SQruZBWEdrSNvmY/hagDmh
cX90K4rwPugd5N98TGrzroi7S5J2oRnEm2ylRJnlYxfskgmSp+z0cM2FkyDjocG/
loip23bhyEqAYSzMPYqHipRWZLt/rdGRmxBka7GMmd/g6gjI6dMcFrwJXYENuP0Z
vXgLdVNMcogHXz4DHlesp6tfwQ5OGad0ZlfOXGrP3IFMVtwbuVq7Pj6D3GDpPZ9M
qxoEOjZiKHZo8qCafjwoH2l/8zKi2OR30LHaOrUWJZ2xrsLRKF3QEVAzHxaXqMoe
009bFl2lcfMVu2SRoX3Lidqhdm1v/B3UG/tS+QX8ZUzbkGkFWr6lfStYeD+Y0fFO
DmAAF3GjznwEUYavfjb0Y4Eze5dS8xB+OwN/Tl4bwto2HRutbQ5ETHFKRRgFtOBB
XdRv584SC+KsVQmpFsL7GzdTCgo5NzUK0HKNhticBXnOe4uuKBWKCEgtNPsTO75p
8P7iCgF8WZoMeRR/P3tjOxeZ7IIXGVkSwfJvXerc6cgUiPXTsVy2BSsuW4H+mEnz
G6sAJp6q9lROI/ydyFPYpzkRO9+y5LPP9Tca1zALCwJvKH761i3N4gZUbaE9Gh4B
KGg40Qz7WuUUUMQLOnrkiZ6aCrwGkOOv4z/IilNyZJhHRy7/g7yITpuwNaNj0CYv
rdl2mXd+5NCozd+HHzIBmZpBubA0M5UKwkGnGRZXG7wtU5+UMndsIX9LD8Lh344u
5I60fdGt0ts71Dlat8GUcv7MbDEHHPtgl6kEbDeNn23N05IikGhkcTFw91mXaIA0
TaplImyVB8s/9kte65LijKk4oqfpN/JMngC5POrrNmxCsCPCww3u9mP6DNWXF4yG
wnAEilWvjubHi347vG3YBgXRuvu0jk5tMBE4kz9IwhjPoPsBx+YBoYGLe82lZo0u
GYl7h8lbNIb0xKUeZArUFkF13bHCnEqGT13yXiBZnMJ/gxAapeGwA87B/GORl/Wt
ZPllRaYtzUDGEYH40s56+WRmwqlynJdYNl/lOjPs/2gigCnzmQmkj/U73VkiLwp2
8d/LToCaQNnL/KTq3ezAXaYnwsJGevvKtChLSWL1QnOFxURZum8G+3UVRIH268U4
YSQyk5GdGomBZL5OzGEpTBOfy9/l+lnQC+GHIVU/e27yq8mZS071rpOWiwX8rd5e
N3F43G+TmeWuL+fAmCRH4DYsVuQUVmnGpXeaXdx+aA2BTaIJ6GJCKMmAocdh+bDP
6XJn9r0Bb3GCknfUN+fJDsWHR1pFxtOBRxfSFMyvhsgl7MJwxmQIkiCHXRtYgene
MiMKo0JZInwqQQaul8mkcYEKqw/XLPcCvZmBa/LpLciP31hDod1Qjtng8UBMk4IF
21r8Y46DMSlyDzT7UPoEvrAbsRIl5nqQ1Cw7eX0v8v919Yn4HPMWliT+uE9QlmNg
zK1vlKBtrGcKRtjQO83TDX70snnjHNTCKCEmktu/euzGzWUhvV2P6oHDuWVCzlKg
kl0DP2nIBjNc9aA+uBXhgIu5HLmBGZMrSWbfKUXgrmJBGLpl818j09s1jbS5LRcd
bWX71vCKScqHK9Mpv8SWbw==
`protect END_PROTECTED