-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PlY5qvDf7xOIGENqRehRDZeslWESHY9m/OP8h34jii/e10kGvL0kKGNOSLjGZH+fxp4WV9QSu7IE
Tt6EVWf3Hx4AB5PDIPrhV9J9aJSQs2VKyygOVYNBfh6BK5aVzSd2QLljpwPoM2g0BCwmKDiMOlLt
kkRyfueoOUneA9yTHNiZ5AIZcghRjDOg7W41KYY2nq50kEpTF2pnJfipFH7Jht/KwiKTdFhnKzUm
D/ifvxiQFOoTgwyrlBorg4y8PMb2r3fI4TPitLCi/et+VAEmjO25+nKQ1dr5H1IdxGda7P44jOC+
v69CHUDoPpDcBNkNcofl9NwIo1pd6gu3DnSD1Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6896)
`protect data_block
5XCrnjJLOm3E2eAB3eMNp/zFpRoSuU71tCMR4hfQQDgD7M8Id/aIhx2VN+RD+SNO+ASb7Knfnlmj
MSDpoPjfZiIlNSPQx4XLDqKT9lJQvsmu+SAD1KXMiqrwluCiYpUTL5WezS1rDFd//L+KmpPAfsWE
g+k1gU34vkKkfMjjH3hJAIXi/iNWCjTpiST/F9YBjx2yYmjbSv7FMyf5pt/cft96qkBhCY8IZV3p
LEbqLN10OV4sYUN+lj7SHYWh8T884KYBy8KTIaF4kBi918bHgGuaoVkAmL74N94PLpJy35Piy4mX
l3hQKnj6pzg1HMYt2iqU96x6QMV3dVlny4f6JNlbxqOFqFIV2X+8c9hR4f3eEGYMXoOuoQAHV5Gh
yY9rwjPIYv5R5+TVh5ChqbRovnh39ffnMJm9OKfuX2/vbyLoheXpp1e+mtMS+KwcT+j3ZDZk9SIF
vuIqz5Ge4p+rcPuGCXZADi8hcpOjNQqct2Yy4hl14tPD3f0LS2XqscA1ESgF1wHwdB5CtpPQnHN7
Pe6i7UfPzSxqMm+eKWZ7wmCoPjDooHlrtPcZJ5GZN9y7AKyC2JGBFJWxaHLS1btB0cQz+EDnZ1DV
GpEhIXqXGj/zpdM4k57BiQ3zREqa9sdq2Z8O53iK6Z7qfN6742y4Zm7bXbWlBq17H1W74svGQpC9
3PPrTZp6psbnfR+UPNLjpGHUkyBRm+C3D0qfOzcNBetfW67QzMh+d/pokTqeZvM6EGltYekCSeRk
vcobDTnTuUu+CORImyWuMsLFx3f04ARRllGH2/3x7UKJ1HuusSucVrXtmpT4qaLRNF9dYbTFLLSp
h7n1po388IPYSIVumfoAo5rRir77F3QzcMQQee0wTmebsorOHn8jelKZRKfR6Eq9A7wIM0H0OQR6
zB2Cqz/6uGRJE9XxUMszuyAMvOnGQZR2MNbevmnxLNgwnBt2cty2dagAEolNygaWEALVl3DYjwM6
vVO8Ibh+mghglAANwlqC/QQIqroraVrwFUKp/IIF9s5XlgeMjCTMRvSZdDrxi8Ylbl/xmXVzwvkj
JIJRJiKFuMNAehbVejxnckv/OMryMfK6wq6lRqFR2LzdrlZWZho2nhY6gxbFHRzjr7Gf6/bRUo+l
9lFtjRoYrdHhZ3wdCtDGl6VEtqQ0ivRvvgG36ybTREJ3DiTRk7PdFs1kTcQ1uXxV436aiFIsJ742
0BwnKYFGpFrMy6RcVZ8KknoPdfmFudl1X1/t2rDoAtMnl15DS1/glcATj3/YWYvKrc8tZCCRw7mC
09KovMXUtTKA6X0m+iV4wweYij5kOFEclpUnPSjoKITKkC+Kcbei7X+XqKT+bkeUyw99uxVh/hOe
EtwnkFiaTUj7wkfiLY3/DzKAIP/Pb+MMQ9evyv/83nrWgq13gQVgSIjyB4DLErpQlS1JCqReaB+o
cbyLWUcmuGBjJuWv1uVctsA0J72g7IT2h/R5RY2pJE1jNTYpZa4kvYqh16fNyhYN5LGu0xWhpD2c
ySrNulmrYyqvS3uWJc0LaKFx9cdyYEdfKk9wZyR06cM4BiWFFHfbVuP6F5W/AtJ0vh7zKA1WfJOr
DWDbv1gbWkRsriQxWh4wC4Nsawdj1Xf7mG+4ucgsM+Dsvp3DZxrHknrQKKSzftQnbTngiHgaDk5D
BsdofBvitN8D8ke9Ui+Do2OR+cImXe6R/6S+RJiX4IvGOX2aZTfRjIQeMYv5bINFlVDUe+4sWOOn
VOGwTW4x4A79Sp/BvpLSwceP+Uv4cc8iodCGqB0uVIwdk2tHEmb8Vd1W39DG9D1bZqhL6B3wn+A1
qm7QBeAnTZZG9Gq27iSdYqlA7DQ0lhsQcAmiPopYU44JeKvz+JwSXzkGL3IzJu2Et7oLaCfdZikZ
BMXhZRB7NduPub3NCOrHZRVWNdxKSP4vIZSxK8C4jRKUKziwQpKdDrH0f57Phd3mcRMyxYZtbxwJ
/fybED63zVM1QKp0mkZIiXKda2/PCdMtSFRfBw8gnakpg1TZD6dUkdJ8GamcTCLcYUuVG56YscIN
Uer9DR0sNx6jXxKOGQMdcTeVTRmAvt8uPsx9LgJKkbvZqh62RD7BMuXb/WrYEMoIhew8GhPIIKex
beVU/itHx0Z+Bh2LT/HTGIXqdqkbrcp6n3fNAI/OA5LBPPdMFTHbIxBtZiNDFlDv2bOZSlHHjRd1
68h/AtNnU1NG+W5UcBg4yyCAdwcXPJmKjsKIVZA6STBBpOCdyJbUOWEcu8b+NH/Xg+8YwQdrnWcO
rMJQqKJI1newXlI87pNZ6yG1LP48qj6balQetEwu2QDpJf/VXg5LSxWixdV2xAeASk4bUwiFYvJT
sb5FMJmmJZOqJfhAosDaTpJG2R/lrbB7NVMbmMsqasYr7w9EizbKzsAs76biXi9Thn29vYWYgJXi
OObLXNcqI5Ys8cri4YwhuTVTEYxl0UtU+zOTgQHesntKshO8bMHIA17HH4cnENaomJqu2oUibCTk
wwE2z+9dNxw5PZG7xhGoPEu5fJ2/xCkAlzd154NtEyWzG/pURM+s0pYYJa5Wr0x/MOiqRf3F8aJW
fJp7d38yNoYOJW7KC98KP6NgeUBk1p+tRt4jy25PzLU6qqg3I+6lP+84CT8/YcjuM75FF3kxVr1q
IeA5wk5takdaMfUl4jU1b3IpV6Lo5OdjC1S1OPXTZ68y1oh9UI37YR2s7jgsC86eEAO2hJqUEoiv
zbnzM52t72pOthr2d59OiA9FxcswC2Ifn6lJU91WphNQ29EUMoPvz/KU9Tyapkn3iMb8ZSm3c5/G
VbI86irWGWPN7W65+ciV/YPjLsmTaxALg1VH+IZuMD3A2tYIH6TPphwLIa3k/1irL07W0h6xwoHg
WEb57DSRkVG1rXTNsKcvRvYsC9IjlzHOaaY+ZCri4T5RRJ38Wn/Sxg0gf5bv7PLfw5IG2yc+IZfQ
wKimqOw/KBA/bcZGBCdC32hcLM4F6maz+eVToXkgDw1GzF0aewO7Kbnc1tjmkLHXcXNgAM+e3ZM+
JJdMsGqT2TPlnOjCY2DIxQGVIPNCYivB1oT3kqhSMUt50ySNr8O7MGAi1rVTqmVWI6GqsFSv3j/y
Hge/Vnoo7ezhxfQnjdqsHvJm0q++Xbb/NbrtwovU6+EGMRRoFFwkzs9bi4Kqd3Ay0FqOpfasI8Er
HwkDVJHG6paHWCNY11RchgRaIHbKdagO7p8cXpVumABLa89nFjoxQhFUwNz7BewjI9AbHKP5pp7D
JLBgvezVdGmuUfipC+ZRXmpAKZk0OTK6bRR1suOLsCWu1ASjYHgEJ2Mnbxe64DNMRBHyd9Ar/r4X
HYa+XNGNFs1gSPPpD1GUWI/4kXmZkmcLg75am/GFRi5qq9B/PDwygZiF32C26Ub66F4hOiCC7f4c
h7IRJcmr3Ve53Jrt4Qhll7V2rFjkEPAyVEVLtuXNcRbPTOonQigrWObis8LQuFiudhMxSwHZg8TJ
bF5NuKfx9U/dk8jV4g3mZNogvuzU1LvJZ3f0CF0iiycDPNtxrJ9uGCD2Vw2eOMzzyp5DgGsM9hJn
Z3ClOFLQAw/Jm5yTVPJCRPKiYWKZsX7JSPFdvjy08XNPJu9toTXYTAabW5ynVc8gOadp0gNJo7fl
BHFxg0+6oEu2UFGvIhQr+oHbIKx3/cSzVEFEFkU9DjrCAhoAtUxgLwWFkZZX1Ol8HRJhP59bKhoP
RsIcOEKR9bRHNFltaD5gMxwTMQ4ZzyOUuoZAuOL7y3sgMaNXat+gVXc0HqkYkElEulDPBkBBmJad
1wSvvyDIHsyxA+NHAOBdMCw9g+7elQL0NLSJ/cWGOdYYYAa/b9hYeqEu0+0xsho7KSlUAv5DnjK+
yRLsz54Vh3LHrquWpWK6Ggu0aBVLZMnD6vaa6f9xWsTKdRV5hfoVbBEZuJWIfc79ovcr9QSDdD9M
tQD1HyN3Dl6sHX+oRS170KLPyf9KhPJ3z2NGLEXtlxbWZo1g9Adg0jOr2qDsjf/OMMvVlUdUAOrr
xkz/jATA3RjPvlXxT+K763HcP68kymyLkalDQgKNESKOp5QtdlwRSuM1LYG2Nf10JIm0Ms/LsScF
RU8qejC+I0DpDsFDqJYsZUm1IFXUZlCbKdp2BAlF1A9ckrrUq8dDV1c9Q6FvBb/cSxKAgcVI56F6
R1bs9b8zuwMB5KVr5Pf7+inCarkO+F0XI0n6sd166Bw8GxEZPYuBrasLZQDfKPy13QU9bxAYcGHr
zrKvSu2wu1Ek513yYF5emhOfg/BR3db1m+xvIqwusX3r8jSSZMna0dbQ0Lkb+0ToG8IvsNRSsa8G
GMMXEkkA7uxm6j0yd07uTNEr5h8YJQHs9G4h0pWKyaHE5rmn+UJ7D4tuAPhKyVJa64OK1agHsAr3
oQdigptxWB9B3uNZIZYHDvdCWRl1OhzfaAlT9CoMAa4k+9CFmOr6bOIcrtmmOEWaZ/EGXO1bBPvU
wgT3K/uGlz1UtALczvYbXq680TH4V/XmLOzS3Ib3tR4u3o1XST7K08q10LzScthcHX2Sg39uzmaZ
2nYGqRcH6HNvoN1ecyITTehkBO6Py0TKPI/Q1eB7jWuptkn0KluD9Iwp9ooqNJF8lETqRnksvuLt
bvIXbimi1lA6wAdXLr6BhTTvzvIFagJp92Y+AhBshFDPxnV6fNXjKdvC989CAUQlNwU593cLd+rW
q4sDamofHQKL7qoTG/O6BLCHuwXxte3lXo081vS1Sw7u315/B54duGQkolQFskjGE2C/+fYzXe+E
1MNsv748nrhAZ3boCe0C42ivZSw3qwcpagkjeVXZ3yp9obnvRcsk2Ke0/2KZ4Yk1AYRpApdedxNZ
0+GQ85nKCAo0z/TM6lEgpTgtZq/K9VOl/32en7o3vXtFdqVr5YXpLm3NgZFZA0bAKEswOWEvblJb
2xIjFjUjPuOP4sG5FL6THCSgU9ylBtORCpQ72pZeIV3/UI5aXwcSsKBjEnT8o3shcYDjm4nBSBti
t7fn5uitptH7gsQ6RSjP/fvgwfr+UcM/KAuk8XgEjNqdq8h2PckbcdYHzCZGaC0R992ii79P+O9/
A6vxi/2rQnGbEllj/L4h+BvPxt56OLW7ETWpkvy1stMtw4klB3eRn5Nelt1VmWhAphe7xqTTrBdG
6ILZGjAaA+O983+H8bPY/UKAtau88XNR+RD8EeFhZZ3YSPqvjwx/Qn8TkFxv7KKEiFIlIcqMCH+d
BgO55eRmSEFlhyOkZIn4uxq+rxZg4C5J4UlEG64H8fjD4xLm86Ss5Z9WcDQY12bhbBpkxEfC418O
sIOGa9FpQkScT6BNt/HFtD1xPI5GI+09hnHgBCNuPGdHkFiZWDbvyJIMvdooZ8qeyU/9vJZZfP+c
opraBtSD7UW/0w/TphmQaCpqqjELOupdlZpinA8fAtKeiZOsE2inULtyoMZdKII3pQrC8q9T/s2N
JpmyLElOVHjDGqqU2xb3YcQ7pPNp8HSlZp1uuwStCQ4iHlesT40dH9soTTQOSn7EkLZeKZc+n3vF
lD/36dVuqUPe/vZ0ndp0GxrsRE4pLAczV+PKglDKZcESFCO0d/r9PdKzaJuVemdEyJWK7Um4VThj
ot2Es4aU1mHWqs04GVZTW3JwihrUtCzpscXJVHmDwNHjproaHnQ3L3g1gE3cSSGXo8LLS9Yswj0T
rBIkf6hi5fJYiYW11eiirvvz6NDLq+0ipSeIP8oifBmG2y+o3Xezh4kg+AFpa/UFjZynI/4B0OGN
fvXcP2pGiW3OZOnWyZ6U3M6zor/4XEflM4Kqf19scVY3zl1fUORp+IhVzVGQZpDd+eUARRYUFJIC
Wq0YsAOpDRudSMPUCaqx0sJd219eBVUXM4vRbccqRqRthCBS/1ds/A5e/KPEJEK+sKEgcG2kPcyE
HryTT1ihJur0U5KtULPNgLhqpWJqv2qw85rAaF7WEwW5CWV9PY2aLwPE24OG5fQfri3jlxy/oSgg
GeW1be9m3/OpdurvWSRieO6BuS5x2mT/ENJIaKLjzuYorokmN/1ndjADNlqjyig5VJCq9R7hW4jU
0BBUmXGnaz5bah3Cd7V2AJcWh0HcdOvYvXAXQhwpl1I4weleluZKqR7jIDZuIw/pfKoEgqvykiHF
LLyM4kjuF12zaepstGViHKImDHWVRAw3TBplSUzaSpc6zPR1zAH5DNKEYVljg1Z4f2Il/+mVnXsX
2BQsRKOh1cb28ulInWNHbAtsVcVF9W4mrwVXdUjj9tus7/OeJFLMA0hWYNP+gHPEY9VvrPTwox87
FRuC6zAAzklczfTh0F9RfJfhd3wOtOw44GIr3uYYKZeUJFMm3QzHRvCo5o5eQpCbTF9f9vD9rTRF
LtAicXsuBnchUbjnxpDGG+cxLomUz+FMT2aQI+SS8N8PZ4L2e24Vg+gmq3AOUljAHnt1fYt39HVE
1yAbC3GQYTf/KyhR3iU4eJY0B2bMc7mjQNPGsWslF6dcArL2C0MK6zxHPWyBGwBlwSs32vukYQ1I
We9sXy5/v/Ghp1IgDjHt6wlYUTssO0Eo+bYtuORZWZ8gwDIw1PXbUBYf0X1pXUdV4YIXSXZxVqtH
rs2E4dpVvacj5TrSv+1BCh+pl5gtJFFwchKeBz+YTqJ34tf4CfqB3cYlkjGxu6rXg7uVjO0XiX9l
wCZlsXcDB+8jNVbCyPbhQSzdiq7GT9qTRyvMlj2xJZJDC2GSbsX+c6vglrvH8LyN3XOCB3gWlaA2
+d8QB9Jf1BKQt18NTk0qa/GHpIki38GYo1JlkK+/XcG3V3FSGyt+PddtzBUI4Q33K33WiUdaAxnC
x1hUT/ecKuCqK3AF7JgP4VCJA9n66f3bR6Aro89PVfY+zx2MMcZixdDk0P5aCs+Cw3UFRlq4CsQ9
XamVN3FLy1MVqfMfVy4uZAxuWAzuVm0mHHIVUY9gZtDlpFtXNdmJKF+mtEMTPPEDmmoXBdCuq1Vr
zI7zSNSQ4hZMqnlmN550rp1yr5IWrx5NYVPaaoWXRYX114PhBoFVNe/ltP2D2S+GWDEeJZ4bXeCi
XRihMkjrOfIcxhCzcx9dTaycyxRh+QeHkgAtgv/SO7cIwHfdoyBgA+6my3Wu+MUce396baFn1cUj
b/OxMc5ezA8LHD376gKRwv8LHyHHMx4CJUo8NdMmUC8QjVkNvqtHyUF53DgvzV0VneyP2nS3Emrm
RYW5DC8MaCoyGQVNyp8Iak+MhGPtp2gC+ANnUZyz4bwgFLFCjEiCLCfyl2K11wQK5sHls0S/16Be
fodJJAHoNfh+9CWbVoG1/9LpNHFceX3yY+uz9/vSAYJS61rMKBgWfogZg4C5KgoPPOvjqXrG0yHi
vklHvMJR9eNjAKGYE7s9UUFDyt1MJfh25Ul1/vRF5cPiS+Dfin2r2I9NkDoLp+l2cb/D8ltKgC+2
vq8aoLOAyLnnMLk1lyXc4qBZroFCUsD5g0VANn5rk0ogzCREMrbW97Ff4Pm6VXqzNYb2wR49RbNT
17bOkdKE8LHvA//PA4/lxPa4hYSE5ph3wGdKDhg4sFk07YBK2FewFMS2NW/bXY67B6/wXFK65y4d
2pzfuWxD6ljOITMTuTh3iOALrR22pKsyl6LntbSSv16g6pKIHfnx9pGN7j1OHov9S6NigGcDHKUk
ym4FfljUrf+AocXaqDAFDP2VQmgjPFldbdi/d55FtvggNYnqjaGIIim7prSLprsmVLJFA4nfy8z/
Ge+HumrTGW9X8eJY+eOhvZt6L1/ySwKtWQ5AM7/MMNkEIPlqXTiRW46XB1y5vKI5VFkYgd2owNJr
Qs5MwQ2QWS7MzhoXNVFfAr98KdWhTXZQ/jCAqj7+Hufi+o3UTJfgRL8ZqEkIgAKxkGunSZ9PZ8H4
7ui45t3YqllfKSWZeuLwhJO2iRvfTA7Vm6ptjxEExe1LFSBqG9Qcx66JalEkVbxkgbUWJ6h9j+o/
cznFIFrbwVwi0ssq6T/06Aq1VqHNO15ZeDlP6HjaUFLayIRk6KDWivqO+39Ese4D7NtrJst8wDxY
TMBtFhxv0RuToItdaMQjp+B9HL5bjOsrUv5926ZckQjPMzzEemosZ6gDTMNO86Kk28dlkAnRyZbC
1gFQVTRcaCpQ6ObWEQnMNCDoMl/I7SHQORw6DIkdrmSqE65bAk79Moo09WwHTgICwZpP3mOlOfK/
XYogqPzRsJ6sytjvLZKhq4ysyqc0w++iF62/7hjIDk+YRqJv3BxWRY39nfupB/vkYkpe1MZKwHpw
InaFxhJq6I64e6qndPu5OTbnL6j3TLqRHgfOwfoK8t16OT5rjRzVS+/tuKE5CbCQtFBznwUB1KCG
iqcW+GD8IhEAAz+SA8ApS7QombZ3KqBLdWrTMZG8284m8+M35rg6ejKPkcWdALuzIvO/IHLCEpsU
R59iA0/MAr1rwKlsiJHp3NQi/Pqf+/YJQlxcINU0rEVHd0H5llQKC2ercWMrLYZpxI2O5pS9nz+r
S/vq35tX7TK4Q5EyC8Znso+xdrwetv4kpM8ocBojbQBqWHU8uu+0Q22Pu7Lz240lm7EM2gwIkmUz
erhkqpoJUfLXhx/VYoqASXqjCF4nglW5EuIh+Sww8ErttZMeSg9+73A+movu6HfuzJKuICJtARct
yfnavOJxbwYu3GoQfdZOxy7Ksr7WO/fCNjnIvuaXD7AaD1gy/IozbYOFGQptwvlrqBxjdFU1LxRz
cBWjvZSW7GJkvpDQYhxgd5eAxu0sGFICp3ZinJL03Hnaqzm2r1uVXf3wLHnGcsxigXct923EV35D
EtuhNQeMvCAH4oMTfQpbgpjAawYzUUW3VaoZaAmQTAu2cHkHQIHhNzRsBGqiqZL/tmav2NscMqij
/QTRK3wlijIJ9SCnNP1dz6DBhuE5hY5HMN9tPDG7nLU2OlQY2wmsVPfIokqty8h9FZd3C0Y9l16N
47kQXk0ZRiP67Cfj1FDg6LZk7nXstYcrZgSQK+Ca/NhsQNWSoLOGkXV5iHRI0cLFBR5KJ+a1AwDx
rSjzMqxFWh7FkeLr++/rZIajqGPdLhAWiyszNHwX03e6GkbuIBPrtz8X7UhDESS6pVsnId+f9IVJ
w0vmUqb31IrchxIhSUxM7BNfRs0YweMoQp1pLELIgie0yhPjBReGfUkeRPecWpW43kygYD95JS8=
`protect end_protected
