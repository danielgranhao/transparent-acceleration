-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1G8cUbTfNme5S+HBQPeKmYJi61IeVLpcvMI7qMVcFGB7mw/+eoByn4XIMQPz5+rS
Hq5jHg/PjRpH4Td8bR54AdTxV0yR7fbT9//JNM8++QkhPHdLwDgafw6s/Tz6xdcc
WU2Uk2YcOl5FnIiBdoLtEaMgH401BhtDjaJ4+dYZZDo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 20096)
`protect data_block
KX/CUOhE/tiwyNGnfboPkZtjLE4A2Gh8QEcU7MEZgniwbqqyrK3hqWrgle/F+sgd
AtjCywEpiMKGc9u5atwLUnqOHyi0WvO69iFN/IabgeINhB0hR+5J0+dStb7jZf2L
KZ3knvbOsLy7ha8Yho8ezl1hM7knibqbOuWBE/RILQZ4/j43GVVS50QlzufIk/Zv
AF7tAecLInLIZCdFRpo/B+Sn4HD0MKI5nwGvwRu+QwSo5qvdHaaUiLfG7y0uNQyK
Fz+eXjDLuAgggVCdBUuEMBMk7c2xPPzNS15VFQ3TZsxrc+HkzDswJY2yAtPFCsYc
U1ZH3tI5ieiQIqhJhArsfp5KXoW5Qopvlj4jRmd5NmWwnG9P7215LRn90z13zsoh
rs4tgE76Ily3myqk4QkyAcM0oijbqlhbHWrqj1mpb1VzdlHZsg5LRVQdwTLB7eQ5
6uzyBtqaP27iueZELutHAB2D9NPcfnHSAb+gBoRt6gDaIbr6S1ChtEt0S6GsVmDi
8lj9rpp3YHEAheQ0ivHfqPYSvD2utIBKVm6U/2m9zza0D/bBuFn3rkS1mc6W5oA6
UcHSi8JVnOz4Gd1RQgXcIqCXzBGR2E7fACzIvCfIoSjAshRbFMkSleC8V1mKk/R6
pgKA+yWTIdiR0yHsA44wGEE3qosfpJaN+wDSj8zcFS6CDXinqdHItdvh7G7iqyxc
qggRSDN/nOwT+Hnk6WqONIZyKOHK8yQiHnwUi2eKAThCTwe1Yq1P4BXT0r3AxE9/
2qeSpIJhk/uPkHmuubwXXO8GBaYuTLJH6cJeBShuTNSBAi39IxVIachQKloCfV1H
qGQ3WBUY+1Chptl+NETPgJSx9Emj2RVa2sINRSxbg2L9gg/13Bl64txvjASWdGG0
SqWxE9V3Zmev6cvIr+9JiMrsbpYmoyRq47p6r89WseXiZJ/GWD3JWbUVyMPm/IxP
9cnbSSXAd4CCR8SatFEJ/9flsjYLWSWJd/ZWtSk9zhFVAwLBzBkwiKNL0eOkU8En
SG2yOFsid0TqY6hY3pF1FxYOhq+x3qaXo55elb8Lvo3ff60Kxe27T2AGGbStR/Gf
WmQKz8Hp101sAb+aNMpshcZ433nu8dc2yBO6DOf43GC5rehk3clS2gsM/Cptb5/t
0kcQ/475yZKRbuzaSkcDL9IFOtq3i+79Zv4sB3JP3uLPWQBuffxhKCf+ntSOATRA
+m4yq/2IsgMg1zjanAQxM5AjN+WmNW6MczVZlmB6f6y7/fNnClGMzKlVw028KwMU
0kPF7dxqvBewyIDAHcm4mXSJgKL8KGX+xU8clljC7wefwxz33ym1DMd2LN4+P3TX
56HajvwcMLj75fcdHV3grw04p1jjFT6E/XKoh1y0/37SwjOdiX+TNdHaIv98WxMW
j288DMkYgM7t/F3km7UhwYnGyIuywSG34bmwhgvqti8N/6S/aX8ai6wpD+74sT+g
BVclft+8jRRIIVWzqtzuVx0ONPpUiRE7n6qy8l2eVj2fALb9xUtxb7DcuzIRe8T0
HYWRrVOoOIjWhDMW16PhNiM1LW5TTJox7CQPXvNEVrbzALiGAJaOClp35Yx/+8nz
7xNdc/JS/W5nghK4O8RmH76PuBM37PN5KxbTTfy8w239RVnUuguO0ZTQ14prS1v3
m5UCMPTt5fJEIhC/vIHudcMB64vpeCb0r9YT23gyKzC4sih1/58RuPnoCkR3iImh
eW79J23p3RRIWQum+0GKq2rI0HbZVhh99rZyidCCCc3NCHlmOWEtPzMmiguT/rDS
iYKHBbVpKj6Ew8kcGJjDikfOTbWSVQj1Z9UhaoBY0UjzcTNmg9AlIuk53HzvfALk
p86rzS9xdSTuBJCv8D17ARt/JX7YoIzl13jbqxTbcln2A/nYpn7sBvkqeUbsPRij
UzSiuzK00lZcgnJkI1kEhm2PyX8eneh8KYk5SBQN7SDXDhglL+0MzGjBpn9dysjW
mrBnHVpHP2O1F3Yp8UW2c958CTc1MsOtVTmMpwy566rKSF3bAsrATk5V8cVBfZ9y
CIQrmsjSyDUBcnmROXbD88kW5rtJGRBFPnRng5MMEq6jMKkfIrQ3T5Ru0N3yMLzA
pVv0HfaIFfEabypDqubsriU89GN0iJBk/GacDENKiGpiX/Gy3ys0YajXA5iZNwxR
BtG1EgRsn2YJ+aKrgX9tEistxSTscmWSvYx2qaL1GAI2AQ2SIUdUbiZd5ccxkErC
JSQLNiOdGNzw/SUD14UcXm25NZOCvvPxf/EbLGjHfEKbgbN17DwN9A25fl5lZ4J4
hKyADuFY4LA5eGjQau5cG/thldvNN0zWVeUsJbBYltCWr4Q7kv+yWFbavHM3k2YA
P5HdaFLSwP2yv893RiQYrGOmeowILe7vGONjf/PWbraHe6Daa/p7wrh38U9fDXuq
YrrXTw82ieLId7f9MGJiRNUktnfwdlD3jgt2+mo7cX+4+oeAVtRiJS2/5P3eNPko
hC6qBC8vlXJW7l6o5h4tZXhE26NlZtxz1UswTLTptwJoSxOJ573wN+PheW7rJnzr
EkbiIEkHeSdocmzPsbfnBOfKEMgs7R0A8xE3iXFOYMLJIwiv02i2tRF3zg4Vuv3V
FWsAPaueBUxOry0qVp0bvyYSxQuZ1FPITLrsIzlMRZrMd44+rUf4UpJlNFtot+sh
geHdR2W0hZ2XpkxdL2Io9o5yp3cOEyXvdqk+JQGX4ilGIKIu0bdiKwGJO7MLhraD
Ubzq8jyBlf5XePxNFGL06mV75blNJdh+pVw1LtEKou0C+oIE+tUO7GhoppmlbOPy
vTXPe2fOEd9QdXZfV1Hx+NVcg4YJSmwFeY3kQdYRWWOGxWHxqG0m4s21W1Ulxvs3
Zw8UmHm9eEdeubYmSa0OCn7L9tWRmB2ltOprF1QcZ8wJFyPR5P76sgh16wfOkMw5
v5Lay31A/z1Zhg4M8vRhdCY2s9FzrtyfmEyfuG6QTb4sOZQ9QJurLQ2oa3D166UP
sYWd9UGL8aAgApFpnZoFDqqqxC6spPX4CcG9KQGe41IOJYbvRT2t6muiqQNQgaP2
ak5TPQAU/EEH2JxGlKKlt33a5swrbONQ7MyNZWCI2kEXNsXGdCyQ2YrcXQmglwRZ
KWultf77fcszql5xNpASdoEDApBnlGGcmcyAGnhe3VjkH4CnG23hLrRbjSv+eFPj
da0sTL3lTy7JNJCatdj26occlqWgs9O1C4rdySNTdzQokhFch8vHH8RCXNUOCX2Q
lnE8+1TwQbh66x9h9ddeL4V9PI2greh2T0dOhDVOfQPPmUenDbynBBOMAt1pzywG
2ySeAaECEBbs4l5kNtcCMY8NHk3igt2F3IQQwd/a67mmoC9t5BQPhsdnkuCODXX/
CumkDjiZz/aFEa/dGOi89uZQUmmzv5wpDrnmfv3bT48N6/sjqBTmGBqRUrWUbrC9
xLNwp9g0hqxO8eirDVIXphpCauqGKAtLE77sjNXiY/BVKBC3VPSBNqRKTglQIQRt
8XA0xm5iPpXY6Gx8QkfiA3Lc9p95/zou5gk2ahofFlBrAGJN+Tjd1+GVoxJa3uDm
rqhUWw2xRfP6QItyT5QCu+yncBZrOiOsRwgrgmdQ42CNN62SjNORdLJpom83KaxB
MG11jfe70m0UkKCPIDbhjUK5zLexB/v2ela4FkB9CcavkTmki13fPQXzvIe57yBg
PIACSgmfsn4JiPJ9Z3UJbCpq7trPU34Yb5PeQXpbynXncNWeUUaGI4ZvyLxthlOe
TuxcgWQ1JPI+h5y7jEFBJw2qsHVWQgkw/YO+1WCOYaXz5R2jcZ3lzlrhLCA6M+/P
2WuPEHy+9vN3p5RZoFky11tZVERQvWNc7zdjjcgWoC49G2NC/tKXlBD/J6foqJXj
I0NqieAZ2RxL2XEzwf7z3jLRGrCSkGoxTodpp+U26SfOYmgy0SRp4PCmvnMHfFat
zvDpmTMpG93CXRA49EqiA4bAXuXIOFy6DAf0+wFioBUgvRpFohZICf4svwyfYCBA
vwUZ5yjtAotWkvG9nNSTll/oNG4pPd9fYq1urk4K5320sISmZ6ExaHK09zhNyTUG
U5hSW/RNeqgO8PwPeqje6cvytPOqrIPmSDrkE3djVZE027sqe3y1cybeorALuhTA
JYQNecoBrvp36Lj1IivLZvNVOyhuxqqbkr0RyMdtd4RWpvLaMqBSdxiwaX4/rquJ
3NWjUKZF1qpb36CAhhZOtTf7m4aYF7l7ZrxOzgW6GrR5vZ3I8T6AFwmoQK8yp+mE
d1isW5HE94hEk8r6UQ97GLjXUT26tMCh2r9ywcpOcrBm8D2eztkS6lEOCicGvtHq
mvgvSI9rThcMotelcggVQNt4ME2sE9HblqC4n8PzlMi7II0fP2o3ABWF/QMlDEYi
xVu4f00Sgvx69ssv/pamg7dsVx5bwe4q1llRJafDeG/DrDAAf3S6zwHj3/jhKfpP
6dWTdW7cbhwkPfjuPTw0cOCc+kWfOr8f7N/gI8p7XEddKUyRXqZW4dBzYVeTkHhu
+21tHX24NeozjXGLhhjRdhewbEVpKLotpx2oQr4Iun6yl26EX5tiK/EmUJOBgMpq
Zsz70MZLxyiJvtaaisixgcNQJ8xpMY7G0jHMUNynv+l0TQ9QJAwYLXNge3bC1z0G
rRKzYhAJ0cq6kDsuWznQncnsaT0dR5kIslhGKFZ/LnttURzSi0Qh/6EV0FMG/xGl
bUtRaO5pJzVqKuOzUMGOfg69L1i6jba6VVsCjfH4y2TBf7eFaUxWjA9Wh2ddTBKh
k4KBCvdkxr8EpLL7mT9anztb80VIHuK33pO1RvwA3xBIEAfQ+8SuRbN7tnWRN6Yt
vpBaiwmlSYpErOi/ACxEwj6FbTvVf/x9fkz6bdg4prcy0ILWKPUbpf3iV90uWAu0
Fd2/bx9j74cXEi5CbZpTZ2qY6sRIbhZgkgLdkImzFNMNDfYTarKw9Q82SYZ4Z0UW
/mzJuH/1d4ehkjCJ88zrT2f2Aq3/EcfwrAnZnKrals3yFq1u1vrLrJjeXOAljoLh
M2nHhSeyBH5DLcxp4DDuXW4wjcVSNanOfe1JRbiCrw995EwTSwUDm3ftQPL0Exra
lSf4xTQ/MTdYM8shhnhgSKBmbRNXZIdLKiB3r2qUmwO7HfksKEUIIuDRJ8s6ZTUk
LwQqGS6lKBzcBUq4FqAE4fUPdp2iRd8+keiV89WjrblkjuYqZMe1+45ECMAkxeLI
TWpxwn0vN1hCJ4ieDeLZ7p7cJ9FohoxW0wjSwHgqXv3SFzsbFGSpkBBa1SLQm80T
Vp+CG4SBuZltANFoPYtjRYqMjcJq/bfAQvZT84HRycCf37JUToNyn+fR/58urequ
f1QM1d51D+OX3lajeLVcHMGnotV7ClFNNTBVjM77RvwIv96Lbmv3gHvmGUs7Eb/D
nPS/OprBLEewKWGlGbPrY0JKtsBGemgwY/RajmoQupgr0UzhiISVadmLZ6z9ig6c
CQ7ZLbYzzxAP2GLup39bX5XLx5zApI1UqX/8Xq6/JuQcTCV2OAvf0KT2zPCoGi49
qdOH9VuZLnoea12OUlB9WuDmFh1zutNvanFw6zfB84cdWlz0ubPVHlChm6lHeEqh
Q9WmPw2yNUE/zssS7pSYzniavqXiGSup7+8PAb7GAUWBiwfxhT16YWxQP4auikNK
RVEkXs2RNEswvGtRuhzNHcZua64WA1K5o6cmc9vU2pTkimUcT1meNfubvdQh3B6c
7ZTYwJ6101seFbUv2ynun4FIGWTbOMunF9xnM02+mZTZsSd22dvG/uVdo6Vd88QV
HBt6xOE3m7NKy+vUrj/jG5TyhmnO/8sjBzupbZZJiHzCchFLOoL6G9USk6HB2Flt
ewvBBcyhpnm5WSa0EQWCbqAlEYgoPAgbXrtU5VmhrQQ6WCfHw4Wb7kI0twyBRUvW
9WwSo1+lseuAR088AGnSrkIYPPFXonOJdcSa5gnPemokpUmHf//qmQBuF2H6bsjF
QNYMJQiCj6ECLYwlydCql4j9kuvJQrH6J1FI7EIxAdoXeqP640ySnPRZ9jx14DYj
UiB7OWrmtciQjLfiRY/XfgP8xRdBXkCGGwS6mnWccWujE2nAp4Gxer8Li6/+V0Uc
ZRf1vckr3ZXOK0P+uCMc36muRo3fQ4s0V7hexJ/u9AKRmdCkzpgGQ6L8re1sMd7+
0XmGF3FO0ocxMNHhCKmql6V/qkBr6Bn3XwxR0RYaGLb+opRjoEhr8a3KR4LOvMGO
RGqssq37aE6GQ6BFW6ew30841LKlm7IKwG4UtBwHhX3cD7A1JyxQQu6eiHlCQESI
AbFW7pHbXqip73VhxGhH0F/4B5xDpSWBScV6C5DfywQ46/7c6peW51YCpuQ11WDk
Jjg0nV8uguibHwIOmu6NjVMDtl/df9aut12K8jgyY7G8M0D2caNyT9oc4eTdOt0O
2mLZrq6qLt4267RPouF3/4lm2ChOz8y6BdFuaU3Dqwi5Bu3+m9lBotsZjgmYDsm4
ADcs9HSRB0JF0GyZ8wPy3Sw/ZZTqaJ0b2zXVy2CAWNLy6Bg55/CcnsgHc4T9zc7c
z406ktfJcG02OBMAMVYDjNDGvDtBRKd2Cg/w9zN7977EhlUCYEw0AsQaJpw4Vn5U
McdL7XAxwdmZyOTle75GBjY7vPsi0jBLT3dG6Sp263X0MXbCLI0Oi4ANo1lcGkPu
oPlv7TFBG3SYVbN9N/7X3l6aR4MsUPNnfZjkb9GB07pD5BOOcDGkk9NQcx+OYFHZ
2apdL/QdcKqrjoBWoHxuMiAIWD8eP6EGj78yhXHP0iZoJul8BRJj1fneRnrXZjOk
TE9hMbFtjX8N+GHf+O8Ax3ppx/kaSog/CMD61QdV1oFtwRnhDJERnI6JewxiiXZ9
rOAYfyOi3+sRw27J9VAp71NO5QNpz5+WbJPoW6Y0hhgBm4sjeQ40pwUFpEpqjQ3+
HYCAO/2qMJU1BJ/nHPoCAk+QVOMF8aoRyAHxYOgMGd4wHc5FB8kfna2QxduRyWdh
NKTC4yucMiCe08GDxIlRVYVcbpQRUwbKfKOBbOszTsNjPtWAKrXsIqMBKzKqtZsC
OzNF1qa4Zas1L9OnBPhsPRAQO5TeL6issJiqXwmqQD1+b88DSHpi2rMBDcXe5mwd
7r31sR3N1EYUerfSCI8bz6U2rcPn70eHi5Co4NJ3oEawnUyUBa4PgIboY9FHi0Xj
iqp84tTrlA226lIPjXUPAZcHAWJ5Q1R0LB7EJcYfni1llIz/SRBJdY7RbtMTVu1N
lauP3FteohfN8icEYFv9dlTnhex5uCGTuwEWqYIvOPKyGTo/g/TqerPb0Dbz/W/0
FpzG0AM5hFLgSQcIZr4nWJXKmyejgp9kFrUSne2ydDZRAZtkUP/iC4bIMVScROjj
kwPmsm8ibGz7MMBzn/Q8UiGUTUvgF42KjAJJ1yyL4BR2Akm8fN+CV8zH/AoL/f3a
3WWPX1weDKpzc5FECSVMHJbn2Tn8tWUXsB9eYt1dAiAMEyByY+xeb/EkkIm0U3ld
obiihkkcuM8Qmlu6Dt6r7dSAxCtTUDWrbBPnKsXUT5yQh31paKcy84knklBiyddc
eBCRiWoYIXyRnYZhHgdir+Zlik+5eIMBmqoOjGLK3L0YDVJ7/Bk3RMGyh9c4wmg/
11BfAs+0/HR23HgcS3Yto1q4Nhwq09DnyNEpfUNahCt/uOzWLsrvZngMYzj9zYb0
WATk2JdC+pDWJdxgVs5bZ6yGYTrey6Z/nRjrF/u60OmwDYq1qVWHZgIZ1oV1Iovh
t+d5TgZ7183BuighYRpU3s5HPoGMGo1DgBwmTrAKGJXcJaNQ9n3P/J9fsvqnqvb5
JJB6zIkp3uhC/0zrhN3znlsTVbIQcSTKMOrno+lIa1yiobEA3n0h8k3bj2QVHw5k
tyn5gpnkeNHzLZr7a83SEqMgJnR4IC/Q39bAt7afTEYwINpkBzjYZJR6UFHHm8eY
OFZwjae5XZcLJwagl+ggLmcGa13u8num97J9in4ORqTHKKgRd5h2xEwQtnE2nnpT
MOheNZZ3omKHtwxfTlo7VeuqPpgmQHX77ZUdD4YUwtB9xd++pcACBUB/s/R2krts
QjT5SpijnrXWpV0Vp4w3KmiL4utpjoMsRx2LPsGU7BOXwDmLoEuOQB+XklqYzmEe
yeETZVU2TQC2ltwRKESjqgFG+8lsm8Ji+0pRjo867kpRcfDki6mUrBOXwl8ohdB4
IuErAa3tHxXcPg7LUwssWpeI3z0RJjv72XJUASsBNQ+gK/BYFh7KpREUyr3HGlZY
B/dnTShJRzjsOPvJs/NZAVkSNncu2OualLo1CzeoNL3OehetX3u6S52YzuIA5ec2
ZlzbkRmUr5BPGpW8AgamCNGKrJ98nugYekBz0zMnu3RxmCQG9zqqdU7cQJWSlipd
xUqUlBV+FWaNiRRzjjiK9IsrEs5vjqYOfaRJUX/enwZFs8CPeo/jf+9J4KXe4n3b
kQjrIx5veLhaBFMMFHHCSC+njHuT9KIZgxxLMSam+ileNd5+Zuaj1hiqeM9jCm4J
7FTAuz/7/qSPUno6Q6R/dsIPCwwniQTlThoHKGL9wuArg/3M7KldaLr0m1ReDyqm
e0UYnFnJG6wk6Q7rnrPpbz2AxG4a046epkdIjQ4SnDOVp/PLG7YF3SJNjiuSxa/s
Q1KyKs2Ep77xH7M0Rb92aphIzK4cgtTHaftZnO5ijOkaqSa4uCe+Q/u/idtPTL0o
DUC60RTevMl5cL5If0SDOETvQkYa0X5/LxeT7MSVSW65A4iganzgcKLWVu5gvrL8
QZut2X5MTDjX6pNLMypx1TPwcDuWoA9JwPwwMLq0VASxmKqLC2KGh52VD7Y8m3/J
LBZBpdIfNv6QGR6yGZZkbv3MzqnkblVQ3rCxjq6CcuyHazoCqxBlQ/MTdQH/hw0A
2O7Ld5lGTE/K34ewWodQCRVzAYju0SirZAldAUn2RvKOk8esSvdbPntgPeUe7syi
RVU+I/hb7tyV6YkoKZuXpuZExEUA//zrpSE0YGXGYaw2ehbxbCiQqlZTuS/KaklC
4udt4wCy1575u4M1Qci8hJm4QdTVhI4saNuv93YoeCCy+fJE02af1X9ZJhpyKdAQ
AUwQ7Pyl3L/7AXvR2+DnT47wWmTIS93phypjw90XcgxsmgW6J+EX+Tr1ylygSPWu
sImXhCLa/kzGgkOYzKh5bM/odpf7HPGr+yyff6TY7kLm2mYL8FDTweIizxE+3MlT
06gwVkmbj0vYYZUSIy3gi36ksSdb80fvVrpH0StPLVKDQDX1b9rNtB1nPc6NcFnQ
9JY2V0U9nflleXwTLFiguPzbV0lI+0fvyz4aaLMGo3WqKLI0mY/IjTQSwHOzbpxz
hTzb3eQrs1tZ2X30Efeac6rIgIKH6+3C7PFxXhnMOdojTGqdKoEquPboDOa3PgyM
NPnkxvJDNywerNEeJrQH+qsNx+1dNZLT0I0AcAkgvzUb9Lw3bDxxMBlgU4aZbVr6
j3actb4lmOJoZny+p+UyO5J7KURtmELwWkqdse5oZ9HM4sb+QbM3HrTDdceqEvPQ
pqfqocm3Jx48SN+CMbU6IutmXJiJeLR+atC5+mPiqtCt/hzbmOCmYwYCtdSY/WNL
e/HDNQiP0XgsmI6xb7jPPsNS2tj3KsPdFV8rB6M3OaSvtoTADP9yjx9R3q9AKM8U
xpkUJtp2pPhx4plrx4ane1oLsN1I/jjYeyAZv4EIn1YW128S5i2u+GM4HbNSlbvr
/bMLmwE6uV+68SelF6/L+ZrSEZIHWTCktV6HRW9r+VGBJTu5Qra7eNq6Q+fYNmYi
r9oAXV8KlU2xV1Tdg9/PlsYaoKO2JZWeTo4kkoMsfyClpniwqH7PQLg8IfNymHG7
4DSuu4v3Hryl+RjP3zEQdQXpfwVyz0L5F2sGwCj1duPBK2KvEbSvXlI3TZ2JMkht
e7fwML86mklZGSxaoMGcrO9EAEqOj0LCjPJw7axzG/SAYDYshvGh2hwnPxPsozqy
Lsw8yESnIgb6HqD09DTgRh5ydRBSpSTRDtCZKU5kb2eRoLi+6DA1cFO8dXOYuInT
WYafQt9cfcF4y42cqQknO2w4/IMQSDDSs9vnQoWvfc27NApg6ea2pD2gOyMf8TjW
l9i96cuqzDUtAV6MzZUaB0PD4ohVKU/XNRbxaElVYBbD4H6uT3sXtIXhnQVcYROk
uUUwEDoCnNtD+oLfEZF/D3AfZBU/TXvNekKVdZleWLUemkLJ5wtKdOFK5tbM47+P
JRs6HM33hfHM7n4iXxZCdH7DRlezCtotHz8cu3RPyDau7wWPtt175aO84VTIl7Qo
BbBGBb7R3gVNl9bL74OXw0qyxJEazgWiBXzIx/AFKQVI11Buqj+pBG4+Vz27suej
fjzHRiFIdPNMscJF2+YD3jAZL7vJZ1b3lCA/dDjO7dMZDQezFyNCSPc/ZzLDIurs
TCT/yzX8mMMnPHvNVbp3ncKr3ad1sIWoVGW2ySDl6mASHEJVuPZsY/mS9t1ZW3xw
TAkk8k+pnB69/TzI94zd7kVvttC5XQ97UdAIeDNJzus8Sl2OHMoBcJMEAgYAnp15
/OEQ2W5feL8mNsSRL+4gU1za4sh9bk7gO/57ROsHLHBn7p4I4QNhCbOqeRW3WkMT
FS7k8TW3y5vjd9o471yBujclHHa2yDCNWdttSZtJJATbLPcDZ66epkktzEFXjd/A
ZisB9EywTiNGoaimNJ5iN2nz9I/7OEO08gJspDD4TMnwPl/4zMJKXK9RP99Qdi2V
LWy80nS81RTP+6gC2nRyCX3Giu8DRJnX5z+Jq5WaGi/xAfLVDxUfUps2i02BAyKh
B5aeFJ4gUDhbJEAO0ZKR5PLeXlMOuBq0tqSTlMMUUZMeh9tOqNCJmLIztD5c95qR
NB3FgMu9DrBz9aIN8Flr4ADn8wA/hJrhKfwrQGtvyD2ed04rj5Z/f1GNBNHC+VEQ
KLg/BZwVndQCKvZrx/ArJfW5/CYbX9LpeZuk0SsTYD4hl4JHjZMyyC8Qpm2m/pj0
fbboteCYN6CcVt2OavhVz7yHAei5RhbjC3GQYmu40OGREs4RNgohHd73TIGfrMak
74sOV+LNoLBLg4w47VzMWrPbTevrJeqQo6AMGUf06P5AFq/B7oT/48n56H7XvsA3
foDmYK/2fS8RXGJaKJGv0AccZXUT6Met2AejvQzRfmDDDXEgGcay9B5sK61i/DWU
1GRtiC1+rj8Pi3lGXcr+GzZrAKh4qyvzZKSvs9HL9pfsuSDfIQhzASDUKBrzwI00
Tae42NNWY8C8wkP6z/26GMnXPiJREiVQOT9YkvXzy4xahGFdPuny4rTq5lhqhp/Q
71/jPlNqFZd92n9x+Fd5S9RJ8UoyQNjW3iImMrCuaAJAMApZVwjbwSx75eybRmZM
DvjPQ2BPbzsDMox/7ccEdIgPDK/6J+SOWckcECEmdGJyJQycEb8OxcfS0yUhBW4l
j1/S+udrV+wTzQRCsyqdDNfFjB1NwVI74BkfP6D7HIaXyN+l7KNybA2C5XuohGXF
0snek8ubiYxuhBhziyyEzThcwf5nuCDW6plMSFFwAVxM9u/7hVmB4eyZI3rzywdq
AmO3MrMRFAD8XtfzWlEgyKcHLMeaHWMFWyhpDCzB4Gf9/coijVYABLwLAqdh3Nsm
KMb1LwRO9qREI+jbOkV3Y7Iwo2VeHeEbpNYTQW7SAhFnch4IEuSsD233H8qmTVYr
ej63nlZNvFeV7Ig84J4JjY7a7pJuhoin0wsBiyicwWJM99ImccnnXe4fVWcxjpTI
oPBpEdipzWL/vZMOD+t6UpdQMe0S89Pz7zOUKJhd4ppWsKW0nu/FBECfRlrp6O93
BmyUQijCL9kvzvBcKe96gliAeGr0vMa+l6RqgswLeb4bVLmY07N4FKLBgcoqjgWH
qhVQP+cbVxVBfZUtXs+aDibliiJHAIox0/nuRMJn469sDnMVgqDm6lI+uJlr/jxd
H5zhBpacRBTmuFQ3QXO8ljfkSDx9U1TUMGa3TgYTrFVDyCytjlIIr0AejHjqBMHI
B2+lgMEzuC/ZPGQmKyB/sbwSjlfoZPDXYk7hCngkiq1amhBKfGh63570gHzX4LyK
TQ0A76ih1ZGQ3bxSPBf26yAuUFH7vAlyOXm4Y8/ELfhh/gfTnlbMRrKK4cFFEULf
yoiLzJqz9HendH44FeNowUzc1rPz+YBzb567/xxVOqujvfeL13HUaJLrW3KVNKyI
MUZUw5N4u9V2mw8/qBOGSbsK3SQHOPKKvmzU75bW0ATDxS/PLgRbZ6tqXuaOxWAV
o3eXLQZ6CZS8nHHtEb0Bp6qlP2NNTzHpxHCBI8Nr5Damez02c+SFgPwTlUVq8FOj
qaOTzs4LsXrjy6arESS4zliR6VStCdn3t+Evu2mi5UtEOQk9TAJ4YrvIwV9C+1Ce
WC278WdSMxxs/lX9u9gD189dKR4kx/bbl+wCH+xotpS4XwiglLAysbTwu7oUZjE9
q7Etndr4jYyI1hx2Y+/e/Hzec7i/cj5Qn6KPP1vUb2sblXvZYgZS8pehiAYoofN6
thCDJrMFb249ioDHpztJSRGWQzGYorHq2FqfhUiFmdIJrCkEaSg/9D2E2DHbKddB
SEOMY2rKpWwyuAdmes/ShPtWfN2qThx6Os30MDUnm51y9txywTD0FGTsqyiwP8aL
xj6vXpQlusrGh/M6TH55F87lqgZL4SbTlFpanX2/SRRVZGzazuzPeKp0RQnu5OUB
SSpjq+8oOP5oq1Dc7e3G42jenAYnxGXvMLOT3ZMRCrAEcOjR1KSrCZQaMjxlX2On
JEpmEKjI0nylI3Ei2FnB3ytmgT3Cs/4ZQlWDBoHE0beirsSYpcmlLkntWvaIA+DX
egrqGBxkaKmN3Xqwc4xJAyEcZHhslpi4AFiYupkHj9wLRBpZUjgLTrORDnMlI/Zv
CtBlHLYnvKNul3XVyCMd8koZGPdBiz8DHtuYabXKUF1EKpDqQ5CVfnkBrtAv1KVs
O4P/eaKw9YyCPgwdeo6dVXaaSwCnuYVtwGezPgyHupUF8gWve3fM3u6Nr7x/oYwR
qBkK2t8M8cR/9AZvo1iBOdebtY0U2Rb0nUX43iWzwnY6VXT7wrhsLP1dHVRTso56
E9gGRsEPcH1cKhNIYpvI9tIKyhcXAaGQ56/wL1RacN9Cd5BODj49o/M2fR9nHXPO
KeCBNwZlDH4fwxtQlgjLDdeU3HgWaPOOcJxnYGoxBhm+AiqJdX0/lXYilq0RvsCY
QQLlh0L+S0E559GT11k2Uf0iM+wyTLgCS6AWMjyOPRSWUU15MA6iS7J98B5ydvgx
0sB2M6VQA0sp9itTtGXuXCnhcKJLnTlX7jku3y4cyx0ScyeS3e1+xAsyB+TSo4iX
yvrlTP14HQhlNjqDt7Hi+sSdLUQ7iiFV4dAhFbrFywHwD5Xp4cXBG23qr9r3Mq+G
vYXgjhyuRNSkXn0fBUkk7zXSlFJl6dB+Ncb46jbmJPqOqCloOevIXMaFqKOvYBAn
SUI3ooYP09r8tUOC2zC3u8E8MC/w7UK9uYpvPpXkA1GGes0lM5ipnoh9FjZiJHxO
QjWfrj+Z+8BCLJvwkhEZthBpgkER04n1k1TUsMiGh7hGcnwaij295EupkKkegKjV
ZbRWlsfepiJbgxZYWbZ0/9GhMdYPOL5jjzzpLPYwHnrm0EjXooZeiogJNzyr/Knc
l2KMRJ9BNivV015iSEe33GCRfX/24buPHKxFRHypuhpzP/VuVMbMco56eMGRKOZG
VJ5uIpqDuNbeVf+gprh9+gE4M+bI2ghZPIzb1IkIA57G7cN0yRruQ9lkkEQulzU9
fNqm9F+FZ2YJkGh9RdRAY2T8Uh/1iZP7lAcucX+YlZEkF/MlySJa8sLvC2HeCvVW
s5xoghDxLhSuE5q8IUnogiQj9/R2ZoVklVL+aLUIjTHoInU6qOJiSJBAyhdd9T6s
w2N1qwmCyrugV2jwuwE8rCJuGuQxbMGcnbs7TYWVsI/DQyi1iSXS+gm7zpdd/pX+
wzSPy3KhMG2+398yMPGO45OevRbNrmPlV+CNxUlVkQgF6aYyfE7PgrM22N6j1i+Q
Mn5eGglcFj/Q8Rc7LcfgNm1B9EAq9Sd/fCjPcFX/NtEHVxxtS5iI/uVC8O5bpbfz
Wpyf5Gq0JRXLejmyaSiedLDf+dVQHFkDrcXvZ9MkDko0ZsdW/51Wm8s348c/0Smy
3Cj94kkKZliFypC/iU97uPwykaL9wYNnbXreRXE5IT26U+UyfDtYRWk2NZuK8EXH
mlTHog7P/tA1nlLUCBTyEz+T2SOX0J90U0xjr6+nDF5goQHr/I6aPV6ZyH5Pe/1s
XZcn2QsKgvhCvWrhYWcGbZhE78Fu4AlkUtGGUc9+Qn5+1hW2WCpoZLqZB33NIXdr
XcLWWtTlqE2uLd9vEmq3Ldg4p64cqKhiA1IOy6R9ZouNzq41gdgZoSzXEamLq6GO
//BUFFR98cJvIKuFwdadWslAZE1i2gJTtyGqUvwbB4VwVAxU58XJf4O/86DzhG/z
eibra3QbnuzEUqlVl4+lNZ32jL78bLHQs8ty1MTxbg1tkOSM6Ju+4E2a97P07UUB
/fl3t1o2dBxV2qCAAp8YDufokwvFmKkiZhKIiaS9pSaX+mGmS7qxj9nqFWH+93gu
fzfRawQaaYFj6PSuMo0sXFn5+QYUCteQcIcgc1HY0cB7mseVG09CEBxw/DhMpw5p
NpUtkstsHVzYBRonXkuxzr4usUFuE0Csy0nnqWTpIAEad7e68uv/OHFg1CEqOeee
zGe9d3fQT8QLH3tvixb0lDEEM7+RSEwSGyCGcL0twJEXr3VhfUabKbyhKvbQGouN
QoFQwDDofPSRKaCAFqUNa90XKzFVcKTtLQHo/dCFEs0QLZowiTkHVQ1sCqkdut0I
oNy4zxH3rK0b0rXCTUpV982gRFdCnEZp4Edu1qcSc0mGCGKH4ATO5vInb0h3OoAF
P7hOkBA8z3WtbDoe2+motLmeQBmYX3tmNp0JkLhKDUPmlRCYlKoREG/lc+IByiyX
B3yiH9loyFqWgG4mPMant7nq/3S8Z1/PBbfA58+0quM0L+lXnU/6BcnKE4yPN2Uo
sDji+XTQOLtYifcjqsnOP9b//nQn/xLW3Rd2PCh3YXyV7ZoIelBjP2a56S7LQV4n
FrBJoVGxDI6dfcEKG3P0fp3bEL0UrYtJw+vI5CIPuBHUXYWMWfYice7j49FGDN6J
n6oq/aOqRiue4h6iLwzSw+pyxgvbJP7RrUDfPHCI4K3g7oljcc5lEI7/34YzR2+P
TLbg1e6YwvhkE2ssJBAh+ol9wEpmv1Dx6e8XtcrapfAl5j5JFHWnpF9U6maT+dSe
HqPaxoCMCsFsP6ey27djrupjEbXw7EHj+k9F2KDkN7p4qxqbLmLTmagc81Wj8SKg
gdWXbnObjja5K9q7xJzWOmfHrJ4Hg21olDpvU6iHW+ohkfbNb6ML5aNaCQQrfhJc
NdEAwPdUDaTQH4TbxmjUoH0xdXpOrMjfhg2G0D0s4hBu0uN3WT9f/gYDMJyFpd3y
Ia0wxq7fEfZyioB9MRLFf4VE+3rPPlk8XPYfouTm/1roy+0Xzgh6G0ujTAo4DxCA
MEXgTD3kUpUHMr5gZY8Yi++GN5EO3UdtBYjOHxl1IzZmp/IYZHlZdW2AdBYU4Qp9
gSxUiXGTegrKbNew11/zcdTiAeF+KRGQByF2wub9Blj2RxvmW+Ctuno26n1CSXB/
tJpRwWmE1DsXzTtbw0oCeMpGVbA1GN1eCsYz/ca3kff5Sn4kas0JVCqOGFqJdfek
GtVlwQ+kNQc+2qofe7C4qUQyX4h09dZfltGVXMFcDLwXM6S/oHjPZNfdHBVhYaPb
8/9rCktLhNhqVxd06mSYSqyoiJnH5kzNyAgT/ey8416mYktLgiPUojYhWtSVA3A9
AizKQGgkQfaS/yxru7AzsiFWd2bHVA6UxdktWNxyN6p3+rbTSnyc1DJT71MoTCoG
fRfTB5DfUdGOYkFznxjXzFQO1Kmi1Z8amESYABG56y0/Ahfuqa1E6mcn+zHXEFtk
m5K0GGCxtaKuEImj9yx/wALxL4PAFJ9BU3QbitYiuuwCRgiNBmgkmLrjLUhcY3dC
XRcfhJOpzpcZvcHLVa5PgXhf2nzsbgQN8dCyfFZQ/OqYGO7STcK2aix2tzNpz4M+
9+WNSUXg42tROfXbKlJrpzOy175KMHtl7YavRv+xs02RKYeZShsWldOKygOsgvEl
l3iE3dYxV8fJGLPeHoDU9nvp6xogpm1NKy51ojMNvB+MaxyZeUbXsMzmKPli47Ju
dX5c3oR4w0n0JHv9ae6tGqDaTc3Ris+jv/ZuFH1Cv2xSdudTtCR898AomHoLKGnG
B6lXs3TIaE4HhMl+GRYhW+HpFyJn9Yp2SG1f62CU6zR0jxIkiP195nPjHIn6DdDA
3AdEIzvdKLwEnXij+Bnw1T2pN5sZ7cdWaAXgHmfOehDYfLiKPuiOjBkv7/4Uuuz8
8jDeDRzREa+Bnv73b35Z65x2ySdHazdFRJzRT+4y82C7YLecB3FxZS/abq5X5EZF
ftx6eFoZsNvdKGa32YPAUiQT2VHB8qJK2g6rK7FZBvPMIgwyQGieSP0hIzLjgXMM
xQU9OXqqpkI6OaZ9CvxdjRbwqezSx0VrHy43WCFI+6nTAfg7p/j7t2CzFmPaY5/I
mr3vw+03izs2/QS6COelgTWZtFFyJ4QgBg8uk32dRuWjASeiNybs4Fjo+EmfKxcA
ZvIT/r5FYOLjRkzZ4gnECBkZBZRpGmjFb62iDKLE2cfu1xmZLpsTaJMmM9IO/9qO
PKRNYnor3F1d4AUrrSAYGbVu7ZehyI0BmQjK8MQR44Ldqix4C50jlFZqW4MLkhC4
il7M30TVm9WpLWp/eJZGUs4+ZdJ/WOS5nYd5ZXr8Yu/96HSjnTgHEdbAoxn8mRiv
lBolAs9z5GRmvdruKbdQ43CAIs+m5BlnC8oXGBqsoEiQWPO4tGKYhnBmFBn5/6uH
JgWZUu+fE0PW7/eRBbgd1gjbduB3Rj1zokkHmIjGw8MgisP7YUJ3g+qyBSDrK/58
vg9vRjav8tkq9UU5xbXknMN8frfu/39HLm5xuxtDaecFqqEYSEz3JYi7cuiVw2Ac
UWL8rYscjj244bTAFR1dh1Oku+rJwg4m4nxDb1IB8i8baIvTm8p+dg/Gez1ZrwyI
QuNF2o9HpdJi9a5mHo0Xyqw3ElzV8TVZZWlX7F0HrTUGEENQaj8az0uD6Va4bPq8
BVSd8fsEVwC7Eqn4YGTMpFt2vrBAR6+jPMULgbVbdioZq4XwDV0HI9EbuQGLBOc5
as3wXKCHAlBu/xc1zynN6Zuoa+arp1Ygn0g8TQ0xp4HEJikJBmkPoRdKLpxyGEA8
dzTblGz0idevU0WaW2xpZBHGOHYsQ/Bvfk8SYSihZrCLMIK/BFEJZCn2WaRFC8ds
OTBEgmMXxccPQfCj8n1Ebpnvq3sekyKH9BfoQQfIY/vl4a6C9TSRQ0YUAmcDTn8c
0XS3yYNV+VSUWQFE7/wkffOQ6GI8mBm0UJh0Cva3YifKAWPH/2Zb0L7xqaXgiPr+
AnQahusEYFsDEJFkAKjpQlm5RGkR+j4vFLoleUyzPaFZwLAWeanl+M8M+pAm1B5L
9X1i6w0TnO5dMqvuTLNIfc2HjhniVu8fDiQ2d2VsDS8ROZEMoVv6qwvoqCbCgsOo
nn8Wo8pknDZUf6wowsnsOaKeMr6gA7nlLFGadNgl/movOvU/39Tki2X+Fa39Ojn3
R6pHn/wmzACy9otxMl2N4Jaw5aCEO+j1VTcqun+PiKLas8nAHtPRl2sq+e6MWJ3c
7AVt5aZVkOp6NWzZ9xQ8w1chhoq1UrqCLz2+sasqYHwOs89O6WpySW/6oyXCdJy0
hvW3xgxWQ6wWlcmq2SiR+JI28mhjqM+ya5yUKgTZfPMAGCpr/VcJG4QSkbCKNDAN
GIF4Fkgn6RAi5NS67RXCo8Znaqz7EuahCrbi0/1oOtUQBAl6/nQcuwcez/ZktNj/
XHacrUyQ/jtVtXn9ONO+zGckTeVyRKsCLq4M4m3qZPyu3Z0tus0RG8mWRIe3XNCb
+8+GV1wdG0UDdGlxMu6c9L3yh5xtKTQ2qO+JA9VYixA2hm16LMgfrSkDsw0g9c/s
E22glrjgEC4hcZW27e95xazVm/zEQZBakrJeo8XY7uQf8Juzy2cjiiz7h5p+rY30
zSNJj4SwvzP3k2IwY42FTUPEGpCamUSRrBIVuWmo/ZhuvJ6pPdZd0ufgXla3D1Gp
O6W6N6OA5SbUKQ/DOp2IJhiRNhiNkGh4Cu0h/mA8wyI/pI6V9OSFomPIDSxRv3pZ
ArEZvkSk1jpMwTkvNnZWroD3bdN9zUX1dF3cND8sN/hB/4HxRKX6Aei+sLAAvyvV
KbmekK2lw8XWE65fkXkPCpfvqbD5aj/jjdtI0C76c6CChDk7Te8+Jmg0W+kv8leW
+rYoql5Rr2NhmliRCLCUkyzPZu4Er1uufAD4stmyd9aBPbOgTyd1K/p/EsNOakvr
6K3XZTwSgP475HamJ1g5bdCzib7tRmwxSg5lEJ1MmhUaeA/4RflNHfAGaN5BMsTb
nbl1w2oUiD7FXT9/YglrdpudiGblPn4FkiJfBHvvcm2emCiNP31tXGgaQkWbnZ6+
k4fFntviTkr3EB00QU8BKtC0cduHJHU7vCuHW10CVNdQR8glIT21f/hpyc9nz8Ux
/ePhSFJqaJQW1Az/WN7/SDiPKmgcIei01Hr1t2yUz/95Rvia0UqEwRQJS2HyA81k
FDkgxVePpoeOBjQbtP3BtraxnhL2qGD6yWgdWq4KIoHYZHOe6hdull/XsUnFSpq8
b54ha1aYhZ4/Y26IL1lQ7U344x9NHznwV4SQw+wKP5IEWyRk4vogukfAtbyTjmVk
Oc8xVlKAjPNcyesYTxHqhBMbI+sx621y9Wr80X2Qr/FUHMUHKZJwvqFCf2n7TseM
lr4+rCiD2BA/Y5l9t75Kq7B1fte73M1caBDbDB7z+pLecg2a3YkVFhkSOeYqOh2C
8hCQv0hWcS7btge33QUWdtGDEy5CUrdNERWbaxYq7Sq7UaSAOj7bNzEnFQXloqw2
lRhtbECTf8nztgdnqLURK28v9GJIZBehhZvkqJIXyVciUrX+RD+8ilvO523sraXS
ngBxg4aNj/HGf8fu06Ys0qn5yyzDZ/fBH2acKzIbE5s1elh4aD+zEGBkA+kCmSXd
GXYxAHCtbQLfH4NvRJnBOVmaGrwgiEVZA1KiH4p87GC8z6hl9J3XaJoTm8Beq1ZG
edBCpVtVF4AXdWDIhkiw7C+jF9aL5ugb+LdHqBwJymFyRZ8vbLGZRgAzhfYE1NlQ
0zNPdxswUlLvmFxJAzV3pyLlYsUAVOCcwcFt4/CNNcj+3q7aRCgPCVi46UY0BjCE
iqgEFi0Uv8GX+pAtHyNbPZjKzfkQdDFIjoIrvehLF1+eED286YJHcCoUBeDCziVO
56AKHWPXcY0Hnl7/CXD0s099bUpTHgAlknmhP8gVfILQRHLuWylXsxoT1zytwFOZ
hKLVjYlbU+93hNvUrU8h4QEpUtHwBWGiSasESIJPcgZ9mJ66BRtqrKYq0KE/Ge6p
iBFJmZYnE2AqdG5Wv0Cz8AOOfLuP25fRBSN6CWC7yIKYy5Xac9WpV86dAbkHZlZg
hbD0smKWEpjsvCPCyFCwDNnKzCaxtRmkCiTJvhmv37ZpyqtCdwukE1HmcFPOHErV
zk2qVc62z8beZKDJjAypsdMWM5s8u2F2LHCW90Jn2EkSfpa3JFerWYg77zxGBwAQ
mtpQsMy/ZfX4WZomtmXmAmPTbMJH7oxRogmoEp3wiI8pNZytPY06hJ0ulBHpcXIC
I7WmFTI5UWDlFloNals3ldp9poEuZHfFzslTl1lGs4McxvfkdkWpec7RX5qqQceG
pUYF6WmbM8Ymh2TmpLJ8hGXDWq/JB3tkALd8OP9GqZYwaE8dOcI1V56xrtNyzaeH
ejrm0+vBPugf92c11xGAqbaQ6X0Wr9E+G8/GLAwyg6oGwi/Qq21u0dWpFbw9qEbP
d1d/qNOp8gxSm3Fa8PViAZRN84WUFYulSQoq5SkfjVfvG/uQntjpruCtZa/L9xf3
YxLoJTQguXPIym2T9Uf8uvGV990l+R14ifj6mN7iI2JAIZxcVv5c1Nql274AKFpo
nI+ZuOWeeyQZ24gjGILAQBHWK3WpcyFTtjgbcFE7Uu+zo8ga1Otr6FLwgv1bl0dF
O9N3kYUCLjwjTbJe6tI0Rl7twGY7qRxHJy8jIiDtXwJHJGzcfZ+WCnYONieIfVkz
kaR1pBiuv48RCpmTCkBir+8hlb4E2xDA7xX/0eaYhCcTqkEUmbwGzn+I1uHb3ZXH
SfHCC61FLRdWOh7RDAm3o/kN9SRudF8Ki4dkLlJilAuIj5uhPTQ8Ot9Y3cF1j3HS
jQawGwtcbVQlXC4jbhSfqlorMkCGnbqCteAM1nM3a/Ux27yw3uqdfjADgjERkWfJ
wI6waIDmdE10ztnu47Qqxp2IWaDM5mSmX1ZbJF4labkhTY5aefBx/cX0PLQx1qhD
zzHgI4coh/vaVoeHR+p5s/QlshzmuyZ+Smi8p3jTIhB7VfhSa+UGAQ3VMhkmGv3k
qIe+v6aeSgj4dd/zUsFwJ0219IYN+jzNxRv45AbWDzqP3iTUHk9ra83UeOS3zlTl
WLRKGb04tgHCap4rSQosD9foJaPfCtEWl7hXtH7kUGdeBc7vNuXvfVPyJ/wIN9zF
p+2PfyQOiGQthRGKswCFNUkC1XFI6d22+s0YrjsY7h2gbm9SvMRSlPQTi5HSY/pU
/gAsHYx5IwhmJH2DDtpIPvzOP9lg49oUPzva3AaFAmO61uwW7qH3JYNw38ZlsVsm
RFVoJBnRPWqhVNosS6WjltsFftMVMhVJm+9yK35nBSvSWsITyEYTzEjl7lyhfQbB
poAUS9nb6E4vebR1dnVCdzzrRehOC+F6Lnam1g975QQBEO/m5HNVxC6YjfUHOrYW
Tet0owpas4P4R4QMhSeF0kHvjFPqV+CQj9N2bc7j9dYwwv6ga5awIiPJXuoH1i7Q
SIBRilz8pcLNq3cm2NQ50cOQSG644u9OPQ0Wxrmmydn/7Yz3bZLu9ppCjDKhoXJ8
gzxlo2goJGEhaM0hOaG265tDDGXSrz8iBNIXHe0Bk/uNwAe611qOSvZ2Q6eLpB9P
myWczPOSBVtOkpVMitHWoPTmTg5qA0VQxECSY9jgjnbq4A41KjGboxfaw+e7oSgi
I217JhpDXKfZcpP3EdVOJnG3Kk6F+Fj+0O9tUvliH1ObIXCOwvlzjfkt7VuXjGEW
PZZwbsolzrwcUgDR4zQ8r9tckmbs/A7Px4R5K/urY3Y9WTfJD5NjpeX45qF5SKYW
njcKOrCYDF4BJx/bQCdMaXWmrG5Sk53kz7iqCi5jJdKBxZtsI8DPTvT8J0YkwM1B
C5r3qtOzoBdU40NxlU0ppb57QLk0c9tEdMhsdcAsL/qR7e6CXLBFCcVxw+Ta25pi
nNxq9KGLEQrquywOwHVtuFU7Ni3netkJT5YyLn3xGfOmfXV/p4RD0styvRxwQ3kj
sT8rowJbvYmj5RP3hwC4Iczz7LduzMI6S6UGEbyyWXjeVw7blMwpnfV1b7NNV9eZ
smQEqyoUZUJuk3OOy4IiZqIyYT3lEpVor8yQXUqNI4ls7q4o+CoOVHH6ODS+CEWl
iXs/a1D2iYzqWCLgbbW/mw2rb8SEeVKtPpUEIp5sgXoFdDesXXdLoHV1cDTKmbp9
qLcxKdSRFbKTXaQka8BKxLvblHTtNNuxCZLT+NIatXHbWjDGaBrf4CT3jM3yki0c
zc1uSsT+dEUnz+swIKNdR+fkDPDAJWQURVzzeDI8OP5ekb7mZTgl/m1gimfL6q7Y
RYvhhcHWp+vFpEnW2YWRYtLWtOEyvnxQVQBgRunbjBRXlCAiHaH9T+xl0MyrPx/A
fG3OV9FexB6pwNkms0apSYlPKhDoNtHkmPaBR1WUtTNQ8wDkLR3wZKmf3FbRatBb
9kJObZI7JnfcNukdQEFYRtkAKYlqvNHHPSCHkXmx9j21oQeocWkhtDmjE66ygf+R
PTiHFNDcq0y3FOjOEQ9ZshqNEhRxJyM0/4oqu49TA2E4R+4Yxxukp/o43JF3r/yt
gMKzjkCmxZqMbZlnoRhc9h4odIA8sa0xhPDfyYmEDyxesJUdtiI6j8OeLlp5Na/h
sqearuGO0w1rJg2+Uwd0sGHOGZmtHpN+HoVyTDrpeUQWvsZ3rmRL0t6L2YGpMAwB
JCYDau9nJSv8+HQ1b2QOLlzlSuDl/hTmRCQ7YWE05MfpweYENt1/fN8KD21mlQKl
YskVJfvKxQxh2Glia3gS4d8YyXmcOHBABHh3+Sw7mJSAYxVKvjfSYcUDbdifCQ9W
YSagDhfVWMX2QzIGzzYS0uIie83cjdHkf6toWVUSo/ztZ3vd/+YVamgi9ZdPd1Iy
7nmzF+cWiCbzfls+mxeQFMPHYRbBBugydPbLVIe1yyvTk/7jnZI8qFwsAwftCUdO
sqEWKWX+FRUy6xy4rF5d2Rn6OIYQxeUP4oI6dX1BpoFY3Pl71kzEOkFXs3kJYVkK
7LF3RK25iC5NQXaJeMnY6p/acs7MUCPEVklIJK0wggC5ZxxYh9UHKA9vQUrpmE9E
GwvqW1K0iMiq3UHrNBIpWmRUeEVY2SFBNAyNVaHTqA8dbvrbCalWvOA3WANY925Y
RN+uim2NBwsVtjF4u4K5v20IuCGOpKK+h5emJwyIscPv1rGFVMUQiR0dP+1M5IGh
JpJhkW7mvyyEHaWIgiQf2XfrgKItin29XyTSzPdKmHDYbMCQtsnvqOjNyMymAdgB
14t4EaAzFH18hlBVmzWWg67y3CxPQ+dSOqRZcAK6CH92MXzFQd1M5dqn5FdZKbBo
OhrIGvaCmbh3M/j6W6zVK0+5wEymS5PMMIWM0tdz8sbOlDfs5Wl7Dkl8YjTCZ74t
qWAbMn24AGF/BFZpolxNgbA9rJJpZDhYqrsdXQM04wLP4ZQdycczPchPDeR3QfzY
2+ESS9olJHhXF2AO/bGu0l4uixeDkYAawj870nTVl3N5a/8BX5+RQyJVZrhxdvdI
/r2iidxlhZQIYk3CLdZU8i84x+NSiYKNY9O5HiBt5uRr6hDgaYIcBz9bwt8clVlR
fC2OA02XiKnGDYzotqTrGfiBiuIxHe2Y4FyVIlEB4Wm12bVyXy23ir112ObTCiHk
wA2X3ZXq5+ZrNE6t/zpaa+Uk1amWwWJx0Ew7ReJni4eBrcjANIyvHd7mvsE80auQ
rzAQ+PeyqGLCBdES8rT4cg0wS1CibH9RTHv1bVCXShpcAV4I18/kUpPNmifyrQOG
WbQY3QQaX6xhOPx6K+2Yh/W+Le5HT6CLuWUd3dwmeeRlmNPFNCcd5U8wzbYF1+Od
Jyljc51FFRht2q/r3oDCnagZ0Z/HwxW3X9Nz2j861SYYXW8gRzTRPZTjGUG7kzr7
r/IIoB32yIGO5b0fQHJzhIONwLZrOLjStJb2K59Vl6Y+/iyPdpwC6cLsMBvaqq1m
eHkYhn3cGnolh/Vut86+yL+by/29iXD/NaEn1okSwWpqw1Q5zYnd8KkXIcfvuYvg
5jNaGJ9/1MssHLiifZ47/vUjn24jd4+hnKyduzc4wEbCUpYGcfLcxyaApYHjD9vz
t3KIGKd6LhfEvmRq/HTEaC7RO+hYx8wVw3GwMUi7Y9VzM3+mFTtDKJJNd30U5koJ
WJGxSH7UCIL6a2/MX8UaQK5jmv5WXmS5f3Km3WK/ASeScKrkiAP4YZbnmw0LWVU+
VxdvM6LBYkP16l0PR2ZwEMNGBdYd1inHDg88H9RhECrTnIR0vYo1XN3zUpybpHI1
avURVtuv1ytpFX67An95gN+s4LKHVxDUJ+qq9wvzshDyh816Lq0mVx6zdc84p+RU
sO6p5I+8I/TutEBxdFq64duGpaw6TVm8s0D6iijXnCzcOWhMdGSf27pzE2vqvs+4
yFYdeU0ZF1rRskMykRMcHrqW2NdnjAJPSv2FBEJRm7BQrL8WUKLrZzqnjAYrKDks
znaUDD77OdgbfHL8+tRCAXpIO4UJUCJZp6mbbGr9ia4Uq7AS+vNcIHAX9ruvwJpX
LXuKajh0oiCIlczUHjXT2eIZnRkIGa7HXxTS5TLdG7OvnrQ83vRWyUa2JzZXzrfF
9jbedx9sSTQa6P2Vpjyv2lzIF9df4WTeV4pxoHvFKD3IAiqNaUhzlv6+lGAlIZ9W
dDJw0JOc+0IhbvXiwZmwockLmYxmtBl693cf8j3mdvBGZSyuKwdHN9AjXCnBZAgR
fydmI390wFx03UtVnJEK/83AXGZubxNvHMnddYQ3PG+GbEer8vibvdeMsDczhl5Y
iSbuMKpWvWeyVVnDBNwMmmMwtkXvRM+n7xkPLvYK6ENqBhQQUsw2Cr3gB2ErfoC8
Nl8wsGE0IW22aY6OZbJgVhBEiRF5Won+S3oqdTvsItw3+NzUTE6O3YTTLxEqzwWU
mbZ63sJLE4kM+xB+4JZErwtOze3PgtohkSMh5+s6XxLwc+RbM+ETDXTVFfvtmVI0
e6ch4CNPnAXLWOtVpZZDYGB8pikPClShvX1mykyXzswWtdQwtbguRjVbSUC7FPY1
BvqHcwJR+a3ARB1LR2WD+yyexJ0lRZSO4NPkwUxQowb7GFcnqvEqYpXHmD18+nUZ
02nLeLpHmrKYZLFNRHRaf6Str3BqiZCWhx1jIsVgktM+jnxz7yZLnMoBzD3Y6EBL
vBSjiT2GetLW91Scu83cDkn49G/aDSPr50U8CTnjfhWaQN6YziGVliSTXlTGLKFm
nhipgRO2+vVLwDG2oWX5RnrEwHZShjy5aDBPdZUl/jBbo0/ijSOB122LZJih3V9d
YB0RDAxCJsdAmPmDWR1rZdHAf8hRmFTMP54mKYRjjbYgULxcsBX5lRCIJ31NgBnJ
IjbZAkQNDaB0/kbJd53hzn3rj+df5V2MbLfNdMdgLyWjFZcsmEoW96JNo58jRGXP
GD6QeiDvWqAxfmBBD0HFYv+3O0/V7oKVkSYH4JhwNeyXPqLJ2hUVOOrON8WAvTrw
dPgtaLZRMHqXELUoL1J33TYbOyj5Ls942meizavkZH/YsKsiSgF0pv3aPIOIF+17
TJo4SCaMIVtbRNp3F5NYQ/h+Ox0CydffWGfx1/ie220uJrQLYoYqjCWIRrgNyg+G
/rCCUcQNMr0wubDfZNGGZRP5CPntqosBqnHWxaGcPARkFopny7deOcXgSQPcun5K
d599a5+AB3fiyNvXL3XqFY+/vzJa6AyvGAg8FC1nr4jK57cxwdV/1FSUgd8HhFt2
vtPFUe8hLACk+pWSUd+TiQJU/nr5xU2dM569cSttxkru8+lql/g9RZbXljZGsQ09
Fr7sBBkw9y43GziMKcarLECv6YD8PIbtQFnmgORZJX73qxrPjMgXKrpVkywrHPvx
+2+RLty/YwsYQ5GKBsoLwtmLDYhlcZnVptHYXsI0DyVaSmrWZfZjZVVIAfNbddvv
oWysmSU6nj929jsLR92Wyl5TQghjToVROafO4lcr+uHpUMF5qwdIWwdObst5BqO9
pi/DwvTyCkGzWOSCR/C2Nr5SAoM3Z92zdiF16Qn5mbBHX8CsW51nZj4+4aBfevSH
GLUeCVijA6HupFZnUAfUO1lsjXkwaY1784btc2DHttUt2dQRhSLSBUG3uFGQu4VC
CtG+J9JT8l8uq2pK5MTsdqKDe4d3micgiVBjCWF+AHb+JPGVjUsafZxbkL2KHgvz
MD6vhU5+VcSc2AjdH/6azhoqE/fPUYUxc5Y+E2QrkBY4zbFC50HsqtG6JLukGhNQ
511kVKUJMzxwSocVzZHxDadwhOqGT2TjI6Nq5OOyy1cVpkOgODhpEiAubgyHoXdb
f6eYy1YZjWrwCFC/SHz3F90pQ7euy1GveTJrfmaLqvK1m7sXPFgAUCXqXVJCZGBT
4zxGF+yRbvkA2MmTdiSlXHLk4pSBQzbiXyWhECmglHF3MfdMuvTOZfgaTZVqxMTC
6GLatAgevL1spTC6mKCZEC353AH4PE74ZQ82XHF1l2eXe8IZXR5GhMyxPkV2fK6C
nC/IW9/VSd6HCrQSXjNfZAexrtpE/bh411hgk2XVRsqd4+a6Il/6p732mZQaGvPC
RYfWRx3jOTBzumZHLsUHQKtVcgCpqs+yj75wvoTB3/ZmkVabi+uFD4NqsePEkOsb
+LkhDI9lQeusLF9ZjDl0OODsotWOc9Up18uz8xQ6xiSx5j3ulEjmKs4+X8Fhj+hR
JzA8xPDidR8Stkcys/yJkjlO7tezJEDJQhslec08idOLiy31kalAvbnGSajuON7f
dv34GUhcg91sy/NjIei9tF/JnE5ADn4g7f+dOFb7Q1rP2Aps0PKT+h18saIZqpZi
NJs+fzb7MLOlIUdw55a7hcFnyZ7SbbzcIopbEeTLGGO1oaYKHlScfTenXvxgSeZw
B0F1RcUjJRtAT69YfqQcyqQQrFc+onVu5driTUPdq9Y1wAlRLlHBmeTEBCK4w+Lp
WsKW25UpF+rouqocVe0wwzFdWt2VPfAZOqSIIpiq8nZZS0aeh82BisC/MVrvOjPE
rDSfeNQp+IbJNt972hQD5DEKMzrIDqC4fKKxn1CVBno=
`protect end_protected
