-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
34h0muTFYZWLmixdbVnLrui+/BkSYRXSISbXVZtMRK/HF0cdB9ce8H+jXlTRi+zM
G6GYhP/lBB5Wd4LebkG/ad7Gcqqxprco5y2WcbhBRqf3upEurNcQB66RdrMB3ER1
4VTYwDVV196nTuf272xYCZqqHKqEQ4l9srvutk73+48=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 47984)
`protect data_block
PRZWy3rYqqWOQEqk8eEkOPrjg8MjS8uf8BhUZer54Isy1j/YREXY7psFqonoYJ4t
U74TSN0JgsZ8kP16zUJ4ZqaKcd8aPO8hOj+BQHH1DI5kqh9oVZWL7jKInvrV2chK
TaRrO7CY5lp4IgbzZ7eq9xF6dQKmBGRNF7P9JiWsCi8t36SM8pWYi501SkA5mXZZ
HW5tqZlPU2fLjdvetLOV4k1GJd48Qk6bAZKDXxzd/S/qxOIKfFJBi3r5G6nSl+aL
520Jbr4fFlHgw23QSercv5rSOxC1bBvj8aRseTNHw/G9eS0jzbZ5Epsoq+jOTrw4
LEzj9/SXdg5JH8Y8OtcD3hVdFe2GgygfsmnRNWleX00pL8dWz6zQYOUeTx79VKtd
16tF5Yww18lxOyw0diQQGgMHv8tcYaXK0ovHOzkCAJ439cCtpmEBD5Ec0661+FBg
3pn03UKBIYoZs0OK4tnYTv9+MSn8Whvq5Ey6ITU98RhH57KHAvojao0M2mcrRJ8V
qw0E/JOG40uEVeD8Nmxj12Bcxeor0ypEWOpXesxzBDQZ86LlTrHSk3w25g9vCWQp
MhujC+mrD8XcrbVii80hmkClMRAQjxNud6TCoDKBbXCpVBCABcsaj5+ZqbP1TZgz
83u40f2dwXNvnPjsSJbicAwbsqM2cj8Uys6NlclOHNDOmw/5K5uAOvCMdkxNKPp3
weXco9gxU7DjEgCbFtHTUvs9iWbEsbT8T+uoz9YDX26fw6PzrbjJvWHYr84mR4M0
jMGigQhrkny4Oj1XR5rMuyKmI4fu4nOm79j8btaDAF/auThwEk2Q+i+x+jSbGYsF
YR9kS9GYex3ttKqF05HIJEzxHS9ShUZI0sOz4dIfgdz+wxJ7hBBqCd+Da7HShdAe
kaWvJ5ULWCQo2S0GUNDVOprpEnAlC3BQrvUPzklaX/QK9X9XIa93LlQ2YOryWddk
w8hujLBX5LW/wBSPAysbqUU/DAnTprXV3DBT/fXZsHXgvaB3VoLWIDOYygx23BoD
NHSm0VXWWVL2YvYx5s6E3y6MHPjPCC+WyBEiKpjub/sZyZUOLSnuY1rkQu6ZkzZS
gOYX3vMcnyBwwHtWVb4RE0qJlIovlY/CKwg3FdlVcf/H0ooy4Vb47aCiIc/LTWS2
G5/1S943IPHQN6iRTJ3l0i2eNc3TnDqACtc60NknHaVZMRGoR/VCbmKhjzEbt4po
dcs6KWzvO9/yIAoLeQ2d2w8dnHGf6HrqAQwBYir4wZM4IKUPEBjZlqYtRYfopjTj
cifMKv1pASqk5cxYi01UNckyiFte/e+pkl7/r/z6hAmDD+63kVsbbbYBLnXit9Z1
ujd9fdVaZyJma8BsfLfInHGIFwI4o9l4OWlqrTa7Tt8DiutlhRU+WyFjvjciKc2W
CEdzMpsi/8RkFEdDIhYb+7VoOVht84d4rsMKzxY0sPNGRqWKQOmeeUSF3jo+RxGU
9Yf2vpA+DTqgLkedNeKht8FMWtdtUnmXeB9IUCPNMdel6jB4umewtf+qYkH6ueOr
Wk19AgzPkXo4PDqDcXgZg+Iwkf51AY15LA96g3Wxmrd9d1kbn6VyZqBd5pE2s+A1
jtCnqxfjTMeUPN/EBzJGKU+XEvW0hIwtjsE+fb/nKvAkL/OzYMu6OqOTAZ6xn5nn
GXkRA2svdWJxtYWHf2k8UpvvuoSyfuEpLFzNoXJvVBzPNDN9hWiXZ3vweepJyA8U
h2SMSv5aY5SODrtjssf7rLst4mavEGhOSdbSZBjcRymuSdUF+DAsiqf7UqMjmR0d
fMgmjVd2jAyxIgGCTAU98q2xxct7DbLBGKFK2r43wwqPE3qGqiM9Co7YaOkJB+Dg
YmC04/WHNDkorbF/4jW+9Nq2Ywcdf5CWjofpFYsobLQYfu74uRXFnttsmpnDeFlZ
2njWiFGNenBLjFJOSlvCL+MSafr739sVmKimPhO19NmqfU2kJ5OzMYSmNLap8G2z
4+fCNr1PJrG5AXwdGRL7bvptWTk+ibXwGATX7cGnaCf+ai2Bli5X6d2SBqmcKVkE
TFPH6F1mgQMvCnHUienxFsnNF6/1CkWCGZuKhsmwO0BzuWfEwsQFQ4Y4I52GMQGC
/uThR2Ssr6hJFudFeBJv/d2MbqTjn2jTxPWKZjaEvKcTciRiDNw5c00l7VgN0OPu
r2NcadfKfAKTJsDJI+PL/Z8AVggvKca1RHwk/vPJWkQED+r66Qcldowri+EFk9eK
Qj7kzkuB1GT4yuh3+23+wqYIH3DIBdWz0QJeJk1N/MWfj4AzIq6hCKGoArDaH4P3
KImCD2cE81bxOxMQ0dG9RNjk7DsF83Q/tylX/QMZO0L/8yL7NDRWXDUWmAOYvP/O
4vbLApB5tUkxqRrgxdBnhDsEA85HwAMpa91B3Jpa4sTN2VfF1D+LE+DH1N4pOp+H
l5a55gjJE9hBJwCR31UL/4nWKBnyVmqcbo3H8kLBIm8VS78ULxYH/Yhp5juwEM3P
g6s5CW7FYfC/JLC4hsxFP5I7/5ZklZFWCJZKA40JvOatWONaqm976ksD807CgUq5
qls9CCrp9P4iB7STFlxQPBWH1ETInunP2/bg/YY1yvFGQYgAVacGRB7cNAk5s0Vo
9W3Ty2rwhl/SgQ0mY2Vwr7dD+eAPwo1HbhKG0uysZALRE4bFfZMC1Q+UeXp0Zsx+
C4W7HZ4SzMSbFYzcAWTB2Pq/6n9P6LAuSCETI1CFdWk3GNpxC+liCdVPy2/s3Dx8
NjuF3rkW4cJeUn+I3NYrmUjSHkJ/wkAF26zsqdg+WezteMTOCl3rLcWKjf+k50at
5VRdktRB+suGQ8x73FcDsl9uMVno7RZvqbt6zmPI+SBKiSgwtibd747sPSmb/zvN
9BheWaP52lUufPtYdPxpPsSSteKwfOmn2XNgFcYP6G8qSLo4DTmYp54d8EY2UXdj
ahfIJKaF306oF/zkjKLJXLix8SaSzptfEG0i+UqXp7NBC5ukCiihutPQvOPc0v0N
e2IMzJ+3PqB5ubEHweMKVbIBxzgQm2qQA3Go0q6/vhfDwQtM5bTL1CibQ7ZTzo0s
0PLRGNZwmXsuOs0t0eOBJq3hlhAJyZqiM1w/fZzLo0LoDPAKRWaf3YPVqvROHgGK
pw7Wslf7baNP2i631blFzfm7V//a9EuXKpNM9Zoz2Jfg8Bzekqdn+h37SfYY0B2p
SJUItpxTrK0+gwtUIFiPfXSfZYcsbNydoNeIV9takyxnziwkkK19xYpeRLv1xjQr
58/WR/4Gs+wBb3prVLgW9BdHfkuTN/hqp3JvxodT+XVWXdLQyZzcSmAJD91ibgCM
pJtn6m7GSBsjBlbfQQuxBPAj53AK54hZVD43nH5dn5hPDXFiTPdlpbOm01JNoNjp
sIfC+CX6qgKob47UCANQTV+uBZTGPau8Gk0kbYExv7sIY0jp6yqn3kFR1SxiMP5X
89qCibVkgD+wnCnw84dToPD01uqBdbrDwwIcc7u7dauDxiPP3snvydjR1aeXv5Lj
kY3CyzWOUKRpv8tHjtkMxGdLILrjeNuS1c9zMkjtgyaIu1PCyglEyJMDyOn/ifYj
Hh01VkTZoE45Dr7u1gxEDbF15XrlEr+NCsNqtPXT78QUyLehjGDHPdzvs/M0mKsc
CEh81R7BnJ5ndhLAT5iWFN7Qp/HbdcU27usHhIXOu77sxBpzrgCxNtQi/9MZzmBg
SUFcqAljMAyfGgLo8D+uYAmhqmB56oc6XJUZb9+Gxx2SNPOaLqnHKQ9ioqTvLIKa
4aqB+YoKwbKuye3TlZAqtVmTC1f0Aoat4LXO4656GYEq+SpP0lsWd3UG+buGbD+a
jsTiVvoAZtzmBIpELdtRPHoowDJ4BnZr82kA3LkvrbgSK1CLp6U/cjkFXR/LEnDh
+04lzxgGE0jDtuHNaP9Wt6TaautIjLsE3nwGw2QzV2eFLJzUNYvUwUFAjpm/wWJo
8/pO2naURU2hFS+TwGDnLwQaGWXi5DebZpRer65Tqn/OE+E2kWce0Ko9A0Zy8cct
n6mdutrlPe1qmSN82Ld2hnnqjxYb5wzcZVjCpRY/C17dntX0o3qZKdseE5vmVzj6
/75gooww5oIvF5zJhK1eVrUgjdVizaGT+6YkePemteGocMK5V1WY1cAfCS1yEg+W
oFHcdCFq/gJk6HkLoq9DCede6q4ugAiS8fl0oFMl+I8CbEYzLHTgAJwvMNoppD+s
Mf8vppvrMNgkVVv6etnReH6ihSSOsFSIqiawJdKopVva8rIon5ChSkXGsjbI1pjv
sjWiTxfgzfeeX8mQLgKXqMaOqk49Jf36gfl+LjJey79m0P4pmE6i3qwSpLG1w68A
bBXVX4csYJq1e60kn56imbEeX4i5l4NEFX45HuFGaYLv40ihFXVa3ia7JCeMLBGf
zwh92d9sYBaeH91YJlKTfPkZyQWGhcZHgvwo/tqVPG+b93NTX/t9hYV7UNFQlSkM
O1Y/GdYA5tGSSOyawBa7O61o795NV3Dyv9oStW4X2SM6lvUgHGW9pWmE1/xMUXE2
c0mqaUJFyQXQ6n8YeMInKOrLNtMx/6xW6uUhGhJzllDX8Ee/QzkQ51C1EMKWLFZI
mmjZkUDIW0vZidhBHGuXX116lhwMY9MPf9fbi9ifdtJLzvXp2R7n2ZWyRDhIojuU
2RNzp4IxgTmdgiJPp8JA5+AKyJEvOVjJx/becfeafidU9lXGklPuRmctDhx1ytcI
/InVzCD9SJcdPP77N3MgDYefcqB0YQ1uFkDUFw4SPEv65r5EMwzz39UcFAYi+dVm
28TZ9rH5jznlJ1aU0wMW4MESddnMP6s+wYkjkdv5KpnP7+Ri/VJZ/JuNplLAx2hd
S/V6uMMH03X9U0Rxj6xMiEqMfuor9D4cr/owVWr2mrP/Nfxqso33vDMxUENxzdNd
b+MC7rS7nBTBiDjaS5T2NKGck/sddAX1Zy2RjfOfYFPbxXJMee+LRiLmMeREc8Q8
xZdEd/tUtFJi82qe+xvmhlRVELY6oEJy4iK2zQtdfXpkQe7yjQFuTvEInptE4bBR
qVicwJhC627uNuInusbP666dSv7PNd0jPKRTFjM2xRDDDoQNfnV1urtC6+6c1ciJ
i/8/ovhFUufDwGKi6S9WuKTChRNniGc5r4SSSSCCbZNNU+ChkqyKWQTy1OkLCXf9
J+bZuhf4L8Hx/6Q/Fbjdq3vR/YtAnsOJTYpkKAte59/carEGi8gOU/hqi6a5Ingy
JqxW+zKJuiBH4madz7S8bL9fMAZKJgGQHp90U1QZbSyrrt7hdMvt6nLgpCpHCI+N
xRhr6LhLR9FvsVeYLayEfp32D2WvP7GLS7tg/GbeOxca8DUSKDgBKMBpiSudOP4N
ANOnF2hQN9YF39j+eYjeWt7ZVFcKO243dKbZHs69LEv8LAO7Io5sBcNvElZJzl2W
WpVa2Rm85VLNIMRo2vprcYcANYZ5t7a3bdqlIOE4jCDOroeb7tRRyx7FBeRHr3DP
KfjaNtJvkmHQqXwaRsH/wGVYAAvBmg2SIfKcECvwWVviz/I9RXcS8OMqAQhRYAEL
HStl+FrPFlGRUyZEv1j98HG6v+Dd6LD6L7vImfcdkboGt6sA7+hqyvYNOYqrIQxR
Gw5zkDPGReJ0p1NcWVEyoiv1D1rKzGQWj9QomdydDjJIxfKVGQrA+iXrBb0l9j11
KAnE2crCcB2wYJT8F0AxadysN+vObsBM3pEfpmRaPWTKWQEkf3JdmUZwhtlnIKZA
6gNBANVT4l4xK+BzPvVL0hng0F4zJVAaqFKCaZ5htZl2I5ncdglofX3VzbQ1qLkw
oo86Rb21wRKBgoS5QDz2v9YpsvCPzG7qPvXgGkQMltNFa6N5hUOPW+6ryMJGALyg
24iGiVScabW+Va8SQtKE0k/j4dq7ZBT3kzILjhwx4BWUeshx5TyacXdFvdjkZWyy
nje1j3S5BcwedeZln1QP1ypCjiqJXC0vJNGwpicp+WDK3B48xNi5355t684ghjnR
fIodJd44AR71ccaMu8t1iE+UwnRDhH2avcyWY45iRUXKObPU7U33RkeTSljDHd86
9baA1f8+tpj99mhX6b1p8aQ1Nh8fNcS5QdBd+jk8qM2pN9Tt+9q6PIRjXlZWGh4q
h0tT4Sn6CATtvOsYHfBV6Lmy6y2Y/7zJPYjtyzrdLR4Qn0MbSdIRRfZ11TetvxUl
BqEb8VuIu+MqT965BrWJGMjPzXtcwb3MUpODfao2iKUkyfQF+/aZlYijzcBOQ/Kb
Q+4f0IX03jBSz004s8lunYKZ5TSi+W20Vx/xpJkkGDOqkVkgDSbwev8vW0+IvdYf
VJyDPV5Uc0PpbCec7fUw8DIenvaUsS9orEhl5GPQsTqyso/N9Mbi+nD5hmgdyFU5
bEwfCd6WmOsmWvF68rZBRSTNzlNFhtJOeeLjYsdj8c+/wz7x4wNyCapm6CnXLumD
ao4GVpsH08CnjluiuhGY+vJtcXcDdB1mML9bwPQtTu8mto6u5xh+0OG/Tktk2UWO
si/9Pxz2K3zvfjuS+blMbfWEPbRV7u4NIZjMRKXaU+WW3CroTj4HkGqvUTIx7TmL
b+KvNMoMDY8isJswB6HcwjCoNmea5z4o4E4H49W76d+HHcIGEnhKBi9/Xrd0JscQ
95Cqhxcz0IL3Dtoj6K5F90wE0+bO2OdjwBTTTDCU72Bpb2To9SlpFPqdtT1MWjd0
1SoqrWrQ5qXd4WEoSlrReiDLICVmKVf4eD6vKzFiBjmPprhYYlan8wrKGXz/2TaW
tOaE4EgdWh/0Bxtk+MJc1D1bqG3Yab3Ik1219Fer3eacuVChl3UFArhq2FgLZaeZ
edWBpbUoXqynUTYJu9fSwcGvigHXdRZM/IDGs6UmHj8nbeJsMZPO7ST31I/mEBv/
j8crB+uA61VpAv+cTHVl54O+VSs92DVYRzB6vOCmBY3EMHcG5sgqlTHxBHDL3qbE
XHG27SbkDKkU96N3TTM/yUAb9Mw1x6ppEXgCTmCIa7s6//kvRu83EPKPbCSp0Tmq
q7+MyuMjBE3+agvr6CDG+AiJla8ftb00SHyWpOB9VRQMk5Mm5KJARBeWXmJLaZEG
6VLSg8HXUD8tZIw4NrV/jzc07n3/sbdkpHx4+Bscnm157gUPqqmRlCMffgtRxWvp
uFHZzYLu8I60JObF1Lb+Bi8hTROatjfQf5hriodsQBKUV/qGDmg79pbO2uQ+Razo
VbLc2VFqxJTCmtkVQSJww09AkTILPjs4CsqLY0s0lNTbWR8nU3pLIu9kY6XPTHwj
mwz2VC/607EIDzgpYW4r5UgCzYaSBnYphkhn0lWHt6wIPt6+z5eaOk4NFVeD5DKl
H+qPeyFk1+AZjTNER3ElzljLog1QHWe445TYTG4cUJ42xLTEmj8RBuprpVCRXJuF
POocM+uRXEjpSFBvtV5e+eahyTC5EpXsuwtKgJ5sLoguQJ1KhY6w27ztiIIXBMfl
6xpqVHAHJNAwfAmAhF6fHfPyXTRYieDhlTdDxlq+OBj+qHwD5hKk0BslTtu7gcCe
w/oE2x3TJ39v1HzlXtpPlJsd7Z5cwB7k5yx1zhWdBuCCmycSr3Ip++pDQGclx++m
1HMCAeQ+y5Qusivw0nUJRQum0qsg30A9kd72vKCsjtxYEokOWRWB9ssx5Ed8yQhz
HQs9HdDMP8xptZeppwxveBeQLor87+zuygvAQ5x76Abt6aAawhLfgbJzS/6bchMs
1DnTmaddq5qRgJhbPSXhQsI3a7nDXiWYSCOAktUA9M03dYUfu4hcOZzEduEfU37a
QWLeYMJ09wUfXNfGNcZdavjy5v7wBjYlHmfNgXHzqpOWo9fkJjyE5hgQm7U7FaDw
OVaWkH/ZerGeoeW77ATO8yNd7ZXB85/yygf+iUTiDmdlo1bbmzjGaBCcayLmDBwD
yGO2yYpQXCOlMfZiCowL4SgBXv8Y6Z7NYNyYe7XbwEK8ltp0p/Bbf+nysKOVwce5
Gsv6P1K+6janUP5rRnjG50TxExTDzC7EI+Ry/S7+Az3y6Mz6bdV4SysU2HYdi4uq
3ny3/mcqGbCcZYw4Nqqn5n5aKyNICb/jDXo3aF4ZH9OfTe9kIqmF5QWLjdETpaWn
a/qP841Qyutl5bCXCwTaOC+UMxl3MmFKarpGFrBn92ryTeuIKgacL4bMjmzBHB9h
v0M6ZmcPjL/RtVd/qUhQYqXMg8Ypa5jjSjRbKlFZjijxIgh8Nr+6wf7NYWBcIQww
e6jWxfPz+2nCTq/CyimFVpITbdq6EAVY36GaAlSeh1McZgE7fJMNzfQcKDhQnHkn
eWD8Lr9zVst8ZTioVE9U+41GEaeIq5FwLoqsAoGmF946CtSSAT+j3m8nQzCdjaT/
fgilxGjAyuhRDBKQKmt5XehOLrguUSGSt5nwnRpsoI/gKRYFmEYijRIsZwAs+AVZ
J3nwkzxHMky2F7QBNQBfq/8DnjejO+6IA2QXx6ogm5QmYEnGLBZRyyinA8kmXXrU
VHBagQO+dwWTJjmmeNN0RinFrBbI2fnsnycY0tPqmgLtfyU4sWVjE80lZu0GPp6M
N1/5Lf0SGaROTsmS6FLhG2ASsC9dYehFaGl1OZcj8LQW01cWu7V++Obdk32QLsv+
EEd6MeOWMfgdSVC0ZgCn1fJLeCDpS4Dsb0UJpKHmNEipEhQh963LODb5fpwB+QnI
li/huaFOK0PCqrObVGNcXhNxDAABmBSOaPM6f1Qf8upQSHEHwWN98M00vVNLjSG4
tz3dsSSiINNxXw+UxB2427rJjsXKmMmIsVAtkEo9od4Y1O+azZBSNmjwyL4XiWem
X86mT+UfaO3X7Snn2IBzx0M8bwA01QC33IlMD6MLFZtMA8r5SzRaGR4UK4JL/Pbf
jlffhZV122X3g94wKlR8U3S30fdtBjwJ8DAXgogH5TsHhvz4uQ3c6eWRE8rOqjmk
c2DemCpffio6p+SqULekfwb0ubvFSDRilAUESDE/3V1c6MBfDFIpSghMYrzILoxV
mHbTtIIntJndlA9etNBAOOKDucO/KwS2ze7smb8aG3pqMEGXhQlWAV4mFnTsvcmV
Jm7hqfPFuQ7nhtHVKGo1EIFztoLFPUtutcjjXrqhgU8WbTPXlCLGNKJxcna99UOK
3L7++h7oZFeBoNo0oHGrQBXIeLEAvWk4g67xFg9XQY2Mb/stMS3JgDyVtD/v8epk
20RsOJGLliVFMELanHUUZi2YuZQJpPpJB5fQZ4cRcMqMp5MfhM0M7ZUtjtFUBesH
y05D6RKsC9plqRWQiY8KtP5EcKbkbLXx3ozbticnNwFRIR01thpBTIuXzQC7P0gf
A4I/SpkjS+EcNG6kFhOiNgxSilU/B1H5w1IWMvrzbkkxl1KQvgOHvRgzuY1yNivQ
J9/XTaqMgTXSou8dF7fSSMfNucB+Y/gwvo7L1zAGAlgnGBndWqlbiaV4KqBHfgst
Cd+vPqjlVaK9H9uJqs4rr8D1SixynW/HL+IXuRmRU+j7Nevp8Q8Su1840fAR7FK6
oxx+prQBccALO/LozQ3U/e/kA0H7ybDsFzymmn4dhow1uWdEAc2g5pKREsWl7jqY
sDZbO6pLdugTFR7sJ0z+mUfp/4FW6YNILEht71QRhE/N+p+t/UnO7HyEQrbw8PGn
bXf7gmWGWG2WPYiIKdai1vxgxiJpUGtW82xa7nMTs+AFg6UZjepBCRXHwG+R2wq+
iwbOmWflHiHCUkjq9rCTRzTCRm1BJbVIHS0yXsEYHIwIi30Xjyh7KKK2MmYf1X6F
Gk1J0AXYge06HLL0Z1E0l9a7X9cdVpvw/ZbNMqNZNw11coh7HtBVFErs7r0hiHNg
TAeHyjMcfeOvVRymgTNzTxDRr/ZN0nFtyp9BLcvkoSHEf/i3vw7kTyurJNfP/u5F
Tpgfn820P6gvT0spVoDYRlt0uDk5HYhuCt2Scz75oaOBCrnxrzbJGUcwMz7cjJrs
RIlSZIbzs95UOtMEwPuBrj5ugJ3J6ito18QaEGX7dQze4RD3nKLnPVdICF77ecj3
ec2Ja2JRvrY+/EnG/Cp3N1/Opc9BBxxuXLPsAYT2UBfqmHqKk35BxifaQqksZlHH
4tcsF49nZlytQYLVLbdmiItGbwwVAmyg5xFyXnfbKxnzdMuNr1bYtumOmGpppRCu
YKYE8wCROncvDLE0rzWRm6vU3c1qLpdjvtDoF7wCqxPKw/0bvfrDTsuTUauj5Yx9
0EO/cSWqaX9HnGWCNDd9Iy+JuH95H3aPpe35jpChMflZqzgZLDPqZpyFxQbsw51Q
jTTO4ctAY+wckzJvAhPUd/qM98G9fxt31QZf1PhopMJuioSsOR4ul31y62OoGZW2
o3kvrCQDvrhCsBYADiLIB/739bfMzkxVfoFRw3p7OEo7aog3GdnmUvkPPVc2CpDG
uLHJ3znYu89KG7EV3wOBFfqW+AUjAs7rvoBYW5BsaJuxFJTokd7i2+jYOwI+f8gx
MrcMdmsbDGh7yX4NeuEpZ35D29/saNLg/DXykN7Yv+LYObAP+AaI/8BG1WbY89pG
mUoavLo/PbZEESgtsM9k3+rysZDLDnKXOmI3BoCijsIg7nSw6xFFcfauXpnY5epF
ennWBGJcTbWlBCEpoi3V4m7PEA0mYUMRmYnTCLfqG77rgQhJuihQdMocyEz/2DS+
8KlZMkNPaAIl8Y8QVwV7s6kb2Tck9gTMG2ii4GedMk/JoAheUgRJTABHV8/4WiV+
YLs/3eLpik+c+auslGQLxAjYIJAe4n3RJqlh6wYek6kRcsc7vsJQAggRj38lLw2n
ZGh+iSFvuU6pXfOsDDdHmhA0jdoq/FlgxjbOOteMIZrdMKieVJOC/tryRTUcVI3P
yKjEqO4WPFNiDDu6LffCQggHpHK9bk6cBTi9dcQbvIp0F6A9G9ioOUv86G6CVJZN
szXq1om1CCgdlX/9DT2r6vt7D40tK4TNecNRb8BBjmF9BtDmEvdPqpXHk7zW920x
ncfnzOlr/DBFOHc4hqeGkJLstTRPlttusJWIrQ8SaS8QidFH7mTetuy17ZtKGP4M
dkhIYFioq8jGw0aSquHdS9L9goeLTH4ExhgzCoDhezQnEOjyep/YCNKOF6ARuaLS
sUKpm6r6damKn/EdOkcJt9BVySkg5iw8mFZbkVFRJqP2llFLrXSamdguoeCNcLKO
/Ggns402jEMwQW51fjhSw+XC+rK08Ak5s5RyQq2l4UwolcoCmsoiGdsM6n4qfJoA
Lklh7LL68oZYetylNQLjvMlZVBg7qQds56jzkjaMzx5XEd67Bs9qGhexAoycmpSC
c/Y8BRDwBSIA+tTAv1vwDWO1ZtgvvbV4m1vaLZ1Gawut7aLF7Qmrp1KofkkRv1Bt
IF88C+iXQNZL/v4hp7SPyUjTT4T/FPt7hYQ4+rwkVy3RgSpUeOVMCXjUDc323+VC
yPHTRgsp6ZF4u0H7kKQMrrd+cPKhdSGbIxQtts/oruNNHVPoFUTtsB1VTiv7Jec+
poDy31c1Gq1NSCnTCbcAZAQ/KtDiOtZHFIVWDtC95QzEBpVTufN892IYoVuzk9q6
09qoN/xcwqpVvHsZTUkSSZFa1palaft7Dl1ECzhuPTbzqHHEN9TU7oWKG1gmwjHJ
qhCzMp7nq+bWK7nLq8dERqjbh9pxHcxz2PV/53q8g8jpyQG98iUBQfSkI85Fes8g
9YHzKX0+R35s8FtGRFt8dZiuaCIWIj7nUSEA2a7EVRMC1c7kUxBuklh4WFpcENFw
C5kvCn+om8M7X4tQKkGbjrFtLfZ96vPh4GDH9PDjeeb/Dz3L0qwVippWPYnuD5qA
TR1K+gq4zPpHnOmNi4s/JulTfsjkqEe3BAtkoOuCLjwsJJa4iG29fA7HE2UEY5xw
cKfZe0WpU7KqVk8frae2+sKXNU0ZSNmjXf85Q+lgSZ03ByDRL0wqbcxA+VS/KVOi
vbaJfCY9/LYYEO6LIDMxNFuI7XN5iSzKB+d5litbycePq8MbP+TqW15MqCQl2Xtw
myLQVu+WINkUQVz4lp2YvfEDK0n66LRrD0lfMTakmR7xr+G2YPr2VQiO640lr5kV
YsRKXeTmUKJlCWdb+oJdOtg87D78akP/zTsNPnWsZJJ2lo4ys+K2Unq/J4JvjuM6
8ys29UNLHfoBnjQio2owVHAJKIIX7Z8zvobEpLijy1LNQoU1wBBUGULO2XeG9S++
5Hp36US0K74vhv0Yr9Fm0L0QycMm9aKsI94WJ3WE5JIlMxw0dJhNz48qG+FUxPGL
NNlgoeHld+bn5p9/8E+jiuM8PUFfqt+4deNiR+6nrKBMTft0c/tUiIMIv9cJWkKp
9nt78F/4KzHVAsHULoWqq/CoQlixsb9gEURDvXxvJPLiCdVnM8kC2Mcaq+boAg94
aGcVa0I/guIHJ9maxQxAALIkxgvy9J4/oaCruEJViSPgvBbyFJtzwFYPIDUDVTl+
lTac6XX3t+l+vODKa8t/xKUMKfZ6a24cYgJcd6S4LzWkzcylinkvuPoPjIP0gsDT
uudrY8/8rwE/uA2Npvmo+V2pI9K3aDX3vS/yW0Zy4/CxdDGmFPbf7nykQdf7lQDP
DcbzHigyACRh5u45FBVxOuLPrNaI8DFcymgz9SeWI/IIYbh/QtHGfE5CKWrYcrcF
s32kwAk12j/SYDoodnr9JDTeiyOYcKaMMQjKmS650Dky3SQGtpVLYeyLZpV30rKq
sjADQge8pgASKYBMf3XXomIfjClX5TnPVuRV9DSB6VDJG1kee0cgES0LcKM0TmYc
MCUGWr7jk8P/sYRJ76aENECee/1XheIQWOGFX13AOrkGTfx5YTxM2AHIWeLGyzV/
lWQCvusDEsnh7W0Tj6gJIEeZkvoHRxVLS0sL3J1jHZOHcBu4xWaE+kZ2siU4++Eg
jHpb+/+oSIHTR62CWMbXBVQ3gIfq7jzJEtBwB7RhZV25T/5xXP+6TfyP0oqmVFvS
Ro/YEJA4gZNBTmRaokTMsKzSIblT4BKL/SJKOODfmp0g0v9e2jxE6pZHbanuHMty
NNO2qSaSThqFdafacReWe/BUFMayvTmFY/JMsgW35KKrGlnYDXRsZGS+1XH061pU
V5G5Pp9PeKfF8lSKRKetnuUtpIhklhiQucNacCsTJkAwz0Mhe5lqqWkFzxJrNrlr
5l87JqoLEQ1kY4pan3S5GSFm2Yl93SCQqoTJrjj2OA0kaK+MVMYBbWpDEdbI3JZK
LzXUCC5mx7tGIovz/OAK4au8sNGwAlrsapGak11mDtngDTu2Oz7c2Lf3aEaJigoA
uGBD2M66S9z0lLhsXnompyg0fAHC3lDzsVxx67Iskdl7B+IBYJY+nd/fH5QDwR2M
Y01+INWA8EeO5Z6phZV7eNqfbc6n3+OGFJwWBm2kWE/FC2WsliTgkLIwfVmIs0RI
ihnwogUC3j1xeaYW+C4Ef6yW/O++Pt2HThTdgA2+bXrXrYhYp0unoZLg7U+QGVi9
GvO8lpVTKv8DQBLvWEGOIZa2yjDA+rNlfaFGZEpYlnJDheRnB0f3lfjaRizgnlo1
wGF06FPkBu68vyeed6aZkxR2iZZne+L+swN3lwRxw0WqdCfRAMc4hLMUkhSQ9M8H
tZwparEzU3qiK2YjiWLNmpk5Q5gsBoTe8o9J+PWG7/v322bRqdO0haQWwe360ybi
h+N4hPw0SmY9TG4Xc9LZxVFD3zPLirz2mUBFBLDCtRfgMYzJcfqO0m7WPjQaWMSI
54JRgHd9qpAKiEz5pHgi49Pq7s6TiUvnaFop45TWs2gku3hCbjzuLT3/f9vwTmVA
CW9f+lQdrcLSfz0DaUu/AI1UYwEXkDHyeiqfPfO8b2nzdYRJnaZpBw/YiTm1i8+2
KUxLSflk3M/X42mJ4rwvE986p6Oz+moFocgIWHLZ9nZqBxd/N+h3EuVEYV5ZEbeZ
jqN2X3cSyUHhwcegRLrQGzuCAyemY11sNLL4mUbHbMgjT5C0qMcepiJjTh25iS6X
cwCEtO0AOIwXi3XAoGzr7hh7mjQR2aj2Aqf83a1xiQUUOnfTJRn0F0yRMB8MKE3X
35ZXIWqm8QuPSytbiRrYb+beFpCzXr/lpv/utAdWdWDzgF8z11l3kkvr63meYXkd
CYygEgS8lpLTET2VSo1pauIQvktw1h8pryoAtTqFxE1Gi7DtT6RR689uEuEKfCIU
D75NqcvmSzsq0AaNSR1EHiaGI3bCX7S+Q69l/50W2Kr3oHqMHvNz/N9x70o1iLds
Wm7E+bLsAxatL4C6gjS2Q6FOwPydma4DIzmc0cyHN83QcBg+lMHeRe+2SmOMwq5S
ro9to3lbDP3JESMkdqKsSqm1KGAFnIn7eRObGb9aysOIkOSbwfCia4+jUAWzM9eN
D55iaWhp3e9p1p21MGs3NKEmhWKf1Pd2p2eWV50pMKUZCXMee0nTxmKEQRqyShRg
n+ZvEudaHyp82b54wTDfLxpLmKil9BUF+X1F708h6Od65K8OM1oJnHHnQ/yzrUZ2
ddvrGU+AaCj1a58WAzmFJut7n5J+UOgItX5UfRopDvFRMCY0zRDsT0Km8eNjz6y/
kUVYz+zT5ScEqrdKl77yDLoxbuUCkQ+tE5Xj2bjCKoy5NVCNFJpwLcl0P7NFiQ5m
LlZ2oSuAU6tB0VhNRSCKDh/gZ3DOjHXEzR4/2kwLD6aYorBCzOQpNWUSFYu/gKY2
ugPmqqERwLTM/Mo28+CSy3HeyeIRVJmlE4iNSDgaPq0gZIPK5sGQMgs4/L2ra7yr
ckAuJBqVDB9c3RYCtrqtCpaXSl1/uP9O1MPXfJ/wjs/YgsfDH7Xh3qGW1bcj2v6z
wDghcAO8s5F1iaFArRx8nFgXs984ke/Co0wpK9UGHumePyY4UdJnNVrqKBk/FCYx
peJz7SY762+pM/K8EQIfaaoCwexQsfjR7ECz+hmX7IeozqEAnNR/dGEY4LdXep2i
pzCYr38FS17RxOlipVmKBeCc8WmkfUwIykD6sKXqpr6ilExKes57a3ZWdvJMkXyR
7hKcahZb3DxhHw57uDXfJQ3hdWq+zI/hBeMP7UHWmm6JxpbepkAm1hSlfTV/azgl
HRp2X0VeeP9FrYgjyv5he90+46D3agNVjxJ5pGewrIsn72eDAmdI8J7rjmJjB0uY
ZLDATzDl3bVhaKgSq3TiNyjK0fQfiaaZlM09W/ViPQvmfdjqGuRVYDeiIg9Qqd41
G6UZ3VMYiMKHEu5TYXWq7V6dxt5GV9DVthrgL/dsigsMFi71jYoSTcllHlh+/nR1
Xt/LssNWVewUEhPCo2bx0YO1x4W5Nu23PFsc7h/4rBNMWPl8gSB9dMaQrNZP9BhH
UdOcyG3CpSjKbdMaBF5zZcTe1fSPlo+1PNi+iHUgnmZCzbsTyjn2u93jdQz0Okwh
Be9RgyZJ2rzazzKEGzwrCBSce1D5Xsg5LiGuoOE9W1OwWU/olpMtzQx+IJsZ6Bhi
1y8L7P0zZqGywJjdtCdUikyTHiAFhm7hyovb7YFC5Frosa2szzD6HLhIoi9a/Omx
+L+7kJjbkLQIYLISE86kVdCmEsEoTSNOJwSygsQMaFS8NQewbBZkObHMD0M956xp
e7fcUwl7ItwU5hXfFjDaW75TJsDx0tDXHZYWOgrL4BxpOQ9sNkbukcNIbI6nDyuz
iFhXk4CLz7uqgmX+28CpyxIChG55j6nywJZLU6A+PjeVWZBEyVK3I3kCi51r8YkT
weibyedYnyP7vZdKs0QqveVOs51m5b5UA5kK7SXBZOVRQvGZWIMTVb+frIlbL5vn
a+FoJBkSXRfMDFt2ub5WW/F6xFTz5Pg+7gZeNSnGWQyIp45sip9j8AWrCtz9yH8z
1XtXSXKj41Wc/5WKgjEtS4qgdvTNdzYqRBJ7fXy9C3vWNocMTWoW+QOCxRna7aWf
0eW24Bn0mCJLsyDTl3oUndHLe7Mhvpw+hXv2EBW/KvOBLWrJVXRpsXJo/vexckV1
ADRPWM5iDy2hGNJkl2EGGGHwclZTmDBj99hIlZjVTjQ9fkp6lXt+46CSS0YApBdR
b8NLem8JkNITsjlhA51EJNfaR8qRzetD5sBJokZ/MTAr9hZDIpJ8dCXLv3Nc4E2n
t7obNy2L37NiqwcDUX4nUkU02+ppGCnTkCfH60w2ZINlR+SOK0LVT6Q5lhitBP1O
1Od9dITZ+beY0I0jVQjmx1xnN9njTphX7wlIiqQ1PyTG5tpW++IEFgk2svymV7tH
xtXYa+wtfZgPxM2wXekSHsWPuL06dO0nr7rjaHgZji2+7rum9+LwGdBcvDZ7uJr1
Y4yqXs6nCft1H4O8E8KWY/BmgvPSbp5fpfymsYu6hRZAAZMWHoy7qqHm9o/MbDLK
WyF4y0OgfzD2m5XBRy35vXCitQpjL7waaC79LmymnBzsobPAGjpFB6yoKYdTdlAn
H9ueYxvvcBv5yo62Qj6SCrComRk/XgiW81Ra0XDBaNAn7AxFTbZnDr4rxtvz3moA
4HoPvN162IOqtji6GfWUMDRSep5IlJDjINoBgJak7So2dTuSt3vtfHfE/lM1Nq/x
+Evk00yflXOXwXkrRQksXJMGgUpWoGk0pu5maxHwMFxsbHnuQwrHGWZxM2poDu+K
v79l0z3cZdTFFfM3D+nhBABVH/9CfuQ5dwhOJzmTVwxrruWntjoDUPd/ka8HUy4b
q/w033x+j5ZQ6mq8eCOnb1Mx4xpiO2fSA0FxQj3nUtdC7P4ppBw04feomJCoFCOX
z0sCPoW+HdWBSEoGNK8ww3UpLWK9VuNnRmHnoSZB4oaU06C2ojU+FrxTAkkfozsY
hwQ43jFEd2oDOpGblNO7fuI9IYO9YUikMg3EMzKdC3pLbRDHKclHatw5xHkER5Oj
Abjfi707Hiz368r9tQMcV6qj7U/yFNSQs2sLJrIcbZvvGyJCf9j6H8ZViiYIpN3d
QDk6yj8wBA4nMuBj+Ytq34XqkLqM+7cIa0kg9kyxaA2wUaZiEI6aCZOZEbMxTAdX
WViV0/mpq/B+G3IRvEO0hb1wfUoCvZVCBMAXI9cXfTEX4UPBdQk8qmZfrugLPilP
awqUGIhummZFhqtbdTpN6ErLb8zFN0LECqSQKm+Qkbc/6QvX3t0qxLka2ElWy3LU
hubH8u8ofxgNBwqYWnF0Rg8LsaRhBfc0vt4ESBXIqwBdAxVRoVPafIX/VFZ+NLDs
FDefqMsrE9AYV02/zoidKb+XSGD2NVgvh9qE/MdWn/xIG8YqI2oh+dKEV7yWZAFt
QpnO8Du8zDUviP9sI1WVvboIvn7tDH8eNAWGke9eqyb0XFX+pBr5h0g3zdjbLxYG
xoLz+uYvSUimEf4zKyH4WlVpvVn/gnXmZbT7Vn8NZSUTytm+h8SRARGzk2sRO+HS
vNG1lO239j4AT72xfbOXMHH59sdPheX2J9/He5dSFolbevkDWRF/0k7A6KoQX9zZ
ZJjbI2YGmOrItYO7icUb827J2u+gA+NGrK7EsPkdZF67T2fHADCTHW2F466VGGbq
3gCxIz7GV42Y7noZSrv2hll0j6Zhdw+8w5wsTMZafg90Q0u/cV0y7LIMvPKpSM11
ENgX350lyn2HKZnMpUOFDA/1R5PuzAFqgPvuR8UuMHPAEuBqXFhCkF5OhjHtq1sl
iAGx2mkyUK90C7Mqtf86WuupPy5mopV0nqIPTANCcc53l6MN55Yyg22tRvz1Uxy2
QkAtumhdcsXXU1DQFEU2n/Mcgl6/hC6kmdGFn3IbT/dm7885WqIzJBejvEcJR555
SssxxZgy8K0j5pxMHXgu6/lwjdrJPJ7brzJAx7h5LUy3PeC/0xQXyEZJ1j4wHyFe
exs8U/Tay8HA8fqyKbesw4jr+49LPY1hMspxyj0V6YdghW8P5nxLXqvF/VISRdhx
/Tdm5kxA+eBsNwXdyoRfTLis+kRfXBVXw8PNLmFzwmbIxHe84FC5UiD0fG4NRqif
GEGFhLKyy0RtfRv2sCLjIg0C+xeOAW+s2+IMrphGH/zO39iRWkbJNgHOZZjyC3Oy
K2XLSayzUTim9eGgOEN77Q9TPZhU/CZBxM6E2kftjJSCkRpjgCgRIY003KncDqgG
ICqAX4f2GCC3IIOBKdYtoIYAR5pIqiyf57JRyOmeGp9qUWmkNcLNtX7LMNmpZS7P
FqQbdkZZMXbdQoZYAABFz1lKbpScopR4RCKK8mIc47pAp4P3PwIbPD13A/+cEQjj
UQoQ6wnfRP5d4EEbn+VU3gfMMXNKmW2S3ictlOUrDeqvtAMZCbFok1miGBLMvXd6
PayFr/cFMKgu1UXAUBGxTHZywTH79kiLMCInF3/MEGyGzT2a2IzAVxy+E212l9wO
5qqfka9nQDWV+7IMQAKPFdzyKpfwNjigUvc0Ru2pbBiSvEkKr5xZC4XxKtZPXnBQ
ueIiD4/JsuK3sN44CnTrzQxKbJCmQ9HhypbLNO1XmMjoIS9jpGW1FpIq3OklRo/t
0uCBXSgoJvVhpHzke8OraMkhvQ9foPKhIfcQbXlaWgeMQpsyfkVXUV5hhql0rRc9
Kz14d0b9XhxpFQOkM9znKeyPgDN18YAYxe29r0GEEzf2EvBy/y2Df3y6gySM7SD9
U/tDeTm3FTbshoq0Z8D5VAWeM1G3h3UAokK6keI2svzvbTuINoqcQoLUtttEehnW
f8XZu3yM4OLR5137L+/eJxkp9SnfNfRwpzH4OHlkCD05Cjc+RAopmZAU9ph+Lz8x
U8RfeRFu0WZeyuNs32EgD6NFnNPwPJJnB4X7Ic2NzrzpY/fCakUtAEm4sfPb+E/i
Z0LDdJOoAG2xhfLVoBdNnbVy2R3BUMY+mx3E87N99xtGPUMCweI4tRKVk35iPXxK
HPz4N9x2whyUN9uCSgR+zI5zn8l82Jdww5Fj48NKl9BFWYZBTqAJqbV7IR4S9b1b
fCyrf/uvOQizYE9EH1/zUciABJBTOSKNDPm2Iao6uR+eWuCSO6d7aFilyGM05c6F
SsbTOzC2C6McG98DDI2dP9ElsHAEsUJ9y5ziJyqKTy74xZsEFMLIBZtyWAqdRU7v
3LJPujj6WgmClLEX1+5I596eKpL+6p2uHdNDC+Fpu4X8Vkaq9mrjlqJU+n7hjRKI
VGQgvK4VaYhIVWd/m3Qz/Rmf/f/dSlDCPEisRcOYvtzLNstnjLjC/rX/KTGI1715
8imCxhxu4xdRvNctdyx0eKIK1UNa8iqBo5VJnLkSWz5yXRUGE335+k/NRVCdDlyz
V2UtYJOAFuPd/OuinAkDqsB6hnIMwI2bC62g8R/cpiQqe3+1oT44QpcMwkKnvdWf
+9wyRfpmL5BKf4fR+4mVES14xNAmjnmkXgEeQf830ZhCxnFwGD073ZxNN6Zao9tM
QWHvkUZ5Af/ESTXEOWNjwSFxv5oJL8ATuSu21cIGgZTfdyMncaEf2Nh/NF0nkfJl
i1NfuvJtDzwuH0UjJrKQZN9MMCVtYA4aRGACVpfpx8xK84CXYoDSHmyK2gZgjZ0C
FvksFz974+HnIPqaQK+RdfQUZknG1fDI6KhNk7WZp2377e8hmgM3/FvTjS81/ALF
S/7eIIUXJap5Z+cm5pgrqE0ElKH/x46qZcjPWKOMsAEX9rJ+T92fdIcVau3/OU5S
M/peNLMKWl8Ywfjjk52048cYqNejEGuz3XYku2KeBxYClq/lgZwG5YBlrMi6dZHq
v+AejKyQfbSuoZpLPUaFTJ/Pze1QiGPaEPxJKVfVD+P0LILwnWgjwx0JY5O1pCr5
mFxnixp9tXYYefDcA+GZSCNb/IuQ11udMpj6+E3FuZ9ZYdIlecBie8rTl9zZP04f
3jJuBVHfW4b6PJZpLj4xbOBtngwFRU3kFYGu4efMa+q1yFfGkRMcAZJkDdLrvoNj
CD2v6fViOOzXckplLjPupFnpPJOALgTuXIRO9TJYgqNyat3vH6TAFVQsedXw11At
7WEWiSWehnJtv3KD5HY2GZZcvRLKpjBF/0tYwZ5XUsh2oaHMj/NEPDFMD8EsJGYh
yppTn67BTOhx5WjwG3rq0HKOZ4/VIR+czH9eUNSIa5LZ9e6F6KqUz3ud18zc/NP1
APcjT+7AWR5UlOTnqERgmc7amjy+u2u1hYvUpneVIUzmSFYonKeUHygAV6KX1OsR
2gdA/xT4m/3PpRMvCrDZ4WFkTeC2No1Sp1WkK27FKcKALCksuSVhew3ada2Wr345
m4LrboCk1uCs61wfud+Jbu7JU5h6T9jm9ggLnkO+gmxrl9YNzLcv+XWDNplJQmHe
O2P9PvTvILTzyLgchFDekOFIQTCqr49zLJt/hG3HOoCRMF/RGN4fgR5OL+OtQZ8I
OXiZjvpKJ7oqbgfSCGH1C+kW4isIgX1J++79986b3qXRFu5SHmgnxqNm5WzVd30W
9u/V88Z/zpzZTysMKMV1MnTmS8qcZx6A02pUr0X0EkiV+EBj64KiVjflomQtsQLY
jAnWLDayXHZhepk1FrjtgHZzgOg5+NQCNCbNkMw9pQgomEA1CBfmF6CFJIpmOeDt
I2vx5ls++tzNEQu+SX9Ok2Cixx1xth/L5NEffDEEcChaUpWd5TN7yfGtpbxtT4gY
ubHsbh8Glu6YA81IiU+z0D2V2tKatEyBbx3CbapViV7Rwn19jBK8PiyoWMXy40kf
ROXHPIVnw6tjqEos0ziYsnHLdcEACrF47iT43VvUfndjKYoXN+gjcxn7/rJzVpY8
a3Q0x0va5s0nd+5YZ59GIefMm9SLvnQHZLvBH3YrGR1ygfKgg3/ACTsI5F7BcJt4
YPegj5ANw5yOtbK5ZspqkZSRKTY4lY2O8Ey9wyxYaGznAlehdSS2X9pQ5Lr0eiGJ
Og3SZcmBJOjVHR+Gv3qSvZEXLfAD/c490dNtRuRrUK0SbLoEcHZeumJmDKifI8iJ
vQbaahLd66iK/o6I0KjA1q+VM6aAiDQk3x+RrTzHelLM3HIhIPLkO+lhbAQd8fl8
tzralzqowTcaJVeCwGJ5UQj1J52OHXOpQhLhIwL7lQJLe9tLqe/wOXtBYQLBZMfC
zcG0Ue88Cuw1qno27vDvSAzodk0is2aBOmqPBj6g933vAzUE1B/p4VlJfw47zk1C
J62d6ER/eBmE39JupqkHP61/siXEm4YiPP911bJOWpg7ZCz8dgVXQ5W8ul3FOSXu
BPqsBZ4c8AD5QgvbM+Nr2Luv6yta8vJTE4aj6sCc7yrEsJPD+hfXeboJ/HjXsaa9
8z9/qxqNgENlAdPHsf69pv4FafUFYX0dAhglK9aI9/b/o3UN/zEmOGrTdkbMTulR
GRVChVxkYopyuTuNW5V6IPfjlmtuyFebWRvBH9OO6D7rJlDuzqr7RTKR0UrnNftZ
VV3Sb12xUzJL7pAGob/sozN8pivSBpFCXa/Dt4hVoXEBVL8pPItZQioK27rcEWmO
Nkg3GLzf072iYvr99Lbk5qTnIou8m6uw9hRQQ6wI3KjX+j/T1vu3DTsG1qu98Sid
FKfl4wBAz4GLqUV0EF17Gefq8B5o+JkaTaqRNbmgtNfzkoRNrS6AXzSYdkXHIluE
yzusd89T8i7shxZ2QLWUReWZHPdMxsWol+QdrbD8hDvmEQcGJaQAOtj3woqXXfsG
5F9j59kwZ8bH6S+TE8jlVnWfofyo7udxgC4IXYn3Nm0i5JMBBELI4y+EBLiJtpJd
F1FP0wZPFFSlyDmPaABSic6IEvVlNPKo0lemfOZ0ySCd1YwkqKd6ykVsOeksgOww
DeicXZVxlkvtqTQH+Rb31fUwM1FeEfv0zf9Y8XhXzrZmSbxV64VC4y9ZTyQ+hpgU
lDtMXVjNYfZ7ZBx3UF42hNB3M3edo+q+X4wLOxcxK/Zk1DDEgK3LJdAsMo3USk94
UmesreVXYnJ6deM+zTlp/vZT0tCRVe6szG0UcT3qSTGReRTf0wigdZmeb+LNdZha
i0t4TIcbD2wsc5tyFnZOXc33cjfuuQ7ELeWvYHmzW00in9k0Gvq169kjEDInzDt0
XrqKT9oqKR2ZXcYZXikzRr3he1bVWKQxFnK5+I+1YzEY9PPIt0MOPDpWIYnZZWST
t7wWFlc/3HiYVoigLa+CuvOrHH/lWybwMOTfsNB1uDhwVj5FNSaxYky3x7qxet6D
w/HNMTxG8XOGwK6gvvabAgKGIWJF0OSH/GNwM+447inC7NRpQw2EQjHuULsotKV3
ZCCTD5pR5DQ6AsLYT01YmLg4w3IaTlxz1Hz5qNtsLm+04NWHTcO77ThSXILx8yr3
p1b16/dXLZpW6qGBgrRNfJrjRoJb5PqrKuMcoBzF8iD6PFgXxcwOBl5QIr1FrLAm
lyqsmbqWIbx+6pvHdoFXMSTgo923M3l8og+EcV0FAaoEA9fqyAJ1no4kZ3tIeGcE
O4xHGmZ7neee/4rBkyVz2b+K7FCISoWU4V/2o3llmoAwzUqMNB55rSLcF0X7Xc5m
/RskGnbHAVgbKxKBXexA5O2WEUD9mDmxTmtyX2svSG+DmTyLufuhi5DV07N660yb
5EZ7jPDnnOFJT/eSu6hk9rs9zaO9/JAG+TOkfQJDd4DnKULhm2PqPAnagf7jV9bu
4MP/cZIxXMjjbcSCkqIExNECyu1nMKd6/acmkaRuRZWkOpU9R4YoBuVs5vRbDd9e
W3ESFsXR52U1e6vcBL7jDu/7nuKehkGnMwc18yRrQGN88lnOAgdkFjIIDRF6R2Q3
H6UEhd8qyUxGwEs6lPENOnqtWu34jeFBxP6UR9/jXkuJkwLKrgfo+Z2KT5Z9dTym
w6eFb3dheN6ymTV+2SunQq9EKeKTBqRaonLr1JMxLKbylbnsatdYBOLQ6bArfgHL
yDSMzWjfi2vTkU7UE/pGfArTz6P28jdUyNqiOAqy2gos67+raOD5BKJlYT2N/zQC
mmFVtjtBSfyvdEXL+ywAH8lUBSev6/m8e+wo2anmp45g7d1tRfZ4Fo8WJgFl9Buf
xcN4GZkdeKlf5Q5kZ2NC7SuoW24diohhXA8n6U18CFHx6HWd3OzrDhPHdvBuzit3
TXert9gQYPcURv1nYL8yRm8VzQvCHtYRS9ohE6fx0RHhqL9ZRpYbrUe9Wd+/g7OM
b9lj0o6bD2YwLOBzDKkys3i9ksVV41Urn5hXvYknhNDZl2kGUJJyIukvfAsMJSRt
5YI/IaJqlFc/sTE2UoLC/8/gJ8GT0bI8+KdTtbFxzDDA7VlUj31gGZ3QNJmY1ctf
5UevSAR9eq0zo45JDB6WJiFvCpdYbaePrXov23cqtO+j1nwBolibBHDWJKKRos9c
0kylUppx+2yfHRrsD4KhTqpK3f8G66h+CIK19L7WDG7R2YmyQ0G9ilSgg8mypo8z
ZY+4OmNBo9MytMWJHs+c2ROSIBE5Ma+/CimAxO4yRlZXgMwlgioDxExUv0jUhKMa
9eZfMTqT3BRpO62ky+q16jjDI37fUH9c/h2iUCJ2JMdrOoDu+to3X1CLu3hDHSnY
ZhBd70WyRPN276K3aBoOn/0tpwEMvEdDeZSxSqU06amINgp8EKZtKQO0SSq0zFfc
5kSA9esle2LiwrJu+PtU9PI5SsShRtvvZIZYptoLAhcgOo+v+lTxER2bUpBL49qC
GOtVv9AvfDPFwDQUue3NUVcuQ4qEXbeLyENCRKnmMXQTOOgy1kabj/qCHbvo2Jyy
bPVXam7/+vsUoPjICe+CgCdO28ZEICiJSqxsP7XbsJkw/MWrPiI7kES6121nIxRT
OtiRNaQNKwcSoNZKpPdm0Mfb4PYYfjC2tMwlbnAVqZkfdrte61BqL7ClDmho4xI+
3H6SIwVHRMKq5xTGFre4N1NAiHkYHLYwEyt3OoHB0oyJcBS06gz642W7/mVgK8Tp
rcSypCu7cE1acddeeefCsCEqMvJxbiJXAAUe9nc/Ij3fWBYCc43xL5/sXR5B7xKm
N67Dq9I39o/JYSTyMy97sJJu/Ld9L7HZpQIj1p5Z6k4tcwz9gaflaf/DOJ9n5KJV
+CCvjCz82QGohJ3Z958L5hbfx27x2it8K9uJPXcnkdURVZKiS+qyn4qH/ga5RrLq
X28OcraWQonL3NRdkPq57nilj6XXpUt++x9W21UacOUxzwPr9VsyjBqke8iqHLA2
PoJLf3mkabizdyJ1POt7oTBIbELKDXv3Zg2V14//3m9ufhCEG9/ht9tuPJthxOxk
PvFZYKRsxESOq9wDKmseVdFepR44+M3BR5S9KmkbnQts0YaTsyDkqHPVEvxM8KFy
8uSeJL+9fcXeQJdq0KutWMOOB3gQ90ya2YQde0nmS2zhgr4h1ddztSF7AEv2i8TO
+PppUL7nncxJJKdt3moiwltJPAzr7nh3ICw9KwAYl/TR/8frOB1h9Hy/W6u97oP8
BVATd88q77ZkwOO7B+Cg0vcNO4k4vvK+RBlqFHHjValnrmzZAYiRbgEwGKhyzE+i
jopJul3wCOcjMydXSlpz8widDbd0OwW4Ed3ueW5kMjheudayEqnTbcruOFDaOHBt
0iR461v81g7PZjYA1msIA7LlpgAIGIAvwD287emJLbXw54zC3tyvzcS/yY2euqa+
8COoMcrnuJ7/tNEdngpZfAqEIIf2KpI26DGzXho67DuZzmPHTsn0LdXGHYZdd5VJ
c9FaVgTIwYf4mO97piuden2aV0GDycdToiWUNdFCQRHXsKJ1Wb+IKiUi56Zfe5lR
ZxIOhy0ki96x2QobP/xnKTslKydmCIknrcT3Z8v+PzwHnizLk0LR1244zPp2eQqJ
xHIZfYT4A3Vd/dniuma9efDtS/BYGok+lO3rEyC0ijwtMt+rmV4z4gDSC9zY6WnM
0KNb41C9FMKxbY5kuIG44i+KsN/hU9/BbKDxHm8XkvgVVYTX34jdWv8k2acVHQ4p
FdOyw3JOu3yqloAtQliRFgzfPPGjHkmwrK1r1giTqf+6UIaD4lLv4Hr5wQ5uO031
Gux+BU6XKSNSiGO5BMNAte5r5X5Mx9OtiHgF+L46qYaHsSHQR7K8E1e1C486KGfV
1pXcn5fOc8EJ8fNGXwnEZNOyLHa67Mo6jrMrhzB04G0PL8DFJGSyboWIbE5SpZF/
ByjKzEe8zTbH8nUe2XDM7ZqtnZqBZ2YHf8WJPWXtxvkwHM2QcYseE3l8xw6IgMZr
wXyz1pGAfn47KKYVfJ38MtLnmNI8S1TuVm87h8tWG9PO3Fy84puCHPgxAovfQ+KL
fmDcAO3buyVboPxDFheav05B8ELPT4DoHeoN03u1DBrl5DtUFgUC0UZVElsuVm0q
3yXX0NplJgnJIZEzq31GyK8uTKh6YQd/dRhDw4J4gKOnHkwMW4h+kWobMgemyyAF
FkTg5HLo3mXGA+dpy+x/3i9rqyULTpj39R0ku7sNiCXVL7ZoN/08UMjvR9Lc87Qo
AJrve49NCEh5q/SiaJew1RyTlbiZMPf6wcHlaPrBFzcOfbeOf2JhlxKpBHrKIEX5
5HnOa4W+Y/a7nLjaZJ1wdzcCik4JZdfb0YfFW9mVQ3TtmNHzVOc5oiS7UOHCoQ25
HnRmULXeGy4vbn57vFFEcA3FK7wViE+01Z7PQhWkNlVf94vqFJo3hWPpU6eRfJo5
otk8HbUyIjK4+3zTaalYk3uSqymMOtMidDdkzUIJ89Ip8SD6mg6Xc2FJcTP6xNAe
ovXdf6WYfb71Z4qItZJZa66uod9m5OPs9uukjpT8YqsmQc5N2H18yi8dFFD6GLVo
wNu5XsgUHxt0gQZj1PRiKNnqsmqERbI3hrwy6tXVbVUoYOPfE21L/hbu/31VewiF
WGtXWVQ1K8ZpjOJ73vmIhU+V6hMKIjvLGOUFKaWAC55mhLgPPFJiANbxJ5uTw+QN
oWIr/B1P3OFl2mztqbFCS1MyWzOQAZsxkQwaCz9s7lwZ5YaUIm9PhE0po9VwSkTV
j7m12JZEtpJgQh3xsoyW950dPnNc6zsIvnqj5poSSh2Tsu0tpeiSB7BPLnsu1Lfj
TX4ANx42Le9HUAYTIkBHKaqH+Bt5ru8aFE+Y1Fz+nTC8H7d+/q1RD8NbLD6BgqSx
vInIONhcrLWm8x4W5+IxEcOyq8cVRUbPMrwCci8k+qlFgn2hZuO97Ro2rXHUw9hk
JKQzXWShlBJ1DGpNRSdLetbaBWBlAggFdYcrOdPOIHgcyMRqPpFwGzDHvXfFSw91
tOEIdVbEyBZEAlkFQk9q2KMnMtPgtCNJczIaFO6wd9NCCejKdK1ORnO8FRpec6JW
wy+XUZSd2vYevdt1CS2nF+ZK5YMi5nkziScSkqAqspp9X/ITjD+T/mzsGpk1EinI
LVTtexDNE/jF6jhAb3/SNYXzErZJfen/OelZEMRJ8lHYad30bFvNcDCUiukGeh9+
uov6ySn76lkfG0x5GGwZFmS3gJ25KB6Y8O0dk/NrKEBLCa0NCqEG3HSesCL1O2w7
S0mC7qdnrmS6hzZdGfuZ0BWOt3XyA8MzhWytGl7AIOjFri6PKEZgMwQlyUW/nHBg
lerFqPuYiR1Pknp874GF4JFEN8AKEwC+tTnJMSU7h6x4gXiXoz4zMRIAcmbedaya
4uGf8RhJOs3F9rpv/F4huEpw3zpNCSwqgzur3gcEAIHn308e8OcN9PrnW9B8cs7p
FydF4RoGflpkIr20pShQ8stq4GctFMmrQD6+7+RKRvyz/TqHUTTpT5k9wq73K9y0
3OEdkAWtxDcEEJ9NjSWIjNvxRzfU1gKL2u0SvYww2CvW7NM1N+zoweG2zm1NihJ1
90RDLLi3JOt1HaF92S65ok9c04jIFP0Vrl9qo6zbCxQ2zgEn0ShIMknUuCOIqkUb
LuICGSYoCpYVA4sU9RQM0N0qdVy4gf/GpMtjoAtj1kpfqpAHlC1n2vr9+bwu1okI
70MPKJD2/lPiXBG9vjC7SAiZ/1xxByzHjsV5DUz4kpR7NmR/iTx/X5fpbih9y8FD
7FsvMIqBdY8oezmQgLF49/W0uRzc0zogya1fz0EnFSb4XRKcyCppPWkVvFQjIkk3
MQV3IVgCMaby1HGZvsiTgsfkvVaTXB1vkiEbzH+Nd6raI8U1ELXYdB1bZDG4n7+d
4p63owYljOHNUkmnwsLbta4sObrgeDpxaewqJBegKILbWP9xalPL7bR+qmtyU0E+
6lQc+qh8AZO87dFt0WZ89DxQKOjqXv72B1NuoRZRFNw7QI5GA3WTVEDoBnfh4Mag
uoytAHVmkxoQMqhxRZP37SLKwWWoS0YMR5EjhwwsASOqcOkfMkwHhn6q5Cg4W+pC
+rAFlg7R2XS2rhdt3+dA1sd/BErFcFJBpKK59PWwEBFlH7IOH13DDTsjd+4LiemQ
x8azseG7BxKHVuuw75DWvdp+tArdrGj8rgZ5UmzYz2I8Eo9ZY4Z5LbfsblNQV+KC
lWp6hqB5BNBbETlFZW20qorspiG2nK1EW/cHOBGqpcrrpWgl21y0QgcdCxzdIZg2
es+QwT3Gvei8gOYFNmJIfqEEFthKJyeLdHj532GwSE128sg/gCsFaccNtGtjdVEE
gvdbRSG2ohCwl3UkUio+UCUVaLcUm15vgzoApHagzaJr6YeqKrfycPXrdjQGvP3p
J9aJ0+GAuU9ApUz1sarxBMUsz9EspBdMBNtnt0N7G9vb6Gw+bi8GduPMPoaLcIVs
iS2S4MyLMHLhnwQv3C4KKrITzRDo8T2pTt/h8v18PDQzWtWeNc3exiQG1hzeIL5r
4/6kgf0bfEC+E1s2XzC5dx48ZvJjRfUJO3CBEtFRTlBdQNy2FHeV0dFmmsDLdKQ7
W5sAkqyFWbaNWNr9ubKwE1Fz0Fxf2kIslUzd+3OatayquT3psd5COhJd3QS+TzDy
IoFnpIxZgK/7XYjKVsQq+SnkSakeDM+g1g3MHFd2UJWmSlof5wflAMQjW5VI0Djk
+mooeJ9wWq5Yf7U2VgnTken5SRZBgB7lK8frdENclEkW3vPPgPrVebevxHY3/1YT
bdQpCov2KgOHbfeLYBiy69MfxeiDQWhubPpng5CFN8LhWxaQNChR9JZB9TydifkP
+ndGVNP4FSdEssHxSBD1HM0ElfXbwnt9mx9p3LP4OQ6iTkfWtWeVwD/1aak7fHJD
aHdjz++uuvr7H8joArzGmN+AtzaBGSSby0wRtiXP1kIHple6SyzjKe7b7pAP1hVU
eN44+Ri6jOZ1KPF03Ej9oEu6NHpo41FhEW8j/nchIotD4EbKaOCiSB6ZuQ5Zvlbq
T1Jy1ET/tHjk0xhSaCzqEdVO2NAI8c2VxCL4buEhN93fKNKHGwmmyBSWAXcBNxyC
7WjPAGDllaMWfRaft65ifP8k0vscMNQVfBi57uC+K7mBJBDEaMLXURKRnTGSu2Xo
yXw7Xman5lQCtLU+SqXr/jGc9jdQgr32gdhQExSZe2l62Wu1ddo/jzxdaP3tqu0/
9XJ3xLhFwEzuAqao1dv80bqOR8sl6APpT77Gnsrv5SgMuG6uOsQr4JMR4hAinZ7A
1tv+OPV/kYosMiPArVxuC2Rgi9+nisSHkwGjIxCKnqUktft1oxC/n1PxFQVdVWWo
kR7V79+Cntffz6EB5RcfuqkV8zTYuE+txxMIEDKBlgJxBrMztx2S9lFTmdH5tNV7
1Q+JlThUvg41HZMeLqV6GlsxOoCqccuC/eEVJkjmLZeqRs5T+fHCzdyTnIQdRXxa
ChEonHuuZgQ1gtbymn/jZ0trLUHzWqfUJFmJAjJ9VCfuKR0aQ9hSnJlIUQaW9Mt9
6lFnUVX6AEPVnFvjxHWJPRzRzUFo2b67Ald+Tl/iwM7fNSAcJj5Avt41R8QhFDum
YZlkOpLZtBUZnBrOKzECkBRZBb4QAaXdbQKHdN7OsfVRty8NLaCgSW4IcMCUCTkj
BnNgIEDcaGifmP2LtJM7yslU/tQIPcWMK7piVQSjIevMzWuPSW7jl4rnkasFzz2+
Uod4Pfa1sGgUat4vnsPtnK3WQ8n9izM27/lygL+P2ZOPWQdUhYyHUFQy2Gm0/nVH
HKT3nPAMsd5tYMo4SL20oAN9Puvqyw3UAC4eEojv58gU9OqivQDSj7w9WYrhYghj
k8b9PVj49XQrBHHMWzLL0pxHxtbV3QVZz4hzrELRV5g5iXlS5ZcjAB7ds6muieT4
13Jrg4e9jtTJnxXS2uHisnJisBIbwVbITi4BaN3dTi13JY4r8WZfYhvwL47XwQ1T
dRSIPgf0A8MNX9pCb2SDgu3JOohbM2m2NInT4yv2/f3IL94vb10RYIcB9bV7e+gy
HlXkajlyQ57kzh9O1qusgFPABwykkkbGTEYttj0J3xzVjynBdG/LzxaP6JldDEXR
TsHdAcXl1loTciQyFukvsuqzM2og9S8wG/DWvtEJtsXZsIHSx5c+B6rFTCPsVvmc
FLyCHOYvGf65wJOhH8QtBYrNGcD7y0ChqAtoRE8hZpn2x8E5BAnzsAb3T6wyMvjz
P5OBSwWNOg/2Z47IhTDeXeVlh7PlXqNAIJiAMGiSIGqwME5ONmnCApRWsok6xVsR
9iMktFCSK7tx9egnFcnpSxKadjq2N5iDhvx19Vvhin0naokLaSKzTDJP9IwgIVwu
kfhbQ6PiIP0+mV4rwZ1m2u5T0X96IPawALzx/XuoCjUACwRB1eE7ecExiC7T6CX5
PsEKWSfM8JPyGcQkiBCEriZcth2m8dSr9izQjPCePzJn8ByzyUgz3uIO+YJIdeHK
LFTEN+BpiTIi1MLNloJLaZD9PwbRuKwoMkTuLPIl9B8hg17IMmcndDOBNCBoJILF
i4ppL0/FJkrWiZhJb1yUJFUGIk/ZIZxHTO98P7/N6HnosAAS9Pnoy51ijaExH2mS
D96PvtbZCwQSBPhMBO9ZYw1azFC+JsBYDyCChjwyEJnN/Db6uFSpj9S3QOSusPug
G1ttHNAVPIGtZiCAL9W8hULkC3pVGCAooFxTEZyl+adflX0mR6ZC2hzh/gGOm4J4
9JalGwOTNgGYoThG1abAeZGZ9VJAouI41vWvPz3X8Dq8bHINZVbKkgjQDrlFv2Ir
tTPA7QMapU/ufT4RNkSILpqa1vWdIRDIw9V82ktBA4QLWywiMr6aKywSc4DFjLpu
BDQxhPheEhPxPpFnEDZM83y/JO+oE1x03uqKTvqrPVxNbWWpm3o1jbFL9ROER8va
lhXgRf5b2GfPZox8ebVPPlnxoln6Pkx/9nK5sJExij4laJwwhVLC8OzXEKv4aoi6
uco+D1N6hMF0Q9voEH5Lm/zMVEJOpEvWfW8HUlQ4IyOPTwmOTxp6TcGVhuY8Le3m
XQ93hZMwaNWVYx9MZUC53ibLACH179NnvpQJd8Wxb21cwjqSJXTScDt4AKibnUK5
v6ts6aH7hXSJU5DxenkIMac2rQIqXQPVFG5nbmx3i2rFP4HQdKMV8vvrgATQwkt+
aTH374OQO14giDiCEAsoMROHFRI8kGQ6RHvzIm4ANkVTN0I9ZSjMfY6IR/JDfC74
MikWUiEep3D4EFb0PePr9hOc09pIOB3v7VIFcyEeavXRbNpUVx5w+SCmOPWn+f0g
QX0T1wmgICKMHNJ5EMm5v6OP7tYxoqhg+vwcXeWn4ZLkcCrxw1J/0OGBN8Es201i
mokOdV1+/N0NsbGtJ29ztSKLJi6OEOJhmUVHJLMorNrsdkSWWuEZ40gmzm0vrZK1
VYUk7+TbDf1kl9PekO4KljQ+i6Poh572fV9/c1sAI1TmDx/2s6WjSSBJaOXpBAQ9
rDn3JCBHjzvaq6P5GEstY7mxsq2MZoZSPcjbJPv8sqbFucL0rqXl2Dp3oYprM7fK
/dxnFxe5PQlv4hgv773M+VAt4gWcfDAOmG8HUQEM+VpBvk2XLfNTbfz6BWFMes5R
4a75lQRkzkofMXNXlC/qgSnBlN+tHWnl7p68tY6NnkdTryjEetj0nDSaBY7OJxqQ
0Z4+RoU6S0FF6PbYB7N5zHd1WRLMAZxTsjPbrBRqiol+RZl7JFeBJORdRaVxphbA
r8a4KAXDRSqgf3aUrlnArugmZnznAmqETfIlDR3hYL/wWKwdvpaphV3+UcAUblWr
WCDwaMO/+k8aRVxCJZ4Jwy6pQ8Dr78xXYq675YxO022wOdB3IhPnbzF64dMsMwGt
0J7/4nRqW2V1DNAdltMz0UJ8YQFIoBE6bvXHiHscBRMYqoR9H6s10BG1ykTcpnKX
s6+IO7UuS1fkoEYZ3Ou5g68rK4aytYMoGmTNUJZpihCgEVIfn7P4GUI8n7qzixHa
eagwRs93ENAt+yergT3FNdI2NRmIwO7DZHlea9A1O6yF2l7TT+Ul/jSc+QsAQChw
Pv7DALbkPX4VCGlZuevoiEwaLdym29sFpAj6VoF2oSaGwsl+JGDw7ZZng+nE+JP1
ijQR1V12jf/2TXpgojtOAB5yqF7pgJzcVWB+8XcNmriJeM24B5gaR553AeRT4ep+
ZkJfNiGOpnMT67tNtr9sRLVIU7OFGQSHA59pUWuOQQn/5W5sv3DT1sGgxw/EFF0X
HOz2x0BdoTB+aOe1Ijqc+3gYM9Ck4XIMW5qZDN4IYaWJbR9LqQ92b7hdlLCIFjAf
OfQ2jQzEOA0F7EOJK4FvaILqTb0ceI8/0pEyMoHfue4GS1j6ch1g6nqICPcAD+e6
8ranAUC/1CmsjiscRjtedmL95zkRdCbUC9nbU3VtLwfBvKe/MP9Z4H7CFzGJUdKH
hXcVloHXomz8zP/89zEWECykd3bes0JZPNqZlw/htf56fwmNiKZQY2/6XZJOary8
jMANdy2ggRdZJ3QZ2hBUDLFRDL6OHa7eY9lVQHCx3FCevEh05sMH4BCXG0nv8kYQ
erfNMUclQfSNyucbMxvV7Olj9y96Jyn3tXNVWQENoS4iSzSQ6q/eUrc4Xjm6tCYB
iP1xBTaJJPS0u4aqxm8Pt4LD4DgdcI9A5hrMeOt8hf8X7P+l1UaStwBbSHBZY15G
5SqrJuMAMy0Qx7m+KIxqlEOmgoAQQtq8nQb9a0/XPudhewgvm2aL4rjq0nWYT4a8
mb/oe78fKPMbloDoaoNhQWIH/Q1a7sop3tQ7ZUZP6iQnWQ3i7VcW67OGKT5MdrJZ
A29mbAxXorfLCeg10Ow0HbCZluPBJCoG4tgXlah9aQzJBRfgu4wC+87ddC66AsGN
TfK3/g66Sccv310EL28Dls7wVCgAQ02opj6k/Amw+wUQ2kW7tHG8xePCBtup1w91
VmGhon8EcUkzVUk7kOzNwRDpjPNCM+MbFR8XoF8Oer5Z1f8M1naQdfn3nY20b5Mf
/2HAW9+09NozouCkbFLV4phMPrADgPIc6qZfUsPaLocVw0Z9ZvkjKbKb3ziiXQsw
EmG1ainVaFX44YRxw2i5VSL2x8BZKMl9Dpwb7reahb5GIY7nzkIxmsO9fRB1sAdV
CfeWoaNZ/xNcomXqwL5C9GOvi9ORrbXb245Tnglotm1CZRT7X4l78VwtpwRItXlI
oKYA2Hb36/SpGQXic5Hk8tTX0dDtWbwFJMWqldIUix7Fs4XeDAn2hEj9jRBGnrkk
f+skD/525ZYLHR0PamP0pF4+hNmwXbNsboETkOVAJt8idfTszWj/JGcOfD6yoz3m
G4XDG7H8VTobWuhLU/WGFxfYIr9arB8VUCUC5pjIZ6m/yyR+lKIAjIDvhMKx9/Ia
RckTiUe3s7kLarQ1Yi1ZyyoVJP7J3I35fYEXaCH3AFDC362/HOVKMqh3E6bE3abn
Z0ERtGbqEV1xfPfDey1eGZTvIKnnmLNdnOOdAD5R5qtNNXXnrkX9OvfXg9NkunNX
T5cn/jyKCtkftxz5ds52eBRmKSgD9bhKdLhAlDSI0tIeoRc3E4BRw7zMa9YM83lV
HfC6DH+QUySB5kGyuLUKE5t3t58n8aBg24l/FJviTgSE/Y2kNS885LdxFwRL7evx
YV1IX4s20r8/LCC8RXoIBNr7Eo8D9wacFcCzMR2drU4VwIAuMe7ZSQW+eag27RAF
k9+i0QqtDbQw4oWBbq27Xn2AZKKPN665/8XUzVhwLrT4F3kwmte9d5/+SybFQTlS
+WhjIh4w7mEo/s5V6tw8C3q5GjDf6ebPEZz/g+Vepcdruk2748cx7cAaEgtDh+Du
v8N0CCIm5sIi28ux06fzjTcxwx7cDFEEF2TmEJl9vxJamMO4viqMZdEuueeBM9EK
pLMKnmHgCSaboERq8eS2SEZrZwMXuuvyXQPINgUj6QKYwWNSh/Y+gDt564yC2qDC
faxdU1xLqFpQSrQj63SmEz4bXLjnk8gIBPnab4QjFeRt0X1pev3Gz9d+siIxg3C/
6xe+0r7jr+HAAzS8ScWh115q/fHq0aR/vohiqL25oL/Kbm3e3f3Xv9ndZ4dRt1Id
xSe9loyXt3B0+K/YWyAiGyRyzQ/ou9G2LaZMIGrV8DWtzarZS64TSW18Bfp7OE35
2nraMzwNPpaO9GLX80L/XBYF3AEalze3hnOgX53mRWMJ4w+LbYDlxR9yhl/wj62g
r9nl3qAws/AHfy70KsyiB6nwyl8GtZrICg3aLPOqELo4HiiDPiVqtBBwxoguiEZm
jK4Yuau8hGOtTjD8GXJF1MVJrZ8zsSYS0Im8ZDjbKSaLF4F4ZV2qmvHEnl1JipZS
lPnbPSDc81hZB02L+tFHC9GY3IHOcpbmXi986PNm7nhmiADsP7y/XvDonYuX1htM
bqbKG/9vji0a9bFGb2rEygsHoXwklaNhn+2MtPQ8iyBtAZuXmaFNMf+Orxv/6R6d
GfOsSuEEeDDN9vwW5vjTZtW/nFu93PYxbTLGdl84TaeWPc4oehQm71oGFk6AxSdQ
LWNRLglJXhaobXwBp1NQHlyTcOBDdMLnCaXjUfOUqv1+kHfiWMYBtrj2czEyWcyS
ERFqTcJk3Xgo9f5d+so79cIEATs/SRevT3xtm0O1xd5am7DHzC16Lgdd8D6ALaQj
rkKgmPo5roru12i8Gq61UfCy98tN8E3tr6jP0T1HNurYQoPY97E7RPC1kGV2Af70
NlL8IgT33L24Q1tnax8ZEoOVAgjFBSJexMp+HrsZ6a3Up0GEN/TYUieM+V+/RD+q
ocP4z6HJZlVdiZh+/d6kBYf+zLz1wG4Zqd8BAVAwo9EYGViHMLq52HnJEwPi0c0K
go9vj2I+VlDebVlnCoCShsDTHDzlUGtLPY/4tQFljonqnpR2O3+cPqSJCYo43eTY
re2mupIKGuLiUKaNQ8rD3bninaITcOqbexauIZEsqO8BVZW2ohtM+U0Kr0vEEPCm
FabxcgSRtHh9XE6MFjDbuRxTMCtm5TZRO8IXOXJdDfslr1TDOrk+y2CHbY7desZB
u/1Jxl+jHVrNrkPw4KOMXE+qLIOpCo3q6h5tZ4RbMEkGDQRRrFyy2c5I2Mo7t7h1
WDs7UBPIFw+8YJXQKfz1pz+oHROxrlEU3qmP7EkfutIoTJ7HG+J2nKXBDNNsSX48
nysDqgcA16kKvdNbs/sRbtxzSEP72Fjho6danr40tfLWoes6v8hXm9OQ6jUvP8+m
wZ6ZkWahwl+OubvReVF3kKHXeyPUCK+0PsjBAJ4egn8P1lGxY/atk6/iK8No3Fmf
6tdNhPcMY9nrESWLBZrMh8O5GbWJ5+HATxI9aXd+PBb8pi471Y9PvNyzUgl73xJI
oMzBra+dXWppmmJUtkV+l2rgvY0sYtnCLMYUXJW/+ttcw037w1k7RCyDy1vu3aFL
BDT2hVkzL9GCvYDFF4vv8ow7mEQQ4+gzjoi56R0z6FpazeaD0VoWv2yNeVTbkXGH
EfkjWobULP8y3TfbeOCdCW0xfEyj+gKLXLuNu/59Fu25sZz8I0Tr1BT7DgYDsSAK
zhojFMVgu5HgOwzS6ZSCBIx0oH4B3aB2urqPyUzfBtQkgVK4F4BiNr7G9M1Ygx7n
FFGtB7GvzCm1rGLzzmLmnBjbY9iGTBDnVbF9o5WpJelRP+K8ADLoW0urVrifcyS8
/qis1439b5yscLECCpO3bOe6nAGV7arvGrXab6PUuuN4a3a28QgCGFXr/eBskemo
LUHBaxpcgK+GykNw3WI5+79As0XwurdWiHwnNgXkrVuS7Xt1o0OVDNiD5hy1c0uA
O/x/g2XM9nur1sDGSMWkkt30lz7y0EpPDVt3rGpgXlkMP1dXglbzybWGVO9TuGqL
o7VquA1lUBKS51JzQRDNAWHGCRpEILWZ7nhSLaBaomlsuxdHCWfeffETjtBhOhCI
GXpl+7MqECwjJ2/a3Yv+lSVTaFoIDYZsABeoe2kbL1tMIal+iyFW2fUPXGIJob8r
wHDFY8WXxVD2ilbVBxDHigLDRLanoKrQJmTH+7sAJ/8UDFQXIx2tORWvX2oUr5+e
x0/WS4BiqUrBsVqwXC4tTkFUAJY4XUAp1y7XXf0jfE0NdQ10ULm4P28vcerPsnjF
MOgmEsCSya6rhuyjs2aV8OqUsuL1fZ1cC20pKxvK6ohOVq+MZmffeCW8W0DNOqOL
xNjCBGrsIm+aFSVTRZh8l+W8mG35NbEOILoO20ioXtRSkgl6zq5dh8YFGncizMzv
y25XCjAArJd9SADUDpu0Lm15G1lB7ox5b3smJOdvkyzOb7uU8XFJDFuZ5eUsZ245
KK8lqbYwH4AgEqnG5XSXIl5+XUbWMnf5k/geD10U5d7dt2JhBiikv8Xobs/ZXQh2
jzRGghkbV/cx3BmDHt+L0y9TFwJAERfD09y/zG99dz41xPkTAiEhAiZZkxMFgVza
OtdBlgT1TloNIRIAZOr10eBO5CpFKKdQPNVymIdjzOiv3McA1gh5Gbnj/NuwOUzZ
VVPbczHexwyQu7mBXXldfJByZd0S+1O7EpyHyNxS5xx1qj4A9UzuyEX8h1ee+QW+
rmIGOl6+eZmX6fdRZ0NXiXk88e8kpcLdPQV+cmuYwX8Bo5CsyYHTnGewBXEypoQD
g8lcM9th/Za0DeVb/rxqP6g1wDlmrkgtpQZM6jjDURE1al3bUu6rMB9sTvdA78BZ
qhHFpiXzViHMEPqAD2yE40AOt+hkeFwBZIEFNxmvtVNs3tF78C6KjCOGURt0qDxp
da8u2qKj4qYHbxI6w9SsCuJYF9OTZxPUFGLp3WqI/nQvAm9gQG/vxazRyzVtYQeb
Ao9/+7RL7zrk3NFigDeHE/w2J+EE4xYdQKc+sDusHbgQbKClPdDfWVKIv+LgBXzG
9wwRHI2y8gGwPk8AnolhtU0YS/zBEptstjFmiiBZ4+NBQNKIkqPSH51a2rMcjL8l
tjoa8zkm1MAz+pRqqb79qWGknjKHrBuTEGRbpGD/+vqsGacemXgtTwpkQHznGJf3
O/PGGWv9JsgHiHVk+QSFq7tzkMxtFpAzfEM2+HVwuQs/4iMj9GnEQN3d25OmfzeP
w1Wm0Za1CxJTkJf5hC8GUk3ks1Gf3NUZ2xnfgG6qOskbyFTije3GKM8WiHW02dCp
HEZH4uUK71vF6lOPKsLfWsT9d1Eyi2yqFPOUM/IDgvaNDhLRWnYxGvsHytFDW7O3
ayj98vWThiexkjj937FbUPbPcfdfkBHGPwmGXLZmcSNP7QMkKgLd3qTWBoImD2pB
Tvaenu39mKL/UuDpAc/1YvLptitDm5BYMNMyDi80b0/mWrdI9pyAGQ3BG5rf8g69
/IbhGiutB33S420eC4NnR4N5pVuohMAqjIoGBGeIYyt3Q1IoEuIdYj3VTbHsNvCN
R6KILldVkz9wgDPc2e8eCa3HgHCZJBJtVZxs9E2n5FTcGa695cWjFd09U7hHjMlL
B60iTHGBZqsG1cqQUFYNpAd3chVNJSewT8qIsPAOG2dB/DOZBnckZVkil6rBtUia
ISLKV2NJc/9JUTpPgVq5DSte2eCRgVNjSHeRKWdjipjhc/V1+9oR52BOjGQf/vvh
ISGULJOiq+m6TLzPPkwPSZts400fIGlPR9mSDcQqOt1+6oW0ZmfG6RleAowBWP5v
8FPDumaUev4mLc1Dz8eqTfoo1nJOxfPY+Jr0VIGw71jlBiklbBP47I7RxogS4Q7D
pCwjGDdFuuyDGM06wk/1EgJ6JfbNJlB7ueiBxoQdiMqiojCV2REhBXrEQ77rZ5ac
1TXrHW47+0jq5ODKTpE3+2RsFHkjQSLSULP0SSTaBxgz7o6s02D8888FW2YQawRu
DrkUYD9M78TsII1hw2pRh1IWmoS8+s6YQ4QD+h3MnTRnKQFitbm/7dwU9kZbbsYX
Ea3NYiCO1sxLYPjmav5X2HOwSOHCYBCiRtttvGi/Ls1z+0toVDXTFO9+Ln2VaUxp
euX9w7E++IlTBMz35sS7K59WxbstSamd7ttaSduePlAlVOR4y8TZQQmZ9GjwLPcJ
Bu/9EmX/2vpuAhXBO+7vzzdSTxyUgITW4Z6ZC9XnnH8cC5SIYyuELekG23cxqUjG
WUJ1+XAZ965s/Cla/LCc7/b1jEegUCuqfMspPfBxCEnxeSxGhsn2AvKI0ZM++/qh
UYfhIoaD0sB0G7avK2w22t3j/cU9oAJ/zTreWScWSw/z3gubUr3zM0aStiGVmmRU
fRJk6Y0Y4jX5n2X3MYlo0r3vvXRepCgtS9cSgPunL1Vx7yBC0oUsXxz5JchDk7Gx
z0gHIrWCQ1A7p/Foz7zL0cW1tt+8F6ttKwzwRWDFeYWk1/fV47F2qxtAc2lWq9wJ
i8LTG7QNflKxDiSdKHhdT72q0lFAx2+SxUjc25pWNN2AkhOnNSdkc4cDBOwBJwOo
sIfIBnQ7gAfkHu9drS4ktqylJjDvJlnpAq0+yXEihGlo9DtVysR/5NhnOeRS+iVN
3tgckCgvp50H9MqacQJ/+sLeu2HjXeG2BoWp83qDgZLBXR5HGv2OAho9iHRSTu20
95/4ktaRSZno7jGEvnz6pQ7vOhZDkGjRXf4rf49BLp+CUxGNBoct1dLDFxvZ28dI
ilPTo2ABilh0ooD66ggVT8qZAgloeNpClTNLLKxAMmutm9Cumco/0h6Tm8SQ0MT5
kc7ciuJODACXmWrXPDhXfAQ69UI0pnaTF10TJofCyjvanZZEUvWtZPJW1rJ6Ksns
KUVIeVwRc90SIgmFjl7a2kSrUuuFVEwL3OmHVMoyC1Sz4QZzyJdsi+ITbFicx2cz
DyFzwdtTzWxnt0ImJn1SzmtvPXmbZbtLpnFK6iEcXsuDVdYOcmd5ajGtOuH+2BC/
yalQhYDA6XWJjYtKujcrwQELz5jxVXaAi5UEKZI+0iVvGbfeX4dGciMu/ASge2er
Ps8OOvAqYJnwmuX09IYPtDw1q86sixJYq9WBeMDdyV79Ia1XGg7w/J2PpcmPXgTB
dtkVusyI6Qs/BvGmEL9tFphdX/LtUweZ+WsGryAqsAG6Hgpl+PK8KXNHqIw9L/Os
XG/Afq31XrrsBwNg0og4dmGrIr3bk03sBKlTbkzvx5x5flndKzb7JlwNabmexJf8
o98PMhyFYQrVZ4Kxhg6T2J3yE+DOF+iRPVbLLnrnvVKoLVNJfpQk4KFKzBPhDMXA
epfnCDOetVNy90sD24HxF6bUfAV4G8ZqSxdVLo1ZLDzwY1CGqg4/TO3CAhI8q7vD
3HnF1fFmBMsVVxsprOfd3uQJ54Y58Z3UUxxsltBsQGxv6DPxwyR4iX3bcdQqHbLf
TML+b5cIP6LX9avcUXPoJU1cgULBbzsFYr69Wcu8TLZTD2DfaugibqyCbZXyQpYs
W8OoJCgkSPLML9BfJFY1BBxDQlh933zT45KeCow+wS5/CvE+qgLX9jmoi9cgkOR4
v8jegyMatcuL2gMjLgM1X6eUoQFB29+x37ye5edQT95K7FgTX2J9ZF30QXt34/sG
4nc8XfhMJ61oJIKNKIn+GlnbBo6gucIIC1W3BIc9t2EZRoszmvpKA1+w50aDsZgo
M6sXuY91wZLKPHOxL7D8gA9Gsopmy+zOqTW4SU3+VF/W90wzGFWgbSF42e5uJooL
MCwxYTyFkPqDRNAAZJEC38orKEzqgOurd/TcatGpjK28ZMSlYwDNN8lXive/taVY
a9lTpBNZNU2auPduRTP0Td1Nhk50juI2J4PBqGXxcAzJHCMkmnhcOuRsca0WUX34
h+8IUPtIYwyXeWZGXZCYDvtiqBptAjBBuORrM+fe4nQij4xpnxlWMfDkwvirrl9H
8ZdlE2Oa97zs1MAOUA+ykuW1IGukzvke3tynQkbUVtXEwrlkT6Vkg+2oOrj/2oab
Glfmum/BR/diko0grLi3yqfkd2ENU2kKxot8xssWZZIvkDMcwJ+c1KE0OeRiuoci
BCXZdpGApcvzTFScQ7b3HLUqHOGG4o0vqxDdZunhh7QenbkbK6lzb6zcplk4FR+4
l/r+DQK0i1FYEyNmia86mnFDh6VNh4NJ7vgWCaos3elv6IrXUAF+xINUljEYrWG3
GZzqlFe25UGLFm4flel9RzmflrrA1/7LiZyAa8kbq7vKOWae/vdk29bhLu8skjv8
3DgJmy7m4/q3kPwpINyU8+WXEWure7QL5P2gikFj4Wa9Q984PyRVki40HSsJHOJF
Lf7NVgAoJ1v+vKPdLU/mQc0XG8uvVnubswQSWY18fOWmpTxYVt0eJqXRSrFiVrEU
gikYmxRj8TY/FpdcZEf4O1PiQCd2ddIGC5Pj7cbEhYdFaZQi/2O/4W4bH94wacp8
78q6mbnLKyWh2Vio2JEKWNrU3Kh6VOKrLzIGlnPubzQxjRVs4BDNbqpBTVj8ebYf
xxO+vRuwu7p1/LEdrGYvlOcYO4rSpurocU5uHeqXtwPm6lUUEfZ+Rcf5GMC176UG
6nRDSUehTBn0tDypkEDFwwWC5ViA2ohTojbuq0YgrMUvnEcEjuMm5DqlEkfKC2Nr
NdyXdIPpoUUAor/7d2kEZ1gZv148k23I4rYpkgvLY9ReDiDjhkoTlQeKjwG2LUTo
Nre5wtnkuCHT+QVSXeJ2W6VNL6O3y+SrRPOLQS+HOmbJRi13YUHfRJXiLyz+txtt
8Pe+A7nTBiQ6fwTNetfs8slRpqaeFv1P6pQBzkvkgtO1LIL8I1T3Bq0KP8QNJzAI
4+RsKBO3M5eNqkxLJaIRyUjhM39WaiCL4M26eXC3GkojRp6zUXM/ePxFo7BdHBDl
zW2bMPFIHX/e8+GYzQs428/Hx8QoE+qHKpfZn8NH4N0AozTZoiPYFReJ82Ks4RzH
QVV+D4CBe2Vk2ausofoNvntVy+lrLXDtsEFkM7EDytw8l2PZLTrGp9BW8Ms175rv
B7j/7kYcgFjTOcM7eVl8Lg360uvHv+tffjJfWSbIv5SP3ykLlzHutKCc9i04YKAF
7Shny+l4RC+bTL8zEGuW9VyjdHoYT1Ac5gkdoak2tKb5wXuwYf04geMYxIrvDEVY
cjM2XIUlAALhjqjDZFDHrKg2MWfsa8fZgVnWTbWrHIazi8+n1s1jRkB+OV8OC1Ge
kI3HVZpjs+jObx9mXSTmXRHry08VH+mXg8VcBJ7KYIMYh6Kf5E+yDApEqXVHMzqp
Qe3EQ79XbWXQZmoHq2CKKkL+AEkvqfCLNuQ2DZp/I/uhHic2gtgiCaDAruF37vHV
wQBdbHpc9sC2zogVbKGMmSajhy/ndGfbDR+Uo3B1CRLInH9TqFyD+kuDU4o7ZQ01
yl5WWGecprlM4cukXVXZzmBup1Cso1cxfKq5f3CTfxmBxQJmYLEPlfNv7s0nInDW
Hc+ZjYYpmiunMLxBqZZV2sBkjnRjEl7VAaFaSaLSyQVSwOYqXdtR2Y89vzTbbM+7
K/+2U7xPgW2tawAoVCQf9SHygIQXdun7S5I65wFpKZJI4IUGMOBZVNC/w6Z40eXW
5u+zgbl394TOb3CPonqgCWNpWbgyDL3WlyZVECSGu+vcOkHsgCQl2PTtuFJTXcWO
plTd+uzA7mF6WAqW8EPGrs9PN4cQOauwiEIWSYX9adBE8n+DmafOeX8lx6NVWx5C
K5VSIfFGLniQ15lqL4diyBAfE39e/JlckUu9TbBe5ysr9BwvxckD9RmgQL3gzrmW
aH9j1Llr9Pp7xNM2rbQd6O9p56pfDMeTQ1vkXTD0D+6+UtNJGRZS4rOXat9EcSIv
nCKfT/g2j+B3JeJGFcgOC2yqTzUGxUb5R3gtsVx+YWvNEeECVJWH1lXOQgP3vSwy
I0v6q/U/Cm6xCEA3+Rn/SwzuMMTnc53XbbRZMpPdYkwPSJ+g38F9ehX8vmt955bN
ICjBZj2Q1LZrtSgvY9khmo+rDJOArtKNw83GZNOHX6Vnbd1KFEmSXuzNSoDuysO0
FJXVGJcVuOzzUOe7OxdmqXKsUKZu3VfCejKmmmZ4ZkVdDIebu9hYLe6jy7oNHdCI
umoC97rQLZf5JGIO+pvLPybvORbpNh2LL//HxkTqZZ2x5O2Nv4Nrpx67/mJTxhpZ
LKvO44+g3q/XXjIKKZiBF9XtOUy3Txphza/vydnUQfadxYcXlJYz0vVDfc/IDLR4
RT5cdAqts1d+M7AJ03WffjTzweDtcGjSuTpF7wXOUugP7wo7cToGT3OVgsdxWbwG
veqMN6tHvrEekAI/8u/ssbOfIXEHXBcIRWNV3ZDccmNBsm/DxXbeplDiDBn1AXgu
xwtYPgXwnJ80gVmsJD1YczFKcP5AEzGfLfqh3qY4rQxcdmzdNYHrgHWMnztyRHdh
HrU2SwOGxYEK9d5A68M33Wx6Jnzi+57yjyQy5vVG8de6WjJdxIq5HTM8P4iQCfKr
6F7uXA8+Zu7s7RGaRm6deQOiOqQCtt0cloU6hM6vllonEIjAkIGUBhaTEYbMmSdo
ijqI2qzvuYGyY1LvvnCZWAIEaf0uDUtOxnxQUbE2B/UcOUsnLv0XQEyWfzOXDG6D
26iOezD4sz7tA5MD3E+L7pmHjnmxMsRwtDPzhkJajZe7pAiAgHNeQbHXzMTW9ndS
Me5mlXZgeulfGmsC0SLTBS6wZqwRvLtxDeCfxFBKZoz9PCqbKpLOe0lDocn86qEs
yefokJ1Q9WCIv54wTq/awfn7aXFCp3cWiXJzRi9SHldNpmYB8pBFggoF8UedWHFd
RJHSZj+/PmigheEMoRl5A7vr7PqJChpV08AmsPnZBYquERdJNZ4ngP+lxmA4xZ4M
fRALawFZzITPj+aTbTTxhdKAO39AC4kDP3DGSHQYOg6h3xJ9gnptNhdSHPxBSOJI
U8NTHL5S3hd0XBjgoUpEepYHgqPmyaDJjvrnwTEUf+fiHctB48t6bzyc3rscyGQL
fIRZV6NdobqOe6kuJ9spu32UPPSphzQDzqfnF7m//8Dff16grmmby/TRgtOQoWaW
BJFp+hZcXVk9xlrfqk1f2GlL8xvMrdEqsO26L346Qqssu7G3creu0hPI5UdiJTgy
BcWEzEJcH3ySh7Gori235m8Y3WGaSQJ3Qr07CQ8r8NswknNClcEu4CbVgsvelba2
ImOkJEkjhFI6Y+d0MdanwCBV1V9j3IWIUzc5sKRcPmZzVOCRxpVpl0pLtbOQGnjb
lDwtzYN1ysRkFt6YEhrz7zFy5RgDphKU1hOTtxNRJMIdt+rBnW7l0oSCNdaDcMuI
GN8VdpGWmsi1LYgK7GEMjfPAPZCZp3KhT6z6hAObjVjQ1nJ6zEUhPR0BkAkXdmGr
Jz6QKXltWG7U+lmGdg/6vvMvAjOVRujJqe18PmxTVCmUyXCd+X55BAzble1tL5Gh
9nODAsvI0ovd6LqsiyVClXO0Ng/CoewlcDoFMV42d+hqspQ5LhioJCBUGpefQ/ZM
nt17CBxHH9bT5EwTdCLUi92nDulY88Mh/fWY+fYW13OYe6c5DqVpKhWHiXATOZhL
XplQoZMoe+Q0PhLQgT3i0LwUMNQ/ctAE8ecS4v4SZ7VU6dEXo0VU5Cb7JFg1aFSK
/lf7OWATyUZk3euuwKAsB0gVMpS9UPMMnmYwTg2CoOw+EystSHaqzvJCJTIPUbcN
f92F+ltJYBqrD78ObqWpOOG8EQH5tAnx8mqOP0x4bp/19VOTDtVJ6023LK63PeIq
xLCDLqGed++gFWjXAEETjHpj8nePoUOaoSKJzbI9NPlSLIqxTB+SJq7rdSK9YcBm
4zJCBUi2L421toZfHvJMVj8zW20myA40WA5LHMfrQY33EanbQgz4boNuC+C7ajw9
j7YqIiiPsh9MC/fPBCfWTIdTC+f14wMZ2tKYYG0HPaCgSBMPbJ7vOb/KK+db35uo
N1skvPoCi9Q3zH0yndkdPN23qCa6wYhRoifsDszw0r9BnAVJFomYsI700KCLKDZG
J8HOb6UijAhQY1iG46hLdbeAXrFdPefesvR+B9FpoCtCjv0Os0DknTk5KRlpafWI
dePWwDq3sNWLCo5jLpgrelleuZsaf9uZstfSDuKxSCMTQHVRL4Ii0P7FGQ/ENWMt
8e+O9FHrn7cNySqea8pVyXmM24edKwT8mIWFm6uN/072uYBVjcg4xayw3kYDNnDJ
AjiRJFkTC6YiIyAVVtnuu2Is3WNCgP6lJaTlpj/8PqlWO0Yfzpf+dCXcOsNuffna
55wm1xdqgb1824aUX3Y2tQVJOxsWTvJOVY8yihrUltOfPqaK37a+Eaq9qM9HnnSp
zu0KlfejKRCvEUTxY1pPZGiGwYc5Y4w11zuRE86N+tWsJ+OBb6bUNXHSl488bmHZ
mju8qVa5emJ+phUiUhyCV7fwgokPz9dOBSSZnlhU6InSCIbvNiKmsN3RGn3TMPDs
rfBd8HnnajjtsJN7KYpX5vJv0ftvZSEFWYJQuWdpHm2byz9fa4rjpc4BUD5lJ6Ei
NPPqFVpiAzb0DyEzorBLzE0kSEn94pGGYyk/nGgLlbuiJHcl+a03GHxfT1kK4HTW
iGH1hiTjbjSqQ3w1IzU4GOoBtGCcrUgXFU1y3kYOwbQtbtNX4w0qw3djcdGugDJw
gpCq2FJDOcvdPlALg1bGp2qOt6ioBlqMp1k/urJf6b5jof2hvF0Kqr0XkR0Ecpqq
ak872JUoiivuijHjnwi4JjB5YBn9UKtBLImkp7IMhR8mUndKujL6VNXfWI6bKNQa
HyGMFwefGmJkMIdpDhZlPBkkPuj6SfT5W1Jh+I58+7VtSAoUTkzM069s647/gBsH
0SoISh//kDpdfTjupRkAYlcjAk9XGmA4YttvQHY3VhWwvzR/bDyuItgd04pHjHg4
5aKJUKW4HxYzl99qcDAxXoKlUIvWlVqekGjF9yQcJe6VzHQBqUq6LQ+PlYzB3PLC
XiCEvwyKcp+mLbyjcbfMioExbGgZXAwaFMWHvmMEDr7Jv7pssRbG57IdC1mVrFrm
pdtogbnLgokACim6JgVNTQV8dwU4zhE8sFtHRd0qnSYQowaYUootvSe1NIAMbzOq
VpbveX8yTwxGip3A7hIqM59Udn7ysfwXj7ngmMwBXvIAfqJLZ77Jus3qvcr9hu4u
vi+Z0JujZkq2Xusy1AmkpiQhCe7/cx7O3DVmHafGV1edIkVwyoTvbO08vlEcUYDM
6+VXU6SC8vkXTsheKtf8yVwm/LhO2wtwKEp3yJFMeE9A7IS0TfpPEcVHqRwZN0q2
2QX2WPeTOFX3AKksViWxE8QvVjBS+siYNPlmcgsA0JFgUikxEd3P8VfkQZa2buTZ
iQ7En4jMf7jMXIBm7jA6CJNgHjkZ2jsvZ3YD9gnPzZM0xgtGHtem4aXOnoYW414g
mwqLJaZWcd4vF369hophFiuD9Ogs2QQmRyftnHAlTWq1u7KyDwyR3sBpvDCYFgrg
JJtPN+m+VucCP1bzi1LPm2dHvdxnzRSOEkGNiAtqbiZzN8i78eGaLePlCWzq8i2o
LQNSt70K471wOMD7cnSJ/c1YzPnoyhf/6/1I1QhCbKs7DYTCrV/BNBh3dzMOHNnM
eCOufYTBUar53biuc4wGH1uMVlZFSO7VT/HXmGVEpB08+JEezqVRfALOlUkU4Yj9
w7qW+oscHLKY+YFDXO2/iC1Is0AyfNtCLh0Rkfy0C8h6KzpOBICpPMUCIgn7w9hd
Ar3qIsLgW+m/TaX8pUXiWGNFd5nL53+U8sgRcWLyUSFh/4jDUbt8Ed1yfwILhIDu
ZYTXeFkqRLOvDvENW2YjQEeUgzOoiLgHS9ZYxI0RVr9gxp1sqHHpEeNI8Ppkpqu6
9DWLyz9uuGu2h6tv98OmRPInKzrxAxK+3s/WxQlAZJhvag6C2ZutuTBxwk/ioeh1
/zq2RcLg/R0HN7/x62RiidoR8wCHrefavckBLb64kDNViboRSo2VJc0a90dLD0gK
J6+6dIgs99bmFQjWobl7b6n9MVdae8TAOiAwMhJPFbadD2tAlSnAAiKKI6E928ZI
0aZ7offfAGQMx2g9nmmeKK6dLDzTWlNS7UIvSWVqjptgYA8M2KwS9WGvDJm3eKGM
xDwpxh2YUPAoHyrjpVe5fT5jj+bb+U25x4PnHo/J0EmAQyryWfT5T5vgs5X4K27E
ifIx4s9rRP3qZdHEt+x4XkXNXhFhK/UHQ7Z3GeiY/N4r1eOFh4ZP1KgYYFV4NLl/
CDRhm9V8L62AiqUXVYXxe2xZ7M3DiGnOweWh2Lf69nwgc0VNF91DxYqXbn4Wtz0E
prFwrnx/Ja9bH0MOSck1XhmtD3Z694vO8eiYAZec2BUBKsJPAgTJvtriowhk7Hgl
XYDkF/2i21xFU4F4D2v6fUs9i8mHOUx8Eobj0tv6v1f1hGiSfm7BBuMME9WBPky1
JovCBAgRlGVoKJ6AuDcZpZN06S1tFSdRMZ4fqZMF3heSPIk56a0SF765n0wVwclq
UYl3N0Smr1EjmMNfRb215IcQgDZpt4p2sOJ30JWKisq9klyLpTdmeIeA2dNfLbpX
BsVCVejcICmCmE7WKiMa6FwmjAHjkaEtk9+SRierLFRSJOOdtYq58XCFJjUt/Ggm
4nuSsQFyJstl1FEmgMA1mG1Bn/WmVSxx9n1u87zOK0yJibeZXacK6Eol/IOo499x
bBMaULaiPixtaXygdxwLm/c1hJ9/d76/LvnQR/+iUvhFaNJUfT/o91bDJQBQBG54
cvtS8V91DH6lNG/pGLMgU0ypGimZWDkdxPusreo2F6FQNgv6kkudRlQ7xuq7V0pz
0c1bn/URNM2nTrO2Y+DciAX1cWU4PSZNXeQTteQqiOGDBZuRCIOR1B8Hd3Addjn6
tNCvADKk8an8K3jtbwj2FytX2Pf3c3cVAMF1BBvVL/nlQfA/WEePTxlNWz1F4z1v
PhzQCcraGhX+pFmT90QmgFJgH2nupWLCOJJiiyjjetl51iKHFC1lHlcdkAtU3Iao
ne965NytR4TjM2zTiDNb4yx7etR/TvP62exaS7plo5uGam5IkFkH6B1+WU/ZaMo8
ZFn4jutqfhoxKVILyp7JieF6G7lasHWTTsAwQqAZ3OTyBg2dAEEY5vgunKYx0TqZ
s1kUHbOHpj5HJGUK0mXHqUuw7zNdlpKVy7JC50e3NjHs/0eu9HzdQZM9l+2PU0JL
NR3lSOC/qVKXrKPNpq/eEwykndZpgiHHq2SEVpFpmlqCwfAq5rptw3REeSn8V9ei
f8rFxzSaQcwpse53ssIvuLYDzcCBY1Da3bBC2zxZjBAttOmJtmNtmTxVw+Sa9eks
x3deQPFWIzD46USujADoUFpKF7+r0aqzeaj3GJs2k9lYCQWCLM7fhbd1iyocgwst
irth7z+ZdxNHHdFOO5oWF4GOUBfBQT3FNkpEjBdSnTIMQyqFixLxazfPUKmKG2Eg
/oZrVGkjaXM+C9sVtFdQ7hoD0s4UhP8Guea7sgjv/mypEJ4OT53vc7WRQLfVHTNU
UyrUgGrlT79d0RcIzw5nMZt0adJLWJx0J5Yso/k4xqSzE7o6lW1IQiFxnj0Ahsbn
qUkRzzz04+ujcdPFFRh/JKFMyWfv2ouMpQIMqLowWAkXgBjudhE70VbzKQLOy7DL
Ius/o16a51Zm4wl7MJUuBhEa/ctY2cCCcbCUe7yBNrla/dCL9us92qFSCLy+Wa5l
1cGEPJzikm843yKo/Cvk6gwUP80RbW69fRItCmmrwV7UCgc+PCKNirkfhnZav7hj
agNO9PVzx20luc4eVisGm9CSMstiG9ebljZ3VIJsAUoJ1VfgmiitXcgnOZvXDeuK
lhi1RgKR5U2XNkQchRhDMLCX3Gt2NbFfWzelE1l8oD8/E4OqbuJNvncGywzCHok8
eqL5bpK06ZKQAJZjJL6UjEtxoOHH5yfQMQGzq9pDcbs2gmqzkbXFNHM1sfkhL6zd
w51JuZVMNT+p5+/+XwEDWcGfUcDK1TBLb6lHsVwIOTswKlvo3q+mAPr6bUiAR+16
SCC7Q7rCrwcgPxY12RxjTxUnbzC55luNUmgzSPvv5n0Jn4wwcc22RFlHr2mCBpiN
hX5OJWiyJVabqj5KaKYibk+SHB5h7m59cU5iv8wTNIq3Dp1tMVaBlL/hsMQurGh3
NDlf8VWtztNwhqlzSPDySiCjZ9+69y/xWVPRZLZ9hYhE9cYvbh2VY3jzF9ryUCzf
RddTsCw6SXyU9vx/adY6YZVO8xFmvTPwxrUJn8HomIDfIztsfjd89owPM6NiAIA9
E2efS1MSft0Pv0ZuRJdW4mS4igXoX0XNgvV+qQJmkFTsC+Iiox3xmvBII1I1HjEC
6Eqaejio4KhIM1n+R6gchk6rwV3jwFAXWYV1PntOYNqnhIMOWsjxPYYNFX4gCwoI
UBDyAw7+Nrw6hKDN2/+59Uu0O4QVJ55ZsXNwOcwLtUfEZSMh8SVrojYUeOceezG+
5Elu5q0Y/9fntkz29aOTby8ngNcYQ7P9MlDqI3jTwrqSVZ7YYbtOYwOO9wDyTmNR
FapBkxhnIkw/35adDi6ILHf8OUaIooIKZn55RdPHrpJrGag0G6xnFaVwkoc/GKIz
IPT2g8rsudOswmyIlRmnRMng2xDS+guI0dcfMf600258PNNWrSX4bZ9sJ/jgdId1
+fuNy0CN7AnzkBhJo5sLDS/P5gyTv47mIsJc9y/CQWiIuA9D+i6o0dO5qhtk03gS
8sRKGkv+nZ+OMNr6LA4LaMywArcxZstZn2+25eVpplXuGbm+ixyS+M55SUhcTlQ+
QJ5qmQ5GTPYBHW7CgIjHjOPWCjSiJqmLJHi6DM4Yd8fzWhkmhUR4SR/Gj7dfEmuM
mzFJTL/WmwEkETta8CmHIVfAfMojQV3G4px3MwO7lyltN+FG38KvpICFpj9wSEgm
wLh3bPRHcGTjTgEWJhPUXi1hIsow7n+erWv7/msDbUZW6JMoIWmPxu29XPb+B7i9
HnFSZjvd3M8Sx+5Jew2CtSG8g782jCmNFu3dcNK9Hljnoy9lVN9ZPPt4LYUhCAVg
rBIvuNZLCToYrltYZeXGP0PwsWNZ2tEbonsaOB7FpAUtd6ofarCWN+Vub6buZBsG
n2coeQitYllK+Dg+U3EZBAYSTD9nwUXbO+nqEj+5Alg8uAbeWXtZ1I9wh/jwahDf
s5Oi9Nkh2OzIFiew6nJbg5H6UqjX+ChVi013ykkUicXaU54xKUPWUWxE9D4sRC0G
+RvoMGVove+dGWLxR8g2szoCVmKvgmAydueLyVQFdpyyETbxzm7Q2FQwXHT19s5h
754KPRiHd6nd0QUncuIrQmPVIdbjS4TMZLuQfQNZcNRzNQc3zB6Ti4UopC6xxPvo
KU9AEdotzP7rVMXLixMA86DuMS3AnUv3hGpfv9+9+prOnNDsagsImTHycoG3AdcD
kNCxuC/NXvOcoDAMb6Vtv5Wgg2li2AWD/soI9lvnxyPnYRi8kEiFuH+llBsKo0FS
r8rg7cRaN/4g+iF/XvGBk/BzLKqgHpgvEEN3CwG+OCsNjLvQF28nZ7dyPGPkOC9G
kdU78ccuNrDlB6v10mjqPD8EGnJNRQmIurUivxtU18Dx0T8ihuwfhefrFXPKm70r
jaRQ9t7GMlw9QvCIiFuiQYgXK6PvvvLuRKJftPNvcicrtVQwWaXkq6X6lKvRCfnw
yryoSMBpi+Cg7D522Fk/yIQyio8e0fij+c+Yr9E2jSK0n0g9w+ta7R+d60DxcD8K
VREZmJZMtH7oiHABHxDXGb2VzaVhigiBs+uUT6YzKqwkI1F4luNcbORG33LphniG
go50Xdht7XCMjKHeC8QBTz3yLt0nQ/y/C2f9/oSuf+qKE+p4ttQW/j55fVm48+3b
TGPwB8+Kz0mn6uYnsZHldGRDGSkclb8d1T+OzwPyFd10c25exgDAIjCa/ARvA3Fg
SO9dLidSb8G8pokaf/0dLhPL7CU+NdO5AhDsYZ5+VV4y1xyjkj2rV7hNS9L/iirE
8JfQl5TKNjWsYw9bMFBbHDF/R5nMlsIgD/O4STFfnBgyL/uUaQ9XBdxfwFkqBPCW
R5Yd3U+wXGJhKu65kMqLtkVIUTgwQJk7+duVKomYLoDj1xF5IlgLzI8XCsUEJB/O
q5XhMatSaVDKlbw4dVn02BTTNARRKF4VER+NV2PeOrYrOMxITCZfS4xUkrCNJ3IQ
I7Hmegj82Xqr2grO3ML1kOIsL8dbwHtRc3ETG3LP9MuWHLG9IJgzXRi1fQ7iV/Ry
X9RyC05YEmv83gagfF6owX/OAzBHhkuBxc2DK8Rh05be3oyUtun0iIYfA8rgoY0w
lbQM5chw+QeZ7JlHami4VG3KPlnDW63+JmHdGLM7i6dYOR9FmxoWBIuuHf0lr7wh
QxpjT37uQuGD7Qgr9ZLkz0xtfqQzkkEtlJn12bYM/YwSGs5eI4yi3y8Vp3CGd4UA
+4AKDimnXGzc0aEtbuBqeS/rxOHedFXWRzeW2VpFc3LdVtkOOFBG2hkQSX2FHXSj
on2/PVOnPyypkbJA+KeHA4F9lkiNmpsozrDNtCFxDId01Rb3ox/EswmtiZwgozZG
+jf0ImWm4VXo0DdoZGwADMfkC81zloPSm1X54+FmmMaPXQB1LNC5zHKe6gd7GJJE
7lYvWQ/a9zLFeVuoAIXqJRWp5FR2GnRMmF1O9DnuZJw1yueho6kfRj3F7eOfHVj/
e1TLTx8//dbG/5xnRqeqE+FY7YjxHbZvlfxzrEkzh9mXXnPSOX9cd959EI4RLSx4
6CNv484KTOcmFMH+o71nGJ8YNpMERu/DUut0iJ4+OcE7Axb0e/W8W3o1WShqcb5p
Y12isgvSGEyktQb5YSGANG6IgWwnek6B0fS3wj0CdNCFGdn/ZTTqu5ynOV41VYXE
VgRhKe4DjrbNKOHXge4bSTeZJ4GrSn+mdCGN8JeoDq7GyIQZB7I1L8J05NBA5MCO
8X7DAo7mUr34VK+KfpHqfmiPO6PKCwWTThV4q4jQ5W1RzjOUMbgkYmIoddZbMb4n
YmWBk0N8FHvWiXypEBVBlZlR6IHW19L58M31Fsb5R7x9zK8ZcLheNKdE86yBPct+
vDO9fGVZNM03yN9JNq1ktaaGMD4Pr0ICVVnuNXypUzwfUpGQwERSM7PIemvhRLEX
2jrWU79NAv8fE/vIx845CBu1IJcRj+ghCF4aEzCpX5ns29EYH91Qrcpm3ySf+wj/
pxxUOIYmG64vJ3PoZTrWQXacnlloq6izMvDzCyRQRFsmrBdTMaDu1PUOqgljCqOM
vZTQzE17P111F1dcOOiPfrWcqxOphFOeczaVUsLNDFK/hJk+8DvXI4b6G73utEru
fTD2SFTZgejpKRUaEnHcCkpBxt7UuLr/AaZ2tvEyV1L2MM4XIwe/+uhePoEIIBkm
uAptILAnb39FUMJJDjQoJ8yxrDQcIx6/GfgEiaVN+N7usEB9yEVnYs+QfG1ObJ16
QjojVWKD3uiFrW6nBUTq1tT0XDC7ofhcv+YFSxmHuwuLSj4SwFkqyRC24mD/ovuO
DXEUupeZaUSBNssw+9i84kHtJ/+OBJejqIYWNNxAr2nhI8ny49GbLr5aXcLYy9Qn
E01idT0caZwwY+9Tb9V5yruhWcP7WYdZeRHUca6q/uBO09GevdzFQbKHzMQSi70/
0s/3Ji0KBS+CNwS598vf4URquwnB9V1wmIuDVa5Mp8Q8ThGSUG5Z7ms5iFQSSykT
HsE9l9sxn+XTQCR9d4ROT/PfEFZFppAFj8HP02aIFHSeJalS9ZK2oT42SbUtiWfN
y+3ZeJcAeIEhk1nYr4iZQoZ/m/D78u+AGmxrfQcqba/H6Nyr7YcZhlpNhUqPF2Ai
OFl1Z0PL4uTGxPuRYf6Qq6O6ESv5TTiSfbJtBLQTjfW8UT4A3SmVBWIp8jX3BzvB
cBBgN6EPgp3D/JZ1O9h3t6K/JoViRAlZCWOo+s6E7W49ww27vidVO28DvawHw0Gm
JPne6AjET2FIBz2AgjqGEWa6iNK5W2mCEMUjR/wHA9XsmoMIbdMwQ1E7Kfk1FOoN
db0KLd+yYRtYx8O73maUOmYotuSXtVkjeaMI0t+VilKPoXfubIaBsrBWILyaaTjF
mnwe3KnqjcjddpbqJLZWtwpOVA3aMeVqJpe9JcF0ap2ZphlGUzDU5GZ5/TMEXcNf
KWAfpZ5z13eaKNccVCLWZ9QOkHq741+FcAGrCjXgfU1tUrSxJBzCbIS6WjiLKwxd
XTtcWTjuJlgD9YQLyf4NkJMHLnBjLrRs4iuOuqfHb1Bq0Rk540upxWKgOhKZnFxr
kTs0NkMJLczq1fjxC5UxJP4QhzOMH/uA1AMxz5oHCRd1BzLZXJwdMrktUkmwORrB
LmXxryvGRGjO1sO+chGjX1M2JxBNthioYUODVkU4mmw6yz7va9OVdi7L05yW7ZTn
q/vGUPtdbYJUEvK2TqbtPSmW/SghEGl9FSwQLtjUTJcdNJxdLm6VmsXwevK6D6VI
oOKHr91wrt8Kbu4I9qhoPZTedpMFOCIwKtCAWPk8rGdoSQrl1OYipjJlY5e4wKOx
ghPUrWaqZKK9YxJB4kS9iOjopmbUOIty68VFayDHYdQZkQ3fufKa7/LjrJQJEwce
vrNEWKx5drFsd87AU7IMuDLzmEhLxAqnU4/s7moSExESZ05a0Uv7fICLdzpY0lZy
pYtsN62qlG0GpQx2klEV9apLDN/9zTOdquHLFbO8u4HYEiqu98NwJTdPzgWGZ4Fw
EQ21AOJaLrFLTHDcplE1cFMG54vpRtp/apGxkuOveMxL0WmyctcOZs6GwBxl7S3k
YtSOK/GlpsJpQsMwBvQJlXNEBOKuy7OSiHXrGjH+pvbmQu8iYA2GWgV5y+3wAOeI
4Nl17QVY924ibVNIC7yyr5gw79/+zVbG+VW8j1BZHFIhBG7WmhYxfXJpfUhgrZtF
A41eOXwcCn8buFC6A+HVSNwbbHjrIYF5UD+4wrny36IJhtVoDlhnifQUx8Pmrtm4
63G4is4jiHVDp/doupuqKhLWBZiw5GuHOmjVFM7c/0i2xH2B8WbwxkZwY12+COzM
nMniMLsYxcuP3o2z0KyKnd5uPLeEnJGqGWY6EhktP6MI8I16K7NztH152kn9GnIL
NK14OYOGg0QOOKMNj1t1GeWk0uHPGrYNzhMpDOjqFOaDJHQJfZ43FJ0xR6wcZOkV
//ocn6tLchcXkRszVIbexIWcVF2yBNpyIpNSxb1arfza1dJOL6bcH0sEkxe0Hs9U
1r5DJMENJARMStPjkxGY+Hgdsc1ONHQM4kOLmWrhw1ib+KjwM2AWVQk+eC+c/zCp
Bjzqed/UaoTUdWRwsiYqRSTOXYopHF5p7vwQ0mGMQsugiMlQOW6TJn7aDNchKA3O
TXLuSDzrxiob9f2b8Ohv4f38wfJNuOQtXkiDlm3bYqcmjzgxKkwuBjhzIZhkq/oX
TszDzr99on+0G4HZOj1WNGEZb2NZvVVe1TNYtvWZehlpeTCZPmDBsJ3ei5Blla3s
iyc7pMaDHEbRKNkcVfl/OVHV68UiAxg7axHyTMPGJFIa+P6kk9Ndcr9bdQ2uT3u/
MxkI7t8Frkxl3/OhqpH97LAVShExJ8jqNgcwc1DX8vQ6TJKN96xJVK0aNbrWtMm1
1JN+Oxs44TFOiPNL2uk7JWRB6kExGnTKym1KLlJejS540ranvfcx+NLIpSNAU4U3
sY70NNgF5eqxqC0ld6/dmc6jQxyoCucivYkbRGSjJbzrtaEWaWDpLJ9K3Ww3k2OK
+aiuUENm/UnP3iQHzvNOWxpCBzYHNGHqgCEczgbcUxbPixC/0J6JFiDZx8FPIOZx
hcFAFCBZlSalyE4SQZSaufatU90yFt/ajtjiNRufocjJeMPKvNTO6WxAaPqP7MSC
4/iRB0Cs7hwborA5VnYUTh4FwHr18vTsgHP8EUI1hGP1mVE/kpceSzM4/Nf8GFxs
/IcPFVqDWcBiVA1ip80ppiKbogGzgWYwvroV2b8vogoDsSyz/ZrV/I4YrHwC9dF6
HElri4+F0HS4RNlNz9PblWN6RryiJCWA7IFzSOKbEAdvoMcHXOjNObzi2W46t4tD
hY3d/sKajbxlL4ahwv3PUvA30VrZxoPOtDXbme8W7SVHn9f12UlBGRIhgGwC+Liu
jsU5TaWdsss88QegMpq+sOnM98DiT5FJebWFFTwnMNrWNqAAGl+zF8ozffbcT7EE
ikS3bd1P90affoAZt+yXMSJCoICEWslRf9LRCITOCZZxIMN8cjFpPpxMvCRiCd7b
BZUw32uGT0KjT6PjNR/tMQkNJjy9IdhdiVY+3cpraSf1plyCWprf0JWKnVplSOUg
vLIa5tAsyHnUHHBK05IJ6zlrmJXXkgYPyRI1X9mJdgJLGAJI/KqNlqcsijMZodyx
8FxdQScbbkc8VQaJx104q1A6CPfhzGTyGu1STh2MGLcbCITRtSQ03x3bqtKN3pu4
gXZQD27P3ufoiwJrre2diyIhOPvXGvl2UYfFuF5zEXyGnvIP+LZtNSkEbNopriAz
+PXhyQFL5hDR/eXKAb9L1i3+1rB/5kxlwaTOk9XwV5VqSFos3scdMvzhBQxbsnef
M1sjMyM5J8UxEZQuVfp9IvBSK3KjvqRle6euJtRmpl/L8/Zd1a5cEbZCIXjLixim
ozlswO1NFL8IyGWjkrFl9DBbTimyLNrw+6i6G2ismkUKj4C8E2bERabdiPR1uTPh
LptfhFUi9ME8vcGvaWSxsqULUm9vT/H/Np51KoHNVzSlubBNuPlOh+EdZL6NWloV
84joBJ3Ez88wAQOz2rB0k8ZOAA7NWeIMhHbfEA7R4AqlAfGQZQZfxnjgZm71iwl1
KcWCYzsGgGK0itBtS/FuF35PcMd6u6K+vxR91SEOV2J7sJiMv2LkRzsJuA764HKO
M7PJfRU9tWRzxOOVjHbmPD0wiX/1AbcfOugrKiA6rGIi6//Vw7i6TlpV2gyYroNq
CCT82eSkJDe6Mc7OCeWyIWZ4aEP0Hs2rqXNYGHgtyNQqVYGX3xP5SZ2sUJkrydkv
80nLb1fAwkv3hHfZnbz+6bq77Vst8CWvTx9yYbV4IP2OmDqZT1JS/Hk20I54wfb7
AF2LeU86Etl3oztKAhO0kaPSYSeAFGKdfMv4xbyjiDBmbczasn+C8mA7JxLVVD/1
rl5fOjdDa0sM4b3DMGQvP/qP3aTLBAtrR2N1nlvhfXsF4E9g/GvTCfN4kNToVFUY
3CmusRrTfmFwLeHTozMvLS7FRk0ov28UMZf1CKAnR3EuRtXXFj6zWsgqUn62CN9J
XkGAa2qeN7vFRN+VojknCW+50KgqICTQPuM1ZlFOviZbwBl7kmunREqta9Yt3g++
hADupS2kH+IHYQtId+sBnDF62gBIva4z2xQ52yLyYSiGnT2VkAKwwUN5hHnvu/HF
GAfjPjYlmwNIjb6ttvDAhNQvTWgz7lVACyuGoNiSch2jsxHALGJFo1FdnHgtRaM7
fsJi+oYE/o3Ml62K+G5zuuNGi1gvV8QJuzNXSXyb9Yqr7Kz/U9wzsNLxv3rmDr98
aqylJF+ji/HDN+zAo9mswd8rM4ylJtaiXHHp6BrVr95o88OfHtD4H3jBzg5hwauJ
wAWFAufaGyHa0WBhR6mmX8xHtHU3AndNc5cpj9C5LC+8NJGwLHi829RVBJhUdtRq
X/MncVAQ5F76gC8G6q5XjBGCQNIi7nBkynm8Y/K1tdhkKABvPSiaCSifMkNC2LfS
cjqKgeIbU7m72I8nsR4054bSMg8root4Hxnhj6kLgBLSqgsPZYoYf7n4KWsm0co6
GQh2TeFgf1X0mK+gvlH6Ecf5JqpWiQZkQqdp6exJ1oQMwXh4itUODWNKSIbMM1LO
D5hvTvVpX3CPBRVV9uRUMY4Abw+lBqLGpOTAvEase4DBsWqOmdKufpihH5/AGDuL
P22ZPqI8ZdFDVnjqVkcQKpUAjWQ1VbrVK/Tlm921ivMv7yX6iCkY2bjKI03KeGih
YIXr2Ui4gCkVHTAyUzhRmhksPUMQuoFPfXt7pgc/YTW9zon78+RmkDY4cbKgI7eb
f8YjaHJadZL5PFre264Rold6S0Q8UILWh3U+ErVUtW3mvRulj9cxiAkyXbvO2qCz
rlQacDPAckSj2lELygbhn93yrjrLWQXXfbji4zPRcnWAdQoKUklLdEo78lW95MWy
XRSfBgCeIVACDMmAqI2B+/8PwwpIWMZfyGQCCxxPeTm/pplZpzKtkbPsjkU480cP
vgGzc5nV2TcavZAc6m04F2DYFIXeBfZs0eYfsGrFnKEqJSzDq3vQGc29A157WhtP
N3Ujss0CVj7Zx3X3eLjGtb7GMsLcP3VwgDSC6AdTfIjzD9Ww7nXdRLJCRqXmVJZg
XSKG4Xkzby3dY+TJIj6EM3/Nm80ilhCB7jkET7CN/M3p0IbydPrcGxW0glw6qk2m
0vrbYXAE6EnV2xq2IinVxOY/o95NNVoXogFFl9eJPwINldJOhdCPtyZCy7eQpF2j
ro9hamdNyvMvNtfTN+qS39FDGWSi+hnZ3aIDTX/nfE2WlwhyKLqzL77ZcH74AdFu
GWjwG2geC+IgteEIxbBKYZVO04MApT0JFrpUeCN1Z51tvL6WVkObWJ+jc1wlN94v
l1fds7X+9Df4E5F+Cdw6W1Mj8k3SZFq/8ZnFWB3/T/DOG6AAtdr4O8spfBhuK8ar
brHJesxD7xg+14Q5pw5nyq7qinsF4TZJNIyqdJLb1PhikzXGCCKJ786eZ1PnFv8u
+WuOGxcZXr+1PDOm8B/6OewG8RWF1MU9nmoALErrk62RcqaqBvlUefBd9IM3uH20
cIrDEZRTtlK85buJH252ZFWtov0L7+dM3u33eM0mckitWwxsH3uUMDOOlPMDW7L6
QgTMUMezagIKKEb290W7fCd1PqL1N6+iIWTjorvBjtYKmsDEVUcQT8GtMHkMuTYy
0MJn1tMH6bE+IsxKXhn34aSjxpM4av0tho1Us1x0v9/j+X3zPBdDhseyljdD/GlN
rziNF1N2AWRQYjPVK8ZqdE65QD+igW2EBuVi5SSl/vPG6sOS7348Jm2mRs/BCBZX
nOdrHDWPEYw0DBPcYNDyz0MBX9t8X5cfMbk+5iZAu7+jBfqpPh11O1/s7tnufod5
o8D38NgBVC87dAMUnR+2Z7o2gThnjvUWUHFynutgDm3vZ71DWourc688+bdTxSe+
t64W7QLM5zj9f+5wq3X2ml5yllPiE9tLbr5rGymhgyNzkvDDM76hzDVOCkZL+I2N
ydi8RC8i2/ZMftDb819AUVoVECgO8q2dRMCOouBPZ285MP40TrT7xLTRHB2a09Ih
OS4UYoymFkh+JbmR1iRuj4aYg8NMkJSlq3NjoaJSXW08zlUzyp/1L/o/+vdiLOfD
wNdiTmodMuOGoGoOv9/aGvhMcTBKm91NFAil891SDl4ooW5Qusxr6N9fjFR2JNPb
S0UpF4KPVffPl9sy30ijb/GILrAl/4YQ3px6VaPKifS644xFxR7aHMVzYIO6YvE1
A3SD6C9i2uiEg+G859boQcCkgB8knvPNXaTq1ewNIYRhh+jk9RLaKt3Zs7TlBCre
/puTzFmIhpQghD5/HWOfj4wNu6j0516WDBHWwnCJXmjNG9mpvmhauZaMJDzH4ryF
yq3wu5+dmrep6fwW9v+gG7KAht3ESVP5pewE8SASPFrNORyDyYDEHgcg9rwnZhiS
1FPEVMlqbtP0wesouQi29PlAJ0msyKNYPrNe64QoHo4pzvjIF1XpCBkxOAt/Rl8w
4crmokJ3dLrVGLEcGCmvBEJEQPTUhpwXW5F1iK0hqNDkE2Rtrlx1DpNXH9KPmZck
6lOnsRcD2ZW9OtOJs6SPPcKBMwCFesRg50SKT+Nl6QlnnPDip0/+g6NWqEgE/HzX
vx1n/tNlr+cKpPFHdoBZ27kaSYQmvzUZSxBvu1jve3OQSWBMDqSHd7w3xFsgPmth
+lpQP8W4oz7+IAUKqQMXazHRnbTx6RSrXzimYUvayW4bxiN0f75SC7Jb8H3PNcNH
EfQ10xAr8ZsF59VTAkr9ykmc7EvYLprPe+WpPvgFmcVAAn97IDBu1NyH/DBraK+5
Yp1Dos05KE6woz3lkoRHZ7DKAHKmxgFkq14n/X6g41QiD1neSmDT+RBfosrWjUc2
05SVrtFezAVEKz5x4d10IE1DMzYTACTjHh+V+94GfiJKSfRWfjDfbcqARqDDPF4Y
XWWrbIIK4sO5wU5czEcbSVBMHRgYCc6tAfeeEg5XQ7WEl3klo/TCAT956Ilpe/5H
yViPRtQDgI1/W7Fi1p4RLdQUmlGyGAHe9jojMrX0ElUP+cAdG1sEDg5B5lBhCJSd
zEyj2MdozGui2L/FTnwlX+DUi+TF3KVxO5G5rABXbX0ScB5EtiqNsUdKUjDmvsZ6
kOWaIdQDN93sAMPJ1z5jZ6Wr0Gmx3dBxtZgIcibgL12t6UztAYzGQiokBLhwB0OA
tq3lrvrenWBFlEfhjzXfioQWz7mhPwAtgd0fvRuWfK1pidxWQH3a6ucCMZ0Du3J+
EZX2dDRxYQXHhY4ckB+gOXD7L7EaAm98/R8ZUBQSi1X0QotySZcvT6bSN/Xpvgna
kYIk2mSD2UAbPv0O54qe9tqK1x4Twt4Ged7sOe1isoRZGsRcj1EoTuMwDupzVarz
r42meooTaR95U7QoDPiiCF3eK5pTrjIzjivGDiJUjoHsZH3GI+pd4emnwLT/Bznt
OukkrFM1yvKujCmYGNuLaDhSagi5R2WrrcKec6zcuTtbeDnTgRy1eCcMR7ioL260
JYUe5W9zJm0GLBnst1t0Nm+Idve/AJovS+46bGD3ZPXzHQmPSOTVDFOYazJXtNDY
REg0UC+Ah5zm6kosa+8TPY3D3Oyl3Uvf2H2z/x3HmKnuS+oFIPXXQPY/ArEc6tWt
/CPCXzuvgqfydVzLarjYOZWiMW7MeZZthCmrHs+6aDF208m4LfUnfCPBTfo162/Y
TFNa60jvUfaYH8BbqaIwH8A9ZX9N7jSP97msTrgPoMweVnXSBMcn815GaN8yxzgk
6DErUrt4nLxE9tEqSDeOJOG9kZwnHVIpYV8wHLbFIFkVT3EjCHc+fkbHqO/PgPBg
SP0ZqC+Q8/zRGwbNtK+BUeilcbukykX05Zxdezg2yS2iI5ikqVKuH85pABcrYr3N
lNN61xBuQ6+xI+XfvyIb/LIdZzbSDHni2zx7ePcQQx3Z8Qr4z7QjDsv3dtsGLJTf
OA8Yzt/Py5/NN6GViySepKk6XzVeth/MBRKXssKP1vGQbuS26PQCY1nti5f6rGOE
3L3ufcGOg6rE/4Kpjd/QpLRVipnTXCnwWdXJC+IAQoAtKFBttFNLyvRzF+bsU6TS
BpX0r/3rUE7yhHdSGyeIsyqUho3q/EnoA6MKjD9RoczER7IrQBvKMJjG7Ube2ASf
mZeXGj53uiZxTOkK1GgXF+MNwnW51ZYWRy8jBV5KBiyXdtu0h1EFxXeN7SpwKJDf
xNYGhMHJJbaXRXn21EpaQDteM2luDsMaW6zrLtzMSKgol1HZlQGsQia1Dh68XM30
pVIufubgx9ksNFeHBCic8huEzgxJ2oPveSZIq2fDpkq9oLpxvSOkSfMJb6POLcSh
AfmSuzFXhEBZV6G8YCdPkrtJ2oT9XAvIS/OaPLLRuFni6XabavsuG1gHzoWTYZT5
0xt4gLNfKdqR+ZWZX/x1S/sU0Nuv4tVSXqgfXZDfPS2eMT3KudK0Z/OoSo5rNxvZ
eBc4HNLXSlrftUXLUZ3q7K9lXDjUSO0WLRnoz+ueagP9ZiEj55wC+D20oC7CH6dC
U6KUeCFM/guf9cigrEdljvKHydJkgVSw2t0lkQ7n78Q9/BapJmXUf3UxQazFuDFv
Vru8L9H++PJdN3Flu9k1gza3xJJTWZ8PdzqH86wo2kl7u+noIlGdIER38hMNT9on
bZV0Vw9au3DWczReTHh7FuyQzPqN8EKajooVH8FdWzzMcSaFKs+Hn2jo5T2qyA0h
L/FNF4oXLw4/Pye/d3C8MVQZ9D84wP9lZzrnIzlKN30vFrvRLSjdiiVbRWqPiExw
DtMuzwWWMkE96PE2HYLyATz4P8W5k2fvTI1Nv/+OyiiW3VMNsdXuGf+LcDJaFmCA
lHx7pnxFV6WD6+1KA0QLVsu4+zfwixjjtao2KadLzIGd07g1ahj9X8fTkeiokd40
uAO3/t0zqbvmxUMpEmIHRy6jILtOGWdwsj9uXwH1No2+9iwozzDdPiKvsxBceNdk
F/9sjA1bwI/MC/W+SEqipCpkm6pxh9K1UUJM/czBfGuf2+iBOuUHnprtCQ6HxIxs
9Wyzq0gxsZBONsakpGYwjNGhaxVqE1DeUvHOCI7Qe+e+gPV2q3SLmLH9C1XkHTer
I/P+mvkKr1xPq25MG05VlgcOEOi/xyUaLqKNG+4VQP9b1naGMpCLQKUeuZ2OJpV4
4XnDNFCSDcAaDcjKLCemRGdu5gCs4zwnRVaCHVK0fOnRFlshxZzoi9PtDa0Lrv2c
OhHAMZMjLV0gwElu+nSe3v3k/xtlsYjaAWgZJjixrbQjX9VnEUb1gbIAaaIJ3x4V
xeorBV6NK5umtMavZ0hxITF/7TDEjrtwSSy31oLttyaQzcNhaH36ZsooZw8yn8yV
w+8eT5L2hTEuP2p+POg9otg6MfTrLCEHN9uaZtZJHXpbplrncDjheXMMj8bIq/6c
JHaVl7iynQoFJMkm4AU2M6ZD2mQTL6qH+5rLjHA1pK/L7BNGTO2CQuAMoJMZ+2d4
0gLWknItQUQgJJBnZZVqFerGvIgnBiUdC3eF8K89ak20h+lroklevCOdL4HBZxz+
3aJ7b/+fgWVCnKJQPzdTZ+Jj+sCiBl5PEVLweXVESmTbo9DhpEetBuO5MYabS1+e
obEt8PGdAArxdMpkuxKy2T2g9hhKLLEYezQPStH3BM49WYozHcIGh7dxsxqwQVef
MJ7GYjFWeOfV7WTvCZVP02sjY7U6W0p1hpkh71EuTmX9jMdZ6DJJQbYMlkNBW4tU
CldlHy3+3rETo9rHIl2iSJBzQVf6Q+T52eS78v3sUXYhA8R32/9eheIMSSmeerqY
dl/9FDmDq7xo5ebxrY67H7p0/l9YQV1l/pTiUEfL2xPMnVxzCtPbY0XQSzIjMOcl
nifQkB+XFuYt1id21XssImUdUUDIaZhIDD31YPehBXM6likrcRO6QCBLwbLiUWzr
iS60cueRqzzxCG7/EwveQjU+Pxqg00/R5IiiiQSPe76OQG9qZJz7053DVFkymZsY
xxhvoU/wtvLZaxLwFosNLMWiKMFe1+MAUY2hy2hCTbrCKQM99gGyaCIthvsxFiDl
oIg/eV1NvKXVojYZZgjhFPHYEHyxgVQ29fwt8obLdpYcpv2nhVDcflACY/jS47/B
DPoiqiLo0bQP/1VJTqli19wWU9kqrs9qJffNtQ/XDCT1+XGBtK86LktOlGkX6LdO
Zhgd8UvPB0hU1uaZYuKTP9N1egsRzHF4g5ayxulb0o7nJuhUCawKpawQZDwKcwCB
PwdfK+kbStNwSbnkhx+8epSX1h5eFIwj8f61W6UzzqR2GZuXRhoLX6xNCkztOlrO
kHtma+OBerw0E0nAEOOQqLBdHns4noMx2bPKkLuyNy1HhF4Psm19N9saVkqGmbcN
WuahxEsgconkuj+O61BHBrMCzlXuYgSRcd9D9/6Q5auE+VqQcHNR986P2l/KICai
FYefTqL22bmWK3ZC5VtgZfCNnj1AHUbCpnQg3puabL5zmQiDHu5W5sPlsQlGXaEs
PVK//YHR3rsSXK5QO7tgUH46hXWleaMzphGjd+XQg9uBZQ3mwQRyVarGChwLD33g
w0AMvTOtEleB6wNs7cdwib1Fb2zdBLxjplWMt3B4JjUy9gyrXTraMFq9eKjHcb3/
s3b9te+c+4ZLeRoyoOhl+M0qUchahA+OvL5tdLzKHK2CHTgWgxwbyYd2XVk5rF+6
pPoM1VWT7ROtxd4x4Hkf7ORsIRkWPwUYLbpfsFncDOYUMgpptG93VY1yDWcc1zLl
rsB86MTRslbPPzqaYy8L15BlB60C2q5GGxMRQi4SOQtIVf/W9FivmI7CnnDcx47J
YpnkP8NVjaxlPNXSoq9zqMkSgY+NRA7OKY6E01KCCRJr4dwaEerAjJ1sA+z1jM5W
d7zzLt7kqOGVxpDi99bWd3Xhs+fsyBQz1lX4hguFsdGHl3eWLmJnZ0lSqtQgApUv
tIttow2gbhSMMPT0GKOogWPGwdgNjfX6efhuR+ITb/+dhRUDxGe5lzHEtBYOEAwV
gxbaWA5zrhTlqqAYdxXIpoabR1BTKPSqHC/ACq3HFaQtD465mA7fdCcPBRC1Klw3
bBpxI4jn0xvK/79X2nhHl/YBXzFvcCmm1aLWCm9ZtF0r15UrDRcFW/m/GhcxIEKO
LgWeWBDgjDUzENpmGhSllE9LiLL0udjYtxxeKoFbL8pD9lDR6qOtysOMfAJLx2fI
tcGd3KK6+X2Mohki7QFBWQ0WaMPlzMpeAw2PDktPSk5zw0rrYxfybOPjuBcVSwF4
tAIFFp7AA4+Q0QB4px4eeSm7wfo9Bu1jZt97Hmaa5VD/Gv8m5/3sHDM+z7JArW6w
ukwLNoELHxQxsu5zXTQrcJLXIAmf9+1N+yklV0+XESMHdhV1jJR28C+r1epof+kM
o3gXz8tDiVqqW1zSToRawqkt6DmdOvMoey/hgLZLlpa4QI1hG3zvebr533SnsswR
2kzKJ3BLi+ex6iSdCyD6VWjz4MIojbM0IubRHS1K6MVQozBpoWy/9v/tFoLNxqOo
sKwTVj/bzCkQXvcmdu7flHBr+813qNkm3z2AuWJ2FHM5NKM4InwR1mhcx3ZPcQnZ
q+1jNHIRUGNwUe03DkvzSYBZKjluNBa3asumpo8Rd8MVprNH3k5nSv5hWSHhFMFi
6yGWM/wf1v12zyPoHGrdB43udabp/HHZkjEVcsG+lECUDSsk4kwYQ8d20MX8XgLT
lWF21byXVVsseWIzKuNDtlzZTLMPFpgQsCd5AGyEdNB1wZQpwxTqr9HjbdwyrXP9
VaAxwV4Gc9mbjh5DCGYUUwGdM63NHwhiN0ScXk26J7VWUvz+ngFfM61sd69lLHV/
dPWIE/VlCIa4tVh372c0MpaG+VBW/H1tds9pVceDYrAWGRZ6Id1c6m6a9usyNIM2
+9qV205+iyBjkOxb0944uImnN5A7F6LTP+q8vaJ9VP98nKuV8i9U8dD+HWkCZ48v
K0UXXep/9y08U+TKto4XgXCmzLPSYSEUN82VUZV/wh1RDPT7Klqcg/J7ZQAzuPpi
eQx4ZhZ7MjucS/+VEUg4euiy2H7dvNDhT1J0UcZ2pmwTKANs8coWJphITZOYPG+S
F9lGj++8ymuqdwe1IpXb9XT7CB77fIpyHr8zxMEIvIDZPIXGqKntAthmZqZNYRr4
GT3w1BBbDUok1f87BbWDm72VZaZL0+CIoQjjzp/2T5JKsk93UtvD5x39vo63Ovba
V3EeyJq3p+tI398eeniHU1s2SYby479bLNuPeg2ttjEQtukAn8lLn5PsZPMP550i
T0q59JtoHEDCyJd6wsBqzLgeNRVhS1+9yKn5Dp21oRo3kZfnz9PyLw9oJAwRrd2H
GptMmBW7EbhnNo/uxhO5jx9S/zRQFHa8F43QWIbGZRAxjkvck8fX+J7R4vkvSEXC
KpcDp/Cpo+06BU5xDeOaFq6+EQDZ5F0xgvraf16/eV56PPjumCAtrg7gV20Fy1vt
DN5FWjjhKmwd2XtNpwd85PoahdANndNUOAKet7FT2fWzSX6pkJRoeHOMl1KGsUGS
7SCGJul+s1O6kc2xOx4jMzVsu4uH/QLMayr5poauSokWzbt/S8ShImJJ7/KoCB7f
vnDpy5P1nEqBod+BvdJnednR6rCTGiS8toe6DUjGUtDNXAAoN1q707iqsAuzVDhM
7jveFoX6yf1ll3ZxCEysgvm0+Jm2/17lwzxZs/XeBvjzGmIlBoC8CFxd2YZ7OKsx
vRg0fZ6T2+3AiLzbsdhuJjAFFP5tpdWAoZRugm7AIEh9L7BGyE2bK3xvynGFbCLS
+Q4HR6qev939h42saFN4WH7wmcELnbwcJfrzzNlpX6UvlXvEp9YvWIYq3QfgKKTi
BUUMnFVC118eR7Ax0rgMTTiT2yzURN/aELWaSSt+Wh4iIW75gKULOdosmefXxiov
SYh+jucHAA8g47jBPbx+G8qZllxTXASbxiN9YHJC2qts6DVLTMxicsdm2yrgXang
xazalCfC9WJ3IrmdEz3eowuX8qH9CR/CPDMC3AmiM9uRomVUMH/ViOo/mR9mRTS2
i06LoELeR6O0bD1aI3wy5mp4nSwJExMid94QmEhtDKbZnuqw15/bKaz7kf1uyQpP
TxOw6MNfLNXmhDHUL62nAgBTK58ouwXEiya1oyhkLoEst17ACnKm4IIPUbsif6ol
37mAkiu9COpoOUlgm+2Et/mRpv8YzW+IPB02eE1yWSuSqvGzCbb/zmO6LXSZWQGA
pRl8xPqr8WH+HmmxTsPwdXyyP5qS/QMJh3j73RDn0tskU2V0c0Aj07h84Em8qbZ2
qBPzZisVbuexBqR12CVzxZ/ZGhebsnjUEczGSCvJBF3qaJXGfDBx9lKV7akoZK9l
CbdYFgNNucDjYtYsMDVByhSrXXdrQ/azrJIH7bj4Pno=
`protect end_protected
