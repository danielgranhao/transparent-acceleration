-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
YUxMssA9aKzaqXEwpMvtBI5vD8tIIVHqoAVUG0f4WeC9Nz9kTtnPkMgSc+8Giouv
RbqpKp2a5OaO+rcV1JYoRBsJ/PpjZhYkWdcS+QGCe0D4B4em7MLLHdkGeP/uwnL2
S1iNsbXHuPIGn81vlqMBqJgApS3jrSZvb+orgj8PJ3emGlp40a5KQA==
--pragma protect end_key_block
--pragma protect digest_block
GWf3Y440Mt1Ndl7DW/msVH1lj+k=
--pragma protect end_digest_block
--pragma protect data_block
MfwdFGmG5eYtuYy5xX95pniZ4xTC1zDggZ9Pxgczgwnu/eJ2YEQMYk2YLT/SDh+3
62xBhKn5C7X+5yRwwnYzolcLU0RUct/vEzFGIQX8a4spnSHFFpLTqBULEwAO8fYf
hIzA4nYk4owbwTQKupj57m57WlIN7stWU6FyCK8Hfk1f3K+bkzJrsBlhHABv+BXI
/ydLsG/CEMO13TrewgW6zP1t1MIgYeyv2Tw4BE6wxfbt/vg7KGtDX/VR8/gOZGJr
ViRiLT3bxYfctnreqbyXq+C1q8gB436X0q33/c7bV09zyDDj+JavZXrCvOr3jrzM
YpD/H01S44rDX/XxpGO2Jvy9h8eePIs1EQyxfDaquLJm9buGPn+uvWaNC07fB3Wb
7bZP9/K9f8+acBlsYbZZFgtqmHYCU1yFIFogCx3cBZRgWM66FepX2+/FbwIgKCC9
HTBQ77IFdMLX2jFd2ZgR4APnE8KL/t4SO++6ZNofU9ybhmU+htRZkjtEbB04b/oR
kSXAWVZdeBKg5wmiRhLlbeisNNwJawdnkO5P7rh6YhC42Lf+BlpwIWi9hPUYfoay
PCzYGGLp/MUWk7HwN7JeUC9scUD1mUU8kK0MZpllp9M8fyXJ6S7IF9R+6mqGjuto
o2L9sKTB2jZ5noNE2MEtnsNkz8yiH6jyD581qJE7oviP3iL6jgHDGPB5gS27Sb/6
Qh0hqec9hAQHh1ywmXP8J5hSmwXlXJ7qPbB56tW6p208QuIAXUND1IAOlIf37bMp
KTTubCgw+u5Ea3QOej0KlcgTxN4dq1enD4tl0ih8B1l14sKPgMUypQ8PMyZlTiwp
SskvSjJWqIVlCpqI2nXztMCWGy32hn2Dx4IAWjW8zo0w6baAHD/1AGwJKCakZoiq
7LtsKfSi3gt90MecbqaUUnvdixILLFoHa3RmduMGlfiL44sD8IQgnscQgIuPMD0V
ucr7Mr77B+6jbTUejb4QfJDHnSBegNVizPHQ3vYhMnfEd4g2qEI5D29YT86k9Xnm
Hw1SfB+xR3p7vuwR4b5cT0BhmbzKwkR4otg/nBmKX0qR1PAlIXYsAIn4039vmYe4
PF9amkY33GtmJqX/RonPTt5CRXpW6bVruQCn/zKjKbaRtQwKtdbAdP2I0Bnmhdeg
Xmm3K2asclzXMiaI+whWY5UD+wqgqjgGDxkMvCPiiRykmmXWr55zl3Wte6GbIRrc
8zb738zkCf4sJQScwnQI0OO39bnVAX+Cw/lfBN3xixGQYu+W7GHrAA9S6U9xGXso
8OhyXQ/O7j2ZX+4WQZLZ7jHjGKq+Dwe0CYW7FxIRmEs4XQ0HhH9pypFRMsFF7Sq7
qv0Rwz9nPHfn8M6XxFpYWLhCWaIwSUxwvLSMT6E/Gg+LZHnsQ/vvOfQODep6HGD5
euWwprwqQSgE/qn0cvHuQJio2tTygwjFXbCBYX7oyi6+P2EBiDP1UfALmO5bn2Fs
ffZfH/NHmjqt69eKZxarKQORfZfp8bNqiQe1TzQd938iX2c3FxradFMRlbu2JN+L
NLTzVcoyB2cZStcZYiu1gtnQ/rPgwqc6dv7Qz6E/NyXReFteSCo3BpmMb/pZfjxO
tukJYNi9E2ruwxEfIe5ilcUY2quf3VRFQy96TzJ1/sFDeTwrcEuefWukpqcVTXGR
b1P7JGLoVFVytBFB57FOnJEFiiMT7j+1RfG7P4c1VxPFVyWQFEymoK3MMHKL429X
m/PJKRebP82hS7A4IkOfxeP0l2WXpCfHLFynwEOpVuHuRHdyGbxyhE8sp2ggbq3h
b8Yr3eN+simzeHeQegvpJJ6xr1bfCiZxCpZfOTFmAoyZdZklSX/lP+9vVyF8gOHh
a9gLxRMyu/zEv4jr/Qe3ItGrj8ftsMpas/qt+TTB0s6Z/YnvpFw7j4RVni0mFRhR
WtrUulXr8CH7EgNR4zMuamTfLqkbVf9eo2cPqPXBQtRcWNHnAQ8TD4JzkqSRZzm7
bjrcsHALPp8aVkBR4bS6k3czOfMQ3XoHNNkIRLbV02KUc5V8ODk91AOjcwX2VAuX
/ygH3brw4HQHVLCrlTgm4NyYlv95xl1BB/1ttVfp4LrsgMKv90fcj5cv5Vf5Yxbe
82dXMpBSgXGHUpdbQdMLR/Yaiu8Oose+xlLsE7uA5N+gsZnb5YwnFDIMI1oO6LND
dUG0kkn8H0ZH+8u1Hwr91JphWsv+jSIITb5g+8BbI3bEWe7rUI1WruSqBQR4Z0lI
vSE+nM9WgnDTmNih9Dq1w53H8XmaBTSwoKht9amYKA4zsDYxi0mLA9HUpQLpPAkn
KtlroWBBNk8G4q7qGCjjH6vXdYAIdv2R8cgVZWkDC8EsWSFlDMrJoaSXepo1KEsW
Wp2cmzMU8qgwh+/aAWAFuCLxSfXxe2kmqKlj569WvhMO90hTcBdCk5o6SmbYRd+7
ZJLCLZzPzhGmovEyVfCrOULir820WeYNMocHNX9Sn1UrpTFF7jcC29eGA92v4bAm
ECLNQpZuum43lbOXQ5BbuepcKH9K2eaIWiQ9VbIj6FtuTcBrNXP0T1+nSYwKrbgC
akJ4MWekiF19GKiOWXcptCi7tN7O0+f0xSNoVQUtEIPRHot8bKtpZfJ30Tc3OuA4
rABn8sPHnKSUzcZfTmNLNVnsnuD2JGr/xZ6jmHFGIhOhCvvhhU3abR/BJ8T9tBNO
xovXvQcVLBcdVtPYHJuE+oDlVeoF6CQjjfkPfWbDo8emKGgnh/miSQaClVbnU/w9
S+c118jDK71D5i53+IUMSbD8suOyrf/sRmv1+MJItsZEFUTXyANbeffw29rz7ZNR
boCA1u/TZoakk471X2WWBS1NTRyuOYsj0UItTh/CqoJiH2EWAbYBE9K8oxHkCaHJ
Tb0/YqwpXWPAoJvZFaXT7ng65F63rTiDK2Mafc3RegAcD4f4hwaqFwgKEZkGo4C8
XRSNW3jE28nBhT0TXjjfvblVh+4xngOjIe4V1Nf3Lig00BhOHU6bRhOXWpQuE6Zv
RR2/2mL6JJsF+DQVgRnDRjftZL68rg5xRTwhAnJpwyl4J9ZjXZj92BRA+9UaYa/N
KR5myPKGylNipcEVTNaob3e8RL1RMxoiV9hmMd9Gv/y1pbhTxpX0eDAh6zTLuFcR
am98uIL47MisknK0nc45eQe2/yRGtTNX2nC5daFr85987cfT+fDTtleIo47pNCjG
ozcuVmCipiYDicKbTD+8rBDoAszLax7IDhV82N4g+IKa8Zdw5V+0gR4aWCNiur/G
ewVsjWuPEukX0IyizYTZvTkzuMfdQW1a//OGX0zDbS5LI3AQpnFEPwVFtTgT96vL
sZTE9Emw+vNNJhn8jKwcxEuRUJosD+M+n1RodLVnG65QdHUKBlOtp1zsnOdOliuz
vnE3izLEysj+N/17H9cIKpowpcPLur2lER6YjqGdnKCh7jiSsTMmjuJY5YIrn/y9
usN1Ah24460bNVXghWAqQm/zAuHMXL1iWznKfxeiIgDpT90vsB0ODTkE0DL1BoOA
WdlvErJxIWV/VgNv+q/Ao+GQcmpTeXrzVTphYc8baMGmJvSUd95IaFfpfycoGlg9
9xZ8Tvemka2iEvFlD00byj4qaF7V/KkfHBuHAlxGIA+w43hjbj1vDB4DvSMP4BN2
4dD+6rVoaLSnm6fjlp2SGFoK6IJ307AW9i07bifSSSJmVo2ijp4BKDwEM3ywkyzm
+Jr0i0ocln4v/JBjwEtX6FQjN4UeSdi24Fi+q8eT6O64JC0sP81lz7P0YfuTIDiQ
6RxNf41RUBn24yqjv9uO3v3ys0tJFXYrtdy1Il2zOsfwIAupwGg5hCV8VI7MPm8J
ymRIoVAHSOKnt4u6dBq8jTbcsC60nq8jTfb2whp5/aZt/p4WA2pBqmpOCdrtUqm/
o7A0CgNaqVBmFqAqHxtp4xTcF+IuqOQqUA05fr4QJE3degmyXoj+4LsyyrAObP6e
GHPEdYjQRP1zvcZGZX98U0SRC410mHG4zFvns0Fi1IkZTgIZU5Ye/nx+1AFWJplu
LWVtdnTBi2ZWLfr7RTLxrGWTWr1waj4DxKZeRKzr3EHDZe8KL36o6K13YX4h0v9s
dahUXK0YcSljWf8ameMRxM2tlG6VjgdJDcQA4LnMzZjLOETMElMW8sJDXn3ILHAJ
V2/yipZtU462Gpv4O2RhEp4azNyQtWyz18eA3A10ZOxVjC4K4Xho3LxI8CH6s6Qc
or1FnZVBua4+lc+/xj29nemxmn3yE/+av8SZ7HoaNFXvtWMB6qiYbYviF9r3Fkd2
8CfSbqyu0pFutCsYWwEx4KF6DFokxSuKnpyY8XCW36QhaQoOAznO4y9ww0qSvoVF
NcwxVX/qAnXzylG//q6r6ryxdbOgOYwH+tm/ArehZppRU+W/M0Jfbf8nQFtlSZ5N
0NbL51mI7jKc7gr4vSLL5+QLhECcKwG7HYcMpPu4VeC4r/4sl/jvVl6PF5ZfusCl
lOgEUeoRWR8d51Hv9f+araRnOCwDawitft3NmsJCI8pCAFqIRj8drKHrTsSoZ9SH
peNdUGbVmzRK+3P6a79PqoZjIJAKH02LqE1OHfs6tcQTkcTjkjLvBmS+lCpw0j1h
Sd/qTur1XGj5e74fR6me3j0qZO8Xl26jJCYgUnRdJTp33YEITHnpH5A5hRpZmcLV
rc9LVgcmxDfk/oeMJU4hR3uKiHsIVpnrk56B9q//2RZlxuZq0H/6nPfeVTnjpowK
nBGILzq/lvZ+40fJ4ilJe4Hj06V3x6zuqbpbUmj0GV7jDEtDzGypbvI4IiY/V+7y
73VmrhQv/Kp0SkjZx4y4U/bNVowkKLhAAqMFfiGH7OikstGiHtwahSTUhJ7vq7Jb
VliXcoxRL+cerOnh1cSgPpC68FZsfLnAEI1y4BlA9zIwyeKO6Uoh9J1HwSArdRHK
7vxtbEF8hu8+qCXkRh3XWwe5ZVHSugOss4oQS4QW8tHq46mKe/NT22NqKuHwYJNa
tIAFoR2n2kTe6pxmrLoXUSiKbPwmHwZqYNwcjXfro9zGNxGvq9qpxB/CUU4hNfJg
oLx9g3HEZn5pznPSxat0+DjTYTnUFLD4+23DDajHwTc07ykWVR5unvpOXtiXspom
Ll5jEW7yXVLN5L5PKMk0gr8bsoOH3eJBux6/u8v/yfuLwCz6hhqBbIx2E+1Cy5i1
5CytwIhTQ8a9FsWJKhL/Gls5xM84serXGaG4pEuRIwkhGIHVud/Dj4n9ZEpCErP6
AIKS87yeeIeBXDs7V6+s73GyBBygCUEbsMYns1xLB9yVo+n+ms8daKq3ko4+r4ZF
jMAt7g4Sr2UFAJqjPkQNrQg12JArLaP4uO5p3LE8NqVHMCvCaHxWeGxmrKTGnDSN
fHavoL0Talr+RADlvc68aDnPq0GBf86VVBaSVjPQZgGiSv9CoLWEN/4TSfq6Vodk
ka80lw0Q6vayBOwMH6x0mhIyJRHqorJ9T/qxFEz9QQugDBGXKneq8bNTnUTjmXBb
fu8epNEqVIPkPe06wLOTKpIsxfmBr4oGxIz6FnANNcYR2ThuFSB0uxKKz+c1NsR0
gymLa8OLcXh2tggF2TNUE+9zgGTD4Vn/eJ0Ml3yrFyDwuJJ5QWu5LfGsIJ3fCz89
anX/cAqvpaFX86C826qrHh524XjTuqP95y/aAgU69asMYG9T37LS5PJNsuIwmIuq
2v7Hdg0W0e0hCH7KNnnWT3dswvSRlsQjlUezskK1Y+coUyJycccFcbhLNJfvZlct
ZJnveOHENoTgTPzR/TrBACAE7C2fsVqFSRah4lgnYT4hpfH7SSIo/sBG5OkrYq3c
XAu3z6tYAg+UyK+o+A7Jse4T+AMVtU4pwo019/AxT8zLpiRPd8YQttW6L+Eh9jnC
kM2358M13Tdk2SGx5r03tb0822XE1Z/a1FyUHZFKVLpJX4G9JQpUqZj5+KmAIP0J
iEUpaHnrecA+kD6mOJ7pjwD71SVE9CYp03yufrmprctl4PuLij7RFtzbSgiilCEA
7bSjOmCVl6gYNsJqo6DUMCQ5K5eQ/7/XsRxDLDrGlpy3J9k6j8cXfxN0L2XlQPBM
+UIcQgBA/LLBcBKRSnhkSqKo7yUje94aoop2zLyw3e0ZE82Ik8w2PR+rBVHdpuyv
J4IbF6mAompE5ihGL5q+6zSpMw9EfsrtDcLabZ7qa53xHuCF4fzk8TxWE4uy1PBY
b8YoHSHYOw9cqJmWfCy5lAl041q3DEwB/B3ZbaEvAVTgjEKKkVit3y1XG6hiFj91
QAQnK2KIVMMWljosCH9+9nYz3rIxFD1yis84c7EbteUjwTN4M1+B33PtOQ1gfhj/
umvWAF3u8kwYii85pJAt7ern0c8z2kOA8wfB98roltj335Sc237CsBepInzVPwAt
9JLz9LxWIFhQVVOXb5Dy5RyPpkUoKbnnWSoJJ/XHH8gA6GDprFL9r32Zr+9Q0GNG
yxgpV5QZojHlBKrl9cVF8Khx6v5B0TJ7tcd3gEtaN0Fq5XrZhLWiMKdDqKC/bTrC
GLQvO8h12qPQ1G4wMnzKDbjHewpAEAan30p4mPXA04Yd9D1pCnWCrVW7xjtvAc++
tQEYSWYKYteJqCCzCSl4qOmSWzpW6qlfnuI9YBu3RdpT5beoTzVc+45EeL8T3Abc
sS5yQbCYTLCKXo17PZnbyhcRWhuplCh0BH19cICxDRM7rfu3OpCU/SUFBFBsJww4
c0xDMJMS1tNKDe5H5BG4Tv9yBfAmRqjJchHqBHi9wfltJ3eWm2OenjyapUEK27G9
8MfVL4UTPeDeuKlZhRECn6t89UK2CmaNm23WC/fFMcr0KZtORgV2scsGZomJ4Q9a
I1QESpBQDHRnRhxjfX520Be1Bkrk85uRXMyUEOBzPOCOfTkq4w9cy3xUbXf/sILU
V8MD9Ya1smGdZ8wkG1o+CtiPHMfuMHSAUAvNnShfXMvJw8UcFYjqDJrR7XauPqLA
mXEVNeXsAjvBkAJ/xA+BQzmOr/Mnp7dYQtB3cfmiSEWSOOfPMf0zkLtE5Uq192iG
EwjFA9L53kiR+nZLWlBaFw==
--pragma protect end_data_block
--pragma protect digest_block
yBr1qc4AY/aAAeQijR4jF9Gfk6o=
--pragma protect end_digest_block
--pragma protect end_protected
