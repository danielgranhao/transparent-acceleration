-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ff0PwLV4izAIIIpUKPCfYn5FdIZfoTzEdRhiHugXRdyvomSDgJzDYpN8uVbsn9BpGHJSp/XOoDvG
3SW6LGFGwP7lzDv8krtxzxtkZuxWb0jHl97dMLAr7CzNVoxT2Y1EIufStFQsoOMtp6k/0wSo61NC
hnaGuRXuY+x1Qz/oaLq+NNhmabysIs8InWWH7aJxstW3UdoXLIS4J7YWQrpeA7g4lGH498oopHay
ISBVu8DvbDHEcxyTearGzMoXLEoZfTiSsvYlXOrfpRHOvdA0L0S+hbOrWqnL5wwHgQgIMj6odQXt
9LpyZTaUeIODj/6iY9AWrNJJe7vRX7UBqaj4Bg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7232)
`protect data_block
KltfuRtkWDCtbZBIVjYJAd4Fv3aGGEqfbbxdp0QQcXU6LhE1jH8wCFhki/UHZRaE5ajCIC8iDYwG
CH2P0AU5OugANuBQxQ5BioMzlmEHpcNceYQWQ2fblZOLSeLw8mMLp+iyiVNU5T8GHrDUbmGMp2o4
M+lZpEhaeRiQR9D4AI0sH9BUH4UKEK6/zwnbgnadsAp0t8e+t9hLGtb/4mbvKeGXmpC5kBRG+KJ8
vazEYvYr0RC6WwJIV5W6sCC9hJRFPmjSe11jh4NRcW2ssaAsxAqifhkod5+OfYA7p2NLUElCXpT8
IbM/0ZChvwvg4JGy9BrcSZ+p4uKO//L3ZlMAl41D3V7WAPSxmhAVY2rCn5oUDIQ7Ofz2RaNO1Q1n
OYcuil9p4HEjGwLBf28Vi2etRkQ06ejmRI9DSKmdlKI4sYlG8TMnA61WGbHZh7bZEaw6QZfMbKuS
y6uPXempgadLmlizkhAm/F4ZvSmLE1v0WBYKaZdfQjSWZGK/lvIiUMKUpkpu80gpok5ETkb4B5rM
4RipUg3FqnFVToDKEVb8Q5lHQK1FrX8bcFpGgyWgkAmo+HlHfSXTxCtwKhAh340MNCbh5Z0TfI0/
DfpX9FlMKRJFbu2O+raoZXsJoauYV8UIwTXqFCydyxnEmll2L2UDb+TjXCmF+RY90xOZNZYV34++
KMLUCOaRMiO6vppPpyBWEdiUiin5vTZiuhLJ7dB243G5WaGXUj56bjLp8OTOxRtMVy5r+rd2qFyi
CXC6/p1oE/3kopcGFNZl1smoDbGSVf0qhMhUEqMs/ca9nhdXB8r7ruRXKkOX1y9Rv8nalR6a6SVQ
6lQKbx59sYEmN0Ymka6xQ1RLsdCNkbmq16d2ovmFR3GvsLq8PsBpN0vH6Hi8YMsd3b2R2Q2B7Z/E
XlX927l+JNEAXAmEGifqxkMxNHelRlSut64lJcH7Zvf2yfvzNCAExvg0WspgwtWstwlRPYDHETpl
yotXps6ypdkHba5Uw+/yGxjSm060Ke91+xrr/GOewzcKxpNY03iSkccgIBj3J06X06ccU3gFYV5e
3o614JVhPUHNVdRR0ytinCETmOlqDhua/P+RNNyE2RyCXMVlSddLcfC0nLoQqxSN60ceZefnZd0u
ptuBfJmMsDoJli5EdUBU2w4IqakROrcbGIx+Nu86r87oR8NXOoeUlOzhSnOHwIZNpWKevRPWTQA0
jEwzAckTBgCMygzw8E5NZ4tTMHjvN1ke7oaq2hQbz9+VvAFc4kXKvuSK1j3VlAnZxDbGKGiyJz2G
8meQjVuXkv6X9IRrsxoyHaJhOhBMoWOKZOJ5fit4FRdMKZCktrtTecitPzKKybtjMg6JuQyUtMM8
GRqOweeBepFcutpuNu6KKjyZEyIJzJC6ZUpkmRL5sEUUJfQ2QSCXxAHel3C7y/0ZNEUKOcqi8YfJ
+E3KBsWQyOEj8EIDUJKFci+/ffH3l99Nt4GWvAgptsLthzKZxTZbT3l9ugK6H4JtwRSe7rFjoLFQ
oPHWlLLjHo7KRuxzgiSZIGzifPxzeiLX5ehs0ttIeIOx4HMwPRutWVq+OUBgXCheHoJzOmZKjVYO
HrXgXmUnMhmdsg6t6uOiLWD9wTOXpsM1iEMNdd00jn0mRjFnh+7a/DuPuQtmAn9Lay4XQmXNwDSL
B4Nc7gQ5r9XcyGD+uq3UXMr5cQ/NNQVEZO56ECvfvHvZsbU142plC4zyxfMKofNmrzbpJcWU4MPe
IEUNClYjBkzph36Q6aOuu8HdrfRzRZNIF03kVOF3GIE4GH915+Ap6psyuA/XawVOZchY9R/we6+o
z7AsAVXdqceRx77Ip+ec6PcNRKJSh6NedoXN4VbNWq8apH/QWjMYz7BhAArEG793+mQix1Hexkb8
dyQ5yy+yHt+OI7jBj7w2HMfp+6u3MGxDxfg6MLnEnbwgKz+05+QzGP5sY5yHNOB/pd4H7NIbA7wx
Ht6I4YVoBwxzFftsEECgfGIasc9LcoStLHjvrFeE+RbkvBFTjZF0JWJgUfDBobvKuEPQRj7klgj8
XiciGYqrXilYadCj4oWIq177kA2WTAvBYF39BAgU3ZVpVYlSXjFpWV7I/YzGSA+6l9N0SeQjdKqy
Jkz37xZWLglomkZzYA0NJcgygEBnJRZZEa4FJ3HUCZPVWIKKIfYeqX5rHz5Diywimr9NJm8Fbj5b
BGhCDrWAcqsOEQY0kmiimbQczoebVIMmLoH6/p+tPQXTXdOR5JR/u9uLfZK3125lW9j34gcHCoY1
9h+zs/vAQJkozkNcBtbJXefEAvSnq/pchCIJrCPZ3pkEYbwIEx0YFRNZPKb80tUBcLD6ywtknfhK
410ywSQEtON9X/WcqLW52Uy0lnw0tnw3qFUx0gQJUpJHAxhvdCqSdMyhai6YCrbcZGLQ6/6fwOA4
1K94ZSGAlt9D/yF3tFdzbJPUdwyjkF2a+IelnyvfZfd7OxNGrBMhggfPq1To72V1fPhKV3lclSva
bS291copj43QhASuSHBedz15no07/xd+RqQVarlyXEXuoxrr6D5F+UqqLuMmMp8qmucPK8M/MOVT
3c94ndD49whlt7YI7M1ceIKXOCUeEtrtYiHRI+jNJqPNWWkFwi+99j0Fhs4MZs6QtcJ9sSGNZgx5
skQxlyIZbQioTcrSdZWMbJ0XiefWRpy/53WG3R+SnaWXMtG63ZKokfNSBP4FecRsQb5/+E+LZTKV
XScwrm11VhlGuOuKA/vWK6PFJP4VkE60eSgs+EYq8qzqBzEqE+ctLceRFt49enIhhismIIgy8bkZ
clg5RaZnc7EfIlSIfxW5WDFDLbMK4DJ642bizhm2YeFi5oL6ccmZaFrDS0wEgqXl0Rz7sSqKlZvj
hFuaaE9zh3vCtsR8CFeBawp2YXGF6JJKaUfvPCVo3Fitsnc5i2jEL5noawGNojZjyyi2sE/C4FKR
Wsem1XwSaY7GhZGPxKmUBRmU4ECOk8hi4ba58vEgTP7E+W6NGyAuFCL3UmdTCyjcjNzaR4CuRW5Y
KE6wqSj+dcMLATxbkVtXsmOvMRe9vuG3/6wNn2xtYwOP8xcnb/AhdnhYP6bS8+FJwTZgkAUc81iA
16Ldf5tSKr/hXRez0EZxYCPfRp6mlZa2mGGEs7XWw8AiwzH2P5Bn+o3hC29EnJqa8ChieT8C9STN
4oZ1RZ3/uWSTecL0FrRbpwBRun6r42V87RlokulnbID8nuDxDRQdWZ5raE8b9wdh85eIWXGmHfje
+HKUuQhxyrkTbZ2Di1lEq2EqetQJ3Pr3l9YbV2SXYF6ZFazwIHpqCiSRjplNQEy7O3nw/v/XTepg
M9eBJs3DapmzPBSlVAZ0zDDsHgRtDqGLk7UmfJ0IaPgaie1/L1tFS44uuldwFY21Kttal6S5H+py
iInjltUUUKfW9pdYcfnCXrPoB9J09DHUlAQgbpXrB509lcwiF60qhyjrJwIFZOdaajbgAXxqHkOH
U8O3FHWkh+UFkMU/DDY+s4ndzBlfaXpcjOxqquUcKfbDCY1H7BgwAa6UYdWoMr9yRVDHvJg47vRM
aXQEszOY+v/6Z0YoOqVILBk/ueR0r+Uztzze2xJ/kg7vjDJzoWm+3z9tHFrURckg5fTI+A/lLqbW
TbIEzl/cTFRkHFs/UibkM5nd5SPWbiz51/K5QP9kdN+MZTUwuPc4zActqOZomCiYoiZxq5vnGms+
lyxOA5LV9JwYpneMu5tbIWhneZwR+G/PiY2NPEWVTtDHQ0ymQBJVFHvuT/Sx8Try68RLoRxeATyX
h7HeYM6yb9pTfUQ2Nhg0x6Zp8lRJEtCaqMD0OUrx1arq/bYG2P5F4bka5//wcNbkwJVjW5vIpHh+
xlYUnSFoQ/SKplJMZPxKOOiQfE7a37SB01xFaLdCiUkCHOE9G+FetT0DMefMYSBy4Y7h2QhGbwng
zs3ZvMF6WtkjTFFX6fAQZ2uvtoPuVC4u9RrnkQzVDX87mbveWGt89TiMN4CQAjkoV8Ya445hPyyd
o28wuFW94yhOTZvCiLd1f6FjCK4iXgwUcp/J6j2LTpRsHxSxwN1N1uwPtVDEFVmYPFZadpCsLxK/
MgqRT5zOjDRQmApxuSvyX86BvSJ5GVgTzhn0jg83X91G1gCngkkjyoL3ISclKBN2HtqLHYOh35i1
6LpLdarVoOda+yKsBWUzRrEGXTX65aFv/JUIUV5zAM2gh2B6WD7758Cnl02hCIZVxr0zC4Kh9JKI
6WDojrxoBAzk/W+yJRK+hXx7NxA2OzIfcBaTBbdgv4PU5iLzU6cEd2gcQCP5PWSZk0JGRDGy63bA
HYQZ3n04IVbBY1SmKy3bGGvwIkU6SwsIkqRUHKvQz4MRdMEmZCx/6Wfg8ordnOixeXtTafssQqKR
jClnfx3r3L0qpNWOVM9zF3fqGfPO8yFjPYkCi2ilSbBVPCrb/CfpKqgrNcn+uI++s9ZTnXqlvece
Ux7Rv0NL8oTNZJpQ5IzzzrdO/FnQZwnCJzJ507znNi4dFRayRYIIK+dwY3/vG4PtEZHqgpTGLcyL
QNHI9yZiJLiLeIeiihkXmOazOWakMTVIWloYKR9IaTD6rKbdc+PeLfX5FDY1VowqcXagbtN7hXnM
TbjNcZVPvvK2eBfAIzvXHGU1Kd3hlx5CkPjPkTvrrNozJ15W5QnJBY2mLfEiGxygnzL28lFH/oj5
z07V/lJKIVJvtA6CopfGoEfklhA7khdDLxqOvy9o/EMHw6dGjwnToFDyFW3fe0fn3I0youvPCLvq
9f31xqFzOBVsvc3plCVoNi29dhTKUSjDC1hxWV3B01ZOBdMZnAfAVBd43Qt4BFtW1lx+CA4JvAub
5ef9rNV7cRML2G6R+LYycniQ8Efl8UM1x+GntC7BfGWq8CiJQCdq/spTvEykrnCAjcK85SeYPgMP
tF93+7qF8PcZZUWzXGeIdUugGxlowffffKva6pBYFg18pj6iL9KbjlvaHtdmHeymWagYzS82NkhC
1zM9Cz959BqyoBzVdRVtKMjmhdomF3vEI9t8f0fSU4efWewurn7y24NtygkYPdKyHcmnhud2L1e9
NkAkDM3hrJKINdKPogsU+8tDd2Te1Zsx1rZ07UPchgnvUk2/8oGGbCdQn/Parg9BAnHksBSqYyI+
aixtT8jCyxdOJG33eGSnfLonQf3Aopv7CTNO0siDiCgfhEJhpdJuF+smI3u2rtn4SmyY8wsDS/dG
Y1BEmWrmBz0FTBPsaDO9L+YZP8sbMGWnYiSxP0DCpgNU7Iuv/xkvqnhXLHe3YSYuKOyYLWld7ubU
JiuBOv7GYK01CUQZY4rwP8ethUXhIFD1VMAI/l3JlL7FwT9gesWDLSUboATd1B+f7IFBG5F+4p9P
vjsJTHtu/q/Ew2nf7ePGQ+fR88ZdbE7gM1/zbSFxeJD/25zIzfuUD1QAt8HynWO6YDnUATbkuFys
YwGjgOUq9Zj+UwwebhVwjk1dwJjLhI9ldYrcSxeQI41zZT/g4bWxM0EchLEtUHKLCpAc5oM6yFhq
/ZrdWDEzIgukbzz5mBQTSujGlF3DWOeardJQ6O0ljvIndP5D3bqYt90Wvy0lQ2O/PyGv/U+0m9pz
2VR4MdlUSAFliZEqp/zf/lRB3rXgtWv8c1/R9aaaR4z5djXpg+FXT7XOaZz52E3hi+qJOVyJCRD7
gtcMNvlKRl2bi0677u7gyHhF27QGecfxR5k/MUiXd2d0KMDg0lHCul1J8DmcPo9u7OY9QM3B1p/b
dAsP5uIerfPYCTWy8z7TbkLYO3qfgy4oGIxQLbAEFf0Imf8gxaqKV3RLb94GQmSgfp0C/7nuq7VY
H2wpi74q5U2zm18YiR5PCEPTfSzcUSs2jBhiDfT5QXyL61MLNzmVta7J6qDIhH7TsxOI+9LbS685
vPxFAJw3qH7IFPQ5VzgU0hd9cndVeCiL9TFFnyCSJS4W6XIUhv1pe8RG7Y+60xsQ+w6zw7qMzuGg
eFN1r2b3DLcY998vHcJkcsnx4W9J5iFg6VdoapmjBKXfHePj+FFaNyyRCTgxaruIukEfZdaomFoP
g9aFVThBIhTFEbt9p9evFBCMEjEr0UPAeBsJsNj8vu+bipE2Zb/KQxmCEzDp0zEs9gV7xtxatH3t
Di9z13lLvziCSRVOX6Ku0eO7y4u0gazrLCvUanpgaNYDNQFz981l2oxpxQmAtqjxh5QvEEgSOp9o
+4Nh6hqK+KjQNO7Ubb+ctSTP7isADl6IfzEYGcf/Zos8s+phnJKMUz4bB1YAkwFIvbbbFaOddLcQ
LYwGtDcPNgiakM0KCDbUSMVCanrurwrw8idzXASr7HrKkY0pBk8tkqtpdXSjQUpg+zTUr71AnRRL
K7QccR79U1dFzPB68D7pLzyLpnQCsF7nVOX5GYRNeJkB/s67b5/UAtS/4XSexWynkqn/Ssu+C4gQ
cPqbWPJmKObQPDxnF31zV18HUNiGt3qkA6n4SCqxiTPyNl7EsYQglCjenyZ5Ia06jFIsRNT8yrVM
fBpcqhzLzFi/r+8SRyMsUjyrjm8xtiVZy1Jyd/xdQwhTcivgzVstcjmAXFiBGClY1zfqRZikF73D
B6FGC6BrhorMOtS4PHdPNgCtG5mOcaETGdzLi4B1zivOLRJBKWGnQTHEv0znlHMB0ctNkMcSpGTN
zglE4TB+v3e5cg5EaYD4WPWEloFQl41xY6DD4uTDqNeA6p6P3fPYVxvnI1OQky3wdsvsyR9XLn9W
lS0lCF/lcH7prAioZtf0i27LYeCuoLuqHXOUIKfft8S2mCpHnXy7eUNgeqr2ovU2BtJxScyrWsBn
q5TqdN49bY9E762Ef1fr5qoM5mYvmw8KhEUd5bFmkRbm9Q1lgVMN98W1h8QQGS/rEIVGgUWYu6D2
jw844JoaAp7tjkRCJEf/zETX/YIeJkpX02xZB0jcqojQrceRXhjl6tCnEOAtVMc6dsChmVSU3PWY
SpywaVNQhEJzVQjlLghWkoRCzWkOkqfUQ6DquUSTW2PQdR1/ab9Fg5fwJoiS3fmZtXpgNFE57sao
SI0eoMNoUaHXE43YrUGruQgRhsXDgOz5KH0xaG1F0aLBV4Km4cgJZjzRkZeSGwcJVhrTVeI32kuW
Wg6p3muCwLxbpG/cMK+bO/AVDEgc2Y0LKNHXHEaeuV5lG/44gNrPquhTBiLJsabBSt64TL71kFK+
MSPucSmkT2j1+ihQg2U06LaedvkdU5z+9upjl72QxCHXk7z4fklaJ7BUSGC8iY0UuR5ghubSZfEL
div9alEh1IcapG+1H2YtFM0jjZ1oSLAs1y5s/9rJzcXQyEusHQBQjAzdJi1EQnAvaSNOSyfjrAWi
TZ3SE/YB9o45fusU3WtYM0A3q+qwbYqdQEwFAnVw824hFqloq5xke55q0UtGIzDJLCYMrW4nXX99
u/yrutCqbed4w+Rsd8ytXLF1DwCnU12Fea70w9sc0UY0R24pB/9onzAKjIoa5Du58GrtQviGPqhJ
oax161Y4GjsvpmE4drCgDyvs3wT+C/5jUi5uq6oBvYhCFc54f7gi9HyrhDBAyNglfhf04ztkHJW9
RB2jRgwhskVwYz0Wr+5cMUP+Dav2qDspjhJg/UND9XFhT0A9pCxbWemQZSjZPagEEulf3p6eBosQ
PEAZFUDubGP37IeySMII5kzFKa/09c4IR3Nr+HK4c2P4y2OVN9F6+E74X1uWUV5aSK+SQyA6X9Of
hbA3pZP51TsM3dVgFOOEVcKW7N2Gu6Rld9/tO0VRj9sMB5g2ASO/6cq1ShvTHeRlGPZJPFBESgnB
qX2M12DKgYHHB9tXpTarL4Nj/0XL/+PcQ3Q9yXw7ZvHMkFLjZ7RMEv+bwDeCbEqa0WGpEk12pC2C
ic3l9OFrcfuHj9Egd3NNh4Xyx67vrY/HQjSxeb5rcfs/YCO4lZIPNKY1TF5hinExp692+SV57pZf
aerpXUW5RPnG92yYmuRZS76STUbdckFVXphWj6rYnLnhVxSxV8ltkLP0hwB3qppFEV2NMqFrGq4m
YAwF51PKLqHB4GH6p5JuuEWl6Of2YlsgrB5KuWM3nL8slG+qkcv2qc56PoaQ+ItqA63fEkDsQwJ7
O/wjp9H6D5QyJAe/E6mRPAFXkTsaOVxAapCbTaqhejRv1W2VO2RStKbtF6LmQ/Xq7l7LQrKIaYSf
1kjIkkYv9ajs68Sb+wzkPi2jz/HBNo0Q1HrTij13GcuI8dcVXhjJLmscWrDjfrqIVrXEU3SkeARh
sTSG5sza29RXpDnt+Xvu52LEM2ZBZAHzD6E2dP+5pwzjuG8kvHdhbo60vLns5bQZpCVLaWN78Y+f
lZd3BvHI7rjd7EWgs9Cc5DdKx9SwOO6NF6XimRerAJl6/rtH+d2Je8ScXz5IyTwl2z0Xz7fmtw5h
lVfOpo502VKfcdYm+d/rIuQIAsJTbOaFgC24e6npGMBoJ3T4yQeV/e1M8wIukrb7B+zYyr4HuQD9
EhYWXxyG1kvynGN1SoCHWqYpShOybN77XjzDJ1H1ixptv8zfkNcg0ycVjfDqm86R+O5kyBIeAaW3
+mOJlN2jQJ95gkeWdR37Diyr5wQ4hZgNeADxymKVBd2GxQZWX1+81NmtFOrg52hGIpZ/1BSk2Djf
aBZJWHOcw80ALefnKoAt7G11VojpaN3Cpxi6dSK60bCv1vZlWGjNM2aRG5HPSapBsoa2Qe0y94jS
Rdzf5G30RqqaZVJIWt5fwGtHKUt1f6yQt3kSHdHh9SdaXzaeCqQt6NT+N4VfSUqBkwlPv51Zjc36
kZ25zNtHnnPQY+il/cwp/7XcRCtwOuXlUa1lNtQzEnAsPk6MvXU9axUtEn13CFRrBsA5lZfZrWXT
YdxNx/S5qLh9zYUaGtU+TShD7oRFczgRtmcvDmBoHh7DO9AA7VoBleKKFnF6yHzMcXXMXBVUBOHc
xNX6ZTHI9gIukdiGNINC396rHduD2hNODsnNOvQjQDbZvMxiUUKPxh/vHqA18SLD9OL7iZtcJ/WF
XWfVarpSbBGiJnxkrDiMXJF/9OLlYQ52iXEKhdtn93313UXxFVrCcexJbBv+WGWAAxspuhwypnbF
kDYp2b2QQVf0Z3UhDj7PGCWpsDPR8NzsssZkySBZKprr5WXQvd9FTFd8pvgoSBOEgZKKfy53nVsU
tBDilK+U3YkisnDuj90dHv+xoOUfekypl6Sgsiwkdr9qUPpkr0oOdixdCykBswfbAhW7fRbZozis
HMPLog2sS2ZFY233uj/x3qX2GKKNhNConOBf0blC5xkA9gVXmKWxScTmOzKcF0E/mCGD7/Lp2DN7
0ZboOUmZg2BJLkyF4RwJNoWqdi7aduFbv1LPH2Rvua6f5G7ZdBq3uWpWMPhJ2Kh8e1rJdqk2XKv4
T2xIbP6MquwswenQIjeYr7PBZZqSAknUn5P/fwHtEfKjdIf6NNbDTc88LmUxXED9/H6Im1MTYqPa
wbZ9VWtj32B2rves5fqZzIxwpWslHPewKUSATVhvRQ0mtPG0TnOu3kQ9cmGXCIpAA7UxetjCle+Z
Ron82Bcqc7FNAFvV+eRfrynayi0gjA6XyjY3NRBnHt8+EpYVapLD9kDRxnMPt225emU=
`protect end_protected
