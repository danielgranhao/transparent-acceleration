-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Ve9tLDPNvk+sZdrgym1upS7grVcFvxejHtmS4o36Zcy91ArV+Y3GjFWrHIdegWPe
wTkewZ5d+bN7GYYQZhV4MU8B9hhVLgMraOegDZJED2UqU8NibPYPbDTWfLslw9Rf
vBGuzcmbHAsVjENxcacChpaHTDIhj/pgaPyQQyNRzRY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 4848)
`protect data_block
g1A/xp5l/qEbs0PZLv7KI3Q120d6Vx98VISkgA5uuGe6uskte5zBaps2hUpQoNd6
VINd08zO/xmooi+gezO2MjVVP3J7YoUNdRMhoWMlrY96tJ8HHhOYEByZlfHqnUvR
JRrFi2dIO36gC6dM8ncGvGS6FtwUFKIyI76UHU3llh+B5b8uAmp5K8MGTgYbhIov
mhPKlEnEdQnul+Qk6BVy/kX6lioz+BqP5z8eVDGuucsKKVKyp4RmlmpL6CRqOCLP
G5lpEuAJAMkUIPjZ97g4LLVZUgiIuOZPayBVDjqDDzAJ1r/UuSRbXzvylVmJxOvi
mv2UcXm6UQ4SZDdguE8DI6V9BvIvkNR0nf/1TNKw60umFFh1fzSqSOPw0MQ9PEqP
W0OPaeEMEl4sf5kI/M35xAAOHXWQkmxMnEbNMZ3brnad+IvWUKQJGW41cGs88JJB
ijvkeZvnsq25TKH+9sK0GVIDDNmwVj+FcrpAIZZ1ypNO6dtNKbPk2wepp2Jpa3v+
wv+4+zGHJuT4HoULeKdkS6nlelOxVj+4YhkTaL7OwKHZ0zz2uTaUG3i/vG7tfyOJ
87ao5F7Omcquw8sVi2EV8UcWUbDa9ehpYm8qp9qrj3rRf7CRj5uZJD+BU8JdrmfA
NJ84/XDEFiv73Lexcp8epb5W8gjtKTAYkTuP9qmbpcTanr4aidoQItmLbdCHWcUf
riq4a+w804lxyKgQ2FrzE4A3Zky3iWcWv0K/6dCARUgkhoEY4PE+EpTXf7fY/Tfp
QkF8CF97z5L4z7U8+skTiX1ngRQ7GPglcbWpvbDLX2RDmOzzI8bBlcw4GbNhqiI5
LCYrbUgM8NYEzWUVUBNsi+4pLbyjNMX+mlv30cmlCbxI/FABMuj66O6AVpGZLvg/
DP2ZoRcHT6JFWXtOCzlxDzqb+yu70oCAlQUARCd9kW+OPBsK9Fnk59Har99FSDhZ
wPaJ3k/tIVdWmJP+guF46G4nl2Q09X3oXmubr5eh2ReVGo0fWpDawpmnkbSfvXKm
G0s4fx6cus1dvkhDxRRYFFMht/eQpPUkFA3NF5Uu9WLYYJWRiLvoONWAmaPbVVOW
xCbAQO6wMrEC0Q6oYUBSfa6yLuCn2y0NkpAaHPMdaHl0eQGTMon9b45WdAURDjCA
L6Y+wO1skSVEMo8uUtLvyEHuHL5SooSNnkj9gMzmYWs7Edu7A/l8T1Eiz2XhpGKp
4gWUGjNZoKwutbc/IlCYqmt/2m88CkpsyS9+D9QLppcZZMZ18fbPbBc9eGeVtONT
sN/wTKlfmfPmoJLknN7P0yZpuuSJt6Tqo6P/CjF0HRf3WVyKUjhtB9ARkF8ZTvs/
A55fT/dLGl8X6RE9uYFKedOoiqwsyPKBnVxtMKfWdp+S5Tr4DcTlT0sGBHFdP7yR
hZdgyVcxhILiLlo3J0nQCaC3+xgv9pRIwVg8Vg+NXJMHLXHoDyvk0zHSY5Se7mXt
6UX5xTQjOVNHl98BDfICOTfXcEh56IFXayq8+eaEZuJdjlQ2+bm97B9IvF7Ue7TB
Y0lCGag9EFLkn+6LTFv5WH7MtIsBfj+3/k4KtSbM/QwhdT14QW0iVeQUXFHhbL9G
F4Nko6gMzsfTkxYk8dnmNvoYcgnUP+7/dUcOuajkEe6hGjApzWR7LkWB6h3/+Mim
G9JkfAY1oWhigrj2Qu2Ijlh/8iT1yDkMN0fpQsnRvPnCj1izMNsOtaGJ6q4KDsUr
ogFccndFbJs03nFPSMq1jU6n14EEhHrssG+BPvxoS1old1ursJTWDcAKDNT55tCF
VpWo5le39gZB6MyduOw5g2B7QfesTYc7kSFJieQUK/1rS1b3a0m1QX8C2i8QltDI
GqhsYFN6bOgQoUe4FeaVuLIB0LCapyrGdPm5Ydq74NDvGngwHYuCO1YgLR5kJ375
VsVww/GBMdZhXYyOKeYv/OyoxJv1zfYB/BkGJmnBuE9WPrM5f6r/UljYcknaPrds
2FBF8I2213Y6Bjxz6jONJ0QLNXoi0i7aC+7Tk5RfaFhWZSY/ujbhHHOsASodTdFE
23D4YSJGZhVPWTg4zcTosjgM9EggYGw7KcF7pXBfCSyOvg48Slip+xlQZmInwc+8
6CfcdAqCz6aVCKkNGNGv8rz41fPgRMftst11xfvNqwfSHP87RxYI5PSttbOEOaBv
sznQcgnKnDKUrOOYy1c3c5iVBUhR165eyOkjAvIM70DMvDQU0O/84wgKOqjR80Yz
Sgfvr34uOhfd/m+T+wuppy4CaI/O603G0SkVwTPFwpYUh6wN7e5frrvJ5FzIyjuR
HoE/NaDUMCt2fzp8G2UVQgxHEEswzcSUMW7v6WzsjtBtlHYUDzu13ZrFyJ0OYHnY
58BvfE/HJOApX6t670IvTvU15kgY2k0xab6I8fEIJw59Jek19u1OsJvJf6DTP+Pe
SH33sNUj7xCb7ixC9FKEzwIrg0xiJgdy65bMth/el8NAkJhVazQK7zrsqiIPpfcL
LVwvFl00OKAzblG2oIJqT107tbDAHXSWbI4M3g6K5VqxowdHPg3AUDsEe7RPsxmh
i/dDX8K8Gb0zo1XEv/7mbpvEivxBVOQifviF4R06eV7HSvMIy2PQFCwOmkc0f1sR
lDpEk6o0zsJPzykXQn7jYGtz6ItrlcBAr7+DKERgz5DD2+dlkn/fo+6Im3B+nvF0
9lnarpb8gRwFlWF1jM+eOhDVMZ6R//LvtGKPUQRZBo/Ryu5lwVyxmq12Z/AW2fU9
tJW7xIH45X8b2fwhW5aEZQFHz04SOniQC3/ITKBzXZXb/mHXugCbUd9j7gdXlIGg
TUxEnnZOa0ILy49qydTzWO2FJzJpm7pAf6T+AqroHTQt9mJVLDH48qOGXJFGyDdz
aRxjZxFlSWd9TF9avQly+55iyMmzp5urwAZKFNY0B4Fl/iClL59DTaZPX6Fkw5S2
E9FCayWOGzQf2xnnQ4empP5O/w9nCvpV869I7i/WvApRtBMRe7B0XA5Egp3Ghq76
4n7Xg6wKesDAVBFtkI4IIWEf/3dFaOs8aIpy/Tn2Y1AIvrOQj953NSZOJzl6e4a4
1x2YKNug9MEo/i+4PR6bG/T+ctInhiA7LE23kon6dYjbdn5MBsSB+IzOGaNJNsIJ
E7xtq+X4KhrEwQs+x8Tc5WkCe1WzheKuNDevAU68cPXuwAuBgy8XELeBE2+UhSuW
jDhETWvvJJQTFFdUwZ48C4nklGDugqjvNIDIqrN+WFXkqV3nSCA5vOis9k3GLX3b
nd7z4ZS+Uxi9jNkpTncqA0RHH9vgrZVpOHVhvP2seJWZZJ9cZok16yflkm9s5rdN
wxjUIaJNCAuEyZb9Ap8rnAayrbnzxyMmTEZIdWLaVJf2gPTvD6p86qFmnfe0VY0F
ZKt/BkYnJGNreYnKL8rhmYig4Bw49XR5E90qTKbvBmchlA8G9MutOiDE5eNpBYXP
IlVQBFbPBkrdv42Hhg9nJ/aNpQ4c3jVFnFP/CmGp6hmerxd3sLo3G0gUF+PIoG/U
QKbj8DrQvcenX0gk3UkhVldplnQb0ZUwRGT4isHoGlY4EK57zc7ocxd1Mu/oUkt+
GjKbexTBaTKFeCKnd1waa5GHjQnL1c5Z+xRGjr/SvH/C+MeWXsjnaym3Vrc9Xfx9
jM70u4NJ04QuF6myXaBHsYP4W5jYLg/2Rey4KXGq2zbz7WXmpkdON3NQTIeCi/ic
LXAHd3skb+U5ntKjW/N6bEagoQ1IHfv9JY1TqbLele3p127gnuLfDdl03/9PDk6J
ko/E9/UnaVgwv6R52q6grZH+fPrZPwz0r3DvBKryqpWOmLgJmILSTdduYyIHkMKc
Eqxb4CAJclIq1XTVO6ikS/r+8HjyCMjecF8NxybrHQuDq3/BVrbdSL7AKzxTLFn5
cHlSJVRrVLE04ZMc7f4lwg6Q8Nz8Icvo0skH2iPj3yivxnNw0ukz7syFKh36mYJO
TXfAvrifZAM0osDf9C7cqdD13oasvHLqwKlIiR2AkKrR8gJhGfWvw8d45md4ss6y
RrR+eZsM0yREChAI7NDVyGiOIuE5hR0DZ8QUDJqCOxIgO/4OW+WNqyOvgusho94Z
355yFrm2zfMLENSoVR+EaaTlIAU7YOng+6J+51u9cD/4aAvOi4CBLi52ZV7EdgQn
lGX6aIqM7tT+fJAyqZIkoFJXoHXM0a8yCeWa4sTjfjrWEp/d/GHpqrvjVg7JRxwF
ySSClyo6r+0/PwNlEH/Vp1gW+sqnyXIH/AfO4Ha0yvcv2RMXUWKJtxlvUMac44MH
qkFV8q8RYN7261VauaUnWnN65E5lNCqqHFl6ZePmJ02o63VJSLmXm58sia2+HCSJ
kspi4j5+KgTa1j8gZ9z8uWpn+DSHRmQ45rPUFiDKhOLnNh0ueUgMglhd793tT6ge
ye7IGIblEGkwz1+O2MShvlhdbTBRIoTnK1uVB20ehszxPzV8yIdmeKDv1lKSGi/S
YmMtP0lb2H2rTogVZrD/f3fX914UF8YqeJoYJJk/2k2BJkVTVJmDuEt51Vs9jwuz
e7FzFHkLgMgoFDkK0aQLu/0bhthMpH539KcO8lqz/TJp4OwpX4o7/fcfaV89Di/f
qbqvMYvbl2GxBDM9MpPmB6r5pJmYRN7FELK7eJ3inTOOID/1pPryfvXm8CdOqmFd
78qde/bzogXOoOC9ZpjOZ3wdw5017AjnYfpdJ/EDpRx1shQJvuOhaHSGIdaBKNnZ
YAdOFH3dXzlNXKOhEaaFUNW16gcKKHejyOezut5IUxCksJCaA7NfJDg2fVkF78S1
O6nlucWV63yFJmrm5YoIT7VV7MKRj2LFUsRYVLeawHNfBlm8HbICttoGzRDbblWp
3cCZ/hBqUCztc44gwQ+v2OrM8AZo02dB+QpmDH+zdcUUvW0WFeFIS79ohLf19P2W
zRtaTIOJdm2MW63/WIWVHfc1YfWoRhHtWYY7KTDOAL7o1Lh3QhqUbwVTtOmBycAD
SSV3TBQC3Pw4seSpIFB1Ss8FykcUh85B6Q7Gc4zJXRD5l7CsT5O/aiZdOYdIRsZ1
KWvWbzvBQUyFyxC5iYkRppCbsRc+LAc1P2ksO7Elosub7TmTtU9COacIyzC3O++r
d3LN8Kziysbq451H/z5PqJBrW6QrQyRU86E/T/kCopCiBwA3i4CjX2xxkVoC4VIZ
QriE42MIIC8vd47T1HULZmUaTLkt9SNM26iDzcPZaLOKnPGxJZrynJUtMCiwOn69
/NfTd0/PEos5d+Ih3kL92Qen7bx1W+FIw+fpYRd70ptAjbBNtrb/u3jiDYzM3fk1
JRhRdANW7DNdO6sS5tFHhMYRc2x/qgQ0qzHZbP2NA9ghzd072D4Wlic9i54UIZfH
u9XCXX0sK7Mn/N2G2cjAkfoWH4e+8aZrdFotsKa19zHlvyYHUp3cnANOvIOsS3FS
tJXEliq5Agxos3OEz2+SgoZRV6Wjb1fA9Atq+nwGTYRdrOcE56JkJO4RIDMw0mgh
/N14rhDpGcO/i8Hp8SCKC08CsFLAU7LKQL5B2jK715Am7cilmESJgKhL/bKBx4qA
gFdvPQr+W3mF7KbSEMHU4CtLQln5mXEWkdC64Z9gvxt9SZ+9dGEj2kc4tCaH2Pj/
VGIvTQO0O8DCnE7Jcp8a6/7JMkQ9DXLFPiI/mdl30PN3g5Ua5grXJlVYEH5FehOM
8mh5VcF0jiCWxuc0bfKdLSFhg1nWGCZypF3uGnn/1344nx4KS3XFhxnuAeG+ZUPm
hvEKM56TFEDxWj0m36Q+FxHtU6gaswUjJcBeN9tZJSPecXNW/KHyXcoWuJuj3Wxz
zXtoy5JRWV5wa5PN9/jJn1QKfPo9Fzoglqnl+q/xXeVEd2j0Hi+AXxakmW5T045/
6te+s5kR50UD+Bw+HCG4fmhbLHT5+YMebdgFOMRCIdM+daFOzHg52ZHfCIpZmPsu
Frwfyd90Ux2aiDTNXWQK15ep6TB1RgJQeYMhF2yO4lOk6k+jcACrg2kBjPqdgiMq
O8cxN+GuFkhlAaJiKbq1ND3/XitoPDBvqNigcYlgvmBgADAGSIDHZdSxpAf3Z6Fa
BfyvOvSWd1VsNig18bXglEL5KANerr0AwmMvh+gKu/x0EUo+dGxOV8CqmyCl0Lyj
nEeL1NAMuE//mE3iEj/hsNP2zziUAKDB7OQnBngXEI9V/2MEgDZ9O3nWfDPkR9JN
J4rcAIUM6yUO8c2emXI+ppXWEXvMxUt2Th7kHjXo/clVEHyGdsewfGJ1a9mtS3ZU
0DWg/oEilul6xng8x8KbuSRgEHvVWzv0pSCLdnLE9SzLzpdRt/nbjFBPkVBxgCAP
l8Hx/DjjxHIKA1P0KSN4uypIxCsRbDJjwHdAJnZcaUDxaJXRa5X6+G76qr6nMfxB
fPGEjV1OUP8CkaiDuEwbnDcsYUtK6sk+G8JKn7PIiUyU9AI2Ns6agQEu+n2emu5G
`protect end_protected
