-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
iviSOkgMhfZeKvJWaKlDgWz2411EYhg3Jj+U6DfzPRb8xpADDBh9hAQSQywgcry+
oyvBXx4YiBsW0NpV3nEBNH+2FArx2LAlrw/HZZ6NVeaW/XSA+NU52gtg6hw0VPn/
zjuTaiDbs00UJuWOdrw2RS93AZXl2/22X4FK8qge3+SYlyod0f9H0Q==
--pragma protect end_key_block
--pragma protect digest_block
M7iFKUDwjpfbVXwhw4bMfG2BiLw=
--pragma protect end_digest_block
--pragma protect data_block
LG5E5WaC7mLU7Mq69fVrqpINzCi+lQtnPJG7z7xqdpkgud+4uK2AcrIeDelSEFlE
lP9Ueu03fWgDgyc0GJ1EVQYPuoHmJ+QMbcp1TmV+vxjYGG1PvQvqo3oSlypcIPWw
YLztjf3CxRv3EVXlSms0jmNPN5NnOibu3NIhj218WpFq/oZDZbrxA8+buf0jGayF
8ot3lZWldGI3Jd2pyeueLDr3oVf0MUNvuJreGEPbVzD+fiaeE4cAwKxNzY3sXGGX
UZ4C9FrgOFIM1Bcx1v0fPmXwgNQ1oKvGO0h3N18OtLD9Eve4llEaIF9ReSlRjm+q
FxoCYm/IrUTaEdL8fMu/FGD4yF6vrtc6Q+B9K7NDs9xGSQSjmFWP0X8s+WAq955O
7zNkdC0WWjbr58BVH1UnVJjNnL0CJXX8Dqc40ZXRz2JmYZAFB9eg+JVKSjZsm81h
DD4hz8yJyvNs2yWBhax7cFLTnaZJ7Sn2WjTt5zOH6o7VeHTWqtvsRQVA6P2Q7ba3
SG2plqUYXDZyu1ECD2TwnWAtPj2ZsatQRlTBJlRBEwTW/9YFHdstspHGCRfWVgyl
BcxLYFPCr/C1tdKa52nPmE5pZ9ZIjt1kkGQCPLkE6Iclg5+9Hx8WJGQTUHAtYY9p
VC5om5QLzg+qJXn4aymXLm1/av280Nmsi4TV3mS1fYlpfZlM7czXJfDLHNLGm2g2
zKJltSI9OeDNjYaN2/eex7R4i9+etGTWpSIwSSekKU2pot4cO4UvtdWJLHnYgcFk
dQ6riITQHNiIf3H60GfEaZ5Yan+6YCgND6BWQsAtBz6A5haW8PV7RAiIhs1O4DCO
L4/0VcEbja0Je+ahDx1BhQjHgb6PLXDQGqtwxdxYWjXn6Ni96eoK5f32wGo/wNW/
QwbsTW5NPpXZBwU297JEw9IpR1bpZ0jCkgTy3rh+hWy7y/6EmkukkzsV4g/w8icF
qvAgbmqizJ8MPnk/mZ4hQJJOIcCzeDuU9eYrQBK8aMZAAydLEWjkSZzRYkgGO3Sa
yQo9dd/pbH11CorHfixjYWDQKleykykPadqYktmPKtfCfHS5wDn48/QiBF+QFQXE
bvqWan3vnAHsi0z+glIOKYmGQVyE9dcmDJoFV4Dn3EHzmE1kag3xFoVZRA4rrhzv
3vvdqJ/cYzH5TZN5skglELNaV7S67dZE7f6tjWRsOqysjgAFSluy0al1fd6+eyRO
z/sUA60j3zYaRz7K8kgAhL4mjbl7yxM4zVWgynPPQxSNsTVSQpm1kFlq8MhaBdH1
TmwXBopn3ro/gOGM8TPBprLzF1Y/EeQ3Vu/3tlW1SkxCykPqhlE0RUDd0lvTR02m
7uahZCzp8iZ1eDYwqkQA91Yw/ODNt+U7vP1M0EXHlMAWWiQHQ4gYrg1Rx72JpAWp
uOGUBQz4XzuUbLuREdxlvSQeHaE4vdO5IMORnHJAwuadWRN1Qc1JvwJHHl4HvUyR
sawlitDMme8VQ17k5r+nh1IomQOjswnYOFA4rkYue5U+6qWTgLR6/HPR28nW2xiC
itO4wbHBrxW5nVB0ikggYBDYf8THmD0n86zO5uRnG1zCjb4JEllR5JQAV1R05rwn
AQzJ1RyZ+NL8L1iDvqzduOXlh2KUvBn0jWpaUFzseXtU2ad8x9ZhMiXG1nD3mE0b
RCjD890nh/ms6pDSYCgzfDkoZGe/nAdYbIXkfCJa1wD91oe+Xu9StwaS0tDlOdQt
9YYoHf3ohNs4yk2jZ+AWk2hiasijDdrTffxQFeOxWwN/CiFvIXhxIpCGsRyesnE+
mqseF//f7UQabS2+Fj4t9SUIA+fTjXpiO9egjNon+J85kMNsNPzUD8uQnvR3hbMH
10aiEJ8rNaMBUenWvYC1oQxl8PuFs2eCarl0KGofay8uOQWIIwKfrHfWkTwWBEda
sKQy5YLXLA92n5DWbwUkanxCVCHOMfd5bbZe0hE573MsGiuIiuzdu+vTcMry9uiw
VDQr5/ufIZNncXQkTSUTMTs0yX2PPgp17waD7gV7TDcMN1mZwR1FvXhbI3mmmGbn
9Pi+Ozes1O/HYTuE7/NlU7qghez5Ve8Tatj/R5zH8mQZWpO/6myCFeU4CmoGzsro
SiSF8Jpd+nkU196p87XvTQ4bKl9+VarXSVgpvmPs7tQep7PDfwNswG56JpGNA9yS
Aq8LsSZNcpNGlSIw4hfVk6osd/LPAhicKki2kXYKU7Bt8+YkIKqZPEaAU4ZeK8Sb
Kx92QTlAitMEsJZaN1XxI5HcgLzimY6Im+VFBVE3yyGVTfoRH/FCR0k8hZRYh1Xz
oBYoZyTRGFsdH8VGbPWTSr0aw9NPfjx0sFfxzobMF61xBB8r9TNtKhRXaUTIOy1a
c3cUK4GGz3ikozuyNW/WM8piGwRCA5qreQZX4AzZyM0r0mhS2wchohfd/OSb+wiZ
CZ0ur5f9E7tHPHZqLLnFM8jxiIkXLaH+GPRCm0cyOfA+sTfXh1aIguVpI+fWI5JB
8G7mR3uA+r9z1Bgv+OyinVOP31ism14P/ERB92DiT7g3CsjKyy0TcjVK6gv27D/s
BJvkKwEDmisBjSfm/pXlwVjObu101x+mJzQDNtzCVUCJTYkgVRTyInCoxvqzuSY+
VrL/FDP/9M0cNTX5vanMFSc3Wfastv3pWK3Fp7jQKeZQbxhd//m1FpCqEeR98n8p
MU7vkSGWyOTpLNFPH7bDA1sDE7BCHAc0HFGwXytNPpFh+Uhgy/+O2n0n1Y8kmbRS
6XsPIYfZwdWZb4UT0An7P8OprDFn115GcBzeDmb6B/M+CPT8WUT9DvSoRlkcv6gY
M+Zc8K/M+8s1cgxRMDsRU8tjkgsrKa9c2wECCpwnDQODDsClAeI8UZB9hUXlQ0MX
E7uBHbqT1zBbJCEJb/EZJcvYn3pFNnmCuPBgwbpSMZXnxRm4MAO76hfsl8tgnYPU
im+YmaPu0XB1owJjvFXJ0OOMYv6sx8r4hqiHxU63vSXx9LgFmPfGkOhHdKzCkcFU
+DGMPI5SeLVlHQZGqQ14D3tKLWubFtHy8EBhFEO6rUDUlO/hPqkDKTSKihvd3nwd
MSb31+BSYyLU76ozdY4YcymUxj4qRjbEinKpg53gfMNSSw27jjAWo7JVrCbPJuS8
wCYWokCWB0i8koMVP1CSVXHsBp/JmQ5uBkwnTHcGJ7kGhkNZI7w4eLvYYPtN7D0b
eUWR32j5P7M0SGF0hBgXYYww9UhqAAJGAzzhxr4CiTvCa3M5h+r0PBJsWwLbR+uh
rx4RWdfklwuTRwVir6EOaukQr4+4D6+wIboDHJb6ABGMpWw3SAiuw+IL1X1Nm87o
kMlsGDkRl+uqt3J6Y8RlMecVIKqcGO3kAaaQtzi2ZqevRMTJkFcp6fQzyrpF8b24
Prfyi/YBdzFo/h28x3AljvVGePvtRc6XnwgR1lD1+DE4wQos+i4NU3nXR3lmNING
uEvRptpLDqqVcMkMJHtNnMjOBQ8jiDswhNFdD4+ReuINL4tlNmzIUnhG4OECIVuk
5UnPk1mAu2NbqMSzHhj1zHjktQpC4gdB0qP7+nBOfTSc+3fvoKFDntkRzCsbmJru
skhWkVi5sC/cODz3wFfSx3hOHOBx6kzTXxaCmQhMEXaY5CWZaG1YmJIINHFvAKJO
w+5JlUBfP/6xMQU5pzZRklAprGVlw3Ys4AZs9EeANZJ7psNHcuy1ZehibI+BvaVG
99DISVbEuA8DdLXUj6pvFV42R1wGqbs3VixMaHA6yRPNr/TM9mhBJFvtNDmBIW5f
ih2LkSuZzeTK8vmW7qLC4UMzQyn4zjzQCKb0/A2ZwkIYKsfTt7bot7o1LYHOhCDH
rUG8HU7P9LkfdD91nVYW42RoSjrzdtiIo47a03XPQC2WLzp2Tszo2XAqc2v51JuM
39Zqm/jNbRGX60y5tajzHdHxRScWej5Xs+FvRtYf5dNguwKGbxFuYEspnn/BllSY
zI5XqITz4KxXM2Ks/7ObIYG9wM3LRt1bGKR75By91RNpAEGGPeXiVG9FTl5Y2e7J
SqtEjvrhM7AEbJGUKl4cDrtrPAIh7c/hvR9hfrNVhRlg8iLTsX3T6hXwik6yS4m4
uNPb9P926CB2aqVTuI3jOz3sRCEYo04djIs3IvVE46uERxbFfr+vM+YNAl/r7GDm
knH+NGLbxk9dW+RPqJdsxaVFySVxQ4Ldb9u3ss0bSpPnZYAw6eDtOjkbdyfBULlY
QF0YUz7d2/ZbxZ9xiHbI+sXdg12lsUHVE/aXgaEsitj9ElrFzZUCuymjHBCdPGan
SqnaZMlHdtrzn0yKJoseUaz9djIBUt5waImMEyqz/lN71gFmYZJPRLciE5XP0w7s
2w+cktgUhIENrnRKRBurN/ef7Pn0RPmyDietg3OXJS3daf2uTCTDbgt9KvNFlLzP
+z7W9Essyj5qyHTrA2fwiUkVFzlAWS6qhsS61bFczaV950gYte3OTBU2IJups0Nd
9jlT2mDvIIMrwUDer/xXbwkiJuu7M9GLvdM4pdgYXhvj0QjJiYt40UZINrcrwSBq
Y5+ndtgEKA/NLditr+aUUwm0CrC11wg/xO7Ar5qJuTvLw16B1DUmdzDxDSUkfGbl
sbXUHArNijvrHz0OAgH8gU871t58x5eRIk+oTzET2F5ql3t2asOMHo3+KPca6y6g
vmh6rbKIQtkQK0uTF6Od9iwYAVynTPuYDs8/jW4SjJ906OqraXgrPhNhEE94Uviu
zB65RdY8pwzMRoZT7dqLznqzT4d9ufwylne/AkYzJ8CCWGlwFTXi+7AVPPv3jXF9
gYE8iNUT4OqzKsUOMxgd35ehzuEyBxXU5TJz624i9PmoRZpetNxsUOl5ZXsNwdAw
pYssJMav18o5LL9PBxN7yQq7Am9tvePPtGZuaanzSMysqwDG9pL4P9tX2tQNIBYL
lQuIdIvsjVaJAwZy9skuh00ueT10hTJCf5lJiSZibtoDNrRSK9m7NQM+3JMTWb5w
95KeCr6B56M+gsMl693eXh++7sHfyciyv2BiQsNwPgnwJ67nL9swXxoLYZad4Vae
kan5zqBaN6j7Tjc4UOgzYYx5hRKO+a9QvLyeN24EA+S0RTuf6NN50s8VMuIiM42t
m1I0AveSqv90X9RPxPWuqkSDJc4lJi4+A3pAG2PEPknzdjge9V71bQ1HOlg+fzt1
0NtdMMlmoxj39tjJZ4gQAtP7nH2OhnZe5fvszBwYd77UAikT7pJ2FEth2b6TXgsl
Ov2ItmT5P1Ai49jCZtP89enfa5rhDUT/M5JexvKSBYaJSMpwrrA9zhSiuA1SxyjI
g1+krIdFxdSPHNh94kovFwxuohh7+dygb2lHqWkV9glNuJjALiZD7wBPL1bj4o4Z
1kEx3xXNErFL7bEaqyT3tKuccoGjBGjI8pLJfMZ1fGq6qHdtnr7XQJrFtsuBNkRV
jF7juZEQTqiWtifEjpPdz+eqGGHGvw1QmXH/rMbgrbseRWCY1KhEEr1ogwdrV+Ai
5dO8rzEYYG9iY6Yh49AvYfwJaQViDddwzUBGyXqaZghgZNslFs33Q4gDzTuYolhu
bYy3WwC0JfcJRJO3Yq6WlKjYGQAqJEPFq6fCNfoXjwpbLVs7wlQdU+hZcGozjRh9
a86e1aOkxJtehRtd4ivf+F+KpflF/ui5ln2WY6Yi+/IrrXs4OEj5FsVP0uHe3QAO
pxSK4yyNbZgXtrN3DLPybdLNWz2wLnl99AnDQ6GhLL+soJjuED726DC5moX/KA8Z
vTUNEnowENTiN1URoc44Zr+daoxdbsz/kXi2hIKgc1kBW2e4qEzhFMefAscK81hr
6u6H4UYAzg0tU9CMDcZRME3raqQAQ7NS2yAw0tdPvX0NYKsTvQ11hB6FREwWQAlt
VNdcNl//n2wRVv7I1kwCN9B6qWi/UD9FvORr1Ms9oW+Z//hATMtvblAP0KoUll7E
80iGpOWaC9/HLxoPH+UsbuUnM3RJeHuv7rH4wYrwGRRxODSvZYmDZ1RndLhSkpbR
MyKLLQ5au6lHh9Sv0ueEyUdF3B3sSxkq6SZYbPcOrAzBT3qYOca76zMjIzt3N4DC
8XSwO3beOyeXdvh8jQ+s1+DhfBnLPQBA/KEm+8kCC0tLR6LhNtElrFdBYZDifrlS
lnkmGTZ+J8U5UGYlh/qEdjl5cHdsD4LxEABvd3UP30y/TV+0Tkc6XxxClbyfnT0j
c0MydVFGnxK15yhPPejfDsJjluOccD3owsXyf8FSIaFworT24WUWqlfb7Th9Pk0A
+kkP535BJd6Nk9/e0COE986m+rTF/IoQ5pOGt6uiax1BnMiQpR1+k8uIXZx0Krx8
k27unE5y0SFqCmilcl8GXeOXPYAGfWxuifzsfKmVIZNoxWTA+bFPe2p6zEO3e22M
fkoVmi3CPHm+AKTwK2tCchRz0QTuNezbjjA6hme1vRtuuNta4LmoqtziSi/Wwk6r
li+gkmSZkgseXKeNyGWKnciC7bXv06ktWEhLXdUTgUQS8H9M4c29eZhCFkqH4On9
z1wK+8O3LWX9dYBNNbQaEoZXMsTesOvhQ7mfpPqSnfqy72x+C/cQ9tBFiZQjaLkT
1bn23NG5tJ5/g27w1QUTp+q/klB667ghOFZiB8leFfLnm8cx17UR9Bba2BkNxpgn
uWcsiOKYRfF5/pnMh57xuBBBUejnZoWObTgon5gufJX+P/hLg715IKzX40sxn75O
V4XMa0j3iq9yAN3C1+VPyF1ezE29XlnG9q2qXjcAKu49DhiytIHyk/aV9MDLlL8+
Bmuop84mucNEN1mrM394lAEAQZwqROgxsxRsIYJGVvfZeFPlCeD5CtDIHqIc2PCl
EsvqX/f23bJzs5rKigDujARKPeHA0gAYl/mQYN2SZxvuApNkxXW8HDBskOPcrFAT
X9ex/zIhWctpURfRx2/9JEdIr/do5h+xrWVw/CIDor1wDXq8oMXcMvsxhVDLia9K
ogAN5D/vEv42l1smoOq+U4EjlDYYsqW18gPDDhE696h39fcN7Ee16yi7mEZPt/9i
C2bFQ0XAsJyINci75cRK0EpOwnKg1wZoxvEWp+iWi5nkYGtcfRdLL71sf0jgoAli
vmblrrmnzmWLxI0wzz2VJn7pERl/JsChvmluU5QXErr3NjgKsfsEUkMFrNFlBdkl
ymgycRxZUx+LORFOJKIsynmVHLRqL2UvkZOww6rDjb/tehvniO1ijTZ84ELGYHN7
mb+q1wLDOnBFIS1aesV2k+DFb2CeQglfFZqldigZR+j4sBnBucfyRPVgvbN9qrd3
i3gQ9X4r28MbGatUEuGNOQ1dD/MM5n0BZco7+GgAKQlA0W//XAZWtzmFI47KCpLX
hIXl+FmxhPsftYH8DJo5xjjGOPzj1HIhVLwv9BXdAS8knuZDhQ3r6AJv2pwOgtvC
KJBw1hdH+kBgA/mOO+HMfCWfeubX5c/BjMh8yShQPVl3gbGPnTGbKrjWngsPzzqk
c/2G7MAYFj4sPhgrkX3s7R3vEii1u0nR/hUCGBVPv2wL7c/a2n+yF3EcibOlL4EE
JPIdPlJ57C2o+wr3OPgidhwCbzLr/r00JHaArowC4EJ01RuxBW4SMybrXgMlkS9b
/rJBgtFNil8pdk1ZGKaWTCec3VHSDnaxnj1uNJX2Bw2vCC8c+IvPutmXfiGoPCEe
bGwmqpuCRaMW8Eso/IgsCba7LxXqRQ7RbXan+knvv3FygEdmd8nMeDGAZwCgM1Il
VT8lXfsvDy25Qdakjm/LPkRmZjmaRm14cNewIPT3KAnCjzYlPcoA7yn3x8Y47f7d
H0UVB2LRIyC0nLoJvlZzElp1LE1KdMyq6kn/TeoqVJ7UFD5vizF3eI4oM46vb+aS
FOBAzR6oieGdl+8qIat4tfyT3t7Vyq6N/bR4rZBnHNyGKgeAsZuHxa7WljeIgnLv
ELDfP9Zjk9DuqjGawCjiP0Kcmtji8y8ceN6Z2FN/y9pWWDTUvHWdWD/DVOUnvIMq
B3/N0mcPYEH5uMqI2Iu4AKoYzDF/5qOWeyZvvaJRXT4iuh8WaRLT9hij7ozLFRG/
sTmREXqYCCyKbDhIQX5nSB8uDj6XoX1knplPNu9MtQZODFV/RtbINjkxQsrFj54P
UCMI2z2G0xD/fb1xLIhPZpNeSSRC/kjMpfqHgciHyUZBl8XPw/6ZnyvdroovXSnX
cJXtjUBQgaTiH3nu4/NPbgRBpJ/pSiNrVLd1tSs9Htf6AO4vOeS3KRPgqEztX6qH
LdpA5dtH+hp+Spvs0Es0c8xXCMa4lUbxpyMRDZHuiTo4oGUu+Gz6qut+OPJsB2NH
2C/vJJQtj4WcdoI+PVEjNW7M4L9+hccS/UOjkW5RfuS4vobC1ziNE8FCnmQ+N9+m
QZW+ZhpLISwKbV13MwkwChRJV/h7g8HI1/o65GPOfl8bmzcFwCsAGMCoHu58xqQJ
mdCLPZdIjP4Bl3yy5S2ohPmZx2H/9mAHRcGx1JSYo3ydFfYwLhdqGj3JlCbnIa7l
jEKKVBcnWzBEmRfp/nG2GaLNlfAsKYXf/UUyGq0F5PgF/JCAGtEpkjikKKBFVL4b
rZkSK46FJ+lJiA8ARKDvnWmaaFdXAa1oSP3Zgypp4RWNmEXrV9MhuaVynvZs6Sqc
Me4CxHtuwMawGGo8thY5fvfoGZOsx6X1AiZEWp0c9IoUDwzs2QjqzSoYtPOmzgZ1
lXnno4AKjwkygQPkN5ZUwokOjH/kMUrtFip75i0A0pVZWavXYp8cGj/0ycxb9Xty
d2tsPCJbS9D9SnRk7TJfj9CLcWBM0dX6CpF0w/kLxE6PYgk0RcxVLJPbjThk0kUO
71vZThC+5TEAbdDSI+ee8EYXoXDY7H/qTXJ2MdHHH0TlGwttKngKkGD82leAOl2I
L6kq/hcyngOHbBbCRmfK4iHXFRsATFBG+YcunSF9MBQsI2xi7rU/JAx+BxPqGb7R
sk9In4pWBHsip0OYBwkAB/qo3USlDx4pot2i9hB+hlCmjjriCZ/C3CadRojg1GIq
M7sdh08i80f65mYLzL/cIuhVSCJPwhNuF1wS1059hzY9rN8t5dXYfU0BfW7x8B5N
nnl31u7r4ix3eIVWXoqVdi67TnPdvgqOMLjOoQPcGP5PV/zXbOvhKRhEgb11gbZg
6nZkacKWhYC+jJubftlX1gVtyWbGqaMVhTPUKdStzQki8YB7vsYRxeqr/nc3VCFo
hgb2fSqnLQrQnOeYJBVYVaMufwOzpl4oAMumVNfoEDQPvohXR8LJ9d5iCkTsLWFq
Zjs3GpIEsOvXbRWPVqW9J9cR/ZWFz9q8F4P792rLGkMkyTz4rt8g1x7Lvzj8g8F2
tAj3XC9TcX5/vpQ3+FG3YhlM+o3yKG0TxbewSGTBiLW5U86vod9G1PnyH+Hxedsb
P6dOPODDi3IGXE+znqk5/lr2iXAfsEy9d3TC9rh2m61Q+XU+WfwpbbJns22qqIZU
rWi8v5Ktx3HxuE7mzuejxepmFiURNUXF6WPj52/hVlqu00UC6MORcoZpFxsIEc/f
ai55OSqBpoMv4BYYTeex6CPGfPO+YW439bTsmoDlz6RylBat0KXRghzo0lwAG+yv
3kFCVluTH3NOEWk5qmUyEVBt0hq2GEDsSMv5pNVWnkqEEbr1CpEJC/Syi/wZt83o
0Mo4vXvtYwhOoLbtmFmRCEtZNvSatne6++xZFcalPM3Kl54jYW/xWVRN9hBbpG0l
pKlj8pYB4NFZ1yLvnrbI9Dwam2hRIVLyXGU6jIvYDI6SJW4aqKbHUx9kdVxyKvaF
hGSk7YxGaZW3RP+Sgz2jgUq24BL2nR1QkatnZ1bye5SsVcl8YXK38Xr88YySpX7F
trJX6ynv8v0iBwR5R/WjrxK49zCJ8/1pPZqxq/mAjgYUd+9gnzQs4rLrc+O2HwYQ
cNhCyD/uoXblrq6A8IShBbzVv8PZXLIHlTtfdBigaCE0tWIesGTAgPrhMs3QxQ4v
6PUoRoH3mysGDHK20QsYXrViUheISwak2pK/fkUXOi9KbvMM4l1v0AtfXmPyYCnq
AGcTqLQjfkzvTpOgcTcM3aU541iJ0zBXf/qwKlYzPZmvkjAB8EDgW5JRbLu0TWwZ
mr+hS1jOZQ1tchlE3QjZceBmejJexnOWpeH/rbTT/Lmv1ufQ7zUxr2/aRELQlCpe
JJzzxmUc/SJYcGQaXMLDcV8cP8ZIjheqiuai2xro7opYeQ0ZuqnaSMUrmAjB6Bx5
JML3z5kUZF/n2XtCtyJuiMBeP67g1d3Fv8t6lIkYZ8okI+4Ox1xQ7NLKQ2lx/pkn
QdUjgzQRA91WwsGC42j/WD/29aUsav1oL9nPme0kAcfnUAOHFbNolzc3OgNSCH6P
15jGakkKtxoRfz8ZaMlknC4rWm9jverj9UjB9pjk8YlCK/GTkPRCnW5Hky2o3Oa6
Srq7z8QegEpDqdtXNI1a3wnJp4wwt+R6JZbxGMl/nRAIGusr7vnsv1qj6WqxgJjp
Qxqsz1P5dte5xllQfRcFYKvNsplXYR825/SRwTaC0w9yypf+DxDS55rLto7Wrgue
pe7sDhfE2JRZmd3bI7vV5a9XGFRObpzp6+4C0NcXjcGf0F2FDbZGM6XiIDuj6ohP
sZ+yWbGTqqzX9hsseokmv54FMpFUb1kYjkk2peOJDdsdliRF765GwChefaKRb4u1
XYde6QOJI4ZYvjXJ4AErTc3y8nuNXLN1PcDth9eHVWaohwr60YCiGEjilUchRHLt
4HkQvic38ACrIVjDOoXwm8HTwQGdWGppXDKZav7KZ2k28idFVAdhQaeCDO2v2Dkp
HpY27NN6awwakmdtMvj+XFwb/P+eWNbpk8Hr0FaUEwgf/sEpQlC0UoBv/f1L04Zu
kb8Ost/B55nZ1YLumZNWlM9wbbT8jtO4tB8TyJ60qq8/WZwbajvqs/RO4nTUhJqe
h/8wUUvgR/FqQNYTgeaLH97st9cScSFlw5AhFvYFlb1HyXbfePTEEFv/vqGcKoeL
HwvsMQjihvS2zWGqzjzu5m61jownVen8K4AYNkaZjaul4bJmPUkuVn5adgKyzvci
IlJvi0OdcQ8GozqDFOLgkc2+YIeBTPS1jWNLY5CVY5Kx0TZWgzKr3JCe5X65b8Sw
+hpi69WeHT2+w7hXCesI5ahwNXdIL5+3wDVjxS5UT5S7zF9dRNX5iDdeIuKxSlJ6
guB0002Mkp28i0Qb5TP0j3hQVwZo809Eo6lWmPBDJp+q3+6KCK1aZbBfkdJzCshS
wvOdZgEqKQaWLIy1oLyaU5N2TTagY2dvJxQr/4YyX78T2rlZbF11J1inZa4boBf2
0tMQ+2uX7SbIJTLdEUvQQahNhz+Jrpw+xiIl5sLLU8Rl5hevnJNiWrml8vL45Cr3
ea0EgtNHAc35TxPaaiLFA3lOussmlrFR14Zw+222J9QADqUBBeA81W5nkV0aNDa/
aSRUX1Rr6jYLcHWqUkqAtSuPyYTVKjesa2jfvRbvq8magFGg52C0+pUxTCURlfnE
Tibs1EuwpJufhJ0kn1Ug3cHaVSmZy7Zfrr3FiYGa1Spy2aU8Qxk+W6C6Xw75YcHz
8HC1yZ/sTzU+f8ka9spOIAcewl4GzCNOhyu8TKcmS5kCW/WqdJiy5dr68V4hz9NE
+MTLRUMF5joY4CeTu3hxJ47iLcdkMUWVeWAnDSGvztgwuVlqI6zEMsoJQNMSqWgd
nklWR5WtuDG7AsLSsNpgSWBDApCbBRNTuDA2zN4XzcsYgaR3ie0y3DUao42zcjhG
8U5tPjmvOgsBEmcGHj0rs6oGx8d5csEeZtzYoU6DTFdZLy/PQamrnYGBMMqolsVz
KE7S+7L5L9cSh9R5BjxKJw8vUPq24wcfN0Hkh6fEcBbNcCg0jWrXbY0ZYYKrD95j
25wOC86XwkpGLSrQHh32I8geGbr5SKxx+LUXx2IMsKhW17AP7sGG72Xh3KgbDyvO
0EqZNk/CBGazDW0Qfjq50suQZqdjtptClfkZM08mywSkssriTqud68n54+b/r0HZ
ku8rsXECSq91+Fqm1KfHtgm6N1BPN7uWXzCeF2FaD3U+Ov9hWpREZsrH6COG1bu9
GXIttXv6ICp01OSPZI4qzIwJ1vOh6TkDwa5MJBaM0Po2CS+shwdktyizHcHJwjX+
lJCsP/+UUVZl1V3NMXfEhRwgeyz8+UrdcUqobYe+TS8NJMC7Zwy7i162Q295XITZ
EfBVQFON/q2cwKlb3m8svcKmP/WKeScHxiwAEIQJ4fo7I0XobTXQgD2JgpFkRZt8
O/3iKLG20XYzjVrG9h04sVV8erKHxfOG+FdnifD1h9VRoM179w1uXguJEBixUz4i
oRqA8F8VjdVcL7WDWJC6GfYNJ9cLtQbM8FCQeuU9Ine4LLPlkAoYzwHHeMqAjZ7Q
HPGmKX2EQuMTZnLTj+MpEq0Kz7ubsa8Ik/NGfQUPPt336EtGUCmKlCtz8FrgHTnu
Z5LjlP0l9SXREnjyCIoLgxT0I9+kSRe0SXdrWxxggngzjVoTnUrcpVBRQ7dzXVXr
+hx0qVp6ugpm7L4sdQbpOMW6VJU9E8UYFRtN8rt8eqr9epk+u4oxSFnmQxWGdmqw
q01HO+S2iwGgUWfkVxQ20IZw7LNFiqEj4/j1JwHFzPAzPUiyKUSlHN2wSYKI1wB5
efOh9toBVpVjZjVjZPTXppPLQT63qlBC5yFXfes6YHPjTLEm0rHsCgCPdEO/hgI/
l4oKoFhMpdqRd1yPiTzJMCG2+r7rYochvIxQwgHi7vPNCLPKuVZLt42Z+rmjL9nN
rDho/LrQRHt+NPVPHsb4W0uiZH2V9bVrYrpYTMJrx4ia5NbsToUf/FZnlehqK0+t
+/7/q1r5JlcO4bnF6QCh2ysSbahs1RsXshyzkPKeRiEjY4a0fLa7eaQQpO/BuPsV
LWRPFqvjtgXhyKd2xMm4ULBzLEfflS94TYef/n1r3KAr3xAuqvJdgwPTXQCZtB5d
lr7S1Hn3CrxEnrn+UhM3N9KilRtWF4KKVEvn5kMHh2IH3vdywQeIXSJKpnp9URQm
M8Sn++Jox/jljLSGES9PXvkPLB4PK3yNla+LiCKUyrA4k7GaBmz3Ya93CocmeMtI
wF7qybJVxUpt3P1FAXWZyrzuJoi+vOCp6hgiPDJ26kR2Sr8ZFPAvxiiaRFsE+lZr
8ZZX16puOCDDJss0O0fzmn4mBv2b7vr3omOJ0Hh32E3tfgQwU7IgDIbV2xM8Rdoz
x2Hrff0WqxnxgFvO0oLMEH0bnvMmqwtytmb8/wfw3IJCUlzQKpnahGo0Uw09Isb3
MQOWEMJLSxX06VCXZtUDo4kwJpE4SQ2ir5i/YRDcva7838TM5Xry/YCy/qLq1aHl
yAfMNMbDz9x4/o+aJi+re6495eToM+KqEHkeh6asMmS3H4kYmzlR8UyXHn/7tGna
jk4AQihwfQaEPbys6gppZiqa+6kPn0nyPFyaKyL/rA7YR2YIO1mXybXGRhJgg9cl
NOVdC//oi3aeU/Q0LBaH2jZhMRHR9IXp/obWaD1yShh45IwV5zLrBeUioZoe4TPS
0T2P2ZkLpTbxgErMvB8vjefYsNrQ2qBKkwqtGfQNlXIGWUBa+/fC2FiHUHZWO8Wg
0BcN+ZNyPUEWmPdrm7fmodUTJ9P0LZshRRVwNIDxhYclByQOfcov6RcdidI5BKIc
Qf19fnuiAMLNHVXmtWlapDdnpBTt0UPMHaFNOMJ5WfsJt1IOdFk6tdTYTgjYcDxd
0hXmrxKGKgsurbrtzJStzFl4/SfNxxhp4LxMpMBAsYSV0XoUjtOCwekgdUDQADvM
TmKZKpuXu1AYDF5JHl/EUNIvJ0hsZjDvM5vuXra1F0eYnBEFeVZU7l4MPrrzFHQt
6BAC0EPyrrnq8zlZnwpSgoyroZyyPKhKBjQzAxeZbaVcx7y7ugivHxGCCh0n2vzk
X2yTPUF+9YdJRuJMcyWu1PNx4in6e91PDi9epILvMMXFm5nCOnQZTbSv0eF9lirn
i2nbm2hsUw2YEImi+oX3CtWNF9xVQbljIX6OEHvZvexpDhPcDr4P+1NqSwjELTZu
Bh4Hb7NgAa0Bgp3IgdV5dHO6/1YCTmL/dxXShFLLJ3GQfZnZRuYaX84XoxNadC5A
yst9+VU7iTpOh1ZMdrsWpKnFgGy2q4M/e4LiXKBWcWnhnoogVPtxrItDR6zKv0ea
yYpI5rfNhLgNVQm8GnqJr2yJEkKjGlqjXUM+k6kDxB/3YTcb1JF/Vl1le75OBE94
DT+lwKfP9T5+PzKHyPtLWMjHIZFptq/K1+FLKyg0hoYfI+4KWEmVUdwGGxoQSNhn
0gHvzXDuWcpIzGj5Yfg8C2DkrllE12c16pq6DNw95HE5zp0PSteixrSKrQgP8eiH
pZG8OUyUNba4FoQqeb55rqGcv3y8xmmT54TBEV/xqmHhbI6krpoqN6UFOYIbP+iX
+X3PSu+lkmSHT808Iqizuv4FaLLOV0lyoJNiY0TAd1ZbHU+QrZV7uG8An6DOs3zM
PF1LBuhhT/b41MrXOJTp9RoFxE5/h2BOrmUuhdewHYVLjFBar0FhYAFmkQtbSayJ
NUIxDPSxBDJNR9S1B9uaDPTQu2XpfhsVQK26EWZaDyni7w8cfm59Y157OzVVrcf3
LP3Qz99ARfIjMxUVKqLuXzvpitV5/iNRU9vqgxktQ0ZeyFhgsla/iSEP9GtajYjU
/l6MHYQ7Jngfeqb0upUFxGrhtJGwHX//o1/3Ogg6plDBhh9/DqaAqtvnaqdNhGEY
tce2i8PvlrWOlC7ZhZLJh951j/jSj5y6e7cHpTxo3p2Z1KPM9GKDspEejjRtuSh+
AKZwrao/PkecMNzkO5O9i72aADgupVDD/ygWyNJYXIl/uKIs9y39EPT7lteEDNUK
IgiqhGEDMgtVN5+yFnK/YjHxkTDSvIfFEm+LFc9nCEWOZ80UFDXPhTToBO3NH/Zx
epN8JrM8z8pjRuWHP7WB5hwY1UYGczXsuMuAkrH8NZ7BMyC1loev/kLZeLxB8ZSL
6U96NlwRdFIKy0Aen2p4kMT7mBt9gYdFGdhFavYKV8nh3dV9dZH0ZEOcFi+nN+91
OPMwQGIH2UFkd3h32oXRYZPRcsMlsmRYJjqPFDZxurYbDB0zxSR0UrDS2s7vBp8X
kncnd0OqFvPncEmTatrQOLUYKrrA7N53wDS1ubDeu1QE5n8UrvK/pcnsa1LnpZKX
5tXvIV9A3QqcrwO1TyBpb6JLeyN3Y6skHhFiYINIgGToOzTFC8hi3bSOM1J32oV6
YNU1vRQJWtBhemcDqgxM974ZQWnn19EH8bJ5BodwoKB6FsgQlnnwide8MgCTOf2H
FxQIkwB4w2OHm75ZBTNFvX8YQU5nCztvNUdJqAIoXKjDKS8fqT9lbkwgLMD0JxtY
rFuKIxixInph3jjBq818zPy2kYfZUxQS6XaZmktOVsmXYdxF5IsLgPSIG9kl1ZFZ
jQsHRKyKYUDTXsvAuV41wLrcqY13D9MlFT1+lg4ry98Ablx38lDUKK2myVL8IAtb
2j1JXiIBmIV97EB5G0u1xa0LttW/HA4x9AFs2QkFqx2eJHW7coqEBMocqGVMCRM4
j1N2a/H0n65Ln2IK1UloSCyCraoYXjFRLUJxlALt5BKuZ0mMUUzg1zFYrtsqbHsL
486TUSCXhAFRKBTvfpjvBJLJyEqXVk6QXQcegpzI7MzCp7EQ2VISwdECbMAw80XU
nwoauuCq6D7qxlncb4+CyPo7eqt6C0GjF051+YogqeSIb0r7Uwp5gXdO6eA+Xxgn
dXOEuOsf08FCp+Zy7AhOk3qZPHs+XhT7Ip/LN6w75oiOgNJXn1gw9N2Df56MluiY
mlIR5Ix9TDqfsyT5aeoeTHhNt8PLEgoY2R5zDwUMgZ7eYXR8gO7sTWvZ2rRkFpv4
cTswOFwgxtgc+IOVYKQ1mSq/G4SL2P2t3UKxvBuqPSEvL4Z0i/vTNyeSxrG6uLJn
TY/OMAMxCROA1yKJrDt3nYBS6KSLu/vglYI1NsdqkjFtbNAxgP/WUleV+FnX3KTs
PYkoOQiFRXrXCH1IPHhS4AqDA1kmrf1aoiGeXmWM24QpuYFGgqFwH5bT+25i9c+u
gFJoSk76P0ahDDRbmXPWnsXXCX9WAks1jNnjZSclKY+IE4hjiasl5/JKNTB0vuV7
YuG/3kDk9ASMPb79M0Zd8PPSAFXz8olkOmPW8pJWeX6+w39HB3jszhuXLTOKr11e
IFIse5rEcwiN3fa0vTvjRhp0ol17GUbMmSUUeqGCkfIhHMbGlak3sGv+hmCZMLIj
U5zZ4OJjMky9k7/t8WckygIzxIfitzXYh9DKTRlGAlvqQDhAVuFqIQfOfzVeS5b5
QNFp9/dUoKnGZA8SZSpw2DVyEsymH63zYLHHirYFusouoqEKwXeSAl7U6GgtGVBq
7Lfs7CCT36mEqf2/nhrLau/dP1R2iTH/kaYBHhPHpSb1C2IODv7khq0I76QTFTvx
foRAGxmpqiMHyQnZeFgOeDYmL4liq+QkvpbF58XGWrNSuFL7Dhoz2D8jLbL6ygmr
JKegksryLvxJTsHAIZrhIXCZngU8+v/jG8Y6Op7MYZgQNAkPC5LLZWLFw8jt6z0M
g+Lb04YPq61rOk9TTPnnhTSF2ESZx6xcn03HJHukPu3SlN066DG2xO6yUmKoqKkJ
SbG1/Fy75+5V7q1Xs7XcCj0Bic2tCH+axsr+0kc5GsLIdsa3GhKfT4Prx2FRWiFb
mH2yM0Hk5wecDTjmETjB6NIKxGcHvRiHsIS57bHFHQDO6EMI2V4gmkkprvECfUCE
PJIPvuM7W+0Y4FVQe10M7dl1GHjyQhKWqIP26u57pryYHQKde1PUNPNwnA38ne9n
ldf8hJz39r4s56Yyjc9864tx+BB65RZc9Im2ebJkoRoLgmQaZws8jJIVLYfJKX+1
qtw3gOwnMKD6jETJt+kN9AVcI1DcaN0EFQ66cy26C6B0k3FcyLhxOoLhk32RN3tx
1rBIbiBTr7OxRqFFwtJuzRpdMHb+v4sTK2yGcN9o+na5F5Dj8ugXTxyGjhQ6urxL
fYIeK6Gls1ZP7iDrXWTlZgQHTLI1NSwbPWBsrrFyrB5Smnweg9JdxQPYwZpVlhEF
4uM3mFI+gx/aGOqVHOB/wEWHNXVGCDsEjbgCreJqONtAMVyTsOPwKL7bJWeX1Bem
XXdicJVOCfXagybxenPWtF7folKPPW3++8OZO3YObpraj4d5tzdRvJ6LASZ2+kV9
rgwGKSoLIgGqWOI5QqT3Q1/l+lUjdDKgKtd6NTkd2RtvtLFyeXFehKEQhtatALW8
vaeKOaBDVpwwUtHzJdVy94wcD7mwx5/v+8q21WMSoZ6nizlSK8DlfL4CKWvnDcu3
I2XO/5p0QczdSvDQHZN3GVUlagmWP/oAwtIJQhEYOMc+NTA9O8HlJnQxiuoNFiFF
KfMMEZ+L7ptjWNmU5YQEbh7mmMW0m4ApYcXDizvJS413j7fsnL8KqdjQrsl9W6dD
sEZ5E0AVqkwsJRB5vgQhoVpW98btZkchE3FxkZTWsTUEJG9Jmg9NATo0WMPjg4n6
egWnVTKavFYenyU4M/JayQ3xrVGLOV+hYLYrkejh6uV1USSFdgtLf7q1YaC0uAvL
r7Lgyem+iFUr2/zuV+pcKRnUMI7YCvgyQGO+9f2DpAI=
--pragma protect end_data_block
--pragma protect digest_block
NdYGYShCXUVoYEiOeTi2Dm55Sek=
--pragma protect end_digest_block
--pragma protect end_protected
