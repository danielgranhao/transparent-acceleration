-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
1Ju1+ePmYaesARc6zqPxyGIKMpT06yc2YIZZptpnLhTuteboQECGvhfinqZVDVHO
xRiHIpWOpRMR/VISsPmGbda09BRs2swNCxQOX/elYQ/gQn0gYDnfPp+0dsMmdcSM
Sxfa/QmfERdeRlM9LqDhvmMcjQ7vqtXLI30QJXeYKWw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 8704)
`protect data_block
jgC7Y0bfAzRa1eL4Px6MywasDj8py9BPoN+k9rQko2QcrXNKgGnsmy9UBR4QhA3n
uXTjfo0JCAj4F1LLD/MOFVnCpGxup6wCtQK2XoAwvBpVHzfxh55wwD3P6r2Jxgj0
m+1YT6Sqs1r9C0hJwKAiPb+nPzsyFKLN3UmDDffQLf/jGQt1dFPAFnDg32S+Hhks
EWRpwojC0+wIjsAFTdgKdxWLAySyGca0xNerXywil6YFxP8WTKeErbvvs3v+/c+I
5uAnMgR0k1J+GEIRIHvH/U7HU2rYrQmtOZWti1mHqUUgZGBnXSd63Vtb1oFyXQfc
O/iDns34xTtR3mwrRanDmCjVIEVt17kuk11DHfEazTd8rWuYqX3Ey2VBJ90kGYH0
8QO+BINCWkq3OLmecuUo3v3f7vnGSqnhEbO1dEskaGDvGcBxyv3jC9Xmz3y5yHyx
40C2H91Z5KUMWgnOvX2U98BxXtRAN3QORhSORhbH8muEv7OFKIBOMrErWPlfYTxK
ZA8fGg6AD1AKf5FL0S5BDus9aPvN2nxFNU16/c9gCZ+sw3aDQDXWbKKEFA4vIk+f
GNI78HU3tZdIQYeDC52tZ07+AW5A/sLCDY+CrlF+0SumvQYO6PfWNLBUpazzNPuJ
MBAJnfLHP+L5SQe8ozTXkrXKHGd4OeFhAvG+P+daRWNV4oPozpgRFYcyvxYKixRN
4B/p69BKYeAGM0/ge1CMZrfELablpuCuBa6Nhj8yzrpNfqkt/iIkX3B5Wk7qymfB
DenclG7w+f0DXQzS+cLnMzEsFjyHSW50CNcLrhkDYar/bmVYI+pVY9tjHUEwc4wt
w7R1RjGtx3QpklYJopYS3fAdc8msWWjnY8eSVrQIxspNf02wWK6O5nCUIwyxZHQj
ls1P0d/2lvte488Ci0eNueeb7ij0+mIIV8mflOBlGy7F6YrPWXpNU1/q77INo/z9
zgAX6Cd4F8SGUvQ0KNA/XgGkSTTkevbu2CLE/L3YsZecp/bcnGe8zNv7jC2HFrQd
zX3OkTiFcDqy801W9BCYcwOZBZR/C+LJbQ9pRMYI0HkkM9dCCYJXZK+/WBn6QIgV
qqtEiXYnswY08uijEq6XQFKhxT4sITPaT5YwQCVA2wO3Kvg4CzDTxKm4Ir8PML23
7DkzHLQQ/jCUCo5SWWdMxho4ahgC7HgdzrYoBe9SEx7e+9DTSezE0RITATzhpG1R
WJu2iK4TqQzqIO3Vb6QTaJAaNQFXaaao/iMu+kxmyLCiXCaOpEeASFc1x7nwZvLr
fyizNzg9oq2PfozJhwhIVTcKpkIQIH6a7tU2gyPuijdwNthpKippZQNh4gYCNjli
InuDeuzuLY0m1mLh/sB+hapqGbmpA09c5JH5m5NPJcxcONeWFYI5p42S6I7pFfWp
TL2ceT6+7HnNPPDmgj03JBinTDOCiIC1FZ3EpfV1up87zz92b2Ke7JmxIMCYSapG
HArTKqIlqiJh3mwMy0Pl0RsJPsGPyCBOpNh/0lU2xULwQLRCJvSBnV+DnDURiIvh
vbyYnFQblJQPKXKR0543fw5EhO/50GGVYJEEfS9/+SB/TdKm0cOlSBzu0jdQWzzd
VdHnSyoOfr736ym9UIhWOV8Vg2ZPajNEFlViRlbQ6KsuIIkNzl0jqy/T0PoubJiG
wmul0bQ1OiGKX6kvs3audqcAJlxT7oZZqrt3k1LTNBmVrNm8+U9j8m2uVOd9dlND
e/KaRRB/u+8u4DfyFAgWH80EkCGQq7s1z1OYUdcvTDae/kEfObjLVCs+4aTX2UFk
MIiHbRMF9C7M0+Kt9idRN82S2x1V1EN3/vZlkCN3YdbOgJoH0WgiDtjcgwvNYjhz
xu71UvxCeyTAn/Z4yFJE+OriFWEFhsksISiQjONs3Ct9zPwq5h2S14+HhScopgpc
QU14arBmGMWDLzjl2XKMbd8+cKyUc1YLGl8Vk4IkWvdtc8T6mZh2eic88fUFPA+B
5q7sq+VbOIYS9nEe6c7mN/5vYEGX8WMRTvHDewmRqcVSf99bKrejnntFHoWUaGy6
zv2iHPMjdp2OnEHezgfk0Mb9KBcitiOEOzmXrBvasYIzn/wJa0ZufW8+TOZFQDGX
/yh941bWuTPepzFlJ364ftpKf0Di3m+hIMuoHpbfnj6aU4rCz/6gBcxjwuBIuJNJ
KgxGutwOAWn0eNpuY4b3QQvVh1fDKjzWWb13ZyObPkCDdh6Xt0wbWb9QGnFQ807T
W+1y8Bv3S8WfQWMUXwgCzSoT/gc5VBPP/KU0pS2psd08K74HsTUY0s3F0uuoeGWg
o4XhJkMzaMOf0eKhONoKzZTSFphehaHrJ9zG5DINPveMUbowPJET9xHTYUxf4tIi
Msd1qvvHLRJfUHsxYNiRWllLmgRep61R4n9r0BgsL6JIOO3BO48LQa9/8obmbKeH
+4jxnZefWCp4N7mS2ZK2QlciMlFoxF1EOs6+E9MY6qMoGzUk1m1DLONhMzuQJLcx
1+cN2LKQ+hwJ8+dKV5zu0j11nFr0sa0mJVFbGMy86yjUgi2QH7kK5H2HW2z29s+2
umnx6pQGJFiSQtmuIWQEO10Jzn35MykDSJAbcKQPZoHtv8hW5HMrUjEywXghQvFW
j5Hoh1VLkHmz1g7R+GxnIbmRPSpl5Cn+u7Qx1ovRuwmPVa9l8c7mdfVUJfFW+Orq
UYQovRnlEFOx3Cv/goutj/RwncOKSsvL3H1lYCFNJwQ3DrivwMa542BtlruARVgc
jOrCICywFBUZlrHGKAI5slaXE+hkfk5XYgCE4pODfuSVUH+euMxER6h2OafCw0Jm
LHvaBa9wz3f5cGfgAorSCLLnDP2buuN0WK13RqnJXQl8GlW9ypxf44As8jvq9YN1
AaMgYyvuY+d9sgUK3tIKtOargMXKT5dL+EgHGNbFPcoLj2CfNdJWrQ2txojWtxTQ
8Gv4IoClCjO7Q3Za3RsejWyS3iPurWR4jgOsRSuf30cBztIww/F0XKsewC2PSoNW
SS2BzVO744nkAU3CrjkgnRShKuTScQju3QUfWBJsJf5jm/o5Gr3+Wb+IJE4YcbJ5
DT2MoIBsFPPUyO810qvO0kWUKrdEPcoOYwVcUnaAgLxGzAR6lHNLlNeHtJ1oCgUe
ogBGwmvpZrOm9tJUd2FMG7U+ByocxwWOKEG5IYW4lsR6BOWbwI3nlLqi51PHZcri
47N4oPuzDVRoqFeITRr7VS6GucbmXBVAZm/0Fomvvi9aiL9CTlZStyJlzF9YYp9f
vM19N7BeaFG60GTCkSNUeVwARn1iorbclsf/wrkkbIfQTPybEE2xmBDQJqhh6zh+
Vs/hWqx7ZjdH6N5Br60JiDMJb9skgh+fSnV+lCTvTGzvjfdUlvKV/4MC1LYcuvO5
kvp3zK9xr32zYRT02O2fi7Aefn8DPUMjwRczvtmjOd8RmoC06SR3r+ePCMTp0t8y
MWWnJ/nGHgchvh7GsuLcOeJIW6LHJsPhNeRQwhGcB8RQedI+NwuKpNchlge9RYT0
80zpFGXdqJYhVzqaNHL3XlGhLEzJOm4HAGYYKFOK4wagEiB8vA1JUaFwxJvy5jqR
TqPq5RL1vT5V2asj+CHggKi4I2Rt5LZTMDnH9uoK9s1tej9JiMJYvuwqeaXeD3uk
dujJDSsIfYiYiB6EqKo4Zplfh4SGaOxqhK7bqkMhpJCTQliXI3EDu/6QZzgImcY8
ZQnQzHlHSIc34psQFV1B6hesz48lORFgXSmVaPWI44+3wvNmYuf0FDWcNnY99vss
VpGfse3iovs2XyrPDazxji5nfyvSaLDVucLgiRDtrhVtylf0bijj335218+eTeEd
E8EAK62Tn8/+9PBQBkb3ZEKF6yieJkpRLd6AYTKtqoteDYXnZNKphq1Ws5BdVDUj
WkJ58j7AjW/npHjKB4hfD6uJeVRbUlbd34Tj0KEs1I3qwyAl8SQYulFkkMEqDyuN
BaCK/pmLuiCGNB26jjneUo47BaPFnNt92fDOD+PN9NHDSx82Xor8S4o3fO3r3Rfq
fTeAYd32OtbkknS0ivy7wrnvvb1ET6uWuqDo3YxkF9o8N+4pbm/LmF1qI5oXKG73
chnyHMOQBQUCVwCp++7wKSbJ3haOsjQNeOBe814+LvTwOXgqrw8YWbDnNc25uzx2
CG1LL4e8Unj+bqCEHQhsAOC6942BF5lKAs68b2Z0iOcrpU3cWaWE+eKmjPzgI2pH
eaeh8431PvhL4w+WPtAKRqUWMZmbwVpQVs4mqtJxUyXQS/CLJduVzkInFnJ0QLBw
g4e1pEUrXwk/DxjWItI2ssZiU4jAABPdAz8v2ipBr2cYA5YyLRi/1A6Dc7S3m5Q3
7cpE2SugNbCx3me8c2BdAK0oV8pHc3Y2MZ1hroc5oLGxmLpStf5C2SCpC7MSQsWO
WfD7DCtxU9+RkBH7Oe1s+uUvY4F9XxcX8Dlj3i3kMQCnWakEHWa5PksIayFwb/Vw
VG9h0ogRHAet+YtKN5KdPSfo0pTcTh1pwDkb79dCQ/kqypNR52ioNbstZv2EU1P0
Oao8+QY1zbhmPNHZnJ2gVd4S52/6eW8lwFLqp8H+BNtxTXb3Yneh0pO8N3YB84ZN
Om3+QX6YTHJRg5840gRRHTqREsB4mYcluCMNJJSTWSW7Q8U9tyAsuhjfaw69gdkM
eff0m9emZCnnILlohG3ceUG+f0Ii3MZ4gMXpoGyjHGVVSnQemXDMGipVetUof/zA
Q8TR7O4xeZoH1YdGNJOVOd67WA5f0OltJeORRA18n0XfZm4r8RAs0f5GUlIIITr2
tQ6GGVCfI+EeqYUYDHxSpI8L21F0xMHsiQRcpud7+2xd5ooEpBbPibLG+YUiSVsq
r/rmhz9rWndMNJU26X7pUpIadj51ceYy/DyEudepnfBfP9z+OrvJ4ahskFFbcXiW
f8Xgkz8EuJUmmJRB70HqG2uwGysLKZlIeJ1Tj0nhFHA56fAEVaXilCbQwh26pKJv
FZSNG7GpKsglWmWfETnPQj+fxY78p01ut+HVT8Zt8Idkr2CJaVWK+YCm20aG79Hq
VnU1jzBLJSL9Ip04d2m+VPvPmOsuqp7n1Zv6/OvhMTrfxZT5j+QmWCCkdq6zMGzo
Op/9tOeZJ0ki/mCj32mfOdNbWK65oZYMXdWggDxNrKtZ3w6R9V0UhG0JValYHMmz
7jypZAUiJCpEGHQelWpfp8YhxGzHpRD8oHSop5iSs1hhOOdLcGRQ8bnKOg3cgNFG
DZxuvENI6I4dWi4FnJOZ26IR0oHYzSB2/9GWkRTxDIm6zb0sRUkSfkd+Q6DALXTr
lLXy2MJgytYkzmeu41F99gPSvqn7ThPAgJ51l2jW0kjJkOpuzWzOY9ENuhOpBVIO
QuIXDLMZEyjcH8JIb1BYkqbwJWKWmPIwuz4LExCWb9ajM2PvahL/JmKOhGP7m1pz
a/ufPeHGTP/pFAi8hSx7AS3L9KrZ1qDm1MoMRr/6zLRONdjAXr2hmGvWHAlNdQOw
gA/aUWUyD9h1Zt107Dhe1fT84VQR6GoGW5BkknE1P8zCBZuqkc/SMWB4ELs+phn4
czd0S2HhKnFnD6DeUT2rAViLZsqAusEL4tRLMI9ft0layckcsadSLF9AjknADDRR
PXMuozWhFpn+i6gyfA01VosAlS3PUUh2DUyaazKbgnEwFqrtJv0ke4AwhAf2G/KI
9nAnNBD/EvAthNgydGUjljINGDqM026vAEy/TR3b0wy2esPo7hGzr6/pbmGgZGS9
Ha1Oioyx0d7kmTmGfzIt5tPk2Ve1YHZJL7BzfcFGTxamgN4qPLrcqk4I43hIV86b
6tSDT+im8PtykhVdSYS5wREsN/awi0vJ7I0PIoEp41KN/+oF3x/UwgoNN0Y+NMvu
JSRCTebX5o0ToeTKaszRQndI/jukh8R+drii8VvvSN0AdjWs7DlYbcWNJ1PIG+Mh
XUme+sS9U429ZY1dUWW41x5SmQV3guhv/XmljN2HXBJfeq0nyRbmmavVYhKG28t9
Cb7d6aIatMordCl4DoOAxdhPWt1JT4eEFBz96Ir0ui9CErE1dxeL0U7/Kz9wFdze
usTrCp2qAGBDQrcw7HjNl5Z8uQM0uaRNEWV8FJBhPrvXtysX0ba5StY4cTDi8hKC
nGj1D/NC5QUluwWXU0qBgIA+V6Ov+QccLiyTjykJyCcHwhIYOt4TUlyuuE+ZnJEd
+7C7oBMMW0EqZMxdrXMwZ6op728bESRYnLG829R0/k1Oeim4/8VsubGtmit2O07w
271IQH57V+H7zXBj24hIiIQAekSjzhajZIQOP/CykkwrwquDCNVdWmAczl8FyAsm
vGpQpW6I2/unWPk6EACevEk0+vS/kM3pkEmB1s8Z/1gXey0p+gTQHUbqWEQraHLt
EcTLS1YCPb6bV+YeVGqwEtLIFAbql6QSXN7JzAFeoFqyT7DE5cBaY/U/gbyxPB3c
h98WDNvhETID006Me53nMLLSbBlcFwzFy4LO09J+AX13MT7O8tXG/q/mqKtd02EJ
5aBTHF4Xx9FH72kcOQd/Xv5CpBTs5knuCIKmbQhL2sXyZG/jDw/FjeogPoBzVFVE
bScqIsf9VC6vzPAhvFPpesVBiY77CMu2kz7oVo7rZK7GcqJCzAnKWvKrVuR4VFRZ
+RQCmdZAO0549u//194G+nEt9ToxjPKCxl8+U7Gogzt//cxQ/FfB7WEv3HMkrl8e
w/2SGG4uzNaz5q3+ATdoy4C+43l7oMddW6FbyuQvOY8H9oha7nZ1PNcsyxqUFzAk
Yfqvz8j6QYSGZ+icfF6F7XYI39V44ZSL2I2mIK9hf/5XtXzr+7O3S7OljNQxUbhK
rhfLYm0VNYkdUlRr+tMO2pkD+lNeL/41N0UdqOXleMCqvaqaoJUbkRxi9NoYq3qr
nPCIHC9E0y8IP9ns8sIHrOq9zmd/HF869qgLaRLFncur091Ny4tISHsbltu8Vrh2
xElKUwMBVoVIQD1EAaQwz76rQrppkcrwNwGBUsfg/WBShEtkSDgtFJZ20qkbgQb8
0yTM/OulCXuj8+xJlKED1IH+Sji2UedJT6jPmkElIzljy8jcMBZ6taYedIp7Fyeh
YwjYLclY7skB8XR3qVV+l79b0SKgAWgMmq92Rx40KB2+Ku/wfWOpCcEl5c+PDN/v
QP1anDm4yrM0yZvUFhZACJiUqYacKIYuqiXJ+h7TlZqjlLuuCWTbK8n1ioHzhaiI
BKYAf1O2XfNwJPlPHIrp3p4hwq6cfTdizEylnNkMYjhOMxPK80kolyOeMccil4DB
WyfuWEusjbIrpiviiGEeITtw8E2eUhoxGuDBnYiCIT7eHLjXEqjMnneYi7Yu1HDw
W4+cbIoXyQsNQ4K8pbfGI6F3l8EAsqNOoXw+G3siOJbZxKHKDK5KTpqY8Un6mcRz
kxA3abcyXW4SbpPN5+MqSI1moP6BqdoJrKnClAGCYhAjh1cL0tZpmJAUmlwfTsdE
+2zEUGG4f0FyNNnE6W5VygjC/cEX4f30zYIYNcFYrukEIROBDwbyCVzagx1oVPFl
drK0HNpPEL5Y9ZeNPjpCm2fbo1qsg+jbqTZfrP6LP6u2gkzaxIoPmzje6Fgwa6PL
g/G0EHl8GoUHd9Vai+Wla1VAEC43S2lcIQdUbjsuHQY9PzJ7wBOz1EQGYYt2PqeU
KYgRg+Qonoc7oBCxOSWTy0+5dTVZiEMPr6YYlDVS2tfcjjsG/e9vnZtFaMH2qjS0
U8A277VvgohKI/Rcd74akzs/qIkswfoe2ypsLai4DFVR6D3oNLHppV6CszQvnAHB
vz0PGonx5k6p1Ovx2EbhGRLUdnxAwxrFGf2jZ6obFKWZC06e0UVatGJpgyusVjuu
fszyy3hXV/pT/iq2ILMr2emRkItvIlWg0J4ZC09T4R2mZPLR+dG8CqrX1Ij1AqlB
+DRmlGNfda3jR+nz2GALPrIEhzAWyHVregIjq33SOh0MuOaBf43krsdEiytaxDDW
YpSFuBdcch3T9XTS6hZOnzj9wOMXs3chu49jU0jEayC5eGULVRjF7LrgdAHNhIGq
oazMQRNzbXZdIMcdMpVkzh/bza7MEcyosDhhp/IPW97kmnycGayZH2HAOioMp7K/
pv5AWbrkIDN8NlLY3BeEMjwgPHRidy6zqAH6Kklsu4nuUUwkd2G/rvZkD7+JACpY
1yzTtag39YkyODzlt/LCjSW+EZBv8HuLjz8jIl0M+mA4Zw68olR7k29g+iHC7oKn
WDRcclN0YPLsCbP96sI2Ty6uBJAzEr8j4spQ4n3mNQsjEavZzuEOLZ2DqowkzmSU
8ZppHt3epO0Sxci51w2wv3HEtf9ZtydsF4HIGlSnkBibKF5m3EFdMjtm6xrt+wO+
wGK9d7hfSyaretpCmLA/u3cVqIkMeBczQNUHXWPhYC61Bd85zSZ1+MqhHbPXrcSY
bskubWhz7mTEPGXufH/1V5BguLO0qEz65pFyt2i/dxYOpkuyLmRLbYR+rzIn7mk0
FvcZfRaPJRk/hZAC1mGnmTUq4+0O9FTX3kKv5Mik3G4qkin1kq8d9ScKW3ft+1DG
Y/pJ2oXOQVrKcxKDsvBbISasMr3e5KUk7hCcc5nOBFZ8eUTzVUr3NfcjXx0Brcf3
Yz3zFWE+D87MZj7LpoYEmGSJofxBk1r4HFZb36WAhWPQC6SotXJRJ2Gv2RiOpJHi
a2yO9MOLelnvygr9Z9R2hMBjxVW9U79szFFXvgU4/XQ+Qr0PP0Q5OZcrL5/HRFoq
7woGdJ17YKOhIfZEf9HwPm/+rOj9+OAcoiH+7WaS4wjeCyBFA7lsYkpkYJV+yXo3
RK3/rRa4DNiR2WWg+zU8Qk6SV5f3FaBpeK4iyn/rExUl0NpjFJhSqW10qDHCMwwC
ukL/oN+tRls1vBFvYqG9e5nLF+SPEW7x1F26oh+GngxYRw8oJXc1HofQFIEzXlj1
MRy/EPeGOosMoBc8OwSY5LoQZHDtNsIcLjCbRJxnGbZP5DGLzLoFQluTTDcpV1ow
UZUhJvTsLhT+LuC9qBH6L1hJrL7aLDMR2Pr9be7mxIMKgXKA4Sc2EMh7U2xOMzaN
9faTKx08EN0xGzqU5hgPPaK6+UsIxfWEnofhijd4e/CJK/vkn8wwxpp941ft9opc
WCaxvKH2ZQSbXMj/q6vn0pR3ckhQnflZC3Yf+aVYfd4v4wZLoYyhU1FB6pgBvSyO
/l2hN6wlFlzNJDvTwRWZgWRc6zAKcMnjCVZjYlXgmp9cYkKxn+sGu+UZs2MPuvb3
ma3S1s3AySL3AU4Bb7lpsqR2voZUMbsK8onytH22zbxJ7xCBIWnOPZlaKnIXlAtl
MbvI3wb3psIzQUo/KlitItnk/OLJMPXZJ9pLQt5k5ITpr9I67vucmEqvnFB3cEjp
pZZz9g8UE6L720mUa9F/IxKF+2JQLP3B5dNflA4GtSRHzvsl3ssbNq9//IAY36bj
hc4W1GtFt1U+DOLSOOsrxe1XH9Epp2ZUyK+1jaUWRJ8pPr2K9aA3x6XQD3eH2sAf
+WZ1AmoX5ux9Ep4NBbcnEx8dsUtB1wT/IYKUdyMb9nfNKGQdK2XKOrawJeXIj2g8
1eG/9vKbVkZC15lEDZiH840sY8La4zEB9XmadLXTZ2x4kuS90DT6Yp8xZ3PoPrOL
ZRw2GNSHpBw8nH0ajeSF9JESKruFUcJzXZbQkpsYAKpAgJZwc6a3Io3cxmgrD5X8
4OycFj1aXOj8Viv93oCHgXdB+MfakMZPJCSZ6szBV1q05UVXWdSGs0aLSUy/BuIp
qj+Me4i+zEJv87OaReRCEfeoR6Z1ZwcxQ/fjKUNFLwShBirb7UV67Jr0Fe/3u6Op
+T7e/7pRI/0tuG5dMeb7Iq/WrQfTGfyOdv/7kmRZnHcAWI7WVPotra2FGMe1q5H4
ArYVh3cW7MoD05eBDBPl4FNpeYSLzN15iJDcLu+nG22iaUxZ/miJNxeL6V0ToQ3I
XHNXrk/GjuU0iCQH5JF7J1AWzJ0YCt9QLMjm8WyPBfJxOQMRgTtqX4xYyCkGMDMp
4FlSdKlWqTxBXZJqtDQT7MF2BwUIxJbu0nzMTfKKZtIg4WIxZXUnOIeLdmGHJuaC
uMMYpYrP5idPMDkAAgv2WV6D5CQAav68avvhlZaoIGZMhX36w5Xn03pP6e7mZW8W
J4Epr5G1LhwTjcsfuTyS47TO8bOOKEuyU/gEFkvD+HoCRZ8sg3YEMBfLEYZ4QKU0
JkkKcPAKzwrjn7C+ECbPrwqHPeWcsCoA8L8KFsfiMN7XcizK4XJHlzm1ZT0Ea2yK
9zL6fTOn+X5SuytNjYgHMLuNjVpKfHtURAxDksNXlVRCZOGAqjBzAiTBxrj3Quo0
T/CCvuSBxNJYjocxthBae2JOQtsGp5WL16dUFwC5bJTt5gix6iwJC297zFxCkVmL
eTNH8iR7dZ94Qt2N6gHo08rmxlK0f4+u+ewkEBPVm4rjaD8jZNsK/JDhMEZ4YHMC
jWspdd99jJ1NSkpvcqn8xttLPkmENqrafXw87a+k6+g8c/CXkszMYmuX/YCHr6pi
4M8KhdhUe/yqn1GUDfWvbFU8agatx1arGSn7KPhKXS50Yi1UBumYGxO59tssHBe4
cydCevtaVAsYYGPfK9j8lhqI5y4a1KpQ2a0DvJ9de4LGD8aPhQKODEhQWRlWQfxi
C1TIf/IQkvVshECU+3QzNHOdiEY81apbTyDGdpkk9sORKXV1ED2T1ntsLqRl1CFU
mQIlQ1Jcyc9m27xbljUvxHrGz9iqOVnJ9xlfQXXWMdKfTNfLV2o6X/lnP2QMXiNq
0B7fMTHLJT/Dz5g94k/RUsHJ+32pyds4HA9rQ1CUpIiQ8HBUf8lek9hR0YCbEK35
XwFF1LjM1Fo34GZILkqY4XJp2QZZltabCN9QZ2SkOzXU+xu4vFACQE+/Lvg1KRFs
Z5URRs8clnFNCRK2f8oTQY5qH5rMgFWmyB1hPp+Mz2gOp6bCaJhyXQaajVmz+ihQ
fXNI4Z9Tu/wVjlfz/dNWA5l/o9bNVf9yfS/t4wd1JKLEkL84meqRtDoJwKf1ILGI
QhODEjvhI+jgPq1SkSvY+yAcOCAD8DB2pEKJKGdjZMIGBSPYTIe68AbZF/xvjSMK
q1va7n4UdnmERhyWwNFIkcEmA35EecYEw7IKhaK/r2GkzUVApaLOADnn/w1Imwln
f0GkLqKTvMPLAOnyew0k2KuLThUbr7bkFIUHp+cQFfd2VnYYTT8+LGQ8mfuTSDhM
obbOFbRvGB25Z9eqZYU8/V4kX1Sbum+k6OirOjvgAJIcuFIiXpWbwJn0IEXQwI9V
Cbd/ImYEzS/mOBRZNxyFc3+i2LOdoZqf+CrV0Bur/EZ3tW7JU5qattfWNg+2gP9F
31BRoJiU2+9JipHzucurFsddN5FCD6V9fbaKkVBG2gbazn/8owy1VntQG3U2PMPg
8bjQMlp0a5JkmnYkpNQdU3V9Ov25ogzH+rbjvxJdyIObd+l5t2RURIbn9xezTaPf
dsMVJJiSDDajuaCUNw/eRts5JBGEJ6rhthgCCtX0o1GiNQTXreVLJ0yBNvFZs5wn
mqPyIEIKBzmJGfqwfcF8/g==
`protect end_protected
