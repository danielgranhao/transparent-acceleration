-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
BCOk3yIMgecHov4fegGIjyLixO5XlAVjuY0C583V02K7f2dRLDxAJ7dsmYfoTKNGqW5MrXbQGDL5
urzmuGDQmERZ08ysrQTuegBvUf5cK+HI+NjkjriTZpSWrBAyvziE/BP4FI7Oj02tPNyFok8iIKcB
ca9YeJoIJfY7FQL4O5Wiuyt2NoAH94MdE4nQuLD7dNcjMhVq4PdbqN4dKnh5Mnonq8Myca+W4XjK
rgDRiyjo0FSixhoEZQf2RvjSfjbOqJnsuTWZpDucu2tB6AtPyPuF9sBLyYX8R/QRfpzRh0m/OILB
8UarYMRkx7qEGWdoMlNxyUVsJw8gQu+Cvs2vSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 47984)
`protect data_block
NgNseKaVbUbBu/wenYfdW6RjxomIFYRTPpsNkCBmasEm1VZVZ5XuPIMl70dI47M0OSH3yW8zJvtU
JuG5GsuuKtUGWstnpaJy1iyKnggE59NBQm3kREq1QejINR+/dD38mOetUC5NcZiQbEVXLximysQP
Q9ypczpOhWkAwMNAd2bIcvUonwo6n4K7xgvBEXNiYxJ8Wh6gaq+42F5FRrJIK0EjVS8PCM2RMP8m
C4MjpINxleqw7016dHxMduB/6yfbOUvHz2LGuKdo6Ww/s3cxDCYS5TsVBQrRJ0GnSwF0Pp01Szkg
udfvkbZ81juY6nrI+8+K0RZibNMwCQ9ESgh/xwPb8d736jyi7j71i9Po1HiUb4blI3DWHoulQ7S1
HwgP4+SPDOThDoiQW9A5QZBUu95EeyKYlezFyf9iT0mdmIGfv+rcUwqTDrBoBTvO/OCh8YsXimCi
2voQmxLbLFoaQAGVGT0UlzjaXeHotLKTyBf4aJ0fh8OhML/5flzyddT9r3wqBBbghrzTTTzjGAw3
lnJKBE/BIMAqzJP1oGf1NLvCc6lIOMsarE7Vec846V84oS5YICA76+Z8mIu7U3yJyrn4Ren35fGy
ELOZquA3O2Z4iZAwES6+b2S1XatY0BgGpZvspXUch81kJa/VI/QcLTS3CZO+1xF4SnyoxjxDith+
4+Wm0CtMOulJOPaJaY0JRvB/5Oquokq2ib3zZqJe4DGWBU44X2yZo4Wb4ybQBUsOkBWoHv/CAdfY
VDzuM5nEsJPVDiU7i6NuC0P/nkfz+rFB/C6hb+PZq2XCrAPN2LvfAWv4p5mQ/c093ihYv2hnTe8U
25evNfF+fHnsmi/6wYbjxNjIjbMttCd+dnyZFNLY8X4zCoF+KKmz5v3r8zgP8hrdRE2XLdBMWtFx
z2+oeI8U8PosRRIcmeIiwv3E3Kq068UZTFzmfiJSm3aVNFQUq4Oj0kPqx0vn3jfjqb6+R1vlB8aH
rnzjgWjvr6/cnQYrN0kGXmYfkRb1u2uK70XF4E+KqBFUAv05uImlx0T5nNbrToLB1sYdlSWzHUAS
pZPIDTOJPL1f1KMyVAKJQ5Z6SZ3LNIae9xYTtN63S+5vfJqIcdYia43lQmwiLZZxhMwFePnvTlvu
Fs6W0Fu8QWAW4gL/x/4JldPZcwdxBMJbzm9xzjxYZd3ZxfZ4frEtCTx+yH9eBCYWf8ncd91tXZqq
nspUl20FqdheY2lpiGduk0lWLcclB53rwBorUCai9EJ5Klc7AJQShHP1HXMDzkEBzr7vZZwWgRHr
YvuS/EYcMoCLXEeJsw3291cWFrqlNe2EWCvGDGgvqKeLVZxlQXt8OGSUOBdJFE2mpERc2ibz04kP
x7aQAYxMDi93FGck5Ra4zJgpiojuXgYmcMSQja2ODp1sO8OLsBhE7CiLjgZ++rtp+Er3NSCA0HGW
7dk89gxcrN2tuTHYM3GQy9uxKQrsmCRtpbZSZJeqqGGcu22CTiNdyqmtIdvj+91Lu47zaE099uZv
QJGjY6v1c+3HY8G4GWa3wmKEoDFq/kwPPMQaz6O96nb8nt506q8m5HIOgMNNnbU6d3Ar501eU7iT
Y1OxA4DPfo87/k9/EvqIeToAxYDVKEjDPHMTuuEHIhwPD72z3gjeGhSo02Ns8PmPvBR90eniMZEQ
ixDTB6g+5YI+4tLjG3YYvcCBGO+cTWV6g4nd0NnqplaZri5LsRj2an3bahD6qmAcxhhipD3hfpM/
LVyAgoaFNmvxLdDsGDuZ9+wloKeI6h7t2pxQeN5pXfPT0cZnWUKGvOS8G43HVGbemVzdFsrQzccq
fYKcfq7CAzLPrQXTbflZTCYC4YiO6qNKye2YVmtetGHc0IWemooSkQhig2srIjyKWPaaRP7AMhtr
BPVuIaFfXfmo29zUrQxI6u+BPuA/Ig6S5cLbaxM4XuPZdlodBoac1pDFlyJQ4fFyp6HTshwRirqO
x4jeSRUWCBWkjvYBPkKkcUlfVXUiW2Zx5CGwVl9hfm/SXbI6VSoQIKGyYMwLAvAU48ufGXn4aq7g
Y9hODWc6TXMrj+V9TUFs6EATgqelKL90fpFeuLedqunbvytLWAGkf+C9T6yyIsYBlWUDRzZL8gAW
hL/Tsbypf5ukJ3KPSvoLUtrWl9ZuGBiL3DhI64PX9it6rj707lp02WJsr61YAzuofeyTn80jjqKH
RihwyY2GiSW+6GakhmaqNgyioKXwnHMVc9C2UfBk3pMuTMofrZnjqIkadltlj8Krdzd9Vnb9nAXs
+2JBW6pIOmAvtXD3RcG7OxJy/1ln/5khFueeC3TR2TMSj37CA5JbPo3MhbNjMy1oeFtRjPPEvEQ6
+eZr5SEjOGMsVLU1QakPVv5BYZY1Y+tyRB+wtU6YG2T1eyerWO4Drr3iyrBj3N8+x7+gsUUYE7VJ
LD4pmIlJZBDiGkgwHVuXc+Yiae+ZB3TWORDGc1uhV6os7Qd5bgaDtljXnNaD7apxQI0pWZ1TL8J4
kWDq0qRztYWulPST1p4bh09KKmPLLqMk0FF7QVz31GWCh8gG56Fd7nNLDAYT0CRKF5VDacfwJYlW
jgi9QcQabZkfp6m3cEiFg915d9bKIGbX7vub/k6/fiXyAKTqnGGEbFLDlo2JKHd1+KmbNNxXe3VI
4RXqffdJxbVPSFS6m8aL76h37YTMqgmfTv1vXl3IaFst9CYcEfkUGtdtOHWx6BN0IRDPmwUtLbL6
cP2XRCYv81+mT8uSiAuPoKNcc55hlDmyfsCajSQio1jEY/rT9d+vUKO8kXMHF6hN5oxxonVuuoth
3oHxCduyxkYb74xmNpwJIiYNCKFDtSfaFMRJR/CaHpZ9EfrMo+QCt1AbWbhcQABlslWDrVVezp9G
nl/PEmjk5PDwEufcAPfLe43cyHyHAZDQoNBgAohCzK6fCRjFrpYMmNmq+8nyT63vdkxD6Y952N7Q
CneCkWD5KVCvdRyAfsjYqTLIjWl3en/P48Kbz+kxOrIu7lCRG/QxRZCkzOMOX8L3/zDhLs63qJL4
d1M70QIgfRSPRECKEUZlm5aRZ7cJB6/mQpfcpmBZCf5WUQ/L8uPD0CKCvwaeB8smlvLxoJqp/H+H
+hIJk9Bz4JYzIKKmyclgY1+k+18Uw/KNQ0ntsG/j2JSUeQ5HvfBFv5F+BHFoqeGwqI4Wu3lIQet7
dWbkcO4DaWKiy7P/MzJxx4JJRfg5axQs20ZLON+mwun9YW2Z3AKEdJrpAYguYdFeUnwIDYgmXlkr
NP21CE/X0sYxjBXeLjE311iUdNpMSWM/qmjwljKebweR5QFFSp/qka+dUOMnl6Gy40KwX8IiR94+
NR7BmzzbKuujpOiwXTK3c4p8nPDNmuBJVQDzRemE6c1gZb8aHgTaIB652xoiC1vIxbJSW4FUbTyr
s5LQMAxXVPGqfsMBeobgosVanAmfQ9ki1QElIY407vrLP+jsNm+10dVoSpwRJaQyJMbK/rQPmbpx
8dgsGt4ttsbYAB+6ComPdjtOdglt+YFTstWmWcDlA+KuBXD1q5EumwOScT9KoPX78o/B7AJyLYBw
PLj4x/DBQeL044cqmNdro+ox2koU6+QJUU3wWRPXwTp5jiyPZAc9+ucgshCm+kbNzus6Rf2fPtbn
Czw8Br1Bkq9liFnP2DLdjDD4kIiGcJ8Me46ESH19lSz3opSttE3PEThcSeL2NCTD070aMkq1GJc/
oVOCPxtnPomRi9qNzk7KT1TaQk5EJ989gBKC2iJvXkxqqq0RFc9WAWRNL8vSaDuPX5qFGxriB1Jk
9/q0VznXK0NzWIBcVBSElNC3A5L0GEivIfgE8sWQwRPNyuROx/5ebfOYUKI/HQU4+HKw+ZNsIXyE
0AdJcPGuYe3hqfB49hf2GvNtRStxSGJr/GM3GLZ7AOuQxHSdKPl6D0wL2cHUoUslQzJIbK+g56p+
kywnhODeekfNxFP+8vX5sS6u6lyvnPvTg2FcM/XcJxSajztAAoWXyz2eZafWuXnFwOwfS+MswC5R
DnM1hV/rCX5OIEeMcQvFdhFQmzLslWPjiTNhgJ7oI41Ytoazgtiek4QGkzxLYlhv4YE16MBeyTRW
/Bo5bcib24MkvNtVVguc/I9zC2Aff2SJsJFCxGDXXISsNn1xhptC0vO9aJQlt+q185B42nBlpLQf
e9FfL3i8dN+kD119O1yH3Qc8ps6jp/9H4R0c2KZZPiASwDmQ1Ov4ArjkKSd/OVtdGgPMFQ/3S4Gu
bwCcJ/PgVobOUGsdOE7nY430n/9WfMCVQzX1Ss3+DFjdrUSP6v0RIXOmJE6m6MBL5E+zZsESAgH2
y422au7tGyOI/tl2JWuoTK9ESI417iztwV82eHeB2Qnb8l7SMxo+Qmmrz0Ofc8lc4W9Z3DTrvNSp
96XHJzTX0hsBjhZokH+ctRmfBYbI+mvMPv9Ne159+gTW1tLD4ILYICWFFx2V0Q8i7m5hFvV54p3a
B5Go0ZRA+6hMc+Pn1AlUhbpYhv9c3zAqZxmY56x6YxJP4zL1eWwvD/tQAAkMGW6uW9RHn3rL63+L
z3rGScI5Yu2WM2dVJq3jK9s7FjIkOqcJuCMx2KQNcnWHEd5JSFwp3SwXBtib5LvwMSCtQoZ/Eipc
fM8neA8/5zzRttf7VU37L2oPgRk4AP1jGDnEBgUIiTdhwRnFiXFLUm1+ZbQu6DWS8sv95CHDPhwM
x10hNlPl3P+9wYD9uSQxsgXPv7a/GfoLzsBWPRaDD83VCj6uqwQquQwqtcD9kLrIJdVRIdlwvm0c
Jl35L0b4grf8wpS2OnGdTmWv+Cn7LbWNUP0ofAvZvN8fj5Ciu1CO8mJmyOibY6dWe+0z5iBsrKpG
lAWAmTHZGLIBjSqmrvDQiZFJxxavxDnpBft2R5RbfosXd7E8cqvCz7vhfGHHSqpM2oMgW/LTXFbn
92wt6A0OMdApdsmNWJxPymzLeQwWWz4HbVwanEvMKT2EOfGU+scYvYh6hN1lE+zJ9vyw/+iIbU0z
LqBOj8wfF/3Wo1HrWFr732Zxc6OF10VX+VlDceIqwO/Kb4ovTsLMD336YwnuJVIJ6h9wMuAKWFy8
XP8BZakGWpeMcDYxeSDeXQige2Paj8+YBJKpLbg2AOxqOsuTQK+m/h4enNatLEvpSPcqQ9yH1XhR
qv/ys2lDiIZyPJA5+2Us8LSEuSJ0yrr0MYZP64Cv6VR99YLvpu05x6KxL9vpKupoTvMDJK/qKnle
elXV1688ErRqeHgs+bfSHLpjT8NWAy2L2ZJTpKRMYwWera/yiZc4RtYuZr5OrjuzcnrdcvZEBhJ+
Kl8O7iElDy233vwirA8rsVQtdj2UOncPM//eDgRC5KDxJmNihN/AHHOq+NrCDX1jo7LOn1X86RJ3
8sdWDcT8H3gWp8Fbn+waAuuKdLYaXq8swTHqXfHfsYNk5kRDx6L1AL4VL6mH/7vTB+SdLUPu2P/9
Tktt7TndbVfB0vcD9RzNZjI8zM33hNALAJtaspHNJxdZOZGPZg0EoR0L8nGJlmE7/VvOk6T+9ZWK
h8Heux6AU9YgzQk5bbw/vuQ0y21jSKjMwgxdgAQT2zbUtQKiaJBg+/upErMyYecTiyN5FDfSl1Ox
pJiKkqwfI3rip+TRLmHpAI1CUYcMuHNoMEV4ULTo5SvV/reC/8ANJtSTLf1t73FhPCmgA2kCDh0g
tmLhru0bSoI2c1ZPl/2frhuZDa027Ufy5Y9wsYYml4M3McUwGOfKvLf8oovt2rvt/FEdnZXwvYZ8
COiM7PjPx3l9ICSipD9MLIe9knTBHsUVVaPAUppeVacRd6wOQEK4VrxeEu/YOfbLBiGJ/z4kzwZZ
R4wyl8u75fjxCl9BFAVq8WxY0/K0zBSsb7ew3W3HmkDQ69vybbid6Sc4dQcZRN/v3qZCZFg7KiDT
+NHB9G9KQLNUtjYotl/aj0XC6u30kMjo5E3AbtsbNeG7C19LuiJbT6/PBCBQXytkYubXywE1oUm2
FOk6pvzhvHBFQmXbT0QFHG6E7N9gZVtDFkjHIs0o1aAiLvl8D6Gf+c76P4My3TBCpes0SAl0WxCy
SX+KqoWHjgAy4Czk7cVRLXNsQchsZyCS04OwwCbWR6FW/R1/xU8M8dvcRKWWoZ1d4yMRqgYEgJcF
a5U1NIUTRIdd0lbtvC9NvRpgkpACHEFYNB5SLsrtKR8LrRF76+0xJmU0wjDIkBBIl5x4SbnluB0b
ydWKPshIl2Ci+rHbZTP93hKted76V7A/NGGuslQyLRw6prSuAIK1ENrxU3kfBp+yt21uAvYmOgcb
VZ7jQKEEOdKG0qdzYqnNrEPqT/BTlFWhjtoYH+fte1RQ55uvSIACzMLvVBPTv4rRdWMHSVhdcXWN
NtXO569Vt4f7eb/6FZiqkUjqQbu0RDUe3hOc+uaRT1080Zm9hz5SyondEl+u88urUIaGguXqklY8
isrv0ichUrTklKE9fsQap+AnyBcWqHr1XdydOKKosFTlrEIbRtJtuv0seiuUTMjJ3Rh+DD3OBYyJ
F70q/tZ31JsJsSZnaZ2MMdmunMFIk9+E96oncZVnOs+LsE5kOAFgz/D7sJApyOKGsGf7TQiv552h
8YAem3+epl9hHHb/FGoSd0uOm8qMqjRulxQRWAuo3lGyy++8MxQ+4tKQelHTOhpyjefVndq45NUe
Lg+s+jj8Hklrx5Qh5YyBunm6gYIbciEV4En/UEO5l+UrE1/PvL87Gq9sMn6lzurQ7Rz22p6gU9WY
jyGPyaKfkkEG66cpxTOtMB8nmabWRAUQNOSIommhShvrOrfOa0GDZUqfBPI/33h9dwGgpLzgey0/
ui1nYEFARsDQ52MDECCv5hy7+IapIHtyBrPw/ruLipglkOYJkhQbcus7nri9/JzwmhGAQJeZ1b/o
AolzGvJy5oSsCgLZxcrGimdtYBzV+7JlLpseZmFSjk3zvDaHAgDhN5gOsHkQIYz7aFxlKbbHJwHt
6HAdm/V55p14IYQ0tftHwlUTZU1tGLR4cY8XGFXChRFoV/G9JMjE5owjMTyCuViPhB9d/D5+sTfs
/vaYAT0MoN8uUjkiT6O1AXNd0fEXIiIOENNoRB29HMrZcH5Nje46NuJRtM141Vv/xWRWYrWYaq9k
LkvvKjSrxDXwBjjMeYubjxWrEZbpnIExf9n/61l9mWvfcxO4HCg5uiaIB45EuMwzDgKBPt/nIRdD
zDv2Jcja/Gm0i0ygvEh1r2RVwR7fc8oS/XjtLDHuk/ExCpRWZ85xlfo6YOa+S5ndscocDNkWJkP3
IvYNkNk3Qx6nhCx8iyo1AjvkrKBXmmSGgCNl1NqgmNra7uZ/bDzpTptWga5iAMoDNSXMrE2pY5hm
J2tdDJSrB2eg7u31/yIj/gGM+DMmYAOER2U3AGOzN43mLjbg6Xbd47h2tkPK9xdyl1wb5GNe/+f6
wJALIizE1r06ZobpQ5IqMOm075Q+TZv4EBJBX6qr0v04AZbqEkJ2CQFhSWQ8AQmjXk0FehttdZm6
3YLbGUWfkgPi21pxMIMmgipF/OQH8zVZvNttGqLoYi498KHIpKTU+6plgds5iXBOMiCAONgGt2do
Duv0AFBQy/vw4c5wsgnT2xPyfPqxS5WzWiokpUjyuysomeIughZ9PmIah8togXQr/wVbCi8oY9tJ
NVcFu8qY7SbbYBDhYnMoZmFY3FUA36vkqXvghV4V1TrUC3KIxe3Nc7NeVdx6PeGPpqmTLelkio0L
A6LXnalMNaWAhyIz6B9oZIZVY0HVJw+opPt+rV2HN3csfxyXvBegUhCsVmYz3qOJk/MFxeUWftZN
0ueBrRfYOuNhFOmGivpS7Ut6e/jYgWjlcSQXG6UVsLFjCqBs/LOgtsp9wsfm/dsjQRo16NcWTqui
ITov39jKB8nppKvQZHPniA5r47SfAw/GhU4i1RADFZRuF6bGEN8ldCcE6enqBdYjnRm5c27MW23J
fbKhFUh6pDBPrVjSpdJQ2881Ps1DapKdogjnuYZRo/rcYsaV7I4CpLFDNIqDW8zkb45ZtNYKwwCs
psTqJAp0e7ObghHUTiIWim2Tm50mBs7xzAzGR/AVYB/mIf/+vEJOrEGbZSPBmvyiy1YURGio2a5w
ymjs8y6rNoBoUbLDQJakLemfwdRuXUzDBm5a5FgghbBCwDcV5wg6/KYeT1sBK+90kDP79XkfjwfZ
4IZ/4tH7ZbprHNWoFtBhLXrh5drMdUilH1mJe3W9BSL86eg/oKiVSMATDeXHLBpc6X+pcba6zA4n
MGnlrwFCkte3/Fzpxd2Fd/zcAwLfipvfM+JLhHftNmcIpgLwJxcvlrD3XFF3sd+nQv6P6wzLJeEW
RH3v0vRctZ02coRUyuCo4Zg03vJXTN1au4ytLatQ7RypZjC4jgzku1SbW5q7geb0JHtGWdYnEb1b
z3N5A++5Ebkn2p0wUKirNTLFkOurmyz6uwcXjTE1DSwpKY7fKSFFm+WYfGVflYIb9hP5Lxb+lnN8
Cf2QapJRBPY4FSogcao83qopGWkl8Gpxbz537OB4dx4juyfSsHVdcD5KRXj2ux/f6fVbQyi/ANHO
ZjbQKMaPXbJT/O2DoKtXgAhJ8BKqv7BSCezJhOh3qgQsX/nqRgkDrjyKMAjaXOcSHstsMcU6BgMM
U3CI0MoVZO96CEf+Vqytu8UAk942ZzMCHS6H7CjS4MA4V7pE68q4VFznjrQO6SrX07rRrcApIYY4
jiKUxiF/QLPYuDVEVEskPcPvWsKb+amao1tNOT2kdRacZ4Bn0VLcimabPxGnf/ReB4KCyEb0IfqV
hTsr+gE7e88EQdkeaNMIMwzkORdYa090CEWLa26vc2mLgudb08fydIBGPk6favi+Ad1aRnpPwaN7
aTuyxpVVmBFTAhyk3jkrgKd4UA7xtJXFL6dlF1e7TrHkwoZnycX73++0VuVmO0TKmtpKiz3W0unH
2cRIdidjh7rQ/9h8fbx549DUJc7XlU/Pd4MpjdPI4dDPxnLc+8yB+GkLruYB8BSD0jO3Qgj7i1Nf
Y/hvHIvAwIHRB/EVmSafML+SmJKmetb672SCzOMWf1nXgJqvamawHlMHkUT5NEVd/J6z2+XRo/sJ
SyJohmnTDRzL/Lv+wWrK3U0Ii+/wEpcAoKjCvDSu4f6TKBDbCNI1hPQiTzdNOBKts+RLByPcVilp
JjAiinEw0tI+74bgtvcHH3VbBHL1HX+kRdP3VxjGi2wcZyalEdPuvQPCzrNKksaRfQEdR87jzuhl
2saPA3cN8nCaBlH8y8Qqwg+3SxRml3zmpCy17B19N7sI1KlyGNsCFfFCwa+p6gNUcJibplgOTKjZ
lR9CvphgtY3244YmdkZOXsDzso4+HCEzGQldydSJV/2hppSi9jz36RG6N1WYcrPXm1jTY+qJ+h+D
3TSENZ4YxRoG7fhbuIRbVL2HdZSeTJPvr6X6OoaDbv5ufDsHTuLMPGZRTh13xjlGohHT8MnoiGKa
z0kuTyS94LRFnElup+5Nk3YKYYsk5gCUAtnU2ozCctJMAWhLBHjX71kUf9UybV5Lsc9BqId1BZm2
9IYIVarrihRfF97GrxUueFPaVoymwVxOx0Jfvda7/T5AEkxJ5I15ypsMcMVfiAITJu6FMGP66U4w
2ix85M46LJJsckw3CG44pqa//u5HdyQSrH+61TBOKPxrAPwcgvCpr5r5s0DIwsNkKngRszOvY/zx
5/OGlb7TO65dB+wr7VNhF1UDrEByCaUOJqVuZbL4p0T8Q0BhqVaiNgLpIUrJu6CWXpJSKpeMaUq7
+QAomDfJWzTjwJ9/smLQdaIf0nqNQkX552Uv95nX1Z5hQVGboWzxI6cqiY61xfCCDuG7wHNQZS4R
Wvnow7p8+7twqChz9xSWqEOFSvgznqLe7sTpzl9gJ941JuMG+OFKos5FSXMTQqncWFJLSaM83J75
wLDHXqsZpOPst4L/W/2MS83ou7cKKeF0krHYA/cw+MoNqzKpy1On4mdH9bNhE+0T3cdgqth2l+mQ
4Xm320y2M2bQM1EoamrqB9laUEz4za0j0QZ15hBgoA+g0bUFiTyRa+3aXUa7MsHzc/6vTKcBfxQm
+hgD8ofmOCv/hgz/wTmbogKZ8IyZfffjx4vKUiZe0tRAmBjsrFqHNuuDEjOBT//YnFlmWxf6bjSU
pYFFxlJIjFulhLOcMYEa4MRoB+Vm50In86JNXS/jnA2MK6rRvOP2ksWylRJ0QhPwDo+FcEDapN4P
DDyDWoRlIcUASfy4+Pl8BJA3s9oyHG16YwOX7ReYAED6B4ClEu0qax88RRkqaCWHI1nf+VGpqNzG
WLxY9LQ+igeoMiNLoTfG9TvGrzM9t+TnixdoDU2y2JsWBR+z2QaReThgwdiYVX8JBUJFWcNdhk/o
KyX9uMGpgwiMKQNDyfBIgGN3UCjkFVt5uIVDJtdZx6Pmx9uNZsqs0u4mJhJREDoIIHXpSowUUjPu
577MSjYAP7PFVNfD6v24LGjb8N7Ryn1/RkQxFlvIhmeeqhJ5e+CcOXxt2q7X8vCN5n8qjO0ZfwdN
4tNKMv67buVWQPJtUkTdYBIECGEeRed3DRDY15mF2Icy1453nkn5d8dwN6senFbjw8exsTCzMshc
fYXFpovpenK+ljiZC2RYZHU1pMCV9l13rpbjvri2+2wuyTjr3Vk9VoL9bnubowSvwXOq/iS+F9lK
+fLbafYvRu8abo/88SHNf3UV2ic0Jwsnxz8E7w42C7lWZvptyQ38cwEeTjyD92LeewDvImpNmJPg
Sq+It3TJqsV+h94JSrnKTgA2BPzpVSrgJfeU0/OYj81L/c1bGjp7Vjv81tJxsNJrzjA2+wiAJOxR
BusA+nz9Xdm+RdW7LJd61yXhpjFZaqUgvitU6s1TxFQqZvBICNuymOl6/OqHlbP6ZOvBvXnPLqZD
0MsuK5bX02XUm4frcbgH/Cl55nAbcShYqwAGxfPnV+7ZbN7sPG4osHoYZR11UdBiOO5/wfA+mtFF
bsfzsFNnclM9q6Kb0MDfpSCttQns9t+xluu0kbkp1HY9yLX2poPVvw3qMQ9Rz5wXEW5P7MzVLBfr
z5srDl4mXZd/zu6jchXChv6JSiu4TWc59b6GpBZPtQWKak76mPaGPGWHhySMVcW7/pJ8TSB2TuQf
acoH6Q2oZmqLqilnaAnc455oGdvn+w2nSlTE2LvmQMX35+iNZ5FPGJGhAz2Cmpq3hnUBy4w/I+QK
8PiKVRcLr0BfYNKmramjbzc/ntqPOoY8ZSiniC48U76lTEfZjx2s/C0KLoBxBuwKAR6mIy4JpMnd
F6Ztpv3fhxmAovATDCCHVPz5/ryy5rqk2apLpm9WNfWbD3rcR4ZBVPcSQfFFMDSWoOimD6LoOxvD
Jdea43F4Jz4CK4k5V+O+pUwJy9L85PyqiJDWoQ0KrILKR+HiALU02JshfB0LvE1kvJA7sDKdO1TE
JkPuZgPC9x87I7OjPM96AT1vQE3odk42ygvfRh5gTAkirZ7OhbM4IGvdIXP41dMTG1b2irciVCXF
aNhHGqvfG7TtcdbQCuO7Yri35DzmQsiyXHBIkD8OfnBR5cKxvKmTYvC1XFtxAXxY+iDZlRigyp2C
YRDTUw4bzztFFf5k5VSMTR+CWwl4ICgbsu2raFsHA2ySEAAEK5bqDp0wgTisTuDM9NhVxDX9Jet0
eFC+M0FgKEK737biztSh3NUlvYZUfcCStl5F+oMlWsa6FcIoq6Q7RAbiYbNbKqYTDI2gZZrGwl5q
eWbgV38shlXtJjRySc4XXvLywXxUgpMItTcW0JP/FBrpm2WMLT6Ki88j1j9Ns/nweNqWghAC6UbS
rvvowpmcm175EVVs7VN88B88ci5/kVUknaovXTPRJyjUtcKkMrPpbdPrypDcB76mIE9B9xobqfp+
pabYOt100Bs2ujW9C7tkrFbXcgm0tiD+qqlw9beJ55gfU8UVOYlpv83Mpjz0+/yGce99/wjt1i28
hNuFLoryWchqgVjE87hQVrWXQ3RFpiOg/VfxNlFdarvzTTgOqS7ElU+dMxU5moccMehcuQMBds4X
X45p11B70GY9hg02UX0HMCqWpTNXIpoqYmySwXUBC+lRJvxzs+WKYU1zsz3kw+jITVaJ3YWFAGpb
Ogoy2vZ89dIT4t2NJZE2KzTiqI+FmIFJ4XsVIkkiURw2bgKAqSZPOFCbpek9bA2LuZA18H2OVqKV
YDDL8ty95KbbupGqYPNKalUH8KVqvIq4DulXQm6yqM0EMM5BBDaBmGAuYDJ483pRDXL14w37xjEJ
dBR/98KPNbHvsDQwZul/1dZGuQVPzfjZXAI7C05lY7WouhYWGUEqrK+WvxLL1HJ7LVUlKo4tFbpb
UYHeJiTXb5ueshllfmzE116+228LDOz703Gn19k24Sho+v66tXTqu11r6ZQvgjLeTt6B7T0jGr8Y
g5glsmTqaYWRvNOktUQTzxB7nfAp1PeYHSuvpVnX6F7m9jS56soBoLNx+eSo6uLVratBxQ11/BRu
vkZIt6Xnu40/1A49/TJJValf9sYUWPL46noCvC92aJILiAozv4K7SPp7YymHPmmh4D56ugOIYqa/
822GIeUlDzf4j0PGRZDawLCbGDTmR7gCR+dt0ldxDW6mnyFrc7wJ2KQSSsSlAgiZ7iwLWEUOVCqN
uvwK4cqjukIXdmWm6TfmuKYhlPV+1DF55M3GVE4G9McGmGu/g16Vwo5k7+z+I/hmBXXpvdCOBdGh
dIwCT8UwDEqtTQ5u1avFnwB2CZfRlW25alXCgvZo813TrsBcLQxgl+mVqkhwGDz4eXnP9NNvksv4
k86//XYw5s9bO9p8CKGQIiQDFj/FJvKw2N6slCdVPxU2jmMFbCTKZaLyyeM7bzfZZf2QUlDHS0GN
yCGmQleQlIJ5VI7q3qtGwSZ1Zmv6xaVEc53HbzZioGk5VGdC667lnIn6jLKBRziMg6dmN6e2AA53
XXCpPTqpzauCf7XkVsMQ/Rk1zJBuk3Qn4DzD+lcOOeaslYH2wTD4H47ECweSqMoWYboZc0BRC9z3
yqm00OB7PQ/hb5ivQBTiQJblY/ugEsbrNUFErUfWuUUh3EyHzd8HxpGHLDIIAElyd093e1IRSmru
2+dzPmrcADTDln1Wir3ut5IfVG75MwGgXD8O6JiPStyA6h2A7WZzPfbSUPmCp68jiIcWomkO6rLk
cE7eI1jadD5lgIYdSYMSIeZas7L0f9BXwAbgmzPaG0hJgwnF1Cz4xMu/+rChMjU47akklNIZMAil
naJtrPXz1Nx6EWe2Jvn9vrtArRMw2963zLfrpv7arb5v5CUXG+gIoAe8SNvLwfSCxCocYEEYVu/F
AjvwCQWZL/lSn/AtCmM6BsImpLbpbTNTLgcGWuPLmTC7JP6w0ynldEkbYwkCLeXCogQwpDjuf6tn
ZGo1VhQ4/hJGD/XUhMxPZz4w1uATxKGq0GnfWm/BnVL29MndnFwGk+XevVa3Yd2NO3xcmkdMAxn0
TRwUcMkx0jRb1lFEXFNKnf/f/jo+SFPfDHP0Y9yELAY6UK1XL60LXY2BnajwJ6p4LQTNgSb+/Jam
vRlW23tQwfghSzfvWkRJ0ZelnHLOLC0ywWMpBuD+wAuaTa+s/Tq0G0AwSmM2/TW7A4rDan+yUB7+
5x8n2K4ozPx6pFtpWJokDLmqoiHyiXiNhLOfRoSVGBz5amXrOYEYMjUQmIGGifd6JCdAL6G4x2aY
TqIr9wbF1XvoZRkRBmOtQ/QPOy8+rxCWM/MURWAT5VFkE85IkyoGCvPjqmj9c8o++mC06gWHIn7Q
855BTczu+3ycR1mMQbOYAqJ17PQplaJ2RrG/h8WJxgNpdpa4t39A4//IZGZQo13ypPwkygTIhG9L
kBYpa1rDSpQqN+JwsaDDOZnLPmClzRb+NSmC6vNDe2eiVtwzvBai9tMBjk1bddL7VMSNMoxasP4z
kzJzaNju92fsk4SBiSEn8KFgw5NIoR/gzOo63kUkARIQUJEPZlvTkA18B3sduG6grjrOOXzPZz5M
6Zenh6V3QO1bwneJAHgSg2TKjRSCfBGzHftVP80PAjpK+2t9ar10xI0xF6jf3iykSZn44TtvdC3A
gyY6AgQYALOWu2t1q0i1XX49SzQfHBB+E92OzSY7S67BJOb2vs6+6pKKuIm84J0hZ/W4UZ9Cv5Cf
9xX/U5mN8veWEvWB1tb+Yr6W8n7TLTDScoFYxnBTEf2gFFK7CaAH56jKFlPDh0+JvV5WjlblBZvT
SlZhKA1O7yiZ9wWPsq5SAAw3qDRnFGGoyDDGADotGPGIjK31bGcoi9tXrYTMkd+/PwzFR5mdALDc
54Io2FcN92Nu+t5kTWrTxREdOCTMtmoI2oPnQ2/jA687Xm/6/oqjcKUT8hzZAklMJDz/r+YQ7SlI
cMGwPlFkNOpl2oFWnH23WAUIFNG2o0qXH6dVd4ftcTZiXDRZ5QBP4WihNxSnjwlCl+7LA+tAyKnm
pngBjsCbo7GPoTDh2n9rAZlJOo7JE/5k2GY27sPzTRg6xDcYQs/9TDzZoW/DgZ2axIJFmzC5uGDM
wjwkediUFVdeiPY/0aaSFyalqkCBNVIo0rUFOiAXi+bmGKlyPqbhTZKcYB1eJ/5OdFmx/CZJI5e9
b04HE68Ib8VSv/8zZFU2/yPxQqSgnsJyi1FZGjQ5AtafnTG+N9wyfA2hOIWO5kQyzQ8YKLtiY399
LVuDx/R7bxFvpyFMna/bFfnvDTQWwTUVG2zfElYAq1uTfFVDtOnMZf4mBLoAXrHJQstbB+m3NtcH
6vhW/R7eDrTYUgXSvKmgowkLxAneae02NPt2NmH51bSdF0HPv/cH9GdtZAQ+uFp5UjUSYW+J038S
YoMu+/uZ50EWeUwj6aivFVlX/r6aWGiX3AWstLh7qmKyD4LYUAVsT3Zu1jKkp2e3vnjI/gMxLHNb
gx+l+icqKa66W8JMXNjKh/UcfedoTUvoUd2JDl0aE8ald65s2Jvyz7PvBAwHsKZxodjmnK20PkkG
QnTjpPNNCC+2e1PCpQJ84igkJJzXkTcsufpsMZ+ajSh0DiXyG0BxI6pEhCXpAWhqeFnNbwlKVrqM
G28eHCM1O3B3+184dnJqrlYb9kkeLkD3a4xloXyYbO086LoqPPJv6cb2PSh9Q1tosUxMmb0W/2uQ
e/h4rKpoVp0or5tah1nCBNb5eseQ8EKHMz35R6T8AIyY3TKKcl2sY0biG1mLIyQqIlu55vkH8p8p
VudMqhMh11xEN4W5gwpoPs6GSR7wJZ1vDM87Mmr4xJD8IvQXHpxveIMRGT9rVJtM8qoOYs8hidDt
bJPzL/4UeJgs2dFntg5doUfQCcrjR8/PtmN/Bq95Cx6qt98ceW27nJ5ww/vNg1PvXJD7C015ffwY
C8DNdnk9z3yL5DzMG0yf7EDxKI8Oz6XAx4omxk1fY2kEfToa5yCddXM+NauPhNOHvfSwh2VQZdmw
5HWCAuzn8l6RimQ5NoJUepoZksDCL894SEYv3avrZagEPNQNUlPkVRrZK+5tblFW1NPThzF+QCNE
w4eCukgYhKGYjVnS0tUapkrG89IGcq1S0nhA1TDvms5JwlnxXD2osfmMjEou2ngp77F4CxFtab7Q
SIWXh16JvwJiQj858mAqEQeOu03H1nHRRP3O4XQwWPYBvL5QYEIAfXN7dz02Yyw/pLqKDEQkhZTR
LzetNPT5c2y8H7PsxDYPGAEp/E3MHRBNbGOkt5lejJsQf2txFFLkd+CzwB4JTjedQxVAz7Wm1Qe3
EGRCnjY9wD62HTwbZN2hbvjQ/1oXJHB1x6uMuA9WLcctPIF/PpZtx/Tq72NaBEoJDROzcxdyb5h7
1qFfRQQBtxa+BNe8B2BOd4MzPKANlhHCYF9moN2r647Hk2TT1P1icTkTG8pL2iz/uAlSqItedVWK
x6cb4uWov1YUqzFxFMAwoES95+CqGkS/B6HqjJzLQ4qUzMWmR8vq5mitWBb8pDnNzCFgb2iolmtd
nITqnaSCRtZxMC9CQHlqN67JWcZrl9/pomXih38dlh6/JKt7JKlOuOyTiwWlKC89lfcxdFiEHnuj
pqFsEDlhal0lbIyh12ZT42KeWrBW/wDigm8tvZVuCUFQFT/O7pyYqsM2Fed8UaD6DPHGpKT84/Hz
Wb+QIhZ25sxJiXszs9FfZ576cqoDuicoZHdtXBD3V+LCZwUKDzNErPdkAv9OvVZMX/EHKPCPZcLZ
aKUM4nND8tVNyyflbtdgnYPOu282J31JB5oFfxqEcaZBYfOXbNPk/QL7Y9sTh0g6fB0tBko6e43R
4vWYuR9ExnO84VxSLGpMGOYB7AtDpMwhQXrWysfMKb6+PQQBFkBmBRSt8crJpuXTsKN6E4mMrjIH
yXOz2bsyrUsG2sCRj8AtgWOcsTdu3tNw33fzCTR6hM+ahixokfqCyBX9TlMgt2TXfz9JQUEJwncQ
8RFUN3m6SxY2ZRWzMhq6eEY3ihVT90PnlTX+CKfwtRf5HXBo2FfYVwH+NWtyiFv0HqziQ3iz0lv0
Ep19nEOupwOEEi6iJcDo3nV4WZFqO2tWyRHKZlpvW3Rg0Oc2emYSFepgY0AVbMzjDq3eE02MbuOw
LPiqJGb5lvoEGziy2TUA8snFK7Ux0WUzYmmZKuTszvF8RCP9FtxHzODfoIDX75IMLymFpKf5vs8W
M9C7MP4Uz2z1O3lMqCCaYWjn3ptVcHSWe/4MdpEUCwHqwi6oDosErnzJTd4HjfoDTnB4yudxMq0e
4Pu9e5+GVsWxlNC9k5TD274/Sc4XLVrMhaLZfHY3zFv+a5EI0l9jIDx26gPSsn7s8zEAXmDq7o8d
xMKBQAuz5EUQiVLbLeF6onEmchqdsGhgdmXofmJs5Y6V+TzsS101g971TkpqdSjjHqghpL6eMai3
jsUO+Y6EjYKSDSYJT0HOabJN24A7ueH6b7H5sGk5JCMNQV0t5FJ1vRRxdmrdeE5fBPG1f651Ib2s
eUFJSw7E11pMGnoLgquVjRuZb9wSFfIAzwalgFP1+tZr6eoY5Fg7m9hxoZEWTWJA7veoeK0hPWM/
W+5up+pMr28dikhz4rdPFhwUAz0J/AQL5VI+mtYLiGsky1qGWFyFIpFVSaK43fAwUnuAqZDS2Rtp
yaJR8U6hJ+wqLe6FZrg2XoHCDhoBbGr68Im9tDkizGklqDwpIXK6Ytgt4dEnAJdFG+Ndlq/UlJhB
lrPvCz7CoRUsGZfRXNnPRMz9UF4OGyXTdM9L7ViVGz2UMEdZXbN/cA+FDFmYmfZzBpSk3PyZZgi6
zmuzs71GPNcUbQJMHLqcjbAZXAnZC6rwIfuFly+hEFsdUfWxAZLK/CRmQvSU4CAPYYWjNmbNaoeT
wXRH/JF9DAPmkjAwng1H8F02s5Wpveaadk9K9FOxU9qxb6gaQCqXyFneYva5MgBA0ge1DSLrPA02
d+tl8gdUg/TKVG09NI/cylMuQQmRRnIgFBEFGQNb/NMAsB5q9ZO/pjEwTaHXIZFeO5ksgeIuckhT
Jg+jOYZldmWXf762vN3H2QtOAevIuy0ENeppM4QUsG+XgB7+I2TMX4u4dwXmZQ4sou87CaUshSHc
CnAnZGyuh90cchWnT3BAz/WMQ7LgriYz5ImSU5a5GVUyk4vi5hdXZrxYeXNYaA6zEM8OHF8BeU/T
8bnBKaVjp2cBBIx8qCl9kQNNQQalP2N8g1zf937X/cbnTojVODZLGGnArjtEpm6zDRWKvFAlJ2NP
LTpGIFcmgpY0XhshAL+XkTfc96cw+7W+mTZ0p42hv7zineOzuSd/IuugBx0QkBWFGRyk9V5cT8PH
2vnKCawDrwmGh+pThY99aHSoisw+bCJX1tGh43qnlwlYSad3QaMNv1GsiQzEjksDF7pM8GifKgBf
idkUbNMK9peDmCRQEqIl04w57CfJagbFUUIlkUNQpFhPZeDwIu23i2irU6UzxEungSbgXXRD6IyS
v6KO3YoU9e6zz4WcPuCCuGlLIXUI5HAD41ZdMTZk4eE4oVlERZs1o9/h6ifBYkAxbjNfBfzobaQX
nA/xp/A4LUWaG2ergS2n2kkzXVkyqKUniO6FVHRwANuJbmfup5VO1SKL4pTmjqAayNgNkJjlR4L5
L/Qz/nJQ2zTfClpduC5Qc4njVaPz2qrbo2e70iuwlSdMFT4mFBYnAPwuwt6nei3fx0VpOWzArxn/
Ek1/csfoKbeDOKAVHF0ovlQ+x0jpMVLQ8Mvvl+lgFewfq1ow/05waEuG36Jxr7V1kZjz8W/Kbnsf
9uPTQrRoXaq4X74TCrv7184XRXlR/Ex3kKzJglUoVLokHNM6Fw0cLiq9MUNHiNJT56hS8hL6lClI
CG6dP5/5f8LXxq59YBOA2S9hFqOVGjvx0dtwvpN4iis99eq8u37NPSXefygaQfo6SOwHIjKd4SDI
1ewC3tOweqIaL8qKUpKvjOGNA/hdHQ5f7IJm0C1mgzPvjbNCNKbvOsKGARAJ3hD38FHjG0ytFPTm
2Vymtdex7JNShofdlyJr2E3LHFvTamVygvfTT5fiPWzqC3VoDsmOSNfMfh48EyPvdabcwKqsGO0o
o7gyoPaiNbR6sV4u+0Jl9tvjhBOZSdqWnNfC5ZvLbUiB5mzTgIZi5H3tZhyNhJYUlsawYK8QUe3W
wScpA5ivxmLHUNVTJltEIof87Oqta0DXtYU3vKZKB5OxNi4sGYE9bhMHqTJcE2JF/qwMG2TPhmVB
LE1Ndk+wyqzwEE2a/ai37kTGXCg5ayKJeLuIzMQvO3idb6jyyRBMBB+lWTJEuOMIW4p8NOBBdsoB
aXaMlexL7Xywbah5Bv4HTJSvnN1yAbBdoPYNIbhN/v+5b7mXxPuVyV2ypY452wyfiD0Pbq/0FPp9
iPeFLpYRATMupAruLfo6W6s2GcM1Jy6Z3b1HY4j3l4pLjcc/V2GRXJLUwt3TvO5YCeTyeD2bCNcW
5TZoj/b3oeYHMnO1604n/8QAfACVY8h5lEkGWV+tKGfbbgJd5wzQmgJRC3+DnRms5rP0vDkgWhgX
ORLQOOEjwnM5KR559MWbxlxqZLYcCelmvsCEyTwku3diydqZoa8DfvTjsncBSqbx80yaVy4y216T
ShRyeKPoQASz9psrdoSZWjDzxf0eMhkF8q82187n6rt45nSI7Uw226qa5IcfYgjJqwhi965//6bd
zp9bxQw+c0dPcZFBB1FWvO7FhfCpvX14C5uZQwH/9MddKWVaJAq0YsvNcrbTNEeuWGpDnrw68AVe
jE5k8GxHP0CGYM11gcyF5lg1fEtOH5Cz2GOW1O9tCCsT1HRjd/xCpN8xi9v/fB2Iy0FWVW+wFW9V
CEIEh2Uzv6AV77MZIDQ3N4SfNJr82AHxJuEq9B23FI6U0IQPkPVFTS7+Qujz5QnIjCdzvRDl5JTS
/qEIAzQdsSxG9183LogUkvt3HXeu1mz0Jg45m5P7oM9LZnBoDcql+na12dHbJ+M5rZ6LdP+PX3np
WSjrilZk0AHfhb50apJtKEEly+B5RrUkTPWbSVRuwlUhPmIB84uxvt5+fpd4z0wLgb6B3002t+ZA
yFfYNv6x+gHpiuoWbMQuXDB3SwWi4tQpwBxH7SDQlr53OHay+7/EtAz4ZnF55P+zvrstbc4P1stD
Hwaapqq/fhV4puPVNpTslwWuIwKYrpVvSyskQGtLvvhQrFunMrspiq2BLiN/cGL4B/GniCfAwFqj
flqbSRw5+EYbOw0YMZy4Riijvv3ulTKY7YrSpvY1gYqv5Iw0+JzZZV+Xynncks1HnAhTWS66IBmK
9/LHnKi2B0X+jD8CA/CrCqdQBm6HYq6cf/KS6hfpje9SmMIAorxMZKC92hnvSzinYsikqeVLzLFW
WeMXDZTQgYz+3VufV+zlhw96u15lNPasXRgw20WhOsFSxMZmc3yclG4DSOmLDE2jV3HdbRd0jhgu
ZCDPsdPLiFC8Yg930ePZ02kEgx8FHvovQgIJZOBJUl01CVFn1WaXwEfYH/gkxLekpQS2JvvwBHpq
yHbdyMZLa024RORAStzKYISqhYFyuWPIDV0Gt4aZN7QitUZYTynadKs+OHQfMdvFO6/aQeFoy8+2
Eyj8dp7VdxCvf/ifDfu/vmmjmC9uscvAYF7lwjynx+z8Hbjd3LNNUI+0mqvX/kqpPAlRhWcCIXjb
duigMZfRHtUsvE/KLren0DEmTlTQYwzuwQQomyhICO1twIRzIxjm12lTO0h/x3hckCcTh65NoyKK
PaGenwss70gHNIXDtmUbV7KUU9kS9ML8EhIbtzN7QYXIuGpOgElA2670I/PL4dgGzYZeYKS3KGqf
W1NzKdoOF9uD3iPmsvWi5O9fDGW1YSoIX/NhDR8M+1Og6380NZKcBDhX8RFy/DsULoRIujBek29e
Cm4jCT3mq0rMasxKP9+6i9BKrR9vufY34wwwSglbZq3HHb24DyGzD/JF5vxSmIvXja3MRTJycyeq
XQgJ4q7cIayBMlQhqOP2XsLosCfdby5b6fZ3dpBp/cFVfKU2589DJ5nL0hS/ngEE7qv4b26rLkWs
IVD1IT3dT9Sq5ssj7Y3jTscg+ZhcNPdXiRFnS9KrisTi1s+yC5yB+Je7niA9xf+ZRCoZbBdReBZj
xYGpkuQYa1lJWaYZgFMDrYR44TCl3raVnC5mKRjWqRlCRG+CDuHXP2IhPQB+A4Yk1qI4/5lXXYNy
aHcnlLRI0UZ0GFg/EVDQiS2tZjMj4uQlf+Y8G8U0J3NhlxsjypLoQAYWDs+KPaV7Njx1D0RsNJqE
MsOrqOqTg6xE9IOlHWqrt8hlDszimRFtDdzaAKehYeJWE3xDGk0IIQthCgnfSdHXYbG5hZ4K5HrU
YvLU/qNHx2bMnZcYYyqCT59mvzCmBKSWHJNEDfuvbcHyAYr1oEFnfT4RNDdeLIZ9e7KguYOZJJg7
Lgt079UR68eHuskKtFsjGWdGgz7aVHk9LPxp23YOfoDOru7z0loa/PwMfqi5L7SzQn4ZVcK3Ptcl
XLut2vHpCk3iUkKgsrCbJFwq0yOMref1i3TQOJli5qjnoQgGVhH1gYeht6EArBu/IYp+PkH+wBAq
uAQ3KAlOH8pMCxyQGmfpOATLcGzYNbOZVng4vIZesB9gaUBFhkJP9ENuo0NUF6Zu109UMaGaMc5t
qcDE+G1/LH7xylDAkABaHztpw8nAscA6N/wsWLfwkloOksTW7e7vQVRymlPZwkJ2AqmaYHAvXhpf
xZHMjL60bQiOPfUB+HGHu6wixamumB5JaH7vSKsqSaA49jNhDeSwppx7l/UuUcHTKQJA1URAeFf+
x3gXk4GfHAV+PDrjz96OEhHHtRud4ZbhW/UJqpxFfqcTIANOKToUdV1mESHPOs5/77tYW1Iu7dUw
brm5gXv4fFLZCqvLoxjOGTmHCtnqcaHZt7JYVQGO0Za0m57G56jxf9xp6A2kPZYaSTd0FFss9r3B
+yfj7e56dhmiUW7OV2rZN0YG+t22fAn9aaaDRCm5P3V/BmyFB1QwHL8pVgNAXvNpV4RE3kX2uaYZ
PPFSDqV0mRJaMTEa0oqjtaJGqrKi7wzisVJUcXSSgmbuIywPN9aaSNQGrh/vYhskFfIeedUqjp2L
mRw2gqA9ePUf6VhkYqMF5yMBNLgsrYi585AzgmbodeTmYRlRDHTVnz4Kym7OnZZ4+74EYmixz3Zu
TDQjIUbup6DfFCRgQlqHI/LxK7s0FJxY+zyYS4FTld+A72NK9Ju+ZJG/XB6G4V0IqbPHSP5mgHMw
1r6vnCO7w/FMej/NhKlejRztW9TGWpJ9CoH2nNMqrOZoju0PjoBfNjLgesEEIMjM7oj7u/J79xgK
utd7f1FKY5jH7VUoDHLDNeG1M4nbXvgdOmcNKgX31pOyLs2UeT9ginvjZqai5n8IbMyGuSJZ8y2W
JmEomDPCu8+5qLwc9Ahh8jI1cnZegt+O/CgPYC6r2nEJAENBT+rUbxDvh+X1pIxjXWb1sLuDuWIN
Sw7gYW7CZkO35aPdES9LC2sQpjhKvR9QXJdXZn9tgzlmN2Pg5PAzimOAeJnZa+gr4wunkF0UyFE5
ILxiT4kUEhXYIO7RHtsC6spI/pef70Ybs/96RDWooIpd9M5h3ZKb+dmp24Or3JIJZzvX4sUu4hbJ
xMM3UtWjjJvslmDhBm/gnvkzNjuPN+X6Hqr7YSn4pUCfTfA+9voD1F3+L171e0+Ikd0darnwrgxM
SXpeVmufdxEMyr2PlqBctYnO5KBTrzCMx/tgH6c7k/x1uMa6GS2PJluFUtrLDPZPN11fQKiV3iJ9
pFlQVi9iqT5HppeYJMx6qPhr4dxlZF2oav6GUT0GxVhmjU4z0NpLjEVGTNf2thRoJsP7ErNjLPe8
44gk47Fy4D3xeqnOEBGuzLxYVgagTiWcv25VxC4wkVwQUQohkhwBapzxbCoaxzMcwTMi6xWm3tLy
CV97dsCglynjcOUg5tDHYgFb/BNNO9jKVc63+mLGeekuASIXiIjUfQCITbhFsKzHH+Jjvgz12BgT
aGyOD7byZuXCBfmXuKN+9By77KSP69bpykF4QetsrR6DShjMpdBuuHRXriPZGJb3EY+eKz4FtDkg
6pPV5uptkgcaBpNTG3yQKeKRcVxj3YfmtX0a276dZTe2wURiFxVPdRlJUk50xmVHemJqu7OGIc/A
BcWEcslLjSOQgadkcd6J8fcBbzAcFuds94RyVs6EeRyKjS77OGDemtHQdRNpAaEBFxH/qQTRPUco
/6qlOkKWWZP+HeJfGm+/EsGDlo57QhwdU4z3+dGLggG7GFD5YEulU8egzLabEB/IVg78Qi9mv393
Sk3UBogapYyjHHLsLBC+DS5qcm0oILsN16xWISlGOvGmX+kCHnaqAm1I2wMEnsFF0D0W0wjTRXrc
568ZSiN3ngkzD1BSxi+iHCVYgKuvbV4JeqE03Ow0fHAeHLX1rylhO+5RFVffWEbOdU2a/ErX9pqt
/JxoAt+hHu9JhB+oNiNOC5OccyrL43k7NRqnlj36lfGARi5mj7jxarpARwUPTJE9HmjkR++0HDHw
4i3q3FnGRrRW51nxKNj8iEdah7ui6SZ8Is13mgMXAr3CtRS7NjaJYEqIc+8LaLa/AoxygP6KYsfD
La3Zb0e6NKLlFwQ82jYDO9vTzn8VJieocwRIntqS04PV9G0VBD+b+SzpXcMvhWGtJUAmbtaciird
qyLiTokT+Wr/YnwG6ocIV43uB7hgk/9NY6cLUlE4ewZvwnHPvkye90+GVE/bcvYB3xjRvxKnt7yg
+TyZ9BqbRHwtqhk9cLj/EuZRUlNMSF1FWOkEc/ZbMZO2PCXUJyp9wnjvjQyW+ccusYiFzhNP7pMx
l7AIsr/Zbe9M3y+n+ryuBP48csE3as8T+zybZNQZDcFfwCFekFLHci7tsDlzwKflUwxBlMzwQnbv
+DN+pLYCnQ5heYP3Yg1H3X1QF59nZUC3Rw3S6eYo+7hytBmXfBkRgUuoIvPXDD7tsHiDJNp+aCQn
1qiu71CGvb0IZ5o3p3hWN88vgr385S8G/AlTATaovlx27DU/LhRpQ/QRs3/xjIoJqeXwmoSuIPCb
RghrK796xdFnJFsLLLsdFih1fUGf+o43oiWk9ilorGlJzNHHYPwW2WPxP0B30GgkLdquZnRnllT1
RIIN/XttW9SXdPFcYpGsjUQRKTSOG7JLfJTxeYruA1V2YWFDmmCPjJeqjsZShYWtZ4IoRh+PQydd
M2+COag7BF8zAwDl2aXOhjbsmYkH0pZbhLupKWniug5hwQaER0pSfRrYgeuxPDMn4tiTwjEymUkd
Nx3eJS9o0K8qBVIZqqvIlgS5LZAGAl9RbjAtU/rPOMs8ne2x/onfrdvvCebzHod1nAcnNsf94tJv
SlYU7Lu0OeDqV4U8A4vlE8gcytsFQbHAcM/fA/d4IvbQoC2Slu58o8aRcQk8tcgI52cK5YJocpnC
fzSn+MyCs1QbiWFIqXUkpitBh/T4DwD3RKbXeXzY3wqrUlLBhWhvap4/lt9N3rQUN+fzS6mFlJI+
/t/VhyWU2/oXWHc65MT09dzUYvkY3CMa3X9dq+AE2dJ/1LYNWsOS6YJIMBBRcI2nqnVGcf4PpC4x
dJcdAQjo0LzMkXzatBScM1PH7kliCxOlHjExk7xvKRHPweS0/3P6tJvp2kECYYO0qI8hyw6VwJaW
W6R5Eg4cpmA+SXSnvhDDn/emHqlWk/QXIu766z8KAPlGd8o8CefR70wNsBe0+84rM22SRhvnNHJK
hvrqWeptBlogXv/dAXtpOEWEBFMzNDhOs5Wlb00I0xpDA3BoTFH29X3X9Dylw8bPIXlk0wuNeOV8
ZFJOxGuKty07hQlbW1Ai72f92UOWp2eZfs2h8MD8kqdx4l5NfNEc728AUXVaLYwjBqNZxYQpvim3
UFi4yisHKQtqlY7Z4W3p4P1PBalaDo5cFnnCRtC4cZ2TV96434OU9mDFmiYLlXHxqLEqKFB9c0ku
eHIrt0bZJARfwEsPnDXrU/x2w5Ah5BVLV8/sWn1ucwb3C6hWPrVJTONpi9CStorNQwML3/bIJrLp
TgIRO8uEABuJqPAha2QefVr4lDyEBC/Zbas79ydf1JqoI+wBgNmIY0LqPq9kP7eSfhOY9NjYb636
Hsoc3qt4+mVoCM4rbjREB3WUEHR7DFTbnmi/oKeEschPjj4eUChYz/bsP7VXEO8Wnza0tbmIxwlW
62SdmKwrbu52juUpQxf8mC876Z/isVaT30yXcyk5Q2wQXrU+3+BRRqRiainlBixbo/I/mxJhLGV6
bIFsApfdji9FbvSff+xAwOkSDLf/dTdrtAw3TMT4lg2o0YSEKapxJ8PNsHxGULd1hydvIsIdG97N
oGLyJp5PzAzBpyzl7i28w75QMQrQhmQNBsP1cttMS5nIt8I5xgAPXGwWNO72qlxs58Zo9t2mtyDw
jJAtih1wwlmIFZsgIMu5dM4v8pX7UTTyUsPRUNqYQ7I9drm4VhkM6oaddWGVS2nulP1v1IMxsAwM
NS05+envH/lIo88ph5+4qLBWYjuNS191yw4QrRf4krzJM7NZiAG66W1lXKHLpWK0IphUeujjBHfA
lCKJR4dbqHasDxEMxmEq78mnlgJzBzwtkHDlTCwp1XOXtiBnesUxXgR225blxv3E8/2sLYiWba7Q
nmIKv/N0V9t5kiuyc2GGydSCW8kQQRDu9pSgQznJJ6LVuJtnkW6Q19tjMJ4/MGvNe+Ie2k76pwXb
dQd7CFZDfFGqFB326ETk7x8q1r4LxUDo0luwrfHdZd+mF7/Qp4M56wwq6NvJ4iqzWPKF4qij0NCf
AzsxkUVIS8YfFefj4eSMReT/XatsWLZJqLqdnzD4ugY0b+vB3q2fMw++xOSoqm6A8Rl5WA2qTCOG
21RYuhGpjlb/9H1hCzWUWr6/QEl/jyDacwO8gbSKlG6gWtbFc3d7NomWpwxjgRgpwTQRJGCXCpDB
FVI1N9X2h/0MqPWZQ9qTUL8AT302EHRUfcqKmcbobO5Kc3oTMh0TYPXz94t0FxWZIFniDaaibWQQ
iiivp3d5eh34IEJUEQ+8CwteW2cTRxQy33CkSWJ+1H0ilkViX4p59sGg1usb2X1B1zJ21GyShfOU
RxOnUp5of8bfPrRmUaD33IaynmEh7+MK1uv1W+H/4gZiJvhVhEC05V+KUp7ZuXHoU1h8cS8Zg/M2
4pkAB8s2nx4XclO3u7kloOyxngvGcA/+0nXkVUoNDIEkh19xNOAIReizECfQZbe0eynE6Xl7O3rw
U+MtqVb9h+W6z2kW9AsLv0vvi8Sf2T09HXmswkgr9HF9q/kXxJcHIzYFygf2yBXrjTmscQPnVVtm
89TLLlepA57wncBeaJ/O1DHI4Wv8H3xW/7tk3FdvhexIQsQFyLCJNPI5kDYVT6wQxhCiJebQ7MOP
N0QcFGteXO0C/w0hWxhowRdJpEkwmJ6+g/8fFND9/DX5hw/Ei3TKrvq1QiM+/SuMLk0XXEjkuUzZ
NI1wv9Doe8zyB2z3ez10nuyPSwG5szeFBG9nWm1jJmTmeOgAa3Bl9Xq5BosZsouT9mHfToIRhj83
JUD24vsQuSnrcRYO79tYsG7MEzuMWK3KkU+WN/YTKueqJAVtuyS1wWTa/m1i1eMO97f/3H4qgGyf
SV8/m5N60ry0fmD6jJ3SvwE7Slkn6IrRNckHUnZAYTuN/kgcHwppIi/puKfL1xt89EwRd+wuuix3
cfnbpPHeTOGZdsWHhxpDGLmSlSxCSLldIfTvpPUhUb/NAZ1H+oK/DQBWyadECMyVYVutXScAoUYp
LKFgDnHRB05L74AHztXdd3yDqpoN6+r7LlvHlj3FdmXgr7+JgwzRBF6o7oVmi04VPZK7XPpuhhpj
AtS9+zSCliIDZIDJT0o7iwIs6R+iu9QJLDgfQF2Sg2WZsWf+LuqaFQ0tsAuzgrjuxUTgu0PR74qN
3n1qFLzSFQ3zfy3ya/IWZvgUTtPVffqSDdhqlJ3TphdRj69j2Wb4okhELLg05Rr2PIviZbzva9XV
3sEcjaTNqvYagmLpYF7wZ9maP/MvkAvBk0sPNj1y67DlcYI1DlIqoyYl9m3S4ecUM/FAMpla2+mj
nknNvCrv+L1budSqwPgbWVuRcFBF9GRF3+9ScVnGXD9QmjFzI1k5gu0SWWR+jj2w0gfG/XoG/Uy0
ojZPIXFxpfuLz5xQ+POSW2hDqi35B0kO5i5JW4Y9xMRX4HQolBaYPq+cHPcb6vcOr5IWVF6HPV0V
LGkxOW4fHxQoO57UUHPKGaeY8mWzrBALCtU/KJt4q3yJzXnrHe5kLBV3AfD38cP6N4d3prCIuQV8
AQUA5/TuknI1fRmnmSzNXPUPY6HMwW8pI10Hfvp5KJjrO7HuXXWuraJ1ewMECHfG9+V5L/sRTogI
hPYHGovXubMpaSYQVKEoMXVQBc8XMHWllQlpRn/NlCctasnsZ62y7Pd9I9T935sNXGp7wqhKSgsm
CZrKq3KAaRuOeqDOYPrlUJXJMNaysLJusZyi+5KC9kBezZxI934FEhwLg0tHYAgJieNPWVtYBVCD
qwlWtTVnadpPA/0cQgBzDrcxd7wyXREbcV7hqNNc4jp5Gqx7Y7Q5RgIK1aDIRM9wtn1vixVoqNiG
MHVq87+NugGZnnkXoTr4Is33rHza6JC69zwwbFnbXAX8IzqqFRy6XXutpCIAeDqeCwQC9uQeL/xM
i7I4nL2hpAZzp+PynZ7vUJRbjLLOBDaDFakXHj2Sc0zzoGZz92fIXrAsqbQrOmW58Mu31CehJEs0
LKBTH9CHMdVGZzuZcvBCyTnl+19uEf74qKjOuDofoDsQjoYA4GU83rfvjsRQrh0t/fRyST9XIa6U
hoxdy9Ph06RZVUaAhBc8wRhzmz2oxpWO967ErzAXQcJWFRKLkmr1LrD/o2zoNRc306njudC4aujb
t3s6qqEzjbc2aEGc/pWfbAE1K6RhWiTa6qVQCPASuSB5VlTp1zKaiEoBjrG+SdCZYs3b/Uw2lTnH
UBcaQevy/BMO9AeH8b/KlyxEguvBTG2ENGlqWd2NW0ZWWGKKF0CpMbe2C4+3VJcmK42ebCUXVHhF
5V0Mdv0FV2xiMoVZz9078iHZU67LJyCUXTBTLtKVELL6whX+JKitj6Qk7/M/4kFnP3buPRvSrH8r
hucMpl9XsJ/uaCSKSPipaHG0lvInt9FE6c5GrCLPWlEe5WRvvwRXNUzSypX7S5qHA9Bdt3ACcZtP
LCpDL7Lcw12LJlSvIEt7Y+mL+dxZS1I+OlzToe9MoJ1mZb/3j6zKL3raRAQ4vjjrltW74BDm+x7U
gMqolwq1Zj6/9VL9Pr60Pe21MroxhNPBof584EE7G5GaNgFszZbgyiaHSWgbBCVnfjFYH/8V0VSK
mHKpZD5i7hVWWvOk0qiXZWNhFXXuLAv3LZblToYQeoURigBBNvD0ZIFKO7O0v6ozUHcqWF0S2/Ne
nmGOXTjIQTSULFa2hhlMuZjqwpNbOOw+QUP99ox9kbHoPXhwRroMzAPptimMH/BC0dopTDWXSbrM
6UL2LY9TRGhh11jqqE7GO3Msa5ntHacUG/9inFiqNhUnIrZLC+Xjm0CuWqIAdOeC5A1UCVwo/zv7
4aLHJSc/FQyvfn72XXt1jhy/sHMhuj7ATUtACwLujcYz8QKVGraPobmnUzTHx6HS5pNzlCkOtWq4
vrv3caydfxuhnAcc30wsGymlAHgtLeBdcnCXTTniJy+Fys3+e80vofU8QY0cYuLT4XgWovutI0fB
fWVHM4raVLyUxxdAf9Rl+HQF5Z73o1RXm+7cPDKtNOKCgMAGnh4cIH31RZFB7kr9mawN0LMUUtgF
IkV4s0/R46bOiBB7NBXny6p0CIYLhfbec7C1VCg+vKtY+mh+VPh/YnsMqU7nghbYDZ4D/LXKhLUn
47a/CVjWO1hP3kJuaSNZwi2xGNqIeKhmKd1VjH8fDw5LyA2aKCjsflcDMMVMmxoMuw6p+PkY2Fg5
KF8yGWUEZLbNCQFY5XnuLBlwxluIppkBTdTGCoxjmUXbKrqW0YbGmDrO7ToZ9mMH8+96+9xKXHp7
LZIJVnEI2S5ZOjkwoHES9jtOcx0yTznoJHp+0jOwzGFD11QmadUce/qEJAbqh1ekatGwnYo6OtIA
Ce1i02xPH6jL7G/KOKwEH0mCEfzXxt7deBJrdNUHW4yXDGW7b05udM1xVY998eALTpLWgZncWF9+
zDLABIIxDX7y5ZLJge6w52s/lftsmphETE2theWBaAO9XTG/3UKz2aJYXYae4pKXORjD6LZEAF54
cXzlClxA3nLN+m/z74mxWNtfI5sITWSkxj7D+vj2N2cA5YwPwor5DQHRGELJoTyzTmNmJHGSYa5h
7zihvRIzVSH6J2ai6OzRdUP5+zt2VUGQqY6h6ihABUEC/v4wX+mRga+xLyqD2IGFvu0HcXhlAoxA
CMZwJl+0LvxeVzeSNh38fKRhE+6LyLg+kZdn6We2pkBpv63oOAo10PJn6J9XUyNKb+24VJr3fzyV
gSV/cncOaOf2op9SwIGJCO8KBVNykPdzArzOgFRIju5cBJT4J3D28R6NQJ/fUK4w5UwHUDkZPw1C
j6DlolaEtMEQCER5ck8mYgVpWPehBTJyVuBnK0/zd6+x5xcmlzpAJaYgunJD+Km3WeX2K/LmHV+2
sVr9P68hPU+BcVPrl5sRKet3Fc3Jk4G/2uZDXj74hK64a8JplvGOu7U0PaPJgdDwDdsEPnWw8sfr
zFyQTpvaDlqccGXM9C7HaJvgNoi+GMTmM36YJWXI51Vy0AD6hXD5SgbkWVlo56CkNgwFFoptjcTT
uocdupG7Km+DfBR/Lcfy657uRiDgd+C4oJMpKSVQfIc51LLGxSR5L/VXk4O0fjUmKDvKA7MMRBwo
0DLsjhAy15tgqXLP7tsJh1DaI0mOb5lSqvBZwFqcqfBGA93WI6VPMo2O8zKLZNjnFZdY97bzlZa0
D3QZUWtmsYXu0S+r2EnnKGc6WBmQzli2mp2l+fztJBu63f2cRlqTpvPtE58resCSTaVVeAT5OL6G
ffegGq7y1VEc4wQeFXm0XL5aG2+w15Py+rQW/0mdaR8PK2YuIncBAungnpxMOlVq6VBIcM6nRVrd
CsMubFC5LeRizHS64Yc5nPue4Wm9jw3wcfaByuNrj2m60CD5ZCCB+XlC60EMp7htnFEmhQh7KQjL
w1hrfCqzNJ5LgGlnFm5xOv78ZWdX4yp2B7ytg93ohbNide/LzsIuN23zfMmwS++1v1Nv4YG/jEw8
JgjEGgQKfNLP+O+Asc2BUwlpmVKs97PW6JPlzyxvr8RXVGgZZ+SpWyqKlB1iG/ccHzOCqzYXugpN
h4tYN23sNrq+npNxR/U4hbvW7yqsldv8MG3QunJ/H+IY8oXwnH0fEuj//M1ALBYJ/QmMcx9+/itN
xWyt1Ptw/n828v9JmgusYB24ptyiwCGVdV7fE8COeZZqiNuRhPW5bhrUPra8EEWUxO7ye3HgQ1GO
Gj3Py3swcGyYBfLGVJzc9UDHkIpIDZ66ko3buIKgyYPdjURFJIR9FHcrfD04njafi7/jE5/TRhg2
QMkhCdw4uke97f2+Ui90v7oG2d7po8dODbFtCZ6jfnS8cC9U4H+rUaLROIuGraUNu3mSI28Es3+z
vPtUnSpc6LimLtT+uO/e0SQRdoog18bU2s4CRCfrxMDyPtBzVOiG74zRjFM1ELwlfaOtBiIWj1xq
AYd1HJgwV4pARtdSFitTR/8zSs5RNF8pOjBP13tqZuRc/+DywN0ibb2U14wD81LOQPOgOtuv4M5V
bmnUTfq+DyV1NMVnBzrwII7E5CuajBg/fTbuOjR4QHGn0O5hg1bu3lZfonxW0SBH4KzOj05f71n9
RgdY2ERp6IXeoMbrFkHYkBL7yRMUHs33cTdtS/R1e8oXdgKsOuxWu3FqSZv3d5sEkdCSsESVSGAL
yMrU89YyZyj0j96lBuNFbnJbvAvkrjB5Rqf9fhExbUJL2pFBatfBD6N+AfN0jgFQEtEkU5hBcaez
yPv602t5YJCNSwE+Zy4ZNRSh9s77cDvDQ+lfqfXCk7iztbNaJ1I1c+p3WWb+V0FlhjCvVBVEifHA
vM5r6hXJCE4eBiACU6mW9i/OyKkGXeONAAwRCljDi7B+G/ayAndU2rru8j6s4uT/A85cGpA1J+J3
JRUFsrdTmgIr4uCKIM73mP4NuDSUrgyx97MphcqCsWc1sERjqKY1uC1r77/HESv8TEbXKqzzW5V1
zNs6d/RnSVK0rUaR0gDL/EMjNoGKf94+I8aqjt7sOM5Y+BVRz3bgODWmQBKcp3ngMf4xF7T3bQVD
nRQHMy4XAL0pLgwxY/lGqc3u47aGEYjvztyTJft7HxMebB+0M5Di+aj9ggxCKWu7+Hmu564QOjx3
iOTv18Gyvg5v/lJkVM/oi+0cxDsCRAMEVufPUmXxpbOL6yWRPji25IwVmCeKAMRZ5+EzniB3DJwH
uQghS1KFfNfBu6d0TNtL4g1u7OsWv+sLBR7SQdpBELTu9oeFB0zgiYVvFV1cp5XrKVggF2zA5n25
Z4HYYKLVRlzKv6n3mI1MVoPFH2zK+lCSW8Bu6VW7j7UaQoY2B+j5JI6UeN4BD4N9B7OvdxA6XEuM
HHUvw6ZEaJ7c9mBT07R9yyvvstFxVWe370vaww3YcrgxfxcrpNXvUuHRQfrMuBauYouKcEXgQ0D/
pFf0Y0KgUTg8+C8BjFOxakX/0lplAGzKtKiQK3HPqw/Jar6C/PU+y8Eu73UMEGlw6+E+Bw9gCEXM
Rz2NcbIR8yNQJlWYiuTZ60YtG/JRcl8pdoiTuOj1tUHdNry6PTOEKu4n9/YmQ4vaKH1qqnATSMpd
Pkuakq2ytYZ4SCnooe/goOWUqEipbYgYI3BMPgM9wS8GwfPWXlp43e+6Zol0rGi+GuNG8AY2S0t4
QdBS53DBUCEnPRUcX+1MoCp3wlH7mPM72eOqXbtfLPmt16W/YxWz1qP41K7uRFGyz7G5ywNtO/Kr
F4i5a3kMdRD1ySio3OBraUIrsBIzl5AHo675wmZOVlI5vJRVkF4zxWDUglFPPou2rFxJyLIP1arf
zHpYcyqRIAK+O8OdPjTpjRcTZvrMNY4VymtSfeb76IfROA1rsAtwbklLkWZMFDoF3wLeRb6xgBl8
NCAlAiNedEkL08NqFgOQdSest+3BVNWNfBmYMbklwuSfxdln9ZGpwcRtnGWv3c2i/sdKIH6DHcVo
PY9Q5dnrdkW/ZIEB3qe/LStjWSc/iJFP2boAY7DA86LbaaOvdaugMq4eS47kLwk9OTTIZVD7Nnsg
aSRSPvUVGMOjhVoMeGOms6/X0zKQncXpxhBLEjt9+VCDIsoSoVaZvt3HhMU7mhPn5lASrJOgKX2M
9LNmwvyfd/eKI9bV44I9FXLn/n3h/t8lf8sby+cYtEigferoNJXeVNktu3rytsWezNaItMqOZJpQ
pnkt1RvMME4EXEBsMJlH/2iP8yUMW4aKt4+i5Cy82PD6q0Aaca9gmk3LU3esBONWtVV67oAVbANP
1HCnfwzAQ5eOvwUdQye1TqaGc+0PChJ6LQbmKLs7UmUlzd0LXmHZSHUarNiFnw4spgIGZPcY/vTB
/QQEUuNSFAfrzbrPO0kdIV68jsbgh+ZJUo2YvZZgXDDN5ymVL5M7lDAdacAp8BRIGb3S65q3wY+2
6A3G6kF/3hHfLZkoL1tL4VSScAKdyvzmhj0HW+oEhr5d5sFMIJQQ6sEu47vR6R4iYVeggbcsjrMq
is6qaJUh43eixFKS5pp2JCfOBU3rkBMSlZD0i0qenKEYdgyt1ST8qW+wwxRhrW82szkOfGQc7crD
vj0LnnmuGGzMIe98c6oir8VHiyqRkCIbWSxI35PXlcLGgP/VXmHXxZt2IaoyagW3U9vQHnWDZ1sK
Oi3MAGHpCa1PmO+8DHY3aNcjVNDle1VKNAGFakz/XMk2Bnm8Y+0yV24GFaGPs/TZXSqV64Yhy4xO
WVS71aQIZ8vMYBbJD9z2TVdmZx1WUNTEGsmvMmIRJoGvOMvK5/9fRJJFHIhfEQ44blGoiIOA4axh
GRijj/1sXEyn5IXzjnDrVJaoBjmPqjRv0SQPKeT6rzJJLh9ryqgMq+2JArcn3T42WH0KjhoT+3+j
DnhkLf4CkOIz6qPk4lTpX+28fmuaKzMIklyMvfWLHQPSYEuJb1xpF3o0ACBjAk5bwZw4ZMmVEV0k
2ZBrjne+sjbb4xG3+F6qgmJQIwGHpMyW9oHdlklFr86hFnGSWkld5eTzygwugkXjRSbJlUUKi5fd
47+heBKQYZxUog83rWa24ZsWC6JSGQX9j+0iY+BtFaNlthUP1O+jNrH8VhfX53OLIcK8aKuwLoX4
XFwYFsHDPQQbsOVVNytpM2q4pDEXZf2udfpRivyAKXqK8/NHeM4FsXaRAWrF4sqwYBL3ZTK6QKZi
ueD3CZaq5KWngZDA3aoge5/5fuP4DecReRQgod4v9LNQr+4X/Lpz31p/cFlydHTEIsRJqJWcDrDY
VJrK4P1eoE6RqMgF+QlOj+Fj/tx6JcoKkgxg8O5LOlHMGsIjuWfeIgRZ5C4MzA4SmcfYiDiAlYMy
sr/OHv4F3qdJXEeI6IZWKJHmLOKDqJeHdYjujaO6uucO7mhgXfTcZfrIWz/hkSpohzAH6qthhEdl
dZHMiiFRTOZTyroKUSGLMnVDmCd+mKMLHrl186LcQMtqWUWY3+AZ2932XE4+ErzymHrcZCMoSzP6
XVG0EFQNQUkvblXB/LXT40nlcJQcAfg0Pqnfnta+/V89N3VslD52bKclYlj4ancXpdfE+mFa9EKK
HW7AJmPTeERuH9ZBk4SeGvxsUQYd/iWYZxsccg6bhHYexLtL2ZX8GLF66jmxOGebuUpiWTGDWWqQ
OZCJS9rpcg0/8B+v49XP9VE2m1NoKb8koX98ft8mK7KXdW6SyNX8WBvnNHnyizMg7UtBxIAe5NEC
X+lBnv9O0DdhZFFHip6sDM/EXQXuvvSsiTy6SGtdnioMSPdWUeoKLSXBA2zANqZRdieY7yqpurns
gzdSAD9DewvAB0e8VusshRmkXR0rjttsxr9deAxFyTDtCEztCYxsu09VycS59Ps1AeAwmb57BeHM
kOTOoZg5CaSGAfdxghpj9EpitlCtzQt1/xMn7zNKn2oacidx1tYEu2p2v6xbo1L4cmTjHHZ5+i+8
mm7C/xk4EChRdJPxmKNcviULB+Ti3qfHpT/U+muYfY0aLYu8xd96nBg7nQIE3d8W7HVtqZNVB0ZZ
q/pcX4PJiuAxp0YqlLiNWEaCdij5tHiM9MUwdyWeBnXUgorTohFuY42SjDC2pd0lBJRpeKaSGVF0
fIA1e5qjgRwGks8M/aNf4Co5dfaQin5h0+CnH5Jr/eth1VhKNrTrtg662vkaXYYBhpnnXUQU9mAB
ZtczQ7WYhTOPTwANBzLtBDq5gOLYPDJQvqiJ4vdrxD2dSY+XOeuZDWj4fe7JvCrU36swJCirQo4x
yjJwEoI2G0kC9/R6CgkEgtNYj9dB8bx9Vef3eIkkNwfoyYjH1oBWB5eb4SOe4K3UHGG6C2h4/okU
+s5ijZusoZgT9XV1IhVM5ms10WBOnmuVrUwFv0xzDYoB7o1UTKtdTq2vQSurz3izSQ9YWBIZlAiw
JWqVbn2tMdXKSdEEOcWqB3XWXL2TKdDRYiuKgMKbUyuGqQyu2Rsm94vHHPWnSyBBL4oORct1yBWM
P8DduLRTtLCyOJ1/MUqATcFBL/7avVotOBop9jVQ3jRUFyNXgFeOqPotzq7BkWiKm6zxK+I/uuSZ
1o2q4owSN+2JbfWZWwlTbCxC+Gvxgejy5PeOY0L/pfTabWDPpKCK7w0itvRxjM/1jK/K5Lauf59t
4HYn6rJl2kx9E+QfwcYELipoyKyHiswouTt3Fp4yQnz3FnINF7m1E4LZmxi3CwdNFtcyMCbLosl9
snsJVnaNu8fWt8EIxkgdp9g58A1OG2GiOIpPEWqfDRxXU9/KRB+7EHW+oNB5o3aa63hl/sxGPDs/
kCvgyaXDO1rSl++9AJ8l6JzyQZ+h/G8MhzWuF2YTjymXqiGuDNFRD+/raNXhQt72kqCWb36c9oTW
e8BT1V9Yhya2tKWGfZUOPg9/BjLE95JSWjQfeKksIgKFYnG+Ka+5KYMmUkVKs/Rxf8/aIkkihUhw
ks1XqC6mUU//0ee8cC0e1csGWAW+hHN7cN2Hr/l2jGPymfQ9gHlWB1Jtpfd6OCCwZa85fYjpdIGQ
gHW39sBBSxYYB3GB3YlCtv8AeBSzl5+xcrOVoSoaxuGPA7MbnqHpG2rXqIh0ER3k7TS4DulsEH7o
e9LAApnve59GHaZdlMUYpv3BHPSagh8364faWw2SGw2YI9b7tEBv0uzqfA6z4aH0Hj1e5jMpPcIh
61uLvwCatoOmyDYPzUfHPhpQFEXoire8vyWwVM1l7J9D5z2fXAtVYw1yi/JDIlSn1BKB+Yy8TiCM
9DmweI92kBGRAg5GAMUPKZon/MG1ZvsrYkW8hPJ0XVFmLFTH1gD3aNYm8GgYW6+tvBG0USJkka0o
JOfxQ9zaOB3gZxc1CGUAgaVwTSDsS1QRRrC4uaXJbZzh2ScSMPdEYUw40CQ7/Sosbd4upWSci855
xrJ/MCBSzgQSbfbW9f1a5vT7NqV8heIZTTl0wtC9ogpz50ZnN0hCNWSxYg8UB/mpqigmOTV580tA
O2mzHQVwmaSZrbbPtbmkOtTaXIJd1ZveH36/CZKNRXLnH6WCEhLtDikdF0Yep75xgZ62rgN32QQZ
OdSUvTatKYvePwANU03xUs2j3vSxYp3kosfoeWf27iUqqUjwS2jI+PoUNfWOjbtJoYu5PCZpDo59
yQxN79tjNGhIqTvm0be1r28IRmFU2R+xDCIXZt2EAW12kW0GmkijzuQBuzF44VE6O70pri7cRZ9U
FTZxPn7MNRRGrTXgyJUuCyjtIsBVUU2fHPV5di3c/Ffxn03k3TcmCDZ1FGn7gOdDrbjLntuHtRH2
pB3gucu5QAyMoZaWWpOx0yJu1aSRb1vfqQVHf64tOTuy9T01rYgcAtWwdFCUMXJugMhMtU7RL6wn
IEf1/xP3BUkQobgp60O0tBuFDuhzU69VPNj09JLYM8P6ZkKZDmvMHiAz4IwKZ5y3mXMew+8QP8p0
oegmOKRrlWliBMb3VwnSyE+I2covEv27j1ENWQzMhA6hthpk8k3uq1KN2v9/zb5dyp49WJdV4mz2
sJZeU0Dri/WtwZtdSlU9/6g612w6ncFQ+V1YM8ge7Gg6E/58jYS1eacfeEZ3gwNal02+S36gmTrX
EaQUdcmcqNM4cSWLG7dCJliMIxMUkxqJgovgn0MnRKWdWVrb5/E3j8KdURLjA1uvHOODfz3cdaI+
HwAtZO9E1m5mdCv/GgTTOjZg904zaevsxCyXDgdquc0YPM5xWIWrYB7cGnzVdN3iw2K/D4izyAv4
dsuu214PVaTO3K9vr39HZbWRC1L+5u/o38+K3VROh9I4w4sOyzp0J/7EHTi+6nGqtu3nlI/up92S
GVN8lu0Uookjon40GncYNfKhAJ6/JgRzB04jXGzXq+pw0OUnzLRV2dPksoLBLD+KRAtjfzlcEe/h
1hjvuIzAf+3QYCNOJ4raUuFnkzEgjv+amS7phM6c+xHM0z4sy48fBh8AbXR8tMwUzNwycoVgqkLX
ZkjXFCE4+TsWLOqi6O4+thhJKAyLgVOHggiqq8dwr+W/dj675YopFCvsz9DX7An6SjXCkJetCawf
j6u7WgO5hE4umXkZxbx686E+VSa8f1Gdhuy2qnKr+cqadfVi8V69N8F+j/YouHYkFj90pyt5lU5g
zcMiKUvHFAV6lKILWgx67HeOdtVNCphGUjzkpIeiNRzVn6aFik0/jWB23qjhcpgAHAxkkwD0+Tm0
YnK3RdaEawNm/yBnqScqwGk6kiUuEG2qK+lY1S8ByuDvmZPpSqmKkX/UuUFrgza32YbAL8JCxVbD
rtuLP0MgUjv6HNEKA4/eN39EzsxBodwbZXRtc2DkTEcOEKDyG7xoqsnw0y+WC8uSciMesaDo/JC0
kVUvoYCHvsT4B0AIMyFjSmKPaAT9C4AJ9rnjb3euuiFJ4Bq/W44B4hk9X2C76nGHye4slh+ykXcc
Tp+jyKvfIA/isE0xAjs08aIjYWt223y3Xm8/bQ4DTfC55WU4zRNgT/guKRQZ2A4DsWJAqLyW0czE
Rc+LKRo15hwSQoUkcfZT/gPEsoxuEFP1sS1U22Po2eRS0NwDBsbnLKeF/gG2qzdZOyLR8tWT+Wew
fIAKTYF3xax2voiPr8PFbqjlcaGR5D0VXmFoijSk1fmUec9TPcazBOJEM/AFe5GxJC7pfQxf4Skr
P5olIS3Z8LycBofMFQG210G6BaifDAH5h0zXpwlFxsvmHZVhJAWN5PKn/VsTuQIZfe21Chp2ft6K
PHPfBHlpw1fKNYUL4bj2+eGDJQOkn+8rE0Rqhy6DZodTwvPiHpaiUO8DlHh8+7pBnsqwRQza12+q
fig9BJWyK9YkOrliWb6HdVU0sLG5okO0sCOyHXhMmGSwGarY+5pUOpKFlvZySupqvkGyhVtntwXg
u2V/RJfAC2bGqO3TfQms7evS2Xj49V/llxSK9y9AssS3oJXkEeQd8tcBmNosVewEPoRpFyVg1Ixd
XahxrEXwese3/UhEYGw7Qbv4FXQgZ1dgfWXZnVDWjm9mEdiYSLibCjMSPBgFcbeocqCdfxBW+9Mv
m07tGKHsDaj01USp6JnfTpFR/dPPvBYWtDZN58OQzCN3osbvD5aRJN1xZFi/WXMlr4/6LZbOcjZ2
NfAx80QLCqeJ0tdV1u6TL21jWmd+6dqfqjjJEVlzNKmhBkAdYYPmNd7WWKqPpAMGWS9wcWsMi0yh
K2ffikaqZDytmVgoQKheQWRBTuWxIdreldGGO1EaHlIy9Q6bKmU7zitJwkpd0pFsdK0TjMaYza52
9NFkBem/DAEM1PulpfL0rG0+spWsTEVzsDv9YnmGsRqREEoHn5PVom9WhmaNvGRUbhnHBsvw+Ro1
vHOrCDcpVM5TyOCDSjNC+wl+LEXmQQf3mm1sCtjImHI3L6+XNRlWtguDyYiLHCMrFsQgHI7T+VRh
FWBZ28Qu9Ytg745Rkuzm2gH03ODICyy31RKxdC1duxg24q7tWar9aAosJpkszeUUA/gnKNjojq1R
fQw2a8IDAhFKkeI0h9Gv4hwa1Sd23YJwBKGaQTVGnfyBKO7Vc6EwVwnXmOgN+B82R+edwIeeehd6
CocGBknqCrDe+6aaGmynxPw0xwl4bLI6iWioNCxiMlcTG+P4W59jOFHHClITN0cJ5oMi9YYTAy6j
Mf3pBTV+GMAhbJBxTDnn0eU98yqtlaMg3Vl1NFsXQoijg5intjUT9zQRuUMlCkBEbpREMKb9/MHW
5vTkpo0iLh7JF8kZYdgf2R0R4pvLfcXJWIy11VOSJf2KF++qGAp2kqxdP5I1vt1qnqx3O4Z28dd6
lmD75tq5VWfXiII17WfTvhHIRrvTqmQfHsHNHeetbvnAajFlmy/1oiPnajoUZyQDyTgKKEzgLHbq
dts3SWC4ajyybHR5E2eAvhSMeiBAvBqW9aqQ3BoukC1zH8gFkeK+NfRE2HxGhC8YnHzF2yxP/2Lg
jp2pnmuoLKcj+cpkh6LSuliJorvec0WX7NekXP83M2vfR6sF6p+Cv/ZmJ3f+vEHcQ+HZ9oS1aUqt
xUgAzk8b5Uo53yDhmpMS5OdC3brKwmDTfIyfURwmapiu7n3LgbogMjMwaJPt7Fz7g2mzgHeYYkjc
7xled443xDYWYsYUyphyjrrRssHwYdkRXY444efCXMCWd8mIInG9QyOZwApk8Eygsr3tDirbYMGN
gbn4UeYhaVYkD04r1Kryc9Yxxzl4+C6bjIBYtb2hLgWh8RohOKoA3DdNMvpvqMhjBVNVrDbQxHUf
19NXbuGShBezCDCeDqbKtzTZA3eJVhzKu4um4KHHtxkiS4znwmtlhN4pJVGKTwlmcYxU5Dqo7jhI
aBNSVCPiCFC2nTzgDXGy+hzX9FwztmQU5v5Qelh8q6uBw/ZQamAexQJDmakS54y+HvaSBz+vUj5X
W09G9WrrpILblG6wPYI5qXCNQMF5AwC4SU5C9TcUQamK1yZnxuhL4xzzcBpoJE+RzHRIyDpUztPu
lJgN9ZL8YaeLWg5i4TUn/U5WYUWtn0FP6N0X/nhPPVqnAT1C/heUUVKTsnWZsHSZHEC4QfXkpSwS
6/ZKWIlvDr8g5G1fvLq1mWEPX1MswRR01Vjugl40dRQW80iQAOe/ZH4fDuISTC+280EsnDJUiWQw
u42qk6xatj/jT6B+fx9XUoB58jlKq0XLEZ9rhBuyb+57r1JhzP9UDcXAPulUw2dh/nI4UczY5Xp6
zd2HkP6HaKNqyRK9YYieFlYNhFvQUzLKUJ5xKAZCr8WaodSP0WRK0YK986gj8Tm05ODW04IYUxBk
KhM+qDy9AYtfYRG4DUG7P6xdN7BNW3Y44dUeyQRNTqmtYw9HSBFXVLkNdLcdermf1gmbSlZrhEix
Qbj7q7W+bC5B/4I1Pv4j3ddaBsvjLpUqZUN1Lv0m3qM0g+oYI7osuoHuXJqwmpls+EL/Wy7si6La
AtLlP69ikHdQKlfpp+aaGrG+g7Uebgg4OpeWJln5FLa5gMdf0reVTmsUnCXNHGt/qw0Q+9DJWBL7
Ys0Oispa9W8k08DfRvEyYZJDgj2m1MhkRdbwYqq+cWrSgCrE6srGWU6Uo/VCrzwA+coVZ889Q8gz
Y/Jd0VezABf2OslvcT5ue73K41+C2FRvIpZi5AY2MOXSupILtGzoEC2JaKvnnezTWmt4YPsrnE41
9lNO7i0v1ZBqtFeN6XI7vZ7DTdLORTO2ITzm5QEMhKpSY9H+Zkw4YnZMzZPK6p4MGy0RqlhQ51Il
RjfYUJ75ezWr8YezdnO6PbZ/PkCpspBcxyunkKQ7DtAEA+IVXnyXpSsZyOYRvFtDf3Xgy7m4l88A
Rj3aJS5ldUSmOLNhX52MWXWjpQ/Cd4xriB9RVD6KN8L8soWISs57UxMEEI2PZZDQ7s03IDsqyZdP
kdRKoBgO1BO9nPpFTZoq0LzHMlrZrDcaHIrGD2uKUDm1a6glg7B4mk/POSfFRkKOLEt7a4wvsE/t
2PVovIn7dIvtpOj5BfRgJObIRFGenbu3OZmnb4j/082skesg9mzZUSpaVTTjonHrQu1D2jSistt8
NJLWwsXGXOw16hu+dx+wGob/wGQyxYifLdpwTJ/idkFRIRl6wNCA0+tnuVxQhSYlLTc0GKn/qoVP
n7pa93Fucc73aJwzx1eR06rHW65/ZLdUYRt3i9DKhfD8FGUicpM4ibtIlwyj4Q5RyO6PSlsOvvXn
NBgWhfZMKK1IXEA9eGNevkbVe56FbiBtzxqwXzqeJEfBXITCS44p9nnyHcZRGNg9zFedZkxcFFy0
HAzrkbmWB4qhluFR9CNahYqqwHnBPX4IO7GorY3pA5h518SdPNL2zJ+ckOybzbzFonsiBhdzcIE3
L4vRvN0mgzEjpnXC8ZAwH/b1YRSjAmKEiiwvA+G/7iJ+xRm06dYQAH5w+jDo+ioTLoVs8nhHn9Lm
GCbqlay98dckY80Mkgi/Z2E1Kt5fSZ5lDxOzHZM+OX7TDTSi3JqVZFSZen5939lmb2YRiXS8Wmca
IS4erEbwkA9addscUB2vTzrkmVbCfkifb1wnJ55dZQnkvGe+ezC6GKRE8ILGZQswQBsSm/eOyBQ9
dkCKw55i7YOfXFDF1/xXOnh2DUpTP9lV7i0f8RCYDTKF7eGhQjd8d/Ck4fAIGFCtL1fg1Dr+ASG6
N97A700g7Z7F/KyW0x8QgYyz5wCISPuor1lAC8yLLtLhvfzHyEigb4SdQ7iFIMAsj0InsEnwhF3S
1MRfDmzSfFtNDcXSKGMlpUHpUjFxqGKtrlPYxmaoXSkO+uqJEL/qAvbWJPZAXF/DcnlOLG4Q+hB/
98L2RBa5Jj+6t3EthGH5m1Mqn3utMg6U3HaWR/35PM94JwNvNOg+G5gBiDkxE3shDwwrYllnzZ8K
CORTXTNZwEvptTRnR6sfKEq3R3i4HPPjWM4p2tuTqcY5npXlzZIy/Ej4IFhVhIv662ovDgDNCTk0
XicCuRaTJrXSZNFg43mNVGVTpkLZtTPefcBhcIRS4D4K2CXOPCuH7sHF4EMBUQlEhq3aNZJF32HX
1h3AHQAKgQNIBd9vaNZIaxGbhNYe2Fok7KEiRkKZrH+URHlvmtwfyHXyxj3vMzuFm1/Oy4V6fzu/
6VS80b9URYN1LpgcRANGk/s1cCIb7ooue7uh9zSZ6wqXCiIh0PcGITrWUClI4poGaZ3coH8qdiaO
NlCuBFfbpTlYsKKN8ONVONkhX5o7ycsH2LSR+afW2IYW4eusPNIWK+amBUefl8S5aa3TyogjTmf8
8oyxrLpHMk9SCXuvkl1IcYDwLEiPtPob4cIM+EAr9vExGz/8SHoauIVjdMRaE2QCFG8q2MwyroVE
ZrUMaxdVxAhVWwHVMq3NooG8UTmx0lXamXcKxOtHL0BQUOssrOijc5RjeY/6ZU/AZij0w8lpkEDF
5g3muNPAkZKjx7RcgAnO/G1dpX+FhOXY8fU1d/5rk61JEigQD/vh2EJaQsBvy6ZEeOU9/fjQGeQ+
N4zXOIx029aOsX24ntG81iACkZn9CHRWAeZDj/25cHrCqS87svvfRO8V8Aplb7hvqLQubsFDi4WG
B30VpYyWXriSkXExzv+jdMt3SLxOC7v8ym/w508eFCQN1PubYiVuMZMCYfXnKsA+UH6Uo+T8oZ5G
T2YozXhpoVPoVYuYifHwGep0yLGBjzkBe5585DPNkOXioELgYOv1qgBhg3XDLxLClPFm4K0wfIM6
5P8t/URi8F9zpGICc8/OeOGjMb0VOixo0722/229plFuyrmL5sqNOdPB4MInQ5YWFQbCqxCIVBf+
kxuPXxn6bAaR26kiUTHz0lTbTRLL6OmraQrlxZE/yjxqMAnreASD1gJ96Tk2CKsMwSTfKVpjWV0F
vr6HQ+fR3A0ngcQhk2X4lbdDD/sPYvijxbaMjYqfSutewumTB2H/6ARWrlC/0YbuV3X7QRLVUGHS
rFaqMh1Cc9rAGSHTE+BRmQe5BpIUlN5wvhvJcA2lbzL5l0yXjH32Eubc68QMwakji8xOyKVolU6i
Xe2nMdQvtaTI8hJSbiMX6QTmedhWdovfSQIM/p2GRrc8RpH6XC6DCtAnAjKwVM3BX+6bTFItgMD8
GKneS0mChdBZ9Jy7lcLw10PHSWXOSXdQtN2mThUnEE+zae56N+BfMy1rj49izltSTpOcWGlBJ8Dd
+cB+CGjC46B71ApwlB0GYuwQ0rMOPn2W43tQMrpJ0+jW5Z04OmrJx87f3ylznjJFg1QKy4dzB7a8
t0xMdWrPIJprMeHvkkJoVWBrGR1OpHTaiH8Scs+pn9aB4iQx5SBiwJR4Sar2eLoYV5A4UIf5llzq
uF9VcH4h61MnCPdf8WqBIqe+IkjYoPt1WzRJnWA3uSONtmz9z1qFu5m0yjEQYTyeNN0Denxvwi95
wCiJ9QPzfW3PxN7ti7RDvLquABxu8V1tTR6gNWTnsTipaDJ2gILoJBXfKvXKdhx8En6VnePQw4Xg
Q8nnfgJaxH4npW713o6axsCaLzod/wf9CMl8nC2ROq9YgV9zatOq7tHPCciMOBVxC8Of7+17wXwq
v/ygXrhwsdWli6zPijo+TQ0M2OeXcEGSZJcC1zaT21adv+VnuGosM6NDZaqujvU7kqkt258WBRT1
ykwT79Fx1olxmzHXVHF83pgB6dVzIfLDAmcnYwG18qrmHS+5cbEVAKdWLf4pfQMD9Vs6RbGf6wtX
yQZr5yiVE9Khnn5jWWnSGaOLLbJIngNOQtAw6AK/b3OuhlmBXvhyhVhyBfRmdUdyiKcbv24zkI8a
6sCEAlNU5w5IDqYLIyYpWJ1GwPUkpvqmaOP66fCEXkx1qrvruqa7PgJIyLYU6fH2aSOvfGm/AjTW
RkZUMhHIY1D0JbMgglmsosu8cRAAeDaW6LtJ3icEMw76xYEf3GhzLa9I2KAu6HTr00KgGQi2qSQa
9P4WH2MGkNjHlRbrGd5fBDR1wFK+/yWy6Iau2fjE2SGGrzJMNe9P5f5ZJDML6L309KCK03HnicCo
vdHCL2SYfsPEfzGZCvFf6LaxLuiKXZbDntpTU7u/fuC+p545wXg0n0XHa/X0vxbtg3Qo8Q2Ry3sA
eCsqOJ3yXpMuR3vLg+MHljRMo5f/C4rWKtnD6devt9da2+Ntou65X8lTSpeAYlWh5AjDuhi/ePXt
TRldyc4WPmHz/HxOcsVC3Tq/A0RHyRSNH5InMjDcxeUxh5+0ylcBB3qgKRrILnUX1LZxfUZ4SwBD
5lSf1u1GjqbVRch2ybZWK/fudKNdNbt7RKR9ncTOuJsF1C32P0BS28GyZJxEn586Qs1RMek12Haz
Jsr64OxK8OSOAKCk/ga+l+wd64iHSBHOj6mCq7mFULaHeUZgv+9d+Ub12rCVCwUWj80Em2W9B60u
01pHw51e+4eprzdkmgnL89eqKeAFmqg+HdAvITIEbAujbVZicWYsdRatmPjoNlKRq1soVO4ysypa
GzSMDRaf4x8LCnTi1NoHAmD8eY7G/PFneIL40Ee0WKo1iCs1U8PaJJSBII0KnL6tkMHrLI6UYAzV
EUNNe/c0UtyrFu1eKMnrDG0JOJDGgt5Tu2KT8m3SQusItZLy9zEfaf3cmTvGg72eidmiUm9WaYlO
yP4sZNQg2jFhS5XwRZctUfyJPsSsVobodMPT8YJQSJRSC2Dq8uydrf9Qprqh1J17PYMKUK3ubY1h
R4wk5MkXX6LWJK2jofpsLgwiKvkgIrMNq6Xba5CeX8aglai8fGHQGW9UXdQKduus+Feirsv9qfub
wvZt6niQQxRws9BvFyN5EKFBC331KwFC+PMNGxgspt6vWlKRDomNEH4n1CoW/VLz7IJwUwKYKc6/
Ni1vb2p+HoSAq98/lvnzDlVTQjHLssD6fici4RtA7CqWQ8rCuUZ9sojEu3vYD/pJzHSsd+yRmSXb
8VOqLU0qLq8+J6BdDjydnmhoKeSffLIYlQYMhPCw7/eNZrfKoZgSDIHuogI60ka8z0qDcYgXS5+a
/JFCMO5R/oxJ4K/wWXVREO/1uQ/rgtgtOH+bWhgv1exOObliiNS8Jp0Jbn6eaq+TuwnsfUYrhImV
S7ue5HsBlSOJhZDCqfq7XRnnpkaAmAJdmSkYbX7YN0ASqaCGCYucRiuFy02fzhKKq+DJzD8Djje3
6EZSbfJOLIRYDCRyHsbR5k/G0SsxOX3nqh2Efbd/GvEOJ4gZRr5sARHl6Yzee6W6hBZFfeviaJBZ
QmhG4VbluNbS0Ivf/rGT8rBk8dFWvfEUnXjTyxWHMlZXR+Q99j1Nyso+4SnMVek1pfI+1OeMFFn/
miS5vkuermvijtNqdgJicDNumr/tkrzW2C325NLMnuShqjWZFK1tutl/aQPzDurmKsofj7eW49LT
iW9zz2fvvc/lWVwBb+/FoZ8NNMDXIDFQXcGYg0zOW2VTCi4ZRY1k1DNxw6GaneM8e+Y9odUn9nPK
v+0PAWPSG4PjLBs65yiZ9lImrt9A8aeVP0knn8UGtqLvM+huETfwY6lh2BcyovMR+iLX/QKDtY+f
B2BZ1x++TJWZy3CHm5T6AsmwgfKbB7dd6q6Rvvs2HEJL8XpbMtEKhTWyw+8Irw3bXcVtuEHaE/yN
BERIxCVHzudQzhp8MuVEcVG9ID8/iW1kk46AQNzSGObzi3Jst+EaMurEQfk/1mldWlLAERvvzMf2
n5fDhqZcHcbt0MknDDQ/KoEMiKbF8HPt3WpUBVE4bb0i4YMVubwLQ7k06rRpJL5U1iDrn5gqg2UE
2m/adVPyLTraDHY8FCGRltU8sXhbam9+rJWFE0AzbMeJtkDCClHb6MverI0HjcPr350ZCAqJYcO0
HfNgJdAoOT2oRq5zSEv6XxgZvkehMpb1+lsJ9oOFI0OzZgVoob0MaBYCVcaHgDznDfRRIQsHawfF
DwdS/La2prpuEit3R44HsmtKQxSEltvr7CwwTgZvKSdUg8IDGywH5ywc2ADZNjeMTmHJx47TVKOe
ylgZZ5V75MuuJ4rz0JaSThIq4smTcgq+rCc09hkOK8p6krjB0OP552uwjSuupCq9ti4IOCpG7+Z9
aZ5CLmz2IzdyL7apwzoCjhV0TBG9evOVxolZvscODgyliaHAHJJmjJ20eDlXL5p2kCWLQycRBxlD
iF3eN4utku035RYYZUhceJiucTnhL27u8UjHcx69JKSUUv8k8jkWrpVnXSNsuCFRxW+5NNAsLP2Y
akgcCWcAbineVv0WvyLHxcb8rl4aB+2AtON/x6xZGdVw+oszvTUAGBEywQ3Q7x8ehHYepvqmkWQx
npm1L/ysCGwIRYIZGeJu0Og1kMdkxnmhVeNVIT+ERpFsDCvVbp6ewEjWxu3Poy+bnrLtc6krTi+3
s/xcQJx3xBO+pbuEYvHupIHk/5o3qqH8xKIUKfddsx4mDVmoVlskQ3YNkwje9yB+iuP1A8y7N1+1
cnVf37O3Jw7TlWszLfGv1BUlb702riVcxUDxzU+u8VxddBD69TB+XnDU0yOLhSTrcJfrnAIO8qFt
sJQsMCsK1PsMNzHQGw1n6t7O2BrQeE2lQpwwhg+xzjGAt1Pz30a9G0LjXkSpRzw+Kk9RDuiD549m
awCh5MXT3ONbrNM+BU8Rku46Y69CeksGHAnpDKFdY4YPNNHK5/h3jwXlGriX5RfX2U9GslChzDLQ
WAUOxCswom4hkpQroIS8Zes783wh1CJSTUZup/0+16TDB3hV3UVat59x5+b0QD/e+ZFW9L+1HI4U
i5dgmKwL5EvXXkST0YAaAa4l1Hd5yDX3wulXiuct7Uiz1JKeWZzpJ7a6nYYinV9qUhHmo1N1v1fZ
Xi96IfdvybuDlP3QOg3LYTxKYpqxad9CQN/3ykdfV7iqviYiem5KgCoiRfPAGuBgzfY4DVGVUp8t
iOWHX9fEGXuthZnZRkd146TlOHg7rgx2LGOcE/xO9VhFMr+6atDvQX+UT8zx2XAQ5V5QGf7HPs/n
uJsKphz+IXkxr37eOHGbvsC6hP2Vx5fd4sxARalf1Zwm655bfBc4rhP9SgPyHc/Nms+e3vEfYyA5
STC5+1lwegVcxWUVb6EzetD1SxRRNNmC7UalcfIpkKqfGDXwKkS731VfOLQjshE8PjvUuMQGjPR5
gjtaSnO0GnUO0JWf4Gs22/IasbMBTzct6nrDSyupc6k61e/NPO291t3f6vwi0COOZEs2MWFkmgZl
miOIDJUEsXwdOXPAY/dfLGnnOe0qYuH/eMhszm1VCWPlQ4zRmQMPeAubOoN3xV7UM+BcB1nDgcmK
4jEpgXhMssKA1cvc8/WxUN7Ojke3LMYSRl5JpiNfOgJoUhQCiTxA6/neXaHyjo9XjPfzXYbjqwsU
NvUbYNtxErcCJOjJdXy6iC4X9ii/wo4vyyZ3+6ePrpop+w31puwIiqt/mrGbRy76s4jwZmqkMTqo
y90EG0B7SjduZ2Cqf0JPvOAM1EpPzX3oWiFToBUgTHl4Ab189FreYTOH7OGrEtyDXOHxU9lgSqF2
5+Q3mTXCZrpsHbUz6LYC2oqVyLxrO2Id0NYiKN7sxmGTLgwyHy6EpjBJi0qsqhiwiDtuj9V+vQiW
uI4EC9q3etdZghS9gko9Slhj+Zmw8Z4le124dOqzuGi0q8KIqfYSV3fO5cVAqS6MoU7t/SwCBd5x
wD2hn8GKyNg1EHerANRhZKxmEvBxkvSyujGCr6FoGyOPXB2ar61PbCbXw7IXsfgzwFvUxKk06nO1
I2PA3XoMkjYfU75JAJxtNQiDk4Hx/U6nD4o52XJoYSMShHyaKXuv7oKPawb5yncb+uwWvBV0wONf
TYfnFsIobuQlrbYcRLVK94w+nLT+yeKQXwdKHNCZsl5o84CusTLT/sBYKNMRzqZZNZkkgkIfeY3y
sUKHOYuiy907TjABhno1KQhxYdYXPACI6PapzN+XFDpR0FnXyNPbpbpJ9YddRxpuEiM6wU98vDNn
o1osu1QhkObCL27CqPrv0P6JLfLl6qyMYFhgvk88hFX5siS4UvRCbxKqd5eL6liEwGw1eK1ZkgTE
TrkXbv1aTuxmgAcbIe4u/UFwKHnVqbZB1WhQstoE47e/O2yIbBSurqt4qBR/ek5vzQhyuUbpvppg
g6eihsj5oariG4fEudqjj9DJ1GrgV8zqp70fy/NX6vht6LUXLxxQDAjS/sEV0l0JO0Q8qpr94bCT
mDmZnWJTWzErvxh8ZFtKvquRgywyqve2Es+nMTObZ6N76HX5Yl6XVrZsxlLIs6Nihj2Kl3jib/qx
ntfwgAP3+ts0mB+PxxLy8sQXwaZ4gcVm0EmWy5BANGc4Uj0XNp8M1UBtAHRAuJrp2Yj+MlgrB8FV
CDWzm+6kDkwqzy+3kjxlYUdsJEN6oik6IddT3mq+KfNaIZ7mUHmGfV/YzW9SLJrx6O/RYp/1SSB2
aLv0pf114q6X7SbDxOPUW1rEZB4ULbEajQ4ZcItKc/W/N71cctlRSFrn4cGgpIZ03jxynYXN2pEN
szKaCGBi8qCkC9Skft9Gu+IW8fkUi8Vyu7biI4fBU8k55s1hc7HYBWWOmCrjonlDLjPv528IDuMh
KK6c6X7Q3j3gL/Z+bgPLPKGMWIaDA4GQaLU5dQGkvEJngF7OJLNbJYCl0fOCACVjh0ma7N5+uZLz
HvHfIQjh9UeWOFIL1S9Vwg/YTULPOCsTGlioqMlFd3TZcLfgl97pO8HL4Gq28/AcXHQi07KgCJMD
hnTRCCzemIfUeBLwW7sZa9iOqRIf5RPWW9PNR1azh47Na2fYjWGdl5NTDU3RrMpWS+LaoDC8ELMH
bSxvjq03TsyDlp4zAMM7plritsdZDVzbF4uXtrwVawJF7brOr9IayVHhR+wb3mwtNQDPfEF7Z6Pt
BRoczQHxSRDDTobqjJp7kEOcl2gm0YT3hTgwa4M0jfCvn4yPZM64u6KVg+bp4dBwXhVIMeShVU+7
fpu7tKLJxk7ycfpRvcIacCxy2fGBynjvoJ8Y7KYvgsRyIzR86PyirHfPa318TOaMej2f92SxeRen
K6jmmC7tph3QCdBf436OBYWqmsCBQIU4cztxAikjzcMyT8nBY71GPEAwN8Qm7Ks8O5fkL5susF+C
8VAPg+AMKGjuFWZCC7ZjQ4/4ErzLnYWgfhZ5Fr5jO607mUKNBHZxY+Zkbh+UJwS87Jm0jl5LBQwo
diTo6PtMPVcmgOiLTlBWul7B3iy7FqEE9/0a6MnDygSntwp2w4G4SNTBHf10rpIYjCqE3j/+yacK
DEaAZKFQVZwFInl9S0BkL6bjSpLH9ZOatvWt/OUGpy9oi/0NW8I7OTnAlR2OMdKEuJAfEM5CdNhK
PJc95jk5JZ59DxZuQ7cuEc1788IyuCpFDYaJEYWceT8cMpMVl9uZdF14dX8zav6xLqWxqREVq/ff
BiK10RizJF1YKE4fREkp9IpKE6PzGpZHaB5275inQLqe61y65ulf/Rt+5xGeHJdiiPZKOlVh5YkK
xRDKEiWc5sK5edZ9pskttNqXFkzmnMt1wo3KznQH0YHzmKqHmoSCPxX//wQrqd7hen0P9z6lUQio
vffhq2qifJ8V4VK31Esqbw9VNHYpbQJn1Hk2BT0KFecafnBKPibj7KnmA62zSbM3Uakxuwr/6/Fw
ZORjmFrNXsit5e//aRHqXWIel3R+CrbDJHjI1ArQjky2aqezkrzx9y//DQvmFbYVrzKRUj5kjFQj
WwsLIYXIzNEX5KgoGO/5iHtRpSlODGJcrTk/nivnXitye+XVoGXvhOa7ix2oRClet4z7crdPZcFu
aoGdMTLnw7R2IgVJR6bk2xuwuomXCrVzAUoJ3jDcco6SlkBFSSjYNElQNSz61L1ogt4uwB0ld5TZ
L2lV/lS2+54EQsfkmOkZIoC7+7qu0EBCthhXBBKafrW0Ikg3TpDkzlj3ZYUvpda3BHetRLR7HyBg
hG7bwY4sWPe7rf/IXI0fP97Rt83iqFe56Yg0+IbsBVCJkRPWfbyMHQhfVF5Cx14sxtLpQz3OhHEg
jYKTbUV4C5ngZLhQ0ejaGTqTeQRN7YLz2ecZOh5tPs8ik3QI2ew138xuvUTV7yHj1N0YscOdhrF6
jlnXFOnBMpmC/ImsmouAWRcxmOmfA0tKG7Uebei8S/bSz31pQd4h1+V7V/UyJOKEOwHP9sYtrVF/
SRrQTk4q2fBqnrdnIVKoJ0siCAUjXMi8CiQsvknTyJg7YpZcOBB8fumoYFoXC9uIMLsAW7rDHmN4
cBF2nkTQW3+kIOEZwDM5WF6v6ezgvEG4MiYv3IPC9ubyE030EoSSZ3ELREs7MCFUTqYpPWhrb3yR
mUGXEHd9vpCHgaxOSaXYXXFy7RkZRsEi8C7TkyFiP5TiIxTiDuj7mgOuqcFsD7uE3f/4fgHeDEEF
iZD+ITrq3PLH15rQUMvSBDUJ4In55Z0og5xbZzuVLPkQJUDqbIKpPN9VS4uPKKMYjkXhyayJlqtq
Zms6tbrevbCMw9zl4GEPmUxvhndCZ+QbC8X3lmrt+cMfvz7CC6Lgq/f5CshJ7K/4LQcBr3GGwq11
Qac4p1Uit9q5GMxHjPbkGGOljyRI+Nh/5UYej5J5AROpk3xR08iworjHQQp6yJ9oiZ0sV6YUxC2i
FSGOPXlz4INWzrWWL+l6dJdyIRThLls+9jvU2CvftqHbvhtlYxUyk+H4TqzY22ybysCTkyvInIDt
6g4TZAve3im3CuQj1lH0MQIjLaUoxLSnN2CxZ5jqKxfj5VaMWfvvaop7T1k/PNYsF3nTloI5XAba
eI6dQwrk8aM3QGg5RmMxfKggCx65Ag9luKtjSNeD4X4DHJU4+uERrXPDhO9uG/lfS0xmESEdTdJI
I3oSl83EqvKOp0HLIz39yP7AcWQsKtrIgxRMxu7tbsZ8zbQHbj/3b/pYYZJnXhffCQjHIm0feapH
oSA7Zu3Pj06wOa50DWYnUV8YYz256+4z8jRIKtsi6rDIfERJluIEUufsw1/+OCBt34n8dxdefOpL
dHq6ajHQBYU6dSPoEAr7NJTgcO8U9A/T6VMv1RtV4nBardKNuJO6jWX6BOAAuPZg44ZMwAw2pDIB
U8coarlO03ZZUnomGjm8TszGO3BzOU7uoFsUZR0/kqVCA9scakmZoFZxCR2ksBBejw8Mo3w/qjyK
A0gpHDqDkIQyULsjjprO3Y2FAPNcYDWZWFs+/+N6LRkAKeU9Y6ywk0SDLt3nhCebM1LIyX/87CFv
uk64Uod0NZs5Qlq/LYTjeWf6dqKtEFA6H0UKLYnh9zb9bWZpQometVwRxnZVwJLfoWMRnc40SDXi
2LXLEuCYYRR5K18VX3fqtjMA/myNT+1ewoKkikc0l2L91ZAQBxP1Iro4/qEGtRWTy1gYKBTb4Xl6
DDfrO/2+H0m6SZi+PIs95vkPHBmx3QWa9qe+eAXIbT+0WUcTiq0TsRVJi8s+3yVyC705NmrszkgY
BVl9cGukluacsq24R5KetlmMwmmvb72+YsUTBNKhuDuxM4ZxNeCZCHwoZvoKq2GWby8TO6EgTliB
uccsc+xe0PojLqLy/7DuyZ5Lx+NTGbt4qsY8kiPS+Q9Ew8F/v1/ZWhM9NX8p775doOZBvt6y9Uu5
39oGowAmkYDpBhTk9r+JWTGPAk+YY9vXcSjfe1gh+CAHpG+4+UNuzxCcLnH6g2+NMXEXKsnjB3Gu
4q1DG91WeQdKB1GNTek4ylh1QUzqeVJo4WBYvGOPE7A+60f+sv+jnwztV0/kmEOO+GQny19KBzVH
SpX2F2RGPuROGj6eU2k7JOmtAT2GGR5OCxJpqGb1xRFI8TOltVUUw/DOKn0sSX/0L1hIYdESK+Jn
55J2ZnGuah/sGLJATKzWsLhdmTW0B08VKHsaDuX/pBMeuGQbfbzdDNFBrJQA8VZUFBtDgPOaAIR7
kedYPl9RNKz9nr6F2aPDv3LN3b3qkr7ND6qo0e/DDTTwFGExNSoAUkljagTA1Ok0IUJEWoxNJEOe
jCgF50Xg3Az2gz4cdM4I06wzBuoMfY/QYhD0fOEDEH0SZJwX81/T3qBFGvv+NGcI4nZf4wJf0EdZ
ICCEttixpgD1cEag0Fa3cjm3UtBhs3nJzOGT+E9UeBqY7Mpe5e976dLJ4MRJCtat62w6YFJNSsvz
Nigg0qaSxbirkuMcjCeexdLnE2EHiHjLdTm0RfIvhpIekHqsr/R/ZAuZpnEi1sXMV1d1YhAVSBAH
Czb28aQBsECd78KtkmO8ODHhLcGW+mdH20653SWwh7PbGdbhCluGlMs3SDRMYzpIGLETaJoLBakU
RvtFromPAHVTShPJm+QMTF8meGxroPcGzEv3FXi99r0m9xTGofVB/aVRDSKC5DuHSsHMcf2uvjzp
RWlfeI1Jfl45n4nztBq28CDmjse3uCVZxaTN0/aMyeJ9H3TiJjhtiztUwQ7G2HVBB+/7YCZNaYTM
pAD4b9ONgk9d0/0cMMo5Q3CyRrYbpeWtmDD3+EBIEjkO4/lYOL3gGyaurfylBV40Tx4tYYIDOtc3
FDoJJsjRfAO6yC6hRGc9b4SyrWhodEDYtZqhbj3ajT7kcWoo8Hvvij9W0waexyiZ723Kc43jnqFX
wx3pAo+gRbpNupnqHreFKM3k2XRO2bWIwec0KDDUw75S3R4/b49rMyIOdWms88cvap15oHlWlutc
C3CWHyYiAXAmVw1/JmPrMuWP++FKyMGM07qc8dtGsAADBSv1I2rtTgc1urg70itPy7lHeSR5g4N2
lOrvWxMsyAIPJQHBDkoT1MTnGjQ99DL0eXVi9CDzFaYclpUkGjXKiQ7ySElWG5ZLRKdL7fkznf/a
rO7LvDhFMAN5ndPy2LAadhU1XgtHvxoSrMSf/REqkf0jXsRWoxkCzoYCHXIwSVyZoi7hYqd0MmQC
MMmLeUcwxjsKJM6rJPnc3DK9hmpG8jPNs7KrrXUGF6YhfepyC85+tAH/Kwkulx3Jl9dmVb9s2d44
G/EtRLAGBEAggjVKZqjD/siAAwfRKK79f8YoxZ8d+dPrNccXddWY+CDnDgAUiFIiYyNj3Tx2oMiI
PQJAq4rj411PqZ4n2QUV2o7ARDSX2NvgJxJKRblKbwPES2Qxk28E5qqG+v29SDTZN7zZ1uEpYomv
SIzrgcsIbRvKOPEW8X9H0JZ7jsIO2TPNrp6iteoKurlMgR+tu9uqOPowQkpTXGbbl516msTHSqqw
5nJATOxYyzGYxLn6AcbX0s3AM1FvK71PgGA6cLF6Fxnr+VNxGxQCXFx3yFXDIKyEMdeE95ZUBYkk
g7f/njTYCwgH5Zvn44L/T/dHdr561xSAgjE41E1CnVW7ol88KQwhyBMUp5J0wHUpkSriPCWr96VY
KBczrTrCC2w/SWUDMv8ABqAHfwzKD1/GeAD975/AxQE4ew0b3LjdL6erBA5eBDELCY8/olLy0fca
3lG7eXTYkha2NYTs2jKjrnwDWqQBjAZ7BXtli6/Rp4Y43seqCRVVtMrT50GDgCicgBUgk5xZYuqo
IGDTpp9zYB4agXxj687jSybsOAxe2Kk0zLRd14fzXOGXNbW1pjOxT/LN2yy6kb8MEwINjyiz0Fmq
2z+dqpFb1OAcn0EYdZ6U1AMJczeToRfBvRt2Q7htPb8By9lOVQq66eARsUy8icqXsHUE2sPhLqX2
XOnb5071K7f5iKzThAQZTGWeJVpqcaC4O9m84d8SHyRsiico57QKfMBX/jo5ecKI50G0iZ8qghCg
MVAwSxsvkn3fBxGy/colssXJFU1MMpBGVFVGvi2KY5sPa9p+Yk8owu3wDcyTi85OF2kRBoLNxVVW
FwEBTN9SfuwFosrLHbuuB0kSSjbX0ZMdHvqt+ch29xD5xczWhxXkuq7NV5Mm7lyRcl9jlqpcdOe+
EwZLS2dI7zBsSgLDKgE1EOgOEJ89NI0ToExU+syZr0cHFqS37heFOrBEstygtU8pkN94CaBHAVyR
28NmdJlPfI9kmjLhk3+WcGDOIV9N+0NFq6b375iUBpNxRS5fdk435rw7ekqU1euw0Wlpd0h/93r3
zAkMmxbtcaPSw2Jnm8Q3CB1ZUdpZ6pImotPht3xLvKWXYdo26J2JiUrx9PgorM+l/OgHxWK24IHw
2DryOSK6LbFvfJeLuki5EB2tddB6zUYM1GnV6qKFm3XF022xn9zCwcnrerM5Faf7eyKqCqjQZK62
Z6ncCWfQGfh2tq5eR2T2sPvE9CEpL0U2Ylk/NcJpEohRnUyyUda9dWdt/bsWVWAPTN6S/dn6dXmO
9eM50WYUFITakKBfdldD1fvj6qcRs0OybWIxvaKFRC8LUk60DtmgF8pHdz+hbxV+5zlh6hvdtpXb
8/pVp6KKxxDlusQjA20jWWIbt5IsUbJztxbwZeRwX1b8s/672TpzxkFxateW8R82QYlY52Efl6He
py+93IxtiahOExkhzUv6X8EB+T9nzB+j8ikPGegrgINHIaWthOkfmW2Dmea5w+hqBH4VLAk1vnWl
G0YlPFaaUQlA6lOFo0fhpVALJ9hjOHPxLYMkBdAa0vMbGMJErBTefege1RZHlcb5tio35WAeBqsD
34qw5qnIQ8UpPGckwS5y0w8+mbJsAZCjg4iqm7JJASIAS9u7MijTfjZGRZYbhdcVzBaoGPDK13rh
JOOxHpwTX6MoCLnS5kXExTYfHvUYbOyNAvvlB5P4SXnwog/Czy8/KDK0nT2SsOYvOxOqtD6DhCH4
x7cS0od0u29GNiCSzR7qSud2qczUo8niW0HxviOJyMPsc0lbD/Q5ZnV75yKceod2+9sAJxMJU+5G
KmP2DMWIi9e/3DbVqYK5iqF1YuYO4rd0Na/iEKzXJMM89PkdH6zDbRUP5yJ3lll6XNpkG+hzHQSy
DrIjf8Pw9V++NLo7horWG7+03UgV7t866zM+5j1ditbRyIhBQHXK8NJP6xwN0jnsIVvBVkfRI+Ow
6g5xzyOvQS2RcfKeBQ5YzQeWNr40d5zUeZWQEKkrmoQ3iwms4OZD66Idenfr8HAPeI53AKRbDn+L
ggb5zSJXYo0HJFmQtpdXxh+zlyX0oDcnD7gXPBuGdwY071etjLsQymlb6lHuAJ/nyRjo51933NY9
GpTesBFwse+Im+2x3b2DB6wgL56e81fYRLq46ND0PY+MDk07LjBrHiRDuy7XTHobNaxGZkG2dUu6
r4HOm2hXYlwAhjeFYB/pb3VUzMGP9Qkk3/3d1txTyHI/+HCa/zhe2RAzwR6mKwHU+JUp7qz/h8L9
Xh0v8zQHksoqkdF/3NZ4vh0nfvU3br9HeV6gil4RTSCwcrRbNbqnOO5usDVQqm5Qt3PEGLpmPUOP
5veNuNAeUi71ju9diKALE6pLLIqJ3Aadzyc6ZS15y2Hqtu++xGMrEy6afgk6jGObf93sKEI3y0Qh
3GrbInf5rrpl4Q+I5Jpb6KJSJ8OypvzHyPZB3QnynAWnDX4zvuQAcJT2Z7aQrHqyikREEYEJLUf7
dsKTZBA9lfTtkt/dDHc7jObap+x4CMnerE5qaDsklDVU4NvwETXx+tbYAGXs845877yKu7TLACaI
42jrTTzLIsbBjWhKoKWW32oBCaoi3y0GNOL+CL9cLuHNT+N/BMskLmtZ140XtIlHcMqppZ6qaRXn
3VqdKsv5QerSpu+dEcf//+aOXHOxeFUnL/euG0ZVVcUoiJii2h4osTqzkymI7Dkgm3UkTI8Mjwmz
4yrngrq/VXw3p4nONEAxuqQJKP+w8j7wdVKxmVwl9JEIx3N/2QhjSs6NiKPSct7uEcOMoU/D2Jv9
uP4fPzwS22+KQqayQIQ89OkVgsn+GXbP4WD49QyXpty/GTkJRn8zpCxnfhW0wDsyW0tj4o4/SzZ1
ona2goCxG8E9nVBh3gLyXa+gM+qqmwYO3XM31d8igxruokWhr3DQa+5Z0OCXEkRfFxAQdhh1rnUn
jwH8QUOTwmtlh1dLXniNBPRF/NNzyRoF45z69myC7EfJf/Tn9z5TlZc2gFyTHKRMVBxxeaSY1WXy
9RQ7bnz4w7g5y9z6Buv6NHpmZoZCNlsoUNAN9KRXYunCIjGbTeMnc2/Lkovro+kQOVapxszmwbvA
b0v2EYUh4007DuEq+AnRpqXKHbndP+PUeIDvYScQzi1Cqss3uMMRj+G7uapD/EChC18hrSBo/xtB
k7gg4TijLMVhcg+/SbBuQkCnaoDrnKuzQv7meNNLmH3F5xhyx8QLO+c8IcKpcORvTsrc0cnKUHmj
0xTs0xs0P68LbY1OXl6pGBvGXeFS59V+H6YE1aHJOiJwaMLKGL/2x3aGI5ggqYqXhHxCWsuEYlSu
etZ6wCIssnX97KvIJ0gi5BhK2XkJLqZN3AhJR394kBtIB0lUjDw+4g+Sou2Nv7PSuk4qx7YwOhqr
/m/FtCVkr0h6BZ+2exBbP/cDmwO4GiPCLCkVEOkGFmi51iwb/zu4IqWNwNp8n9MWUH/ztcjKVp5N
Nb7WONAahiTjORKJgSsBMshzy6HIBuks1D6R/jjzp0GbsFNx0dMEfTs7Oae63QCqLlBqe5AmI1bp
ySsG5slNCz8KAvVL3O++e8ULonBKXP5ZCPraP7bBnMVvSu12NceG8S/hqPusJHYzYuJIOakuL8WO
i4OZjUe6A+bN8CswKNaL3E3DWGo6dBLxLQn0z7DVwcwnLEhyorOfa9SrjdXTcM5Z6RKu0CiD1BT/
1Z7/jHHhzbTs9PPWhYsnDGOUZe4uAZnRUwIZXmWE12XxdMpPt5SAnxB0Hm7Yi9cxNiriz4FvjdgE
pZTAOtcJrONQuvG+5ipL39/l/Ok2+X3BRWcBLvnCVe31uhjemgykvJZt53Sy/6tLl6cW9SBryGYK
85sBkqPXaaU0ACTR982oMDRPr/9Kx/1kqDF25KDrCvHNoKp5b+aGhmDZOBlWMMCy7PGdenyilZlQ
td+w74fElIq88LxjHBlCmLu+pB28LPjQqiYR77+Fmo2bdraDQR7RomYunNifQIXCp6naRmz/KaEo
gMVx06OW6WX3SbCdH+VXbDvOr9ytyhrxExwLc9NBE4U+1veaUFSmPYnNHvDjBATZwSxjqIlr+MDv
ZrQnxzNtGCb1j6F/pp1DMtBaT9hqj4ztMrLNBTM1KjNl93NnmveZmS2pqW0imlsIGW/lX4SvltOG
HDuAW4x4ePv2pcmTnl33Mqp4vJnPO2+fnJ6jaWrPWEYvsXcvz8HDtWA3Oh/eUaFQU++PESkTKQyx
xYWeohh8nkXnB8V/pPYn98VKala6t1TYbCn6D0BPi68SRajFk8Wc+O+qE1AtN5/Ko0Co0UuCbLgk
u4MiMwsB94ZeJ+T+poB8Fucy4FqzStQFZwOQjOwI3ld6lXKyhAHlHVwfDz9tSnFDBcCC6kHtsDcF
31PpRwH0jZzDHaJnUfXcINJSdlNg3+ijSks2WT0fpTlWUG9RHTusrmmnTRYlZANRHLULMjd3E2rb
/qbWcgo0yItnVy0RrR1MSHf2qXWx45QlsaA+Vx2JMwu/CGOwBrwFaetzlEthVtk1JbHzvzRT5LPs
tYyZLyZIZk+Ctcs8aCc34tJO8vcs3wxCQyzy4qJLRT1oEzk4vFDYBv4VX3JWpGDUTvshZ+IqU3sT
6TzGr8IoZYm9uGOlmw5OLk5GPiQBla/65e7ZjcXo3hqEBE9Hz0RDHmPTN4nLwKMJK3ewppDouHM2
PHxcNNXxjBL5M6cpyIR4MEXwIKI/MtYLdWHiX0ww6uOXQkNrvqzFVloQl9hRajujPUww26ZpBjgE
pwVWs7VpaSwDCu/baeuaLVuWnakhRrnByDZOJUma4/8JIUqVvfM8IkVSoRGWtRW2eCD7KosYVeWH
TJHUU5BHjcCa4kCm21W/AhhL0Z19urchNvYQ65zWESZRdi6qAYlQmanW7gcjk3A/Ks9I2NtLc9lz
PXzC4SnBNZryTDTCHMBhI8jMAH3VluF9jDnvWXnzn6ypKKsQHFEl7MH6ufOkCrH4L/KdP0UdE+nG
+64GFWsVSAPjVMadhJLVM5dUtVNyYCIU/eCzs9wuH63K6HP89wOm3b+xDDoTL0fBKt/P81CKDDio
svW21ktwSIwmup1ErVCcKXjkXRjL3i+U/3hEeLLU4BqOSE0jpgeOHzGj0FNzqEwun0p1f9IQESBT
ghbsujXHY895zZ0V1f//2GW858Pvg6p8ar7pBSXEI8uq+tCEsdvsGu9conyQa3HPJRTDS6eVNqJY
bbw0Q2OMGypnxdNzG22uuvK8JeT/Grq7A7cR/3IxDP23/lD2JeeXK4ow1TEoh1uNNKyZl6xmHV8u
uzkvPthm5pi1iL7wd6mT12Cv+ajoVVWwg/2brxbcOhKDL9ZkFQBgmkV4pKC1/iwFMoGxV21F0Lv3
Vi/+4mkTjypya82b63ujeW6F19VXjJM5+WYrzrgKVTqyb3JSEqdcaLap6/A3tk02NFP04RpdD6NU
7ukObBDGbSbzhBsqzX4YiTPojwf4YKK0EEOpueuXCp3pKoYMR0sylytjvsaGDLJx9EuCfYAVJiI9
6FNLIW2sy4ndFAHKQUKEecU8Z6ZtbXE1pzyKNoWkXvpuMJ++k9Uqbfb+hnLsSDDvv9G8NW9BavzN
CUE1tZdFVRwf6oHOLaOd+9Awoeg4xWtAMKxwYmKW7bzpUljR+7+N54LVGDIsXYSnrqJDMPpFndFf
vkJ8Lnw45MldMSbAN0PPv248R/8WNflJHSyG5RytpnZqthUs7G57mpWcVLtbhVCfsOm6Wsu4udhO
qUvTotIqfZDNg0Em/MhAwPSFQStaduRCKudwbjrT6Wq3ZvhSpvKWlLTZjPn+aIzxy67VrtRmhRtx
LY1xTwgvKRwAo+Da72TYWcI7W7pi2IjZVzsx7hY4RtL6gYNxYlJZVWfrKh6cbRB3uIDfcbaOKNmF
O/L9fMDscbvtG6Axct7oI55f6oGwyLjM+8NsGDYNsn53VLH6psgBHB4rl8g8nflmrXpZdN2oYBty
7jdVVCAl+GAGLXTb+Dhh1Bh6bbUoIfoI00Fpyk082KMowQQDHHfXvABh0sc9e8xQpycSVE80jYM9
Dy3haXeqOFbp4356SyaRkaItDQveMlDzWwSW4YLRmo8glkTnJFESmPzrSqIgG1r6reCvjs8eAZ8s
6z9Gazy4l4Nr9TwUJUscMHfTMGiGU491+RS7Yj0wu9DFNTTaAzKjCKdN2lk6zB6yFucZ2L7+gT48
xP+KiqRys+VvWAs8UiFyASLAhp6r7woZx15u4EMqYcgJr6GbGs+BoulXFEN7Nofuj5WUYA/Y3VFQ
IiM1+4ww6gRdyIEcawp025/cYf67/NEsLx75dH3L29UNyCDaJ1Ywu0S74K220xqRxZbP5vXLu88c
F6DDbkD2jClzbIyNDS0W3Ap7nMf2IRHB2J2tLWSOqDwBdjd9EqzCfHF73gp3SH+VIcbdM9SMCcYc
PMZH8PoTosStRk0ePFTrgqNTBplbt8aD2gRXwkJqzh6cd0WjZ8bdJMRx9awdWPVn2Ec3cVuUgW9w
d9rfft6PYP1YXNFpK+aGBm7457mPL084NdHigA4g40HjjYy/PjBny/GxVmuWFlzn9awMDa+VEaXv
u9hkHu01I26jmw1wxmp+k9r4LWi/SZn/6I6RQdEp9GNGRHbdmgy90Y3jFAfmJ3q0kKLeAL0L93fi
n2281u7HZLgNPiAKVq0LP/JiLZaXrlcW0Ci7MNhxw6ZAzl/+5Vp88/opCO52ZodMpFnakQaoeQiH
R/R5B2aMAE09rkyZRfBzeiU8Fm8dqbtbF80vps5dmC2Cc8/34QJfZB5wWsCqRkMpiqxaQh18Zx2y
1Iq/VJwRIJe6O7EVDZceTtH9AbY9kBlAphOLcpQMZM/LiuiVf56Nkf/htOD1u3u/obwlkldCjLsU
yYo8A29LJE9GdMi4kkn4wVIGI1vpL4J1z8aHbVgKUGyyl/b63yBxNn+vmuGtnLQZSB8SNDkNurzk
a8O0vZGblJu/E6BhVxzcmf+nhvzxGeUmKE1/kU6ihuk1EaIVyt2gvdo/HVSDB5Pl/xWmxlIIbyAm
QtNtJZUggla1cKuRwdOlws0LLOCO/VwEIYNsT4eyxCy5G8lwqlgUPQcYsINQMxQXJJrvhAFSAbtK
UYNNkyLjAiVZyuIOfo1ne8ERb+S15HXpzU4iiF8IY0Zv5KIKU557ynSRMOndG4FcYkAYNVw0/uDM
WalMmqD0Ji32WMgj8V0n/d5DZXP7N/VIWdm/ujdpgyIuhHFlJhTEviWanTKZ5mTHDYeWkOaW6V81
FofMCLvFOupTWWqtvHJfpUQq75QcA2lwwycIzNRbjlPiwEVJ0qbxMOAimPHuuaCnCRwJXoD9Qpp7
HisPQB6pZmW2Z4YfDJesF37dVIdNWyWRQprQXCXXFZKE0drPaDeUKmizqG6JFns58YxyWNZhM16R
hVCfluDVT3DEyZc11dIuHmOtfsN/dByx9eIhQvGdq3Aip/ugL6SXtMZSJOksTBkRxk5EDZcupbtB
ebF7qDmoUtR+4kBvEk4UymHFydJDmhXqcxcHSe0dStbM9nHV70q0MjaC1ImmHBSo5XV7BIClDfu2
UpIItRzy8tvl0fHj9KBB8WeOGmL6cJbRKNLzmTPwCG5UVqZK33/J0moZMfMg1fVFsJQqP6WTXU3e
RLKcp8go2ie1dmOTHs8T1TePcNlglc8Cm6HVTUQqk87hNhnKykGPg8eTBuJf+bLDQn52K0h5V/Sn
7sIqu0UapImbfTWL+egA/YAEdKeGz/o+KrU620qP4APZU54y7JcEpqSAji837rHUFaSSdWzAbKtW
A5al1DUT3ojLYGdDs08LmlcdTcSn8+Yx21Vi/oqa3t9Cmqdt2EEIp7U4VoaVyh97oSklADPmE8ko
+n79eOEu2ArGriKwGBxbY7eJf7PWqS/FyR4ITVhxl5h1ewUf/lhaeF1nEqv3f9MR0P3MArF4XiHE
IR1Utfyl8m/8Nc5AiQrMcksxafHGYVJ4TzrJggyn89ldkoW7t/qbFjv/R1Mwe0XLt6BsthE3xwyM
4iYvG5Y3R1p+zcyc13g9ZjfwGztO3a4RQEf7NfO+yH3xjojJEssMcmUA4aK3CK+WK6Rmy4uZosau
2rNz8LqCMDl6mmXB9SYcl3a8RJEvZ4ZyEVPre2EH/kz7ecDkjzYWm5oFs/SJe+rhPr2xxPo86NoK
u8ezVjYgVpd7DKKN8RzAfqtyt7qosBtkYPPyPWkjJYpv0uH2oeT+ZCAy1LpopqfX+Jdt6MSXmzXV
qq0fG+rJ8ZW+YgsuatoExyF3NgKa+erJovgVfV1OqfoqFY51bl0jkqCZ9B8M4gZTUBnuwJCQinlk
/3gNjiyyBKO++KJSiK/ctdryijUyntm5Lo90+9d0DIN5FZhVX/Vx/8lNoMcGn9aZvkLP30sZEf/g
rKAPI+u6u39eberIV4hfsXJgi8wMGYlZnVpupQOsyI7mcsyaUijSfOftGW9cZJ3ZxW9eW0dqXm/F
sv/ldJR0l73M5R5oP9zyEtHlQ1PSQEIy9KsHjJ5BMpDy07FsQUoKjZQ8HPgvume7AnnMwKb4aMRn
EIsoJWMNAjpAH9sLQ2480O8L75jeXUX++t3UvKdDhW7u9CKUbJNx4ww4AxMBYszSeeB4EkXTXCV4
V9eXMBooB3FaIzcGcUZSYzUqWGy8WklUKCKKYtP/1a8pGXur3HNvYV9syqeUxKUVr0fVRFm9bc10
NC0HLhwufT9T73LPm0reN+PxNQnZCrmQNHQ1R1gOwkc5NBOOtVFWggVeP86WeiM0wEERksELwQgh
AyS7YAUbZVEcDEnSV/RUmPIuyxbki6Vsi7exCSSb6rMl7InumWhDeaDXrQJM1sYYFyzzXs9XFwYL
taXh/7R+qwjSX3NuW/muTHBin11SMKbGswFPwKZMGNUmMI5uBISt/ZSZ0KGgWYyVzXZQSlXdbaLm
L97ozP2RGoXTv5UKrHCAZmGAfql1Cb8kUaKwzY2YlAacic/vAXkQzzbgk+j2muphYllQblut9kOV
z4a4pqegO2uGvC0eI7GYG2RUauiZjAKn5EHvKsVB+RVnTnKfjxKMcdiiUHfe6wz4tiGik6X46BsQ
jI4/ir0xgoZ9aZ0KQr5dIjxV8E5YucOQunwneMT+KBuzDLoYyHS4aB874ITrrh0zFswaeh2ARoGz
PTu6xvPMJU1yZAUWbOYm15ldvOzCoA+KXAvAekm0l7Ma7daE1UXGC26t7wVF5//ZbLhPf9C7NPeT
OP3YUeYD+lXalmeVgDzRlfGYZrTbC4Z5XGZa3xzIWcdCAWY6mHUuqYVKP+x+9d9mrjXzbL50fjzS
T72v0G9ZC8JN5ln/b5uxrEcSoQx2ZQlCTN51GS3kQLAdjjFGxf8Sv3LaZF4JZVgF+vU6Tcxis5YV
UiJUDf6SjopLCE6sImJQTnk/3rnLTckezqazYkKOUNF15VpEL1831cMof79jfwooDGTP+aXC6wG1
tD4AsImFjnquN2GzVqJjuF1JoHkKooNB5kuPGgtZ09d7u7M9TmltXfsZYpFY0mQvhyYvq/p6bVnF
ES6yMunXIGP/AosepSe6KXIwAMAgJEqy9X/GwWHF/mvj3cMHsocJP4t8riEnyq4OMYOp3NhSzsHl
8DjK8zhyc724Q7kZ1GRysyDjYoOz1nu8vLSJVyHSYrqtlkGAZIMYk2PpNs1kkAw5QPRiVK+IJjfX
7NyCBYaWHD0YVyF/t85PgD0ePaHyBX57jVG1ItRLBv2ujuBMr4ALJRytJ5F6aMqB1wdTIPpQGQl7
BqtxGau/Kl4Ca6/MvPoWNwVNinkRx06UR/BDB/cQ/9c9OQNioz49mrzVHZaO4yHjN7ofY9zC3RGq
Q9U8p8tBTUvrVznhFJjDm4vJ3g0Hi1nPMA/7U67CwlcSo28Byu2BjdCa7l00UTjRggEsZMx3oNVh
xWBJmWkUKpXBvv2/J8eGUFvJ0gxwm+qETW9BSbSpW14a4oifoHen7rv49vdBxIy72v3zFMXytyiP
+SNwEC52qlq9rclEiWrI5hwtS9mbX9paLk3BoHB9wsyJnNmI2G7RmTvVRSA1h9ruOPbRdgVnUA2n
zlHmGLeGV3gMcJvfnqYJIN6Jg7e3m+Kx+1gMIx+XDYr1SdnF1Xl1GI99z7IHkqcTRRdWRofzpY3p
3sPaCHC3vSyC427j+t62C7P1QrBtpeUidzNQKaDmvT7psa8NoMaWMBdwHpfhGBLIYy9MHERsj/OB
9jUtMn4jXdOPehCqRqhvddfg/WtFiaPusQfMJ6r9L1vOlfqcK7VuNeazV3uMZvHk+vxvQfb+5hCu
3E3ZbBy/e4HpjMNOgtQLn1PHVqzsoi/g0A4QCI+h9QJhBZqvkF9ivUT4VgF1Q/zeJ4VZOE5Mdrv8
6fRTWrDXkv8fpx58AJ0R4rdLVW222VHEqbE5QHAbIkzUcIkaiKycPyjOj2IiIv9OcyvQuu/Z4XcC
K2fINuDj2PFZq7fWlFTXq1XwdgL/AvUpdoQeB9ApTmGu4xnAUDmEenGWho//N7hediIQ5fE7ducF
vgiVBjdwmWXrmmvtYXMVbmgKcOWStUgpQ8MV93/SfSuzR4G6TEN+8ZV3WYZ3YtZdZXT50dMHxKmt
MEJIVA17s1PbL9QOy1kkwdPvQU6qG8nrohXTOdfBDaomIW+YN3CBC+lmeUB0Kxilc++k4olj6rif
7wDFCbf5kF/LM+igVwMewkPdCCq+UuKpxLdL/UQFxa0p5XG4BoyuAHWjkyEZCfAlCkHRnmt0iaWI
RtPt4jztI1pZ0aX9D5x0fmUNRHTmM/lGn5LQqXXmQRbNrCygtFAeQIKfWNXqJgjGMWaA1u/3Wdco
mCD3aAaIKmv79Nk8AcsgtFM59IyNvSCDg0s5dK8f8iV5wfW9xx5X2F6QcXJHHOCcAgLvRyk2uAeH
y2lFlTqkpv+PXaMCZBl9qUVr5YUEmvLE5etBICY0d6QaIEvzMhp29brKwsPU5dxn5Aiiqh3bsI32
GmSWLY5WZT1BuqNyRqAPJuhO2/Q2ngHBU+k1LsjxNBMbXGPmoypyQdxu9o4V6v/eHvQKksJSaSrC
lw9/78sNhbfJFRMPxlZOMxnPX4qY45ZQXmRxRqlvfMrXIgCuKBo/FyviXnVhkpLbQ0uw9DkPJvcF
kGZHFs80Wp0qyfAVa+Iv6bEWRB6MTCO0IqZW3PWRwzA93McF+dyuHV+nElabMNxA4qQ9qfoF6LU4
4g8OCHl0gz9VtXRl64xPbDg6WC61C4iYz1ZDUHCqDrTxO7aqyvZS69BuuBab6bHrPDRWB+0iseLG
8JVXd/BTUIk/x0+DRVS03fRJx2CVR2aie67Va7g7tWVAL469cs0jaUHtSc+0bQuAaVKNgidSCXfs
zxaaD565v2GX5DHYFyu7GQiSjuw8OWhC9Au3CqmN9j5swCuwp9/pxH6Gj22M8uCAfgsduZdoa2oI
laq3v97q9U6HdTAtgU0jvT+85PBV2uN6nU5h4undf1xunU7qSxPKWlLVhCTIbPY5mSNwLTB5NyQC
gLjFb1f4798jXcjlZog4oMoQsFRbEoISbdKBavOz1T5/QsJJfnkg3hxx8W3RZ2ksfonAuajxkgw5
IKMU/WHWBNKBK+rtWgxSAL1KvLgHsDx2BfMmIpMcN663GAi16qx/4RxsCxRnwNIh6EKpwWsDmWjk
UFGDGpXJWSGiRFxjHFQAoucq04MTjBjzuVeeVMbkaX2Qx/Za828jFYckosxSi6wf6TZUHBz9zpx5
jT8GRp95V4Nadi9mcqeOTfDHoeeW/Z5wzFbTreDl5COdOz3Zy+PfFGnYrk5MBOJmuMSu6ayF/XtF
ed4MQT805iwyJ3mrx8anNwFO4mN8k3SHTTbYmDSmkrOaXRgpXl8IWuMrj6ks93JJ34EHVg0f3jCt
LHA69yL4T7yY62kX7Db0twChbnhkDCayikszs78YeXZXShcMNAM5GRS58X/r+Bu7JGxR64mUBFuX
a4NN63+ilAjXd9uXlgPjBAM06BhmH+oJF2EGPIt6wNnL/uhESTiIbqM0IxiAqyVWXUlqTV+w1afK
RAmJhkkir4wiIl6TKt6JuMWE6+m5MiU9SrdpDLvyyd9C+MMWUTbTdDwuMI0A+n8=
`protect end_protected
