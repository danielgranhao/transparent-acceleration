-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LKybQ9O+P9JmxpgN9HTQ4TwaRaTjKu3CyFdxnJxmm9tjLW/9zkpkOtRIUZ4RO49/6DA4k8PxZJkS
q8l1BcoBQyCf+yc5F4i+uC+BGB4U2UB/vDwGELSclmGQZqJ0uiMVg1gc/HPjOHlJCe7kxCesGo9S
D3nqLIdJuWkVIScdNMUsmtqJRGXFwPYMVfSG42nOsRj6u8BxSWpN0d9QoXF04YziQR7sOwyIZ1GL
oAjf3qf6OcU6efRkCrMRLdwfwnsTTaDB6OydGTeJcdduAqIR5qPRYZWeywgy5GhwOkf2PhxPHa5i
B7z1ucwMkkAwEPb6SsCZlDuan1MkSePpDhawDA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 20608)
`protect data_block
5R82zj7ME6FNApRcBrUIjQY4vaqvNg4q++4iMLKXA8sZ92y00kqUjNxPp+tTEqSbZGOoL6bp6mXN
l8FoqwyTrrwM8BA8t3/WGMO2aRKqViX0gd9RJ3xo69IBpQEaNHH+MJmPtJy5xeCFa/BiJrl6YHXs
2Rh+rmVmccdqzLDiV7oIzQsaWXVc9H1kNcDvqs//jLqvVsWxNj7u7MHUyGILrMGmVprtS1IbBE2T
GrGCdtlNIMcpaF/jFEQIx9Ezh2JKklOgE/WLG5dj2u+DDeNVekq5ErYd9Gmn4GGAW76I76KQFGu0
NCxOGZeMXZSnsAL5CiY4YggYwDsUyn5o3iJvwUzyu+nM4TIlWuoqc/CeZZUi80JEL5h6sG258I/D
Mlv08l1vTZSDuziaJxmP/YhT0DiYKNNVU+JaiGMU3PF4uC4Vd013GyJQ1HOhOluQLMy3yrP34Js1
lxt2Q/UaoGF8IdHJNJUwywLpkoA4lwJR5L8uWrTgg/ehbxyXgUbCZrztBcbnbR9GMLCPU12HISM4
V/OzBJEINjCeeot7j310dmr+YF4+0io3gMQlKn4w4ouCA8zfzyQmFWyYJPU1PczhXQpBgP2vWOEG
4eg87UuTiSs0Osfzwz3nmFOny00NQJ32b5nFqUpfNh12nTY1ZN/Jzp+FGdMitCMqFZIHJKezp+Ds
gRLpWFDmbLFpQyaL18apBbPWn9wl22Vv1bUsG/ZVLBRkR+ldZuC/VsbJj8li4YPHn6ycwgmkqxll
si72TEU6Z59/zjO5I+S9RgtbKvhFStJesl+Veiovr2tyZsW57fyz8wnC+MvZN+o/qOiTUQzB+/yZ
IqNb18KziWJgh7zITBWk6zmofwCpjOfpCkOYlKYtMYtBLqaeXXWiSXXeVixlJskGsuPho4Yxvz+G
dkGeDNOJghhptKI1uetqLkSI5B1KPWStv3afOstRBCEPhd04JdwQk0ZnZpuHUSPw1nV7eo3hCrt0
BaQK+LwmSBQ8+0hl/tG2uA/b23v/4IXNP1Co/A88DS2cKXvXwYxDOeOadErk1IzK5R6UPePTL1Di
Y/+V1W30ZspXg8OO4Je3UgRTQ25wfSQx/MC8onUSeklS5swySna00fX3VM1fXqx8VrIFD0XfNmDJ
nfwOsKDqvSQG7BY87t1FHjAUmlyg5GDiS8eCfQM8E2LM5j5uJMBAJlYDbofjn9/VVN6I+Zfajz9j
vdFOBPD5LfN2q6Y4ZMueCK9jGmvTzl1ZusmbIBEZ0V3wBMeyfseDQwlLEYe8cOeWx67Y5bf+EWAN
MsRlB51jyJi4KH2JI5FDllTL2rJHXnF8D9n+d2dU00I10WAF8YSdz+uDJ8Rlbq/Z5GAL5o2AnefS
+NDBPHPOKhsuVgAooDCeZoiG/la1Lq57HzHZNgXq1ffvBlpQJLVBqvcVhzRenCMf8/KRIDdjOujB
jZOLDmxFPiMMgoJ6QsC8mkvQNBOGP2j7ZR0MlZofDlrQvNVKirc7W6MU4MwsQGysLdssp7+oaKmD
2oKPsjkm7fGyFMkptW+co+g73fFLE+lBqp/AZy5oE2et+23+rowZzXUuVx7CIuWEhv7IH6mqaXWI
Pv9tJlbG/n2qSi8eOCNXbgDCrMLzFpZMjj+/pr3LVgBRwvJseayZyqMbADhWFje4gB8b9MeCqhDO
aF4eeX3AcPTrMdXKp3RsnTLGJM/22H3AOYpawoW3c6cj5TrSUsmKDthXpy1cgXbLYbdT90Q0e33L
eFuV5HRUT/rqSuyslnBKgUA2ObzTxS+JbXWyJDLSVTGOeduN48Tm1gTr+rpPr4ou/4x3X4J0sJWK
puvCruDH5ELhko6hRLHmD2eSEw+zuTUVatahUUVhXNDDKzDUGciNM3UqB+dY087D2M0B53ubvgod
h6RWVeEqT6MRALgLvj8cxE3y2MrDVZQoEok6d/ddst3AJIC8jTpJzwkFTiOFViRRie1bZ6oFz3NB
hc+1mnT3JAJO9sunZ9dZNQNNWW4h538Sf24FVoPo0YxdAzQjjGB1kJMPBjvKj5M6BQiotuggh+az
Ju4vmmuvnBNV7oCDPWf+CAvClFXMwBYVuHV2oSkX/IzAfk1/VBhvVM7SA227+YNboN/AqiMjXnf6
l9cnKQdYTQzFGLpwprd9/DyGuGS6LGKETaVKL1xYk+FGxv3/O823SPGkFFXT3aXYHh4tNrQRD/Hi
FlgN6aACBPMzCOGDEd9K8DAmac2U+mZRDVFBiy5oSBYoyaBtfkcRsRA7n3d004EQ2iOgc/778RxP
k1+uV9G66asu4Kvz7ac4UG1Sz6rCnf9kghxh4Cyc07RpRL3Thzx7LtwBSmQUdHGwT8TyLpZkaPA8
/vT6YcUMjEomkTNnoWaGHcUtyGxcRSq4+3dtOoz9uakqVVarr+LOzGuI5xWDG1xKQGZjzn7CW3TW
iBJyg6dNQdQ+vAfUdEyD0QtohGIp0wHn3rwH3NbwvCxJRaojZ+lQyIm84aVJIJptjquzi/UucJz5
1bwguq0ffpK1YsDvPLfCnPvo35+3mtCZn/DBfhNi1+yS+iZhuS91I3fFIpiRtbeIcX/xnjks6q8+
ILhaYXyQEjnDXphK89SJs3biLrPkeuJDnzvIt8PfmycS8KkgHEn0BjOsv8VQPIASVUt/jWVRGJWr
abiBbBDrMvNsUpMgia8x83S6+ikW3MY3Q9+zIiqU5OYJNxL1zkxqIbR9tfB0NZ/9Klf1eJ+08piC
sh1H6V2jGyiDS3NVa5FlkiNkkXXbJVW6X77lDPW3viOUKd9ip2vIgfaBaX6zKPxn/8ZbNmdkx6h2
Q/d3UQGSrirnmNgLlsZDpVv3bLeX78Q6p5qNS2nPfN+x7H0oyxLks77zUCzplVamWH9J+bpzIhpn
8H8tMaNRaLrBtw4iPE0vFlc7y9ZH7CLgShtimwHWLVGjaQJ/BHqsV+LPGzKPKGLdzHGUgJnQmKOh
evPpMlJqWIexejyLkWTVgcHUFEK1bTZSUwx62KDsDwU0VIHAWbwMp7s6HNFReou2TYfFfwq5/JLX
PKLimIAu62TVdEpR9b7bvCELrTugkHy3oMnTBR921NR3r/wTrtDuaqmMm7a40SapkJdwjurFDCNl
7YtDjgbDNaLf5tPmD72oJ4ymVlCDNGD/LNeWQJAmsLOAP6zW5XQSBACgaFnk18utroPi+U+2ai2n
sTEesSqa5LLIxj7TdLjYDI/W2d3J1vDdOtEn0+Q7LzWH1hz2p3yTsuOe8uym7PP5UQCuZwnnQp6k
069BQpmuUKfxzqM2NF+YP/xw0CEpdsX+vIH4tJkpmvSapKhOQhRx0Z6wbyJdqJgeI3ClAq78PdeZ
jREpQupL5UwRIS4BsM0qnEYMp32cwphWYh8tacE/SgqqpAy8Lh03LCqxYUHNNaNIQTM5f1/HLHnT
90sHisB3POdIpN2daVraDwWZZtSfRaveXOkOtjDb1K+CnYnn2grkKXy0l9soJnon+fTZU5tVC6h8
AdYp5TjXwWCBvAxuzMw0NXgf2EJMxzBBF9NZipULPDcr3wdTNkhNSUmVz9ahlcZNLNavgVyez6SQ
MzcDuTF9tjqKLvH/xXXQoDmF8cbi7mkoiIkQF0nvHn1KrYjfvU9flVniNmFAGEcJGhQg//IRUbRp
5Hrl3mObQFOfmqeUL2csmPxdird4lVyJN9uptVWKnueLZNolftioT790xZHQ54Qky2PdvAyqkQes
vzDj+AQEp29asZsGZGlreh+kFerd38s+sQK7wOch6qvniQeqgA9ARQQeHHn/CbcoouC8IUluX2Vy
oBLry/QpKwIKnnXTVjkBeJtNXnJeEXGsuCF3uaU5So/Ji7s8/Qyc7yKrcZlwkjwTzR3YFlgmGffj
OnkWodNrF/uUWeaWJW9M0WwxILXw792c3UraLh+nU2ilCeZCpWJ6jiZZAg9Lf9n1zY/oCUkUgg6S
aOgpd7ljZDyUBISPznMuCr44cwUTlVjNX0apn8SEOaZ/2Zi6vl+FDOJ3bdgqtanPvsNS8OaWwiq4
IBRRv3g6AF0CtdVLwqWCUqPO3LjBl9BzHH8+DbFkDojCaD0H1fS1mf7k6Ky31ZIPdnxlr7gqiB0G
u0Lz9WRbizHXjm1DgtA9BQugR+nz4Q0QyvXxe7i8mb1Z42rjedlj8aDakgSZcMMXR3vUhCGQPAya
H1/hei0c5e5zKzvp9zgjTSlHPZjXXyFVytzdjIgWM4d3jvIOgbnMSkPeVkKCsU+bQm3m9LrrpWoA
8gHKVQkoonYxv2IO+c55sHX1mXgalgcwm/P7/BF9lCui+8r1MeK1TmGcfnxHzVPMwb1MJQspopGx
I1hgSGk+qlFJk616F7+U/94jIy0E2PFLYAWVA/M3clWci6qmOs7AfN3vPBE9igcm7N4a/aLmRH3q
y4oWwjJWpKco5wPanhxDMZoFV1xs4rhv8UtChlekYCi3mqPvjLbAZM4OnnHGeNdA94TV8TbmrRW4
iMO24klNp3HLj3xCqCthz5AnReHtu3C0gDUH3GDOnbniTuvicQUwhyGWlEQRXSMxf15rgrremfeV
2AVGPiCRwJK+//C59EBRK0xlSuw3f1zf0OCXRUWewNCKZKCuu9q4cUVYATrQT4sX8azjgO1E8lo0
XVLVvaDzoViTBceFT219NVuqzne0lhYiC4ofrwvQ0kAdBGtAaPWe6DMx0L1kTB3hz28aFM2nX2ZS
RdvKqJcDTIVUxlJj0kJfisVAFHHXKFmcYhQnSjf+fNtElGN2rHu3h8S+bIKzhTIWuz0qRQK2qg3S
HORH+mhllZmrQKFGzNp0ytWMMmzVZbEBVDqcUh1L56mg+yDObNm4zYe1N1tgwD3FICh07FVMM3CF
kT5D9tWP0c2BRpQa1PvSG2sEUuZRM1mFpejSrotvqqEzI2c1xBgLpbNTBv+x23sx/fLBTIy3nv7q
WN/lqmtQTwaMFXxtTrZFNloCT/IDtDTN+PxkBUYpnh+87Jjyevx6s0YTbkHQuzrg7Bx+0N5Ms2gB
k0MG8uyXmI906KPx5k1CA+SKqTNPCg1ybvbOkVimBDF59NYkb0Y19nTQQ+TEb5jLSuVyHnn6SkCx
rItMJfH3se0AtE3ZDyaJ7OUaZow7aDCaSOwDEWOc1MtjcohQ2W2IcDPsOQp5StjNK1KlyLdY86KT
yG0NK7wKP0pdal7s1IygQEAgnXOjVKSGDEi/scisiWkIozM6en0FxmQNklIVVOk3Uo7BwytwUSIJ
wZprqXqJv5Em/W0VKpU/oW8+5OeUbQ4iN0Auz0OxCl49oDFf4CMkfIoReAruhXtqxO3QeHz74Pr1
7pUN7OPY9uSeM1YFerUGLUDL6F1YRxfhV+v+zxYeODUWGL1z+ihHXSfmSSoo0ALiOY6trXJZy7h2
dvr05Sxlkrqz2U4Zes8FdHNZTM60zrolEyT7drMipbXu8WBJzk0UUYjIjYnBPDbF11eCetanS/Hw
nl/iAjOPOQCaT7UePlg71SNLsmnEpgfsonqNu4NwiqP27kcfLhNEmqnZtrZUkIuy3fh1QipcLMZo
el7Qh5P9BkpvKfZh6ln1Q/JU9/s+ZQ25oVWVZ63Fl95l6oijzdDVEjkEkxDpzO7vH3Fezvg5hqml
WQq5BxvA9yPH7lmXcF9pmBrkLqLu5J9wanrc9QsJWxwPhVX5gUw5MQOOx6IN/+9Z9/CgkYC6vrO5
ZbX3Sre6DJD3C5SMXVvxSIr5uviC/7/CARioVsGlsq9nINwULaEubFzUFClCmPSBsylHyXPcifRv
0DrTqL3uI6jwNQw6/qL85B0xbhqtq/z7UXKx9iC0Al09RVbwY9JNTN/uu7ztqIUOEuccdOfI9vma
mo7d8LAq2mwHamtTGwT6LYsdiMVQrIU2pFYA6sP1LSCDjP3KHL1vQwPEk8/oQjYaVo7fm8ni7jdF
hge1o03MRXZvkfTS220TfTgs5PAvKect0MUXghQ4su9fKFGg/98qd5wrYq/uTHC3rCn/LlIJirNT
vwSg2VYzRSQ0bmfIbA1VLNQYAB5jUlWNWZSfOGn7YZGtbYav9VwFin2YLNgbdprAOtm2zl2MI97l
EAeNWit/M5DYw8Yoy1EZZdnejEmeY2jf6MRSctt8J8cwchZ5kE3aZfqvtaUKBS/Nzm+N73q3uu3v
H87aqTRHouEdsnx8qRn+jrIy7E81ULasIq5GgmIs69vkSJKPXAUsaI9DoGqijRCYg8bIPd0ierTO
oBapB7h3FuUf2sS+UTOb19yX0XAcq59gzYumOEKXusgJrkiKLIfY18AQXpQNwqcrJ+rc2ieSc5g7
m+06ya0LvPBkMgXLCXYy5eU6wxuEz+Hsqc7sR+pNSy6N10Xhtws8DPKbdYdekd/UUw39Glgu50lv
vDVEXVeuiX1dfxUdI9fGSJginWQK59DA6mPym03GiYb11tC7HhUPPIT+onpdpOnyTvGVqcn5ZHiU
gcuYS8YMKTH7T8Qw9mD8HUOa+Jqv+i43qYOMyTrCVDkmemjsaDDVOs1HNF7MNkdcOzjbsbzHq2PS
ItvFRSXArV4ToPBCTKJdI+qj5uwhbk95OmkbpSmTPJ+aK3IEff4+Qh+dYBQkTEUfsqTLJ1WCE6X7
HsFAcqRY6M6IsBhfjYIlzCJWS0Lz93HtFBFH85qdmirF7s4LA57jAjJ9sWE1VyBkAWQIVmCR+KyD
7UTj9yiCbMXRnH46+Bj+65q7RL2j2N/Ix45Uw3juEEHWNZxqU3Af5cXtMjKQs4JXmOaSoP0MzMCe
rq3rlf73rlHLiT/2khSzJpaV5Uvnh7aBK7xWISu5YLiLuoWXTfLW3an0SwkMWIODGLFWclz0+WLl
KgBJzXe6kDfC2aoaeS80QigMC8c/0wbEwyGPbpt46+iXp4IUspjqhB1M1czwStBjEGCBWyPzY8hK
9vVcSKyv8fRTGabFH7XSIsBbjkI9kokM8lEAJP1EA9JAHgTxfWsyIRWe3foj4yGs1/F71AZYeyD+
azglwhM/CW8Q9HzYfLje3cU4qoFEVDZYAkZoP8U5WFy5CpYodyXEOEXZUU+8o8PcDSaYASLytwQ/
Gy+qfo5GaDX5ssXy+iJSqEleGF5gGTaQD4SbXiuAHo6eb3VGP4hE9t+Ci3PxuM0JoLP8mawvtgms
DHJ8OMcfptwWGf/zKyWOYCZ7BdmKBgif8WxoZbizO+n/0c2kJT1s6S1H9bQVblGU7oL7wGtn6VRP
fewo3AUmhqHLDlq9TNcpNpr4zco0opBcEj3S85ysc6C2woXpKXRD2etd59T3AaodnbpgORjiu+EO
ngRDrJ6AogoB92I9Zk+CjkaCurJsqI0DPja61ttTBl/Ys7mmoxk8wRG6suC99STP22clu0uzbNOg
rVwtczM5838wYfgfKs9pVUC8iZfTvycuaEekvrVoWFdmWPc6cnodDz54gYotS0bQmsWMQ5EbNJGK
aE0I/mKgb+A8T3x5Ce9qdc3nEBiTZwPx6NG1u8fy4twgxUAcXJ78MQHMx0F94OwW86M8UjZRhRuD
8f9DKsvZbRy1mKkFcwxGu4hkp4xI9r+auFHtQVAIhwZx2Uf73edW85xNmuKgyZbk+5QR1hCQZ/KU
E5COLTjtGkxRT1V3CN+OBWJDspv72A79fnw9nBsM5eqH1s6K+TbLaZB3Yy0KRKIkv8XEusCSfno1
CIKEGDMMDaJKofEhyzcWC7ScHrRBuMU52ewNLNAhwE7/x8UQKpQ2rF4v71ZWwC8ikvgAsGSC8un4
3M3OBOZ9zNtQbw9EAUj14xBqXwgCqP6T+cHiS9DcKSKRFdcEgtaWRPG5lI5X6fGuSLECn90hiyLl
XN3LQt4TnNuMRfa8FFovst7/yO1YKPnU7cfEXL1638GvRwkXc2tmLBmW9lcmeJvZkNN/FTUx40BY
4ldPRsxL3uVzuljzLbJQ+l/M7V+ZgvgmbJUOlRsHjVvj+4qFf3hszIEefqvYFChCb4vQCm9WS0OL
GiIUNLGAsb0jLWZ1OuotQ0FRlij0qFnyqMg56xwE2GcsMwrxcpu1Cv0RsS5F4KAGGkl/u3TmHeT0
ZxkMQ8Mg7Dp4Ys8iw9eAcjsUOXAEfyU5MceB382Me/DFHpbQ1HV7UZz+jGgnNDPjoEIDVGKofKWD
kV8T8F27sIkiLshtE5yvoz3585WXvgvzQtQmTSHnMXR1Qol7yB8+0IXTbhtXyb4nLWvtTp4cgBON
R3d7KlAQxs7xDuEnkiJwOhc53X+ZZDBtNSbSKSAthrJObzBDs8E0KOLQLcJ0BetElPt7OvQFWm+G
ZPrSbSSdGIfAdsXz0aBzYAKDNR0ss8Z6xHg264OKLVLZ3Np8dCvD9V76eq7Hgb5s1e2EU0Xa9ejm
moQnIFP91B2922B1TZy6coqtF5P97RrRs7SH0MFfwL2vPKW5I2+FUEZvj58GyvjKo0fb7rJZatMR
SITc4ggC+pm2VT8anhawTjybrynmqbOq203O29I3m+HKNOZBZMmCI1gFJWnbnuYrR38ZncF31bm6
npb1/a9eyqGpoWLWNLq8ujFDuuYsIUq0QFY74fLlYf+NagoeEfxOLxB/3Ytl/p1Ddj1a7aZ5cdMP
UgDThVZ1pL1jVUHB9riBH4eRfVet/iWaAQTVxCmLu6RH78fTUsVWUlCN/+d+A++ylPsP4XhLZ450
D3UCDnsFZOgeTDUTtkPLBKE7gebaqnzSR3+1O9AblvukO7RNVguH9PTMQ0ghV44jkcX9KkxZa9bF
uqqBS8c2xdkjaOd4d0aRY+wSUIZCndn5pIWwDO8N6rkL+u7QNaJK0M/WiIQKOOFfWV6oVdghUb7X
D0MwfKZ5AjLQIbeTB3z7e1twQdSBFwxF8MLJ3A/XbmJCcvv7xz/j3JNP+CphzPTDV5Ln62sJAfYG
opqsUG25vXOqbQQqFtg5b8+r2tIAbEyamPINPtK/JAH+SztqfihUTMqSIGOBWhPv2Gl0JHS6RajZ
o1FjTRAnUkrLr2kG7+dtydK1X+q4yij2jTHRRCBvGV4V90csVYSkZfknYyaq37CTiL+0+3KQ+nAp
UBKpKaOvh6jYC4gwmdNbHFZueWDYXWKxPIeP6/o9DAvQ8DlR2uj2skq/MOT8/X5ehA6sV3rhXCtT
zK6afYlTrW2PT7hEbJ4j4dzdvX/XSaRycHpan5sNwVj2GdMsr1t/Z2UU0ljfeaxPmBEgVrxF4/nV
RTO1ZRnbLhxj3g/XWOjTBQBPTlAIbLw9I//OgqNnrm/jcTIlA6QBs5aepXkoCNmlQSzeKrICu7uH
8VbI8LW22LSCYUVVwalYooBV7hNu0g7yS4EArQIZqm7luwEfE8uz6xHxUaoRL5lk5q/3+GRXq9ll
rF3i6Sm+9ub5BlbRh9vH2qY/X46YB6oOzLgXDNp0qlT1vWY/2DAI5YC7P1t5MZR+glYWXJzn45oU
9lNLmkDrta0YsRiBq8cHAqpWzqB/+Tmit8RY1lmtGDxieIBUmk+mhRqHFf138jyZpqdumvrArLDH
FlTMX5uy/+Ev4Cf4GfcJFVSv9zY+rgMhrrQhDxzOrHJ9Yv447HlYwzs1Smv91qehPkhAVZ908tY3
+uEMTV+QU960cvZBSH7c/joYFv3k0zuThKO27LnxNbsDpg7CFQT/1VoBzPCQT900CZrHTRXRDopX
toRQepp+ZLNvW4B6709SMx9QGQW0ygH1QBbsGBb/AI6Q7UavMlt+qJJlbp1z6xhO2TMUgwDCvAvw
jo36/PxtAdvLwWMMaELRrC6p3KbsS0CRqPoXemSe6MjsH5KOj55bo09MngJoLfn0zDp2HPCltNSI
zzzoi1D5XJHoiDRkje4kjECkbEPF08ktXZkt91c3acvkBpId4kXiAfqT5hLMQghto1PvZWxVt1RU
AIBNvBvSeJHA02cbij7SxOrS+QpcZIPIGUQ8cowL1zztOaXncYCQi4GPjB0VumkJWzRGzBuLmqHG
+LNGPyiobeJCxxsICqqAUE82qqXNrLfV9FyauHROjMl9UFtlI/12FuR4K6oF9jWTw9GqYef4MfRt
7FCzGl5DDzf5/6ALjwACbwRG6AJYeUKrGjYaSdPAeOSl+GhIDhO2K98kIclTqg63JkkI1oI86Mp5
e0XeTO7xGqbMKEdIpzhHOt/pbZZrl9JoyED0FleaJBIgDK5VF3Ah7allboRGCwWOYSggWHiFJzAm
bng5SS2nYfUlbU9q/qo3d7JCU0q7URKPmLAdrhu+mJiCFPANFX+YoXDVhCufc7zD0CQ9kmlOG75H
UiYobScDhHO4yH/Ekb/p2sWRqBzMEQmXO3TP/LrjTuycdVTIs/r/Po2Bhe2cyNO6mz6yJz0LuI7m
Sfk8U5GCnrUyhfz6LMunDCZzDNoXiQgSpyDFiODTm7eCOC7fjtvT7k6g4TGfOCQBQfpHlz66fTOb
9++s+N+EljdC9rv2CCbC4xL/CLsTj5g6ajObRh73ed/KaOy2Zoh0DQBhwJL7NwhEE8f1nv2CxT11
SuPoszIDCl5RtnoEoTffxGuUkusXQITVUnTOeoEQ58kPXdn1pL4frV+NoqOaJojETxDT3EOTKyxi
Mbi/KrLE94fSwHZXOS8pd4134ApyfocaXa7WjxALfV8hS9Vp5drw/+ONGok1tfXtW5MnLcma4gn0
QKFypgQkPcpuSrlcO/wMQk4pq42QJ9Vr7Z+1oUbGlE22RyEyKIDhQRAUS5XQMxjmvl77/rJDw2/Y
QrcfJ1i2mJ0CmCf9RQBr8Vrsamq6igERQWtk9p6smNGuOnxU8mmZ3o7OCOwMKmjgZ89dLjZQJOSz
pSu398ahfVp8kMvbDZxxltBVRM3ilTAw8aNqZd3Ss6srnw6a0WMCuiC1ayF527OGeGl7sq4nFI0Q
kH/FSKOIx7Ar+1aZGoIg7KKqXz/kFemKW8JleghENLlvZw0xvjeYBqBjt1txmQjzJZIKmHPXLGfn
J5mSAp4HMqeFeOeLG0XkbBz3RpBayUpX+0sZ8+gnmTziZfxfZONVyRB+Hr/zsdCPYcp8I+QSEnZg
AbehTgAKJQrw1OECQlcO6qDtcjmrfG5/rmVR98hC4M54SxAAIAr2UXqwvR9WDmVTOzPznhmz3Vjx
ZPZ2fXQ5s8wvcjmCwYjies2Ftqvhp9z8m3EKfesefSo0NFmjEm6CpqJcSjRaxA9vSnEKIA8pCAmR
qGJkzgJD3GRJ83zjxMTrRR2Q87ss/+AJAq9BLr7Ce8uVRRspab6yxq/cXw1gqIOsCI4elAARnoP9
yobGwbWdNz58uJUjNIW4McqOjQFTvuQqexdG8UEPHaqFwKUPhO0HwNY7JfY2fEdWI+vENfmVubyZ
DKHa0jijhs1Bhpx3X0nOZDSXf64UWbAzUWx9UzlCLlJO145VPHQl/w85MxQ6rhqOIjAsZaVCBKHP
5Iqcr1O1/6H0fu8aKq7ttsMma7HN3r2bBPtYGpcJitvvu3Hkmd+fhKD/QoPLddsRK8sIK/YKVgZc
d3LTmogBh5JdjEa+KKmeSN6B68w+lVmy58oC7vjkoeuiCGQ3BmP5+Gws3thCEgskbQDQbj9Q0YQz
YWoATEHNlAFjBecq+kvlPQY9feF6qIy1PRd12JMzsNFG2RJGP3Nxfwqwd45RHhMc4ikVJRyLlMik
bLqOjY30gIns2PNWCfGnlcSSibM7cnm40uwzvO9/P1Uwm7N054dHaomOTl8ZHziqk1T9TfGdZkE+
vTahn10k6SqJU89mk1WEdTwF9Ggzea2blrrBbYIaGktVnSa0/b+WToJlwdpaj904VGdchH6KZEDh
xJNdPdCVLlMzxw6dA7jprzzSmeUt/sOGRpakL2ThFldKzZSUuEkjOPhgW34mWGN1GlmC5MyblvJ1
THg3G30rgUpMR7DWm82pd3yJ6AlXv+1TqEHxNpGFqfmqJUGvaubpWvopfyO2BKmAbJTgHW2J1c80
sTwQj+SyzchjR7kLRhyN5fM+jgNYISJ0q5ULV5pKb7H/tqTLhuaTzR42UDKETW824FgKiY/Owu8v
8b86Byb0PPYH+I0t7YoFJcprzBWWnjRJwXoEycSb9ZCUnNWUIHgNOkFxzC/9u29exUSh3BEORxCR
bchZVrSWZIMPghuJVlVuch3LOhk1+FM5pWQILmcpHFRpIltLTkRK60lKgB9+M/UWJpb/6uYhkenS
HY/Eb2E1L9h07reGSjccn1+VxBhgjzIkfnOCAQlRrjUSdCKm7lXlfEBIeOjyCjV6Wwztv9y2PRKq
Q/qenFIAPho893pMH6qQWs947cxbW8lwyu0kEajjJWriBiqDoqdVadG3p15OMaJll4cvY6kTF4wm
yP1xPWuApNn/90tJ07FQgzI4393TZ/GEL/lBlKXTuD+IuOqC5BvyXMShIDRX0Fp3ePtyM8LQBQSW
gFvDvYfE5VmVNtQmyvgpxK65TLIz6Mf1bz9SJGYcqCfQUOz0xZemSOHhtRFiBL3uSi8Zai46kVuG
Ar/Wd/cNcBT7Y8d8iQFsF464cc112VzrV0ppD87HC6ukcThOHLSwu4q9Uwh9+mhp+xV9l+XQkj9Y
IKWNg1GkBjhF3Ui9bzC59njhY1sRKX10lZ1iJukmA8J0f3M8KL8yQXWEsK1EGw9BfR7zjvS+9dmR
JQzlF5KhCIW0COUb1fR9Jd7Sqr5JGL3O78nZTJwydDqE9mPlrX0IHl5PRve5+naJXQLF9B5fDw4c
x0a5KWd7jbMkVsCQbTI6IMB+tL8q5/HGzIkrWlZIfcpUjHF3imiEJDV6opb1m88B70cjKt57CtX5
esupscm9vCisqZ5c9UWvlgxXZanqqEWOW0hcWR2QS1olJHUFm60+deHJwdTbZLODeXuk12MObr4J
PNvvSHSUvmrChMY39tm/P37C9WPXKgfOXX4mPjit7B45wpBdeCRzSJmqkPOuNRNkPCK20vbFOBNW
nMNsNSqUPVMURH+3yw6O5Y/NdN11Ji7TfDhSsQKncWCeuaseTkd+mxnRwqvdXgEfDgyZdD+uuA2R
JH3pl04fcpO++PCi1V7ZpM/Fi0pjkM/PQVxnPj5fSWZVVpDBdVgYk5/4lUD83B/590fbBjT/HpHn
N77OSeQPe3GSL85wRjQytyp0aSClOQ0ijj7wHKiWJ/kvW+CzDoxIQGkaeUX8bZvl29Kd7BspkgJz
yK8vAPgeIl4CmLP0wX3rBDko1Kk099Fe42XProu6WOyIF3zody89xHvUA4Fr4ZYwJfpraeXYR9PJ
faucjZ8GQzoerk7gGjkgZ4bPtchq/o1LbYzhsJn9stUUhQ+9TKLOr4gRqL7EgesEfsLHnZmEaVRA
LrIPDDlS/v8N4kU/bvSBonHNAfxphYoEmh8T5KXxw58K8b2cO93QBb3QZlGUVqJfVkhcKM+xUqqT
wTowpKwSynAS0RM+5FMa+tgUg6h39Xqtd4ZwA1JYFHZ1KQl4CHsD+Gpb+po5vvvfRL2gKsscQzt6
Bdw/t5c/zXvhf/9SRU1GXIXAf6KWI1P9J68IJ3E7ZKMqhbLiKyyMh9DYhmrgPyawUwEFwVd0Joeb
Qm7x/uIFItzL4mu3PxovRlzDX4gOl32WRh15ein7k01YCoAd88SUryE1poCnsJCGuDPQ0792pXYQ
2FErIxxOcptKhoZzPKuNLGeZ53FvQwdpM661dIla542M+SYjcnBn8eZTr2ZOXJyJHW90P+qtZeCf
9sBv9M0hi16iwCWaW5TyNJSfwUfasPvVu6j6JikeFuNxrBxQM2QtFgUj7jxbnZVfyMZPEdz+0z4T
cWY+2CNN2Vn8xATO+xVwM0eZE3S+1y6C5jMNJZP++I5n5Y/nkfImvVrIUgiRp2550F0ske8ASEmi
KR+oZw2hWmK13KHDYNdmOgLJFo1VHMpcbdtn05uRh7zxrOVvCmoXQGWJowjhZ1gyP+YSv+Oit1Ue
8f29T/Z4KzvQR3KrGrLiWZ90yJvefrvXuVqPGaEv25BcvGBuq19j/TnBirYiRPH8vw6Dhwy3uBVa
WfCJNIOXsi8rXfNDhmMc2jkgmrVumdwEQMti7VGKYb6TLM8iqbHdFRm/xwqaXTyBaHGypomfuWy8
FigvfdyMGcskkk41QACDvJKQ/h1NY9MyIE0eJuuQMOQyh32R43wS3PFuITfj9Ha5daXU/mP6m0ST
b36EVoVyiEfFps+G3vVPdaeGdQPJ8hIBeBHmNEjBq2OspFV5K83eIy4Qvd1SFehSrgGKxeYeK8bE
fjpQTv84JkjMf86aV2ymvOaqwDMkRJbGGz88Y6kCiQd9ZCGmHdX5mqmW6iHCB4SsC4JPCdqPLzcJ
qj3fcEPB0E1SG6bTQbc2SkMS+CzREjqB909r86pJoMTG7lGGnt57eiAkwbPPLWJ3mXr32VPqEXHJ
XHCWnN/JfY60HFRacgaAbREa1Gm5+octA/Q+4ISRBYUxLnGqrYg5AbBkv3/+D55qPaXwB5dzWyEs
YGWw2CaX8Sj+lbRfvw0ZP615tigxnQfm++ULAzHVvVXAwFq9skMouESOptA/LmWqKfwNWQwjkrIR
TBG2Ug3iN/DGhtQYLT08jja/G8/jBUWk+JOD95yDcdRarzRAwCYojIXYCU+71T+lA3lv3JWVtuUj
rCyEmUM0iu7Hyl3sAkSb3MXiKhzRxx74nZT0N2IHz249PoONj96vP6Os4pf4zohkgtlIwioY/iqu
aP0NyQECmjdbxPpfQy0VoQofHT/a2yb59YDssHDlqIUw633jV+XEPGUvGwu8JxMwvLzqBwb8GWwb
nPb4Zz1ifP7UKfTmKbcwuriDa/uV+H4tVV8A0HpGfQvmcr2UxDNBtMpGkXXs96atwy19xL9qhDzZ
kWLZ3f9+T/AQ8O+D91nROS4NEguNl6wMbBG9lM57VtxwJenHzZbWlQHF+ugVb4YteVUMW3uIXaKn
Yd9TPaHCR3XtnFlyyd8zb191/a1z34wwbxgU1XM/X/+MqcKhVwIcuq1tTPoj6NzP4vrwvS35lC8c
TYN/3oWxfoC2LZDOuEBArzwT3VS072TOI50yxBjKELgU1gF2TplsQmn2HuMJh/eSZOf5S62AcJ9w
D3FU9GTfN7zRRtbFtHeNs8LrKKzeS0hkNl+6bIb67vHsMN01kjY7v/J3wZEK3/o+09LJyzCf1fux
BFVzZ5i4RlsG/SF0Sg3yzXHdzy0G7XRHXV/38ABdDzJVhU+ZHNLSHmboG4kMCgb7VvzEZOPPvkgM
+GHDrz3SV2HWIvMCf2NO+dkkQ245Trd5LXG91UyFtp2E7hn2iL1gM8F5RB62N3HDdYknRY85JjsN
Slu7EJQnL6jihuavULWRZ4QvOltWhZfcpR+zpcbXsOXjv2wvApE+F0mCaYExAANgy2EJSk+oDpZI
9Tz9GYr0ndsL4VEo6D8UHsCCgOWT504m7v5LO4SP95n0dp29oIoheo0Q8jl819MGM3EeXJ8pAi3K
N8/GQVGRonxGYCGfLcd8AH3l2WPb/XqGjIA7VnMso/8Ju0cetsLMtLCDkMhRpLBFrLLRvj1vuy54
1m/QiX3hl+vbmaoqaVOnv9NFSn5VDKl8rJTIxEKwt4fL/3kUDyTdTIn/rd9Y1rTLBitHYmJodkAt
bG19fe4cIsiSPUrIvuZAdICUjNmV5W+4g1YFzFPT1qVlwn89ma0lNUGqdYvcw5RW9XIvaq+VR7on
0NNbtC23yoCRNDYRUJaFAmUz1IirvlaK0UGsbd5hgdOLDMKzeMmxRTEdZ1WE0AhE5jaTb464iIvH
gBwyGlb3xg5DvEqFC3GFQDzzI47/7NS8LY6X9KyoZv+qwY/jLX41rZqli5CmdzP6qzwzfZjm61Gg
VRDF1K91+OWaEDY8swYj18Fx9sM/DLU+/fQPjjtbSKHFApIlIpzpL0vGV8EubmAXBk3Rxen/Q2SW
nc07i6F7YXEpztTywDe9r5UvAPFEspschN7kd5DyjHw045xoJ+i0++E/2szaBrxSwe6VOoJEi2F9
tMAOpjpyuxaRWaHpS4ghEz4HHxc7OxBJJ9NyJP4ULsKEeJ0Xjac3WCbflNJvEgHI1m77y0zSDLvx
5EXksNnTkv9YdVYKoWksfJ7+WRugOECZmvYEbrNFX+jsuaaC1SOl3FNJLs6yM/xsyhBgzvsWa/uP
/IIPlRrYI6HIhalA1bcVDj60p14b3Ny2PyNJ3V3EKzm7XqUx1RWAjfVBeY/79LfRr16QxqL8n+3Z
r7pM8FhocclTxy5eytK4fsHAxknySU44SorNk4AjGH32jFbZqzEzuTk6qxj2wNkReGKcXmtcXTsP
XTsLERUxbad4ixdhEPrB4iu2Jmq8ADa1/IoM1V9rSYgvYSRDYLMaLsm7brI3CsI44JGGgPnih5qu
Je4liXUlriCYnS+yLmtM72VNSXAmYvvVZkQBYmWZyG0Gt3DH3rVe2h1WX/Gs1Zf8h++yKEwmECUc
jyRTMi18VurDsVat6e/7NsdWHOINyeXjvXnCSNqapmoOHSxOJN3jucNhUMPdVhDOtakFJcvzmLS8
4a8eFZrJ466SExUOasBJndE+iX7x7BrRMwmvN48Jl9kOx+umbHgW/mGsAxdjCj6sIX3tsJvRFns+
O9RMhFzRZ3C7MU1l9/uFTyY7SsTzVsZcuiWk7SoDTXzzwVP1/cC/0uqL6fPEBDMKPRYs8YHhDi0I
L5CKKTJ7DVPWt3N0LDXSOQ7X07aEHPn5Nf/4M3WqIaShjapkX0FRbPXUuf5PYWzHX8SwDrW9Itoe
UuhR5EKNgS6WIG2IjjAbH0CQJ9Ne5oinXYg6V90TqwYfBy1bbqPsAmA3zmLIwU0eeHZ1uGlSgz5y
poKrnDTb7JuQiueWQHGlkjy6dIOcnjKc+KzsR/R7pTyVRrobe8mMLpxIhLGjwsEwbspnj/E/MyRQ
D0Ngfl2IeUV6zXYLvSZhmqrzsWBgp0bZr/D6aNYwVTi1F7FWVdF6MCnbw4xo/SoKA2NLza8wYOju
YL4LG+tUWAjyg7dcjk7P96+WP8Gt+rsCxZmw+B6Z2mnfB//TYiU6etzvQLChHh4UDdTFfFUxMdmF
cQOHlKj8nDfpbNbgQ40i94uCefJnW30jsSFxHAcF489lvhoG4EpEjKzyj8pOpDxMI9xhAlR0mJU3
jwD0Mnv2kcYEwYm4MMtdZfnY9yYqusZvp4+Th/VoPqM/74I+DXaNufKCflWR+RVE8y20rVH5zzsg
Eh+zb7uATPiiW+8wvrkH3xtTSXoi+cU/SahDYnKAUN1HW9hBYbSsxjZd/gogOnYSOZA72y+LZ781
LZVVUNyxosHz26iEjyI9JU13dl6p9RZz5XOW9hOJFQ3XuBYyqvRYQmcBdP01798sgeeV5ahdyDAF
aSoqz+/lXt2vGqTB/7AlTBSi70ABoaon3CXYiFgHoxmG2XFg0eh+rxjYV8opmmxj/C0iG8IO8THH
LqX+S9YGFcDJKiGta0bTb+85gSN8RyVigxcfnZVx0w6FGXn1UickZr5qEXKy/YCYZkCo7F6ZShtW
M1hnYSH0ynUdK2GXAxwi/nNkCwflICl+FBtZhuRKWFXvGAq602FG3qq5fv3BrhDXCcVFX+bBUf0Z
0oHgB/8Utt6AVVNg3vEjEk7mKu478Yp4tNgFI3S8hbLpDdEF9ThChKyV9CdKy8s/A3j8Np2yLR+f
Yw5YZHNAGufsUPwzjkkRaRjiGdj2Ap2SKj2NBIysH88m6HlZiXU7SlbfOT6E5l2HwoyZKxFF+srp
IvaSO1YsaM31G1392IzW+vkhiPgVoxzMik0CcBy2yopiUbEBLE5+o+i8OjKdJik2h6YEop0A0b1C
KmTgstUANGNWS7Sji+lAAjx/VlhsknEwxYaqqtfQsGIP0xNKmLab6mNocDaxmqdMvy7GxSeXCzbV
6DFp1p64ImWoH+IuLza4OOF2ll7wyfjdUiDwPQyVZbwP9cGqTfoIaM4V4+5itZyuxIunCGddWova
mhuZPti/aar4OUQ0wPASiSAhuByw8mdGk1WHnmbEJ7/Bu9wQmVOM912M2COnlBLa4/YZMaF+tsY0
atHTSg7WEMiMzdBKGY+LM0asfyC66ff/4O2Jfuhg/vMmFytJKsVIlBM245Ne1Leep8aW7DrUbiTw
Nfsgpyvfi2wzemmd+PWnKTkmJvhJqXz5VG3IT+xDNJ7r1GCdLgZnQqsIJ6as7dSeXXYPJ91faVLu
yTqXhKbdF9l/t3G8JN9UtPmfBUsAZJOWfML1vebry6ochOmuN51bOevMOWbV/1zjyrDixf4TUUt6
LMpIzyLWEE+PbE0CER311CJQaGffu6evSzsC2tmDu9W/7qT1itm7qttOu+CP5FCPbtUwQNGY/ShL
PQ2b59POEpqlRh8KajKbfpogdrXt8QiwemHR8KC+d7+LlWpT8VJiRjavvFESk7nJn/h3SEh0iOPa
m+yYwzp4gWccjE/5MWPJvpfPcxD66NfdA3yHaJTZPJVjh/pXBBBf9Iu5DX0dOscgpdwKk7cPGFtu
woTuVvWA7WUU/RkquitdMyLdUFcA9Ls2rMkxFFIoMNptHWGtqD7phMCJr4jxWkpdIYZmmVI3IU1+
GCk7B88qKqsRaPqYxdg+480CC221qFRzVk8ChiDvtEVeIa5/Jejv/z5lI2Y9JbiO6Y+5e99/opVO
v6Ur6ae37R/RdK0ssPXy/sKl0JOhp7pN0k1Vg6ZQVaaLzcDixa9jbyD7WYF/ghiaCBd8lx2VmZtA
kjb8qS2kY+rN7It7FTIRbuIat0hkMcfWyfG2MX6I9wSdYZAYbN0fnom3aX0i9gOEEBwPr04Ro5KM
wnSB6+xrW1DHGy/4XokFxYntin7t2RnAwIWvHZMT2Iguz7ydz0sz7skslZFPb3Qm5b0bClqdYJZJ
1zGebS7b0HDYpX9Oms3eLYrsCGmX3BsYTeRoVust0H6WoQuSyQ1DvZFHC+9CWRaQW7mOxdQeuRwD
jtFMDjOiT/mh0gOU2+R52+UdQKMAM7NqhMHeoTuXtiphDeRefKrsWZxKycMqg0MB1aUInaFv+Kmc
b1QgcqKbELl6NUMt5rh4SlECjB/5aOsg+RV+j5iiR4F7gcYagEINnRgmcVTKTRhV+4VrdlU9ywtM
/2UX82V75lk5bQMcnImMsBF6CahvRBSeo+nbW8PUFMBLul/Nt2tevv0qtpMwcrMkG5tBrKaUPWDH
bog+IHseBBSN1oOJygwxuQUB/YdUFtwPYZ30igRm2Mp3cuZPR1ffs3J/CXdWlnYdgC68IpI8ohAL
2BCbIuTAOlwIcR4CjbUbrU+OK6QOl8eNzSk9W5AiHskt8WrBlobGSGeqFMQ+UW58RNzIgC8gmUaT
i0+f3LoEXJ6eg3w7ITE35AZ9zXhzbMf5KRsJzCRP+/L3xoDM0O1I6xt7H9i1VWgeLafFMMoPpvqy
aMtqGe+zaHCDHg+aMeg3N55+SafUjFjJRPoAzX5nGflWt1b9FDhhkiK6b+C7xhMk9x6IaskDe+J5
bzObmOHHSyiMbLDCA3ll6OdzyK63a37RQg3eQYC2CIOlykpWAZSlouOPupkN4z8KQ8dNtrfAmvRS
Y5whczgvSr8bLn/ovGjpmTEZ8kWXjuI2rvmWSqMlicENH8Yb8i8IGDFhIilPmnT8UzZyTuUPKxnc
c1OPmAQZLQDnzWWnAntp0pb5qEJN0IUtDMXVM9CjobJT8yyACFUJVZJR/8MEatonPJkJ3qQAUbqB
bNjB86BCWO3sVYxU3fFF0s4vimtLmECKuY/xN9RXZOZx6sn/YBE7oSPWU97seXukEoRzAhbDB2JL
sT0joKZi16cKmC3Xh49h7CkXmMOt7Vqzk+CgwiPdVZl8XVRdy9n/ACrCTjPIh6osGA/eArV2zVJH
RU1XX+NpyBzbS2ITkyheMmOKw/csk0BGJjL3d/FpS01+1vcVASeJX/bo5+bbe+QQGKLpQdXlgdub
ZcOu31AsN8OWdsSIreA/RZ/pYpuJow/OpUuO6+IHsUM3ttvm/Pzje4JBz9zbj8lC2VhL/oON4x1Y
ujHwvN3ctUHuYgYT2n97lEj9IZ6oTRFYkPFPow8U9COEswZhpx1pHkdsvqZ/Qv9ZQSVDukKe3Ns6
uks9lMyE3KxD3rRsIEz/n09Ybj3fxFIC9f/QAIL8bCioyGCmRG+b5uaqouR1RSv0gTt0LjU6Sy2S
8/NIMFKToQ8WtknH1QP93XXzaGjBoeJbQri7h6S2XKqvGpteD4/eYDkp/78KvoUI29HuJ2Fvmi49
8t0YEowjvGjkNWIH3bWFDoSO+8hcuisAlZ4BLxP1lcpZBVOuHVtiH1yxIfvMn7GDtttXoFhFdfnI
T5eFq4saVTxnEiLUosxL1wJJoJyCXCRF3cjAHjR251YGXcTBek4o6Z+xtzR2deh3jPpw0l92dqJz
HhL8Sv91ekNQC+EjbElFNlL1g5RiXVAJJcLlbPz7kn5llJtL8eOtfwZhZocDcXpcL4DNoV4N4iGb
/M1dMCcU+IB+vUNAy60wU2/QXZ1xN1WQAMvW0my2HLW6O1O0gI1bidhjvzU3FFSlSurln8Rp8iSW
wB0NIquFzfIEkD/0rJ+7YoTTONAbbo9q/OZIHU0aC7IY38lY8ZoUBQQ1LGx6nU7iTDipsDmSzp0p
+AjlSTEz8X3OENwq6k07UMzT98TmY4b6AyRneRti5vpJIAoMU+k+a4ErG0TAIurTH2bF25xThCwl
dV1zWykuPYRSn6bQg4yIASULk4O1tYt0v+l8fm9w3qKzVeTe50v6Iq0RWTnQXXYuUm9rAeStacbh
WVU/hWf3NWxQhPDawcpDr5bkQ7xbguFcgCSR2BDxCkh2+llLN1+EvMCAM3dXL/VkHAMMbf3iXmDm
2Iwq9chYY5hk3e9gxl4cCFYeycQu85gmDZU1LZlQvRuntF8H0/xMsn0V5gpCGLJtWwHQDS6c972B
WeKr6qxOXDCIfAwxlrbb6SOl3vdTDe3NLQT69lYNGP25xl0n4oOckoH/4DWaZ1b7bZ+PsVy9eces
y47/CIC+l3e/0oKuH2jgzV/dcK9w4ywez+17iMhpm78zXt9JLg+uq8i8ya9+vYLgO0OPMVe8slBp
2aIBSTfsvlE4Uq6i+MKgUadDujaAuGA6fZXXKncpeX4UnXbLki/jhfmhZpB6vu59AvKyFqm2Kzfn
7OFJ7kpi/Ij/uAecI0ECIZAKKJDKlV8sNu7McqOLtTwafLVbV+Y9n5nyB6loSXY5DRKNdhZ7+04B
9pROHH5NMgrCIzCAlfc9v1u03fz2Vc/+jVhW5N20mBv/SSK/11PzRqrkiQ8uWy92LsCEgrHoYtj4
QfpV9q49TsfNVW6PYYv9A+NL6Ep8z5BE+Ebdw/PYAByZcKrUIwq98lv4hcIsLgmJjtKTH/6R5GUl
2ABgRTJ60R2ZccuLCvAISESPX1xM4C+7dNVEAujKLUwNpJ4w0HQtDZJew0aXZijO/sXTaG+2Z9vt
HNWHZJWxZ29ebcsQLRag4DEm0V2F2JHYmrfMVrG/VMCwJ//SwMQCcTzCEbgid0iG9Hd4PAnvrnW3
O5RDqTbERgwZ8AZTEdfWzEYaKXYxiFD2Liut44GeOMd3+isvBSCald/PeYIo/wvbNoYc82uS8BrV
1n9a1xlsJvEUg6Dm/Q0h2c6jIUALndjkhM5ad9K58NtFInECbnyruX/A+j69JBw1lZu0SrZIdNBb
h5vjtcCifBpOH9D6Sal3Ur0VX8w8xRxOQkSepT3ZdXyrKvm0Ybe7CEEsM61FOsbRVlzh9dHXGAQ0
06jpEp47bBQdbGIGsR+VBwXCKVHqoE3gxeG3xZNX9jJqn3VSLIlbye32bEs5YINcwBYuFJG7kGxJ
yozvdDO1ttZhV9VAcaJy+j4FuWJSXNxlu0fg2GPv7Tqh5k3WrfBXtaH8mSULbr4RB2nJyjpc1M8F
0mabBO4wSUj6jo+2Y6B84H7F8Sk3Eqgjc9/fc4ey37gGFn3NwIbX5h/zNqVrAI4KgPfXB+DuUSkQ
OHMjMpniDFZqg8YX5pSNQ+LDU2+/PzFRZV8gNce6T2Z4zY70oyPVX6DC+S1uVL7WZc8IINrOyuNg
xVswkW8u7emlrGvFbiPFbdvk3nq/c2XANYe7pJm9OTcBa8QNN2NHJKw8NaDf0CIXxJZr/oqJrkH8
67xD4+LBXhdmu3cz8ZlmQK0vk2NZ7NvWTp6XSL8/sJNszunlElUwWVGuNvl716eOijrfMzezRboZ
UTZp8qDp6chuN23I1ir6nGKPz2j+mYc4eRubCRsczVLRFgU+UKCxqZa2iXcIcfRbt18hOhxB81T8
GRMT5tQ57ZZYppVwjxky6ykBBS3bytqViGzAM1ol0Y3v0Pb2Y7Al1PAvETkj35aq5wQPR/XDA+B7
FWMKqH8L4udICFT0wKBLE2Wfu6uWfWmzbhR7xMLiBLwWSzGcXxgyTLr8Z69RuhBAE0EGVD4jnwoX
/swXcg3B9rHR2vQAQvEessgvJ4Ydpg+Hl/GUhcngsvEv76FJG4BhtHXNDR9Y/MZXnbs3wg/n0rhf
IQpM4sI7WbyjAIlWapN717HMZLM0XTLgws4pf3sAiVWdFu7qcFjC3HIEgnYmcSRLc8OyTDJblynY
lmNrtPXWfxOLn3j1mHMzOvbbBg+N07D6ZS91OXv5qSkIbxLmxZD3NUWs+IdMD0xYX0pS1yM6RZED
IyugVQqTe3qgnLvLoNAB0vSjGKNPQXyXCYevJWrIiwpNjVNCb/nxB06ueVOXLh3iCsxSflwbckb5
Qt4Zfamzrgjn+vlhFsniq1a+y7Rdw06Ht4pTX5YXpoSGU1TRlztSKj5fLElclhyax53BpLzQ04FC
nYyVJ2px/OD1Ak3Jn9w+4zHYbz25mS0vBbPQjHd+jBb+QAOS2/RE46mTOEPxlXy42aTGjfcOH89L
a9seWj0xKh5WHFaizffzy7lYhm7IGmJykvn81ScCImoQqCM3KELV9MkfSAti3vzbuWwHVUqPBCEm
7TtigFmt/fTc0tKxktu7sOxhuVOUappVgDP0dpuHQCfrMt1+A+5pEeKSQBYRZYqvoECtSQrwRWZR
QMAklYhH3O+FIdxGzU/rRCTIpf+/2e5UylG/6M6A7J+vGTmKLNY3wrIcGF1gRjg27HDX8dAOtGyM
8SqYzzfF7DVTZEOGATgnuD8pxHZiG6sXGAhqwKWiYdEWvsYaLTXmZHBGKldg3wKZqlisz1BUZVkO
EDeF+Io4lu5u+69vt3nOeFWfwBdEH+biwtyrkBMW13XEVeSPk9O8SwJm6WrAbeOn4PZnvkDAQKHa
9vdgcNBoSd40SE5uUqKf1t2S0gji25ivwE9iUosRlmbuJQfAUs9yA6HTQD+Apxuhdd233pqYQhII
9gI/9xLauSiIcASHTlsn6r3iEH2IE3gT1FqAKrn6W8qMbLyijC+J+ZjQQ0CeMKelsl4tXW75lHPA
oT4/srqW6R9GXUlSXUXshpyUtqCeUOzKcKBDLUeViC7b6x6eZc/WqrU6sCH2LJXCrnUz1VWM4y4F
8YGvJ6N5u7lBwNMFPMRKLjhmqvCUb3jQktfcnQlFXS15dA8z8UfO1sV1Gfg9ei95WS+PgoQPF0nc
UI4XNQY0TORB113+ZCwFbbr3Nw4DF0JzB2fzxM7EUQXD51MckudxWQVNliUMA3va9rDSPhGK90y0
6djUqZWpkE/K+T3BJEP1G/xhE6Sdse1/XtNhL/aBUDC1kjPvYFzIH8TfLLQoAb9hVAey1dzoYW6u
TjmIOOGUOvAcGzhI55FhZjdkLSMCvhV7xHQRGAG/jpjplw3KHK9s4oSJ9ELnAcWHdu2cASEUei3s
zinmLApFV9eBLQ6RXCd0a7IfJ/Z+Y8ykQpXGdFnWt/grlkjp7AAoAS8FtHgiTwNaY3Di4JuymHn0
wkbJOXct9FqK00Wh7konE2fGexNrI/MIvKuOjXu3iWI/64fp6D1upagXv3zZJTYEc6BIjb50/gFy
/+7JV9JmMBFhFIrr7N8JH/q6q5CmY+ZyzBVS+scYNcZ3aap6pkDGfKXcWWlJHRgV4CRODDiWYCLe
i2+sRxgPGIb0VVUOFePLb8t9VaTFcWTRZsUR3BVXVa9ZtKJ8aYOneRXFaEiOCL/OTPo4oJB638Qf
MeaxNE91KI5HIu4E61QxQkJJRJSLee/C9PfxkRq+CsjmeTgmXVZiTBeoFYXmwu5BNNAE631xhwKJ
959z2sLwXbbCAYz4nKk0GbqhZqWnd3o6dl6x1GoHMSlo3Jb9sl5eHbtNSPt2eRswE2Y6Bq1gi9td
z3nnAC+QO/BqyuT0o+KI/HTYBBAfhS/VoNbXZ+IIGXB3+SFzLsMIQ8Rwpg0xwLN4xihYN/MBYsdT
ibZ0Pe9pcm2KH7k8vtRa+vv00Ep8u4yVEYMkgyBWYZwKDqEoaeGT8dfu4boB5S49iTJlO0frHIMT
JM5wFV43nPfiSnIhVO5G4xRaUrz528X67vdSuzjaMmT7Lgs4oi06b5admziT/oPud1XExvBCxG26
gXNqrab8sZAG/DbMIDrBNgupl/77h43ros+eYAPzSqT7+WV0s9zVRA3ypHA2yaOU5TtRPOfkNPC1
urmVzusQmzXUtlaFp9r/5dgJkgDqDqVrWJ6HEU/8y5z2bRWK1qfzqW6oYl2jwcLePzfeqmPRkDZ9
vZSdz3i93EqTMOQIZkXqSq39UoG0pwfYT5o9FJ2X2tfFQari/HtRv3Md7KxTUc1L6YrQ368rtgsb
+t4YEhg4V4ZPaX5tfQjkPjQdmCCGppZhDWrL8dEqPvHfBxKssSTttDa2+OyMbG3O+UhSfDGDlpfo
bi1LqRiiztnV5SKZm05gTXAN9Fp04OrqSMuqvoqj9bQAoPz5ro4e4RHQ8/tT6OBqWq+2jS3b+Dpa
qvh0kfNECXMliJItApJR/seRtZquB5F+nKeL8mytV225SUjCO+LrizhGe3NSOAnwy6SlxVRqxwr6
kiWSsOTPOPkXAv+fKE9NU2R6RIPDODGLHVFz3o6mvxI1iAMpsLjCUQaGLMwpaXwgdO6CYtzcRqqY
jsu5duWtK8rDJImPWlVLNU+rvf08If5DydhrolozS9rsIWRse7UjWylmpSDtP4b5HsJ8QaYYiFPe
XJza/pzwvSS7n3sXLGZj/+fiHfaS2pWrv/D8tVyGgrrAe1eyxScaiEkzHHdeWTeAgmmAjQVYcGBI
6f/YBOrF/+ql18nuMzK6SomK9+3VUC4z+o1FjQm4PdLUZpplhn/UxgNJdNSP2rGA7PG9q0vWLhhz
Q2ayZHcAVveRd/TGekjLX+nsKFcgyEvdWVkCJJPfbTXRaKlI/Tv+cMb6+WqnrO9mzlq5CG/yhUIy
XKSepMdyibTojsusaVGo0YHqbzUVTqIS38XEq/zyMR6yQ1wqt22nZLyxM6QICuljGly03RX2SR/6
f6RhdTyuSr5yDw9fRE4PyWcxZQX547pbz0fLoOyhOMXLGYz4hQO8QrDFg44xgxIxUaDmddR2Pfv2
9nT/TMB1cRhnnVNkZ0TqKtDrvMYNylMzaQ4wPxK9H0wNNU5kwfJADNWahV1n76cHQy8uAg4CFUk9
c8rcUkW+lCcrAG6TIYlRm6aojtCR4kTaoEv9UczQPo3Itzl/1Sg/PbKPsKWoxhGNlYZ9KsroQWHk
YlJ0cUdZvNXb6oOZpiECoRc1RlJe6M0VGcSuLh1uLJNZrxYxEEwP6wfPQlp/r0oo5ylx0fYObXpL
PTfApJwxwZflsSLfJ0GKCUR1ZV+dGt9ey7CQ09W0oFhhIIW+oa0lCouMJ6B2jAL76IlZ3anAXfXP
n1FmNC6/S0c7zYun5stdq4SpPc+HFcaMzb6K/zVNUOZ8x+ioaiKpzKEH8elc+kc+trLEHiDvvsep
Q7P+mR0KtY5oBPT8NWjFb37WJpJwMcDOM6FZjiWuStlKr0rPjjsvN1IlRHTDjC+6kXvuwCXe+IlT
KTc8HtaI8F0AKNv7kipImiZP+sGyJb2hml7pZ8Z6x7sYeAOXYrt58gzFLUlv2F0uf5Zh7YEkfQlp
I8j9gjQezSQeXZix8z4RsCY+nDgdBTAWKuNC7Af0sgEufVtUrcWNKHiksIakZLgagN66qL+u8eiX
J3U65SKHSLSm4Y69VWG21z6TVX2l3cpfjDmr46YhiLvNZLh9I1Ti9tFngj94ip40BiDgGhtHo2Os
wA/uUvSes8djlXQTFkorRQZx8Fw4Mv2LCkIW+fP8B2rmLuv2QH1clIVZD6OTfLn3HSPhKijCZd0d
yb3u45dD9r57LXpdTfHhyZHB6VUOe7OE25n9ZUb/n1PU9lqRIgluJRUdy52DGrWC5EKULDMRoisd
eNDm0Zbj2QJgTteAyKEaxbsp2cyWJrKsJBlnmNLmUaAzwphlj23I6dfI7HuCJRSjMbT6SXmPFazc
aHRV+76he5l1hBc/FBIAh+3hOOSybcZgZ77/713Rg4xL2cnabLdpjioIX2xE3Gm5gI/tuedSjtxl
7lBErmLCt2wXNI3Kn5a2MzpnUdZtnqaarS1Rch9eI1RaDA3xkUYvSOgJsJdYLyJ0V9D7eOnsowYc
0//tOaQHXj1NToUiHRB/4wWGjJYD3+E1vlkyby12QouQIg052nl/I7nCw56dPquqRcGw0CJCu/j8
HepTuNhwQWSpGdvJUjlPD6lZF2DceExXJRNVyoro1BUBbHb+7VavY7QhJAeSUDoZ6kNcB7Z4pNwh
bCvFZdyq7JLaWsrG1Bgff2Nuvmanu6P3lM456Z8skj6vNuvXumUqXIM//J9EJr/5IXvXZXQ3AAFM
un8MfiRbTWFcp3g0dVHwYJOQ9Ax4tu4Sv+5AuUMK26C6lPZTNZSJaOX58Uupo4soFBtYGgDb8FQK
v5iUbe7pWNCRzSQLstM2HRlXUIT+DT2xqxw7AKZY18OQVwxhRqqcnxc+PquT1x0DkNtgMXGz9LgR
G/P2x4Ij+N+4YAbw0VzTPlw1xlyHFW76GyDNWl4iXcG0j7ba7cS9MaqEI1P7aCU+c4AXAutXJd5v
UMk+uNQ2Qing/o0mw4Co6qy8Z/lopgwv2VSribmqlFBtfd64YVQV2XQDylBCPNt9tEGgUCq/XU28
DL2tyehNbbRt/0jnr99aMqWK1e7LY/asdUpyBmPSjZVxeQk1lJUGxh20KQk/NLi7bBXidB6kSm9J
whbru6aFKVrTMVKSN56HR8qH3OszrTOo8k1cOQ+2MHqT7CXMqTPt9Ssw7mR/w6lTXkNteJGuu8a7
GHCTqoLrzgZm1V9QAUEjt4BdObVgZyu5MC7IEOwUQo9jTb1VI67eWh346daGn6Sxup83NKWHJcdy
oTzkW6pPLSto1GEP6EmSQh7tBBB8DrsG20KbCN0oId8hInFYTLxiAQD9X6ZydF7ZNmbhSceZecrj
wIgDZjxGxMhsF86ZVHvThWD3SicoqMuBbIwgY7BcvDH0Hqm9Y3a6ugPvQcfHFKkAXwtTiPpwVQbu
LtdUtjb34Ro1D2lJ+oyjcilQFnGPZKFMERF3zq5hZQ==
`protect end_protected
