-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
i3swIZ3VDAqAjOxJrDRbuZDwHMd+a1PbNxAzxaVa1tm290XsTfczi1fqOAKHiO9qHE4rny2pbr45
MgcH11OzeVrtIPIvw0hPtQSWvTmj/ZEpHEg9p0MQ0e+0twhIP8j8hnAi6mS5qoCjKBXPgAqoBUba
Wxk8l3soCyW2RKl96vkz5hIIn8vcXKnwDsisPbYVAff3RXpsDs45COfQYLctdS/T3k+1b0mlBKOl
OLOl3eDE9QW4po6t+QLKRAt6267I1CcUTKFtJPP6+AhDTSqAlHmHGXktBmVglb1UEUNV44f+mGdD
1UN7uoeLqkO/cwUI5eTq+bqKiWRxal+udXEAqQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6016)
`protect data_block
jj+k9RFWH8CkN7c61Iou3nRK9dd1XoQmd3E4UioBDXgYWojn6ckzuxD3hUFecpz2F54vTypoLwvF
f/ZUHgvJA9OYEFXKY8DtVyykWmStlXQy1f1bbJJio+748yHFeREj+VkpO2VP/gMqJM0q/Gxjpw+d
5JcN91y7STS0e+Hit1Z1ApQdp+wq9ZGceO2qRNbStnsy1yY0TozkljvOxayUU4VfTwxM+D+hH6/f
Ygn9phCXmlp5LOERhr8+XzT+EVCbJ3DUabiM8vJeP3QJ21C87gBzB34UqfP5NubVjDPuiz7GR28X
4VqQEQ9Xy4zKg7h3UYZSvy9CrSKO8Wn+eD0UE6C02kTBMkOweGGJrHkf+OKapCExA4law3/OD7N8
K5Biyk6mxpQb4qOyKiuFSaSpBE3NRCprUhZgBYCZjDJXDmKOtwASakL1tdORfzbrWUaH6aHT7nwj
7oM5UXL17ptLEW3PHi/oP796CuB8tNc8LN8RjzG0YJyddjs21QBVT9TzlI4SudmXGQiJldwEF1jJ
tiK61HdCXEKyzfqCcdJwfJbyS190JMw06HE/b/HRw17Rq6Pn/rhXaFGEoivj2nROn48Z1ygl2NFG
KPu8y0cABS4H4M3pBSdqW1+IxmhGBR5U8Z52CbMlIv/VbGqw3arg2ibz1qE1YjtCR8Su2W6Kr0rl
C3MVRwkthM8fs4WU+w2cF4JEMrt+cPC/VjsiaLhKymfxtK7WXg4jvDq2rjecjxOjyIm+HSRt1Hcj
dGeMf6y9/ZnlXguqyvhyVJH7UhWH4u8xo2EhYSywtwJkkegRLmeWmDRnae5RhE/tKR6sVijEZNc3
FPxu2kjf9Zj8WPLsAAKfHfNGIt877jpFftYGgnGC0arLMpP2x+t7qn9ojj9/Etax4qFAIHCswtWP
WZb/Ca4auuLzjwY37dru+g39LXdu3XMhQm9ovFYifmjmb/GzIQ58z7/avDeFwtScQqnFq1Kt7bsO
cfk5pxemKGqIrsm3XF/TbXY2QYGuZGXuvKpjBTq58zuU+0X6qlFX4u+g9o43+SM+tF4WCSDv2S0L
WaiTfQk/1yrN+J1hbz/+D+vWqLO0xM2599487D4OExCHVygYbP8ofirzBVCe+xvSRAQ8ThR/9iKi
14eUijxhpj5WryIvLGjDuHqDPEDxcgogOqceWHFHljScMmgCz1VTab0pFqfHeuwBQp6Kb7ZsRI/M
baW1hQ6mcwFvuCRsV1Fz0kRCWIvnAImpBTeiCK+poCIIPgk4cdtOfK8GKaltIGWdTulOHiN/9RyH
+noFmrOVKlCFL6qYx7d5eLcPYaGVyjd9hvVS+Q7xgbuQPc2MOdKrAqzg90egRdauvEIVuVn7h7Tl
vYl4NVrqzIgjz1bDuRFrcTUA9I23ETy4nm/QnMNszfT+gNJwVrQkvtX8KZfkZpkdhGrr+urUWpXp
Oise3XGbEHVeC7XTZlguegtAoQcn2QGyZu+nI+hhXQUePnehPkksx3izKt0lHgx4+sxJBPnojyxm
+lWa9OpuBrL0K+76HdvSHuUlN1J1OKYk5NdG6uhykloFxX2UyRSXvbBQt9bSeVIwE5sAHwHlGCwQ
piLJEd1eSOoRhnMpcqzuwN2D0K1ewUtkuWwE1jTWaK4sejWjrvRo4kyXXW4O0XQNJhLZ2w2BAOhx
VDsoxMeZD1KDfKV7rFh4tr7wLfjHiKEGI1kX1nGOtObutZ2NKUP+W67AppXRey+GTK7zcRAhZLn/
VUa8AhGv/RduMkDrsbEwXApGWiACfuad1DNFlN3txma4ZBkjfH4GvSdq2C9DkJCIhWmQPllX6SRA
3v6pVu4r+BY0ThdcVt1cBhmyqBFDRJslwnTJKgh/Svj9qn4FIQCid0D++Sosl/Hw0FQxUHMUrO/V
P9P0JWCxlj/8HxCPNrhp5KlQhPSGnW8LPbwwWZAABT9rS6pEkg4zUQU/to+3LSGng9NwElB9kSSX
BXFEVTuANvwLZWcb79XOnr/2c2lQB6Fi2sqgND3gmFXVDfXdYnb9ge9O/r2AjQMOSRuwuoStPFnN
26MjvK+km0MC9P5EB5oqYHy7c+amphhE6HXhHCgr1Kf6RpWw7fWfxczBs7Fn4hLBs3Fu8yUP7gJh
rR4WpeNrSpbjgsopmyEquHHCErPk2vI3DwwraSt9qMi0wtroF/a7YTxUXaPULrV0BUp33DJbodn9
awgEIpIV+kfa+JoENIL/rlhGhgFbAlrKoNBuO1pIbnL0Efb8QmnA79cS5J6qaOEvTNhTm5Akketo
K2cw3ltI+0jrgTNMNS+DOxtN8i9YvxJY/uEFdzTCC1sCnPOytRSL364tz4U9Y32K3+U+teDNHSNM
IapooUBFYEXM/j/hknbAuj8PqCIO+NkLUBWRj54Xz8eBKhIyqw7lTHsX7atikt4x56TB3Pe4pFFy
3/sO761RkRi5oHFWJiZ3+In0BQzUUU/rQjTxUI0sf2K+9+x2mUV3TbBmRBEIy5zw1Vjesm2tz+Lt
s89CdwLEQ8tXSEj5z7kp0lYVZ5HEe9EdGHgniW87EkX/mC233PBp/NXAwOF/D6e11QmqK+yhsWvR
lALoaClAIAy6f7j3qrPKP2pj+ErpDgDAu+YV2c82hKj/QO4Qj2eC5b1xUUpehw6UMXgeVhxNT2DQ
2foMdvBfszgGbnsTDonsgh9jh0JPVwVQVcOe7DHI0+WlR4CaPyX1CfWFlGvz5nxFX2aWvFHk8h7X
qYXmMrmIX/C1F4i/pJZSUDNYSgnlFAg2pbpeud7VDAR7uFOMckSLEbknFuy56jq3gFBe6Lwd26WC
dH+BRVcNw6XMu+8ITHeFSqQZ232+ZDZwoU41MfWtys9w79B5wc7JbDJhLILyTuZjQ8JaKbZsjpGO
tkUe40jjFLksjCVjrvEgoSDEQpuhQoBD2JKr01LLMQanil7zpcBRVZrJ3TgWG0C7JPBNjoqz9skq
jQTXCZbhAZaMLGsI5nFAWbr0VOEz0ttZ6QOjmCy2YKpNno9KwaGqTsqnPdaMh66+kP6qPeHZ+iWS
J5tWFx7b3yyT/XnJzqGyf8PSWwXWcigThE2ASVvC4NaQTUcceVJGIcbWWIFbszuCC7xzgFwB8yvL
WGrMxPeWFkf/KgurzA9qCjZ2RpKwiITIYQ+vzYi2U0nEnbhi+qdkwOk1blAQU7ghClPJDMrlyA/j
19EgY/8O+qNXBoCrvYxN5jZOkMSR9MIq41Z+hxy0SyxLh0TBFVVWNC48oihTdYk8WnCzq8c2nfGA
l3rwtGzgaS1RZbEzutGvIYfdQA8B+QROhsVOOkk+P8RCthH7Ooq3wbOdywN6rRjzXY1c5FZaItR/
UO3YeiTGmCcMrTU7DBFS8UbYs1mjOAlnynZcOD013KEU/t+0HHKNYCEFSiZcCMaW6p6KlH5cdIdR
upSi7hlq/uJk7LlcSPTh3xrhJ85rLtZeREeKed5N7bOylaBUBDNhfL5cfvsRyxzXhWD5xC/2co2G
1xoMKQ5raHbEKnTNbLl2l05ii1g26DyJF6RUyqsE1BB9ybnGwjIxpfH78ehc+OGiQGXBmrvdVi6M
HiOd+nvuYqxKLAyGgTsTaI+V8NRUGr4GWGn8+TS5XJaObmh2/PtKvT1pPXywgABc02wA8QVXuLI5
7Hhr/g9vAAX6T9vYHRmM37vDz7JPoIYbwsAekI6FelCvkKgDvZQRQd7w+mygENHmU2ioAz4Bol+g
DVPVCn7iENVk0fHX7Jf6uhdUlA5FHSEBuPz8ugyk3oa/q4caou2C2R6ofQqTgC868PFPoRvf1XRc
You+lr3VnvuNr3vfJsqDZDdCJadmsAybW3ITVvnMT6GqFcnudwSnxxMFUd0an82ZkxFB9AcPjUPu
0gVBiQN9lTTUTGCdf/76W9ofa579o0/BjTBlUXhUVUnAWi2wSrZX6Dl4UEY+vMB6VXvC41LjWu7n
amAb/S6TCz9Zc1f6gJlBsgwTlvfe4K02rGWbkWF3DuoVD3/ZnSEA5q29PsFIr5D1vaQ8yJovSqLl
WBgBePpUPDWq5uXxzbagcuk/5fqFD+9xqn3YcKtlv27IJNvQ1q2O7LJ9zGOZ3zJt268zwuAn44ME
yL10z9wSQBCeSWoWf8lEhm04dAk/5F7AAJtAnxzi3kL2MiPQO4IoQ6wVfrPJu3gfJ/4tduFfYe/J
qCRMAM8PuJk5QJSYLLxuNofb0FGnoHyBddVrHwQRD9hoV95TxbjJFhQvRXMhlieGYlPTLkC+d6OT
9VNvkF4lDlVOV4Ta20+K2dd1W6PEPWiDQ7/VM4LV8/IIP/FsGRVVQ+hleyoKQ2kvn2k1uw9O0ouE
oYi7NLuA3yK2ZJsH6bNoVMvoEjlKxhrYWoDwqk+B0ccfSuNUaoDMkf3FmFGxvLQNmgsGQnguoing
3JvYrEy2R5i7XPegJZ/3wvMKW5D9jMByX5NLZq2aOImz3Fee1EFbWu06eiVA4pexGP0iiuh2t291
PRzm11/kPPoW0aem0Dji3+0LK/4Tr2ptrkx259QBIqPM6iC4m8bbAS0czJJdKakAX45iuM8c9Zrk
eHJShz1497H++gcPnrjS1QzKuBRQzg/9Py9NaS5itP1TSJM+kG2DWFZ+LT7BRlzzeylsPYMemlbM
iLLpJ+qPkRmfSa7gPd/S4fbm1Bq/i4ifvjf6rmRgMsy9p0PCLo++LU6yGv/vW0J82OVWvfx9bN4S
qLbri5qVzYHEu9eueStCB5aILNOY7oP1TsQt71dXIAO3drSobJ6zcI+/3red9pwW7LGea3maH71l
oAVgaUcg+w/5ujWMxBAu3eP9jAGgMwx4Y9n/sZzDxXobBfGWtoCCyxzKkYWltp0LOotCgESQ6cVi
LSG+IFZmNR1L9zTCTJf3u1mJrAGowJn/M9Wb4scNo515uN2ix0rtv/IsRfYvZ1KwBDsKCh8Fd23e
DZK4PpYUjmbJGgHcSFtXGdo5IL9Q2tqeMDvd0Ml86s+/Li9yE1wGRTIAbEz2gFGJyvc4TXpzX2wm
Zu+QTxAtF7A0/28mTjVFoYn5Oi3/ZXDeD9Y8iT6q8AEa/0x1vbPg0hrNfGlO1N4erUu4o0oEE9mT
4o1J3lYp9HSahvRnIZkI2Qg0/AqT7G1DWqA8leVX3v5drCH4LevK+Dtti9xva1FTTO3XbWdlUw5I
kFgUFknim5Ol8bHDdXpvRkYPU3q6wY6g4fIDx0lRq/mqfROzFc5akIukoTSEtME65LjdqufYKukO
x4kbQ8It3OEPzPQmP0NKzmWVDYv7Aql9ghxqxpu6fuDy8L3rUCJ3kkQn/7c9JBI5VBEClM8ko+41
hpvXuY4WUHx9ajoc12hbnr+g++KbS4JsDLMkVdhljUJWKKQx13UXZ58VphAmGMJbIEMBGuWAZPzm
5BdV3q6ytb4FN7fWFqXMvX39xKdlM7xBtPfuAJuGPE25hGFSt11iY36/pHUwmlf9gp1YOM8SffVV
++5sDhesNF795zjUFFRhbEynTlUxhPTJcVBZWEyliznWdle93sescdH85gxc+psTgiPo+ssQ01Qk
UZ1H7AZ1+BVHljucwuzHWEVUL3Oxalq8CVYWTuLhhJAKIXpcUOTibPGpzZIGLEmlyb8mwimIsTjo
wZi/fMN90YJ/lnEyA+r6g6d5s5h3R3l5QBtFHL5gUcTeRdz1ZJXyK8ExBSuZ8PAl2b36SmAUfC6t
XyglOJXYR8JT2T9RH+I0Gjp3azjX3OwRxI8/kbqYx3JDWjk/ox3Wgfk2P7uEDiDLd2yJL3/ohjgO
bpsZeA1L3IZlNRVvb7n3Svqm09f5sthOtsJBByHdcvMcvvc0XqhOAcjK45ZHVdoqRsn3TWBhZkSG
cdQ3nlYBnVTcKyqM3JtpkKb5yb99IjABKnuIOc0fQ5aBEM7PDSpws2ydODe7VUmox6n1GJH5P43r
Af7kec/QAeQRciMPjkFhE6g/9QpdLZLWtf752E1Uck4Ro+vLNIznRforPTMBpW8E0YNhiBB9jOUQ
P/+85oRtNr7u4YP4uP0qUngDEr7LjmHh/JTLKQxzQpmRLGqLiE49wehBzYsCM67azrWXVuip3zj8
LJGS7kKtc5DSUd8UN+JTwnV1aTSCuf53Y7ywZZnefGnp1641p5qKT23qSjXYiDWgcTalttMotYOe
w8xku9/HtgaN81HmgRw11NU7/dsNO0tuX9922OBfkQ3GIIWoCGws474oxzYsvRVhD78x0EUOi99y
X2OL85wC6nvnWaQK4569irl4zv8ATYPdLyt3Do5qdrdlKVEhkMifj0Ffe1/9e+M9oXzivh2f5HxJ
wnxMc02FCpxtj6d+Pv7dtQNyLV/3yO1GdFWHC4P6OVjkanjd0S8R6UUg/Vm5qJBd/Jegu66hvPZr
o+EJqu4hxWU78YRaIPrmOgEHuxVsV/GB8yMc0pjOXWS67EkbxRbrC72XTUY2rrAWvPBrIZQXPEo/
2Lgvxe/dNghA7Bnp1RMYKvL7b0aIRaWVwCysdHiMxoH5+wBr6zsnHhidLtKpy2mMbb7hJg+0WcOd
pC9TAbQIRGnnuarb/wnwIZJUSSjaz9DbgMRsEYX0EZ2RR7v1nnhCuOJYtuajAwZ67OYaLcPXIVyJ
4uxNCZyrICR/eX+viNR/mEKv7A7wKnD05YYZHuX8QaIGSMSJdQ+czLfV5zySfM3hEKasvyuzV5AS
W4OzEXzizvIsCRu1RNpMmrDnGxjkQiIYmW2i+cQLLzJNz9dkgqXvnIQo2XeVV3AxtaDI1d7NJiHJ
ERFsNB0Td+9aah7wJEiUAjNCXrXeMUGIIDfxEl8zBlq9k1r9xJJ9/SikMkyeUGqYQjoXv9ksvKhU
5pOJUBoSj5ASxC5L5ToQb56x0m00Ta77favFumALB2WnP6snsko3riWRq0U2X78ye8GrBjPpx9in
RaxI07wKw++cDos+wX7oCuk2UplkilG4ce6A4ADk8occ+tl7qBSbb7C4fiGTe0lyGV4g2jeVzo5b
otwK99XE5GB4yvS7oy74Hv62YSRUfd6P6EyZleWHURPsoYEdmHk+UckbqoEQdXQ/GP/xgfmIUbCs
SazUCnw2LW+newQBsL2fMOWQsqRrrVq5t5rqME0WeWGGqWmL1pXnbKpm1JAIUXqnVa6vWkvW12EW
pa5JnERd15pCCxa8FGPxsasXE/8PoMAd0GzxWib5mfpR9dJHPyAf3rkgzr1Ypnv4zuyr0xDD8QHv
HZZd9frByonmz5IQsPOdf5f18wLNWWLatKBiwTyZLFBDftQd4cEjGiV/C2925f5vNOmNKhYBcZ2u
lrpgapJoTUTgY0dhR0JfjNMQ/ffFeOTzZ/946KUpIkkxyAs635vs8Ixd6abEY9DzzIaP6sDDq55u
uWXNhL7y2vyP12x3dU5Xz4tAcHjvf+YmSzub3P9W2cDBJ1u0NtlVNZy64KSeNlx/DRHi82FTepdN
aPZDImxjTOTKeKmVJP08BN9JTl2fIg25vL2Ka+hP4CtIQWO47rOTXdU9QqYGcqekvTNbWJwR/uEe
NxxUqMLAttr80xoJQTCwWCeh3pM6rbUw3gj9Od/Bh/dxl4fxDOI/9/hEmoFEl3TZcl3KQM98AdJo
K2eYY+ouDYBWAWLmfJeYOFs8zygxjN+Cj1T5G0Hez24YWW3037/LUgh/LXd3mf4ErfX14AxFKosi
bi036FgH2YbZpasnq/peKNJjqa8FwyBX4rHN5GanrT84uzEfhVKQgs+za6VEKPdukmlhaMyUTsO8
bWU0AWB/onxTIHUmwPNQ8UdIVA+gMlvRM7tUcvRzpGIWHFQFx6Z0h+2NFjkKckFS2pdKZRzBguA5
Fdvqh/jBXRb7gk6Cn79iLvbnHg3SFSQOGOgTt/zKwmOD3TqaHTTfzY/bgc8+NqcuMDQh5vU+JkKs
5alp5FseV8IT+bYM6lVWZJIlBqXDLvZPHVtWvHQqIWVu9D7IOYHyA6JTKyGotDdua0HQlDAeDMLv
VcZf6X++rD5rROh5lIAaIDlkZKcca8oXKILPyN1wSA==
`protect end_protected
