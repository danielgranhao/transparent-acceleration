
module fp_mult (
	aclr,
	ay,
	az,
	result);	

	input	[1:0]	aclr;
	input	[31:0]	ay;
	input	[31:0]	az;
	output	[31:0]	result;
endmodule
