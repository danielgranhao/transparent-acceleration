-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
hctktk+qYgwJn0dy6XarWQoQhUa1ym/GwJ9kvI7voLC7ufBzaTjGpeVUZ3ges9gU
ovgmptj5JBBDbP3MXYESM+xOtO5ABmSuQwc4AkiVBPOO9w5OANaoDVfWTzQA9Muj
W6Ut8k8JCP2YBF2fAbjb3a0d8YRGas0vN+POqb2Xj7I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 24944)
`protect data_block
xubHj6N7l6vOXOUhvaVoDFjsLzc5MtZcvQ/MLftifCyR7LumDgMVQCzJ4ImQHO39
G0bfzfFE4pfutcI1Vkrt6r3EE/iwlVBCn4/oe3VbCHdRw8mmOXrZhuRPKKjig5EG
F1sL7vW2MbR6bNfI8ncH+FepGmQI2WTdnX98F8shFA6fzoud+DK26rYT9DmanRYg
Bvsn/ps2rjMsQovMVWgGoFYBBR0Pi9U+5PCsDe4ZyB3O3fVIQq4ThB27p+2583ex
lmN5KHxlAjkPOU9JEOniIj4U+3oBtBbSlXeCVVBzKEneCsTyFuHj3rWNtXR6wcNt
xB89hXa+idouvkFj2YMDZDX11arOFvSuzqX6w3I3xJn6MGsA5OqU51PJ58p4HpJq
G07c/7NcD+6G6wL95dCm1Itxt/yLOA/FLY+OujNV2xUPI3MmsHc4EkfVu/lwMkLp
unHwy7X9mYAIgdMZnhO0VPLi2brWUqvYsfG8FGCHSbFtUUyOTcUkVFTlLablF4Kd
wLVb1SR8gYVbKiWzKNJSHKlTWpv6HhDXFWN2HhCKecISse6g+S2NvIp5ZE6anJcC
TpS0KplwzM9m+f+5uRigufdrnyfdpYqZM6LLEOmtr0fdrmieiVuuUOKMX+ubke98
wSHM5+MT9+EOgtG0sghGWGrT5gUZt7DFIGtYZ2Yyuul3+wbIS9e59iCXL2UXQwQj
II54d+4bNGjf+dJJ47IhbJjjMOX1XNvS5XDKcqw0Gg3BjxCN4KPfAP+5IBV+V0wf
ImXMqDg/lHWV/pq/E0rJWZT7toZ2uNid87Jo4KlVt8dzS+WzSDdeIh71ydjoPejT
6YFnyuzR7Kjyhf9dafALaO1VFQ3vyRq4M71L/kSOyIWOH1U1t0/gWJHnZRH+J+Xe
CZl4Oyg9aEzY8ftfYXkEm2Lcj9AQrtlx0Y+EnD5OOz7/RL7IKxZFcuonSqxE+DPR
EUKAn2Oce+4F3pvzQ1x7qzHdhF23pu7TxEFkeBzQasuJzIximj4XfQqNZJaZv2f1
qQnmXo6rcQI/FxZBAaUtj8O7HjQiC6Rhsl70zjdRz5GIB9Fxt/B+h0sKH2Uzt/o1
Ol8N6ZHNzHFcw8ChprGLta96Vxl8W+8y9/OtBZyandawxiQLYlgVhxxVQ4ge2UCq
PMXjw/kEplypXlwEiQTzuN5gQDx8ZhEVg2v307qk8ZvHYuxrbBwmokqWZgNdz12a
2bb9d8/UP5vpgKRuI5lTtPFSUBj5winkCX7osMICHZDhYSSaIa3BCyWdblMJb2xh
Wxa5JrVy9fV1xr+aPbwHoBVzvAHC9cqV/Kh6k7xifKyX7GWZyI0S5o+O3+HOG5VE
zg87o3RGD9xTcw3gRtbWbPkWJHKyD5qGsCU+DTWSF4smq4dYH/wNJ2t+KkY4hpcn
Tk/0im+FeYi42bg0YrXzT9oScgDfa7Vd42V2h3/PxVu+sDY+6cXu0PQuUFYfQas0
9eK/8VJmJSEznbMJvHkSNCvcIWApnRrYgzKHjsyWyamek6805RWilekHtk9HhW1T
hg20bu5OBC1kQf3Wgq6Z4gbJittKfR1+pAYunmhxwfLb2pwBB37EIX4f6VlX0MBF
ElufPWcKXfJQH+qugOh5R7pkVE7n7/bipF5DswkM9V1Mk01qga3AU6eRXbQh4hXS
WPy5Y325doU7ML2QtKpv5sXiTkfOhY0hqA5LC93n/77QCE5N+uNDFy1yn35f93gY
iJVAA18QWmAdfCgy1C78qv6zrgBsoqDWY29AOvYmnnDHnTkQviSxPlFbQXXdC49x
qpP+geZSQy2UvSbFcl8wUWDH+qyp8CtbB7ihw7aD+qhuntg9WkUCuW9m8TcY37dS
VWdsHNMEK2iU+crnJsHULWF5ko05kn+i+0segCsM0yodKPF/lsqOUG3wRMMs+jT0
3OzFbGykzU/qkLLcv0az0yH3C5CSVieSnO17S+adon9mxHIAxw3B5w8XwIfJGq3S
JkcsCrk/0FXAEwLCJc/dCD2teicSqf2E23cxXN4hb6285GGTYUCQ6KhDV41fPFUZ
GjXZw2bCNoNJiT6N2uVbtkOxA4FJZon7nXSIc4k3MaBBDeQYUpqH0t8bE5wS03dY
fm+ty+Zur6T4WGJJSF+yJOZ2ttimzN5jrKLRWbYwPAPrdWIvXLfD1au1zOx+yzPh
cyNDNa+FfSce2oO8++S2Y1YPgkN8d95nitK3wmnfoWTPLKb7PhE3gnUd75u9dXpz
LI6dyGPBGUglSJaXgSCGM1JxgvkxUO1iaqpMHa9AHD0/GD5fQCnkYTEm6LcKpPqD
7/K6v/FMG7ulXxOhl2bOVgLlGuv26RcbsdJWaUn9fpPLatFh4bnnrb0bjcQ6QVA3
/GWwm0YNUECTiVMzVYBlP/dsNDMSDpAL0riBVBBM5KExNpJo3uAW+oWiLh1ZPVEQ
ZuVrgcK7yV7BLyzK9cFQyj70lGHdNo3yYP5WzpYr7scyUdSrU8U0IukWOWmsdySZ
AEsZBZ6u2MEc3hsMelZ6ADJ9icXeDL26JfajGpYC3xFkbTTwDmKy7d1jkV0NPKPC
MD7WKgu9OkThCLWTHjzLtQ5sZmgKUba0gSSDNRvYmXWXkCR5vu8/Qxu2ymYyyMWR
nV5GAD8h4Fa/X2Bxmb3hOhIbdVRZLOz4ZPTxGiPGAJJvXvGdO7JqvKdAkBG86CI6
KLi3RJoUGsy3loO3D6SQSVa0iQl2CIgOz0JtSpuhjApJinv0dksMLNSGAqnYY4fO
3OfFOmt6VSdmsG0H2xrHjv6zZ+pdjUlpsqgYU/q4/w4yEGX/hcGvXzOSej01PpJJ
AF1kyJMF92F/S0CGsE2OMZaKPT6iVrPwGEdKQh4Bvqk8uX1SgznluhMzWh1T+UaY
N5vTq79HmKptbj9f8UXInAUQvXi1A/LdpLJ/HMeAxA/3lmBQMmC0VEPZD/kmaKta
ymxQP2FQyrUM8uIJpasvBlQkSOHD47ZXLAseHoAWYb8jeRtXcy2kKKC0wK97Dyxj
vY08gdVRIScTUbDSFphqocS/50Ve/qpBxivr4pPZm0J2r4ybZgzhVd3w0oKZavfd
BIYmLuqR4ef/OvTQKThIZF8JiqWyJ1Hz1+qcgcSVLLmCT9ozj8ylO/MOk19us7J5
S7jGmRJAYhFcXR94dgAnBSWXwuxDlXlvRjEzJVmrdOuro1ZVqw79Wq+3C8NLClyA
EUwHhnyp6OyVpFKRhHa0Kgy7qWEv33o294v6+1eQGTWw2QgjgEgPiiELHKYYpuo5
ta9ldrqIdIGx61ODouBvbl0s+7ov3xqUhUp7ClR0Vn3Icz9fnTUqnM9IKiIkJgD8
6m/ic20jlRfVwehMsYrgqCPS/lhdSbWxBE9VjLvZVB5Pqu53t1ltBWxpkKlVgVsn
oiwokJ/x7rQJ2rt9IYS/5JcQamjE9vpSus7JDvbb1OTghkzmPDOM48gS8a4vA7Nf
7UqxLpRUEezHTCrmlNoM9bki4+2gyVs1iAMjXBznB3C3NUslZWGRVeb0oLLh9B89
zdV5yZPCreYYOLWLEX/aPFCnlVUtVnWBeRpQVyBWVyMHxO8AymRlmL/0yclHUExM
9q9PCsD9Dtz3N51c7KLqNXNnkB2fSoHuN3jeIAw5tftRTcrkXOYfdeQLvnsPIr6H
IfA3zPwS0pJgweagj0KRBFrOG8MdVG/tg7mlog8FyEvvKW9qNs+tu0ncOwI1/0xs
H08pSQgO+zkKqvgFWV0YrVVpunWtjrtvBEtw8aU5wBnB9K5GOsgEcC54WeBAX58I
/cOBC7QABDMX8NtAyw2epT0SoRUSevlXmOwUH0vtLuAb1oBqG5Yz+iYYuEjmJ5YK
FXOYNHG5zBwA79KBO0ZIkuxGpDVV7BWPLfsZT8VfVhCi4KVhf0Q3YMg4UvTEJcAF
kDOIQmzPEQkeL0qx0YTrMJ8AQTUrF9Yfffk2hnaSICPBkvST6loUwsng1GFRB6SO
rbTopD1RL9XYpygAl5vJGqzVjIJgbdeC0XZ1Y2/5Qk2CFEeaLYOo1jZ8bJs1cjhv
cf/CM71AIvQ4xgivtaEweCviedJtJ4cIzIL1bHc5yz1RO18S3p0/Bp4xx0g9T3g/
macibF+ErfvK/uLS6ROD5DPE5y/DTej258npotplIufy6Mk4xWm5RQegfD/DCFEf
/d20/CpsMXKbhIGUgVVfU0Y7hDWwM2ae+MG1IrmNqzfLFWwPdQNxUXN0Jl4OPvOs
9GEzWTq4NcYlXuk2pk+8fOwh01RN3s7Bjm2yzggOyv+PQ/b8ZDcfQyJ5VDzTtshX
wysd4AbVZVjfXCgCZ51kRyCVw68PQ6su+rwjcU3HYVPGvCCW3z2AxmwERtiJX/vu
HcumKXUPIrGR2+OYo0Xw4S3FPCBwcS9tdZptXpeleb8L6cGp7JGAO7NoJMF0S9cG
B9UuqjFH7OWmEuIRkMhiLFmK4r26nB2SzR2QNVaR5I0ll6mzVKFl2CUC4SSQmM7e
w/KUSKEionH6Fsk0IlXacjoldChqzUkQwC9DAnRnlDrfpex0PWf5ZOPAAt830h8A
5p94/se0Js84KLyRDqOjApuJw9m6gqY5NTmQA6NdIqCpIA8+O7kQJi9785bptnxs
sEKKHlNtwDZBk1UFmKwPby1+iSKmtrOnBJqWe6UcNL3x5I3jcP1Zf520+upK9j7z
NqNNFJVmKWUp0jhgPk6SHdEUNqaDY/vhBcroEEMkqpYmXFyC33t5yVbfWmGUnHtz
jy7AjWUCxfy5DQxHilBXDoTEm93ULuyLAYdw1tn7ZIVb6qN95EwR2R29jEAoONhb
DIsx1TwRdMz1a3uqAvtAVgyo48SiiTDGtO2ph4uYSnMebBd9do+d0mozl1Pb2tUQ
nif4fqCmG3lq5K/ZokZq3lYLc2stPqkuq1J3pNiyFu4VVIn3ri3oCgZzrEhuL2pp
/Z9uymux0oFqNktiAIeGiZ5xyy99JYQS9tMSM/jrqlISvHcJdatQYMbMoKzw4YNA
lUV0LvV2KC/8WeMIzW6RAMFIv6WKpSldVTJsdNeIV/GXO1++JMOQPVuO2FIIq9h+
zNX9xnpgdpseAK4eeWN9QWyxSImPtYA6bRKSwvIB20iUXRfTKZfRfXDSO5uDD/wV
WyahD2OhYtPpe4aN07iKnhR2NFf5fB8CqsyzabxrCU2HrdjChsqVRqv001CgGbr6
9OtfUUm6pbyHRRkpnwLomSwrr8uHgc9T7aTGnZMBfWTmCte6kFwEZVcacDqyZR5r
Mn59jAO0tXUnD//B3BCjGNmrlXPKleIC40SN5drE28ByWOLIiyBJXcibxGXvlAKA
NERaOTv3RAx2NsNfBe6GzL3DNUlN/5ZpevuTXD6GfWRK/J69DLo481X5liq4t8j4
6QhtXOV2cN14Hj5ahO7FiZK0iDP8/mKUJTuU/FgL7lq4IgKnkug/lRmrByMjPfLz
RBQETn+kG68Qm2NRV0R+kulmd4Z6QKPC5WKBx4oHa9zk0hx2lM4NuCHqS5BcaUcF
EmpINKR132s7csKAMVTsyeCYex3B3IsgTa0uC3AFWS6P587t5cO9JTrRRvDa1iQ3
2KI1x5tPlM8AC4xV1q6BEfr2/gawrgeqOmnglcnKsW2afi5IidzvSBcRZWrIVweg
S2+nbSGGQK2Lqd+ATj9qt1VCspwP6gD9mQkVPvUt31KxqjOb+N0cYWRMDklz1ZYY
GXHx6rEPmlx8xmFK7BiQnc47A9XfG43+EsoIybltbmMMtB6508PlNK4c1w3emggB
9ir493m9P2/xJMe35LCPMB6c2Z+1889v9ZtB6m/N9A0QMhJ+b+oxQkc/kQCAdRxD
hd4rSM/X9hCRw51beJS+bkNvFKyizCw1iKpjzBZ9qW3wDSSqGe7lWNIVA5cm5Qud
Cjr2jQp+VlHDo6uvATAo1W8DMzyySs1jIIcvaEyjBUgbWiUEJt4W8Rh8m31ExI7Z
wjnI4DC4a5lB8QdM7wu84nzMfc0VJf5YNSgRwtFJIwAAcjPjoo8ha+Ci0mJlFhF6
97IlE2BDSRFDBy0aNNhw8ohM1kX8Dq/tcnkKuSoyXC+zvXOiLaCZr1rATKhIFB3M
aa79d9Cg0dkj0RvscrmkGtjOzgHlOQW33CPqMcUt+t7tK8DrDWojUq2Ap0DXf/ru
Qjvi2ndk2WZMCoLrr1FwpbIWttGI+UPHj23U979ebZLDsOZzQGzWDxCoNUEbn+FR
t4oDxF6CoNahCrN/EzMf1xljEUTIanCgw1ggeLkZ+WYPd9BQKa2agAKhTny6/SW8
IaJCfq2BnRv+99EEl+0Gk8nAt0MTCg6sMScAFB/DsnppVjNq506Yp3VDr3hoNuyB
MGTeZ5GKCP48pmZa5fQ7aBGS0IBAcRbbU3hxBWIqyfO/ICYqA7M3z3Yh4qDAooIM
FgscdvZ/i6X6CL4B1XJicl1pnWdEgtZ648bV6var8HuKhT4iXsLWg3tLGqqfSdYF
8XZAsa2k0EBOTd2m64ZyCjSUdrE4Y6/a+HbB7NWM+rrtoDM2sNEpA6UH50+SqaDr
Uz+UTZHbSlpettjKet31RTtGCfvgTSxJIH5Y0PDWJ3KjMZQA5ydCp7mt5yYnI9w/
Z0fCyC4pwhamF0ByEBaJ9gSFckUZB29S8HzE3XneRBdjG5hcoaL5KbeDllZbFqN1
7KyaP21qWllF14ZMh4xWqcNXydMiLF7kZOiWkfWzcqEvKAsLMBdxjWlaTZpPInM5
LLFM7T9xLtyEdoB0Hv3X+WfWg+w7ePxGVdXnZDj5/aFq1CQOHRxViaOykSbmmEF1
LzVXtjD6zJsoPSBvG3BAPwRGQBd8YXqWny6pj9Ws5woagpgsQlzwBYM0meUjxTjz
T59kFY+F7fabeFGL2NWQJsWO8hM9SBiJmiz4ToYz/NKhse4MfnsOIuS8BqI8rh7a
HXLbStRUGHnccAlTn2mc9esEhLJdRdh49mFhRjiL2R+x+4wgkA/usBKJlAheUWRt
66vMYi0N4cX3T7GqjAAG7eFLBl2OPp64VPofvcPPhcgHykvNATSlApsn1WkoxXCm
83gFgSrXedHxYPpEFHoAJmstr0oEb4d4c2jfmY8BEDqP8IJ2/bJ+etaS1imWW4jo
q1AtiT76QPQ4VsixTMxNAoBD2ChOQfAQmb74zitIz2u8+lgTpGH/OXuTTweyY9DP
NWqdC6q+r5f18rquOvHnZ3WYy8AeyQ7FREnvwj6+kzFRQvUwfPo1ayU3SztcTZLl
qzRXGNqaD0D7NmvL+EKxgs6wTzxC5dgDo9m+gaw825TeAM4UFIx4tJo+4DulSCfD
gwdqlLX4nfuw1JTaQFKUR3NL9vPPD5QfhbSePlmrrYL8htYSya9jN7TXPmLTW5+m
+NoRLpbRGTYCLZ7/zQJu5BT9EIapfXJxmox26bBRv+lPuxStuq8qe8DC+nfHJWtO
99c37u1jRY5I5l0YDdzTTc95FyoCg9DDfOC831pDPqsVE1gSMSWkI94HWI6zMgon
SxaOu52STFnr2vP61p+2hkzKlkdiG4sjb/FbCPb20uAXsGVyqMUHPs7G92mxl4Lp
Ggv2kruZnfRwVzuMCbV/agunnF2dSPkKc1QVXhdvS2PUxGfuU6Gk6SRNDlpZ2Pc5
vgfg3xitqK+tWuQElJOwE/pUpblVZ7rkFjkl5Np9+5PQWUpCG1C4c5r8F7IyC71v
NC24aqUvh38IftTjqs2mZc4RTvEN5aIoTUk+HUlE7Tn+IYzpOl6v9U9BdK0S6sr/
oiOx6zK4fLofVUUo3TMtGqEoHwitT4ZrbHj0iyTUlQtb8f25RrTL4OL5Yej/HX9C
wI6FjWY6jdGbGgDwPPISL0tsakfrn+mo/v9qbGotKoWqF+Wgd3RoRemsG4QC5cqg
KlkgActLHBwWaBlvB+JQxQbgaaYP8bA58+Wz4d5g5LVYl0hBCnMbRi5Wy1erU5Yi
LjglBkE+5uwVM/9OxNEDu5AOOyjE88B6EOvpp0G1zn3XY6qgWxOnSThgG23rhrB0
thNgl9gi0yrVnp+SZONUT0i3fZktRrZMFHi/kQVVCuJkxOm/2vovTRLutjfno+dL
DRKcSDl9BET2jmsy0QamTuFvQBBX0fenR6JJkBlbziMK7xKsiPJNAJ7az7QXN2N+
IA/Oa+6Zwu64eFMY0gge0SM50j22HFFsdYZHbBUOuoqatok3XAqC4/Z1a0NUDyEV
69OeVuehKQlzUxvjm8eXjAkAnUDLJj8HfXXbzXUmwGq+vR+pX81DwZd3EIE0hUcf
V3wj0fD9aJiTKWzpXkAh3ufSAnWm14pFui1BoPPBfb+awNOS49r1mLSafR9wIKZz
Qf//ebPFVpBouWAgjY1pHQ6/0uqyUnUiEabjuSbrIg02ML/xM3wgLrgB2PNrZ6CB
cOV5wlUhYQq9Ek7msnU/QnrXfs3TTmrFrlsvTMob0B18LS1lH9jxYwZTezcB/uaq
+meHRCHwf72KnFvPsq5c6cZFCKv3vFjQ+Cvsk2pFH40hZGx7EbfalUPcKa8D3e6H
T41r99bfKVhQQh4yOf3k1yahsrglQdAZsPZ9OPFq66y64AKjv/G3HCzJOMQ5GFQ6
rTxB0C5LFw7RRLDGGBn4qNnHnPpleE3x3EMe+ZKZRGoYjzGtRH3rr2x6WQAoeqOf
rS5p9lrA01ShbGGChzWPF+IGb4ybOSfrVmlQSPlBpVfcCyOWpwTp4/g2N4Loe2Vz
9dGDQyvlZUnUFq/3SkXjxDXHruGnyK0toUNdoFojqILGZU7vGoUGBk+JmyhJ41qZ
iBror+oeHBalbQW8qoqTj7L/cHrCuO2m/RzzsCPY/LOKQnS/dwoHp7oRsIIlzzT2
ucNCJt/ALc38+tfjw+kclfEZF5g8BW8oH0dWuYqoBFl/FC8caCnZ/dhaa2zGNkDG
DQYqOB4RM4x9jgnTU2mewYHlVpB74G7yZaIwYyFepDXwskfwkQUR9/GCzLnO+uwY
Tlro/NUvCIE9qXDTgtWn7Oxb0oUTmKEd1Ys4ZJ2lDjKcMvCDsO3H1gh1RX4eFE1i
8MiGYja/GygHvA2eSBX4IOHWRZj7zqD628iEPG9lm1mzNtzWTBjo1sj6yvc+y+F+
1ii6VHrqjCPidOJ8H9QF9+rXhlfau4BF99NHwvpSTa6BIuXCpCR+Tr9/8Hgr+qfj
QdEqj40FsbCSy9F+ec7fg01SeG8a1DGSYnl2h03D6ICsMTlMR+WmxPkxWLAb+uL6
fwYE7pXyxYkqb7HmdmnDzJU6V0ZowrKxRaEjoz4/V5IQG1CR8gmxbBWwvyMS4Zmw
hawGVCUVQqjXMMfwnuC2O8Oa1mv9lWudU5BQuINJ/D2yC2GWG6zsA6jc41nR5zto
PHpojes5x1gLOOtt41ugXpiMct8snNtCS+jJA2Ky2RufPuX2cSYIUGo5dzHDpuuR
/QpoTYoZGX1Uj/tYp+vJzV5N2VCbMC/3FQyfVsIUOdUVTtH5akJNKBenMA3rRZth
jg8I8yI7KSRfwIxO0Q69xCM/ekLSHQ71VvkRfWrM8U4VolCKZprIIlTW8e7NW4Qe
qJ62mffqKlsikEDt3Q0eUv6OTkAbuH19uOM35oFxncbJlSFXJ+s2qYvZK5VmlcsB
cOXRnEgfFsndvIzPVUex9uIR1d+TaGr4uBzozPGS6mKDrV7DzyWb1JcpLX3In336
sRnSR7s4K5OSaxQvf3oZVAGxR59kUIIkfwPqcxmvIbCdPZyXuBVGgfLCkQcovz2R
P7tAbWirQEHvKiQApaisnsF1TI1wXAkX0Q9vauhWsYUZfepAxGTQ+2RcHVZvaxB5
/2ivD1PaoAqKvkz+N0V5uIiEokVU6LgjAAfizkmnE3iggBxQ1hiF95KsgTRKz+9x
a5DcsjLPVYt11i4R2ZtGskDGl5iTTXA8KZwrmUcRyj+eG3RKF/FR4Fx7UE2GuDtF
XPtuGI7g/Awv+5jhpZqi9d+IuQBAoMXRSda0RbyBEzjLzv18yZmMpBtVGpHv1RU4
88aoQJKNVL4Jwh2B8mADyeFX2XretP8B32tywBWisV8hNiG6oepfoC2Oke7QLdFK
c1vGwN+27n6zXmuNuxUvX9EnApUgfW7q1EzxyNGnZzRFfGU23ruERg60wuP15i+5
Wi7irouNt97gGgCAm40IHXxZ3RNyKoBILuAHIBflYPhzDyj9GG1KF+Zu2BlkaHJp
auZPzq6Rf9nbHIv0YjzdoXlJK0nlbLbOeTMESDZgprhmKmlMsdVkkGQQPJddDi6k
YsbjZThv09hYtCRLUb550SDe3hddYfa31NVQ60Vn8FxQHFlT3gvfQqcnd3sGIwF/
Z2mxZuZQH7HkObclqhcwia/yB9pPvLzu/69vBHkJs6tSNHFYPnIayvC48WiHxE/w
9VFHnoW7Ci1ytfS0l6tkLqAlM81/RBjL4ciO4lsFgWd22XkjoEX0qg/mBZ4e+JgO
KsGXQCjyvUnWiBsP+UuVZk+hnEAlpfw8WXniywQvuI0vSgX13Ad8kWzoP3B3PZeV
vF/l5No9KTLGIuS99/DNqHSvwAMlF/LwpRuyiM/mcSEV1zaxUuhAGxctbpnp5q8m
hwpVZybBwiGdEkdNCDD5LRcFNTNI5xD4KaQR/WYUDlzD+ImLUSdxU2TEM1+yghfy
LBXnVoJK9i7U46LEbT+MTuKyBsCYnPH2b4BoHn2hSpPkgjwt3bAzP2FCp7LMlsde
8EwyBFYeCCG2f8+0NmqucWf4NoJjyWtHNnZJDOFZ3B8QvO3OaE2IsMXv3wMQydhm
t5rWS0uD+LSyxBbPkV2W5EXwQSygf/z++MIIk9e36Lt/jfgG1Qe3uBMVU2tVwHTK
yHzcvojGKJp9EoLcq7OUi2gpdMaOEXzU9vvPGLDIHdRwBrRyhDPw9f69eQrgc6HX
Kg1BqcNKMH7vNdLMKfYdtZNErcHFqYoUziaa7nyEMwxBfEOZgBCIoLl46Lr0oBon
tVNBzVSJf6IWnHeq+m1rDoK9vK0AoJRaIpgCJBraUpJzlJTDRJ+5wG7V1S+c+yMo
8ILCfEp/iH1GIViIqIp69mz65uG6MAhtUtk5apSgMbw0zGnKd1wwl9gx8dwqIxAf
ddWVrAqNuLYP2JJ+77gGr64xc9di3c1DSOesyh/6kY2msHJnTQfHxK7h8Gps5QoS
yrQ2zWPBesXhztegJN5nw6E2HQ6xHpRdokzJr3s/lIe3qSLdwFFp/zan6aGFzwjf
bXqgIReWY7udBrnKIsxPpsSkJcYqrUVst/cHrL8T4TpCZEUMqjnOTPxpVvxZ6Y4T
/UGOwF6eibd2RqIr6fZPDpHZRUo/nZdaaUApLZsZO2Fi6lX8m5/CznKO1XmiZH39
wugg7e/sXRu6zSxqYXHqICbGuLoz6ZhQvt8oN5ifoTsCGBD4qncOBC61r3weoiCv
cdX0PXHq/QXYNWiAEPbIiuvd44iMZuMGWAtq5hxEg0eocBA4R+lM7aksl8+VbmaE
I9YMr4fiyypQv/0z4/Nk3D918zNbgLJMvbCV/nV39artLE7ejiPrVECtp1aTWBsX
FMtP8oJL+R4/Av4jDO5a2kfMytzVbwZPmXJMPo/Ph853wNrM+OAzWLXzGTUf/uv+
cb6QLiaDz2VsmC97LMooyyqtYRMZO4ZUz7f1LWmBrrJDTpk2MJ+TWRpASULpjP+B
0EuOy1ZorDZ8Z8CXjxIDmd1cA0zqDsVTIs//7fQvJ70Ty+YDOr9qWbn11ENEw7BK
idTBATRcUKZvEQueLu0Qn4blE0P1Eb2LFfch4VLr14uRptKUUi2R1eb6SB7PJ+c/
RIK2n3u8XgpxSxrWNgjblcDA7Ecn55dmOZjYTZDuZHVuLRF3ze7QF2h510oFk57S
wuGiukGmBoL5ZrckOuTQVqmHdvZS/4OBPT402uI43vBTmTKrGkCCjDEWJOAJI4VU
VyeX+ivGEm+CZ9IWz6kEZvbkNr1gL5vRUBBZKWYcZ0KjAwSqnIr6SiCpIt9UhsKr
3sg+UrcOagdnCrINvOoRFn5cpjmWwDHmkuwyGMabmMLyHFrZm9cakyJYsRyLIHsU
TqsKDEpjb0N5q6ifzTClTXyvNrYbNB9DNm3XUBtWdKLGkzmMZj2WVbGRz9RZLEpN
/PDybiOxSjEBdElURbuLlHD9WmwMW8FRGQCFh2IkkRzno8LYvdBZGQa2vpFokt5T
rNzH1SJetYZgp2IpkGUAzjf5mLpcIfZ22EebwMmUVyN8V+FFZn3iFwOX49YKfJib
1m1a1jXfhzBhqHVronaifkDfRTxDNJOuhQJY0RttUI1aKZIgXAxyLQ4HTuuejHJf
JPtBsx7a8SPKLNA4TbeQIV0U75S+NU3d/gw2rwR03pPFLJLjmlmVz4WPIwq8Cmtp
yf7aOz4v22e2BuLe3G6X/R4KCgx3CL/DJe/KlwS31+EJMiFea8q1HiMbcsqUlvS3
TlFnWv+YcI+96HcBuEpBpvAjRluXMnxlSZvZvIO9kNs52qBithLCQ4lNJs7gMtFa
rZaXcKQkhVy5N7fP9hCSIC/YleqNc8cJudzY22Y0OWZO54LroqxhQuZhlL6YnO2/
OAubyct8Ta5S/s3sZKfPlHItm0s/dHli/HxQ76XecRzt90V45PHoZkrumPESqMy5
o0Hl18A2VVKasAYwf5/WWXhtOnPfBrTMT/okIO1fy+rDjwrezgUTC3oELFmYD0LH
4/y04WTT/yhKQIArNuhV1dsEY+HTGqrb5ccVPAaW87IF71q1FPN+npa1g+yLb5Qo
pbc0YBZ5B878UFV9RCqZvfc/4cu3pYxSrd8LnfP3oLlHU8WeJP3CKe+ytfGv5UIA
+K13ZYz+vkgm7Tfmu+M9Bb1guJLH84FgrVjbZorHelSs9EfvnB9mSS7wefx0WBEV
74wIFUirK7kbmLBcriTZcSa8511Gu/Bn1+AwkI1PzmJ7neLfy2ldSSzZ4u4BNF2E
Oxqssb2nKrOS6Ihz1cdOC3K0vJrN02x+50MLJf1vE5zQ5VFu93mpxdnLwYiTvpkW
v/M+ZIuUP3Nxg2Ub9Kt9VHn2rdLC+ssy/HWOfOtiZZWqiWvuJwQcSzvn5TF2esAR
o2XZABpGwjAzKg6Bav2DDPEi3EJKuPGxzfYGOsx/RvMf/ml1t4QCgIHT/Ga4xUWH
x6iWXjfq7Eit8l09Xc3ucZ0cPLL7ckeL7xGkJNX7pQN3puU2olDtsACJHDFB8t0q
drYWv0KZBs8icssAOt9GaBDcH55AhbriDAzlv5MdBPHstPxKifROOmED2g6su+yf
tvm+SqTHyGrWzJCHfGQp8yNZ4Ft49K7W/7Aeq46HJfq73ZqGguyPdxbOOlFrLEWg
QVZE+84g0vHg198tYdrIg3re5aEPpiL9JBltiInvND56uf5J2kwOc2bV7bJ9PEZu
hXx4BEEf323aO6Zi1ILHMFY8s9TeqhH96mnl53z+h+vqUs6yF5mog3dG8bHdMAG4
2tFUg5p4NOtnKcIJluq83zX03O6TPhtyh+mMIjhy6/YwZRxtb5gLObJJ/Eqd8091
hLgxSluIRT/wDn4i4wegt0RdPOOgpO/vPY8yjFnYQGAhOKlsLnNtCkwbk/OyWchx
4+1JAAswM6LGtF2g2Wm+aaFM9+KRaCUKB1ANWgZ4mgmiKS7D4CZWR3YdAzzZp2/7
AzfpjihPOMkolqT2YOWr1s7Yxe3SSh1MbtywR5UyKZYOG0PARANB1QrQJNvnYGsZ
m0Pk0YESlz9VP+e1+ud9JverLefkKboGUAk33qDLtWdeNlR8BTjN5C1Aq3xxkSar
bJPkIQdjTv+zPUaPuu3yVGGUmqsFk4u1vRJ2TpE+07CY86ObpzhkkGKD5si2IiSJ
6qVoaVPMlWVOWhI61LMykzyH+GNZ5DR1XMR5r6FoyXp847bckaz+2nz0JY8xEDlz
5SXbUTxbMFL3qBTSKEE4E0JjFMo7cPHe0cKzn1a6pr4sOBvz0NzSXJQ0KQGNNMyX
RDxpZO5kZ//5nV5alUjFOqxPxFhTZgOEid27LV/Aow3ytH2DniUPNu7j+tse0A9i
BXU+NBLFM3V5Biu/hKDt+wgRcizO0yfAM2bYHtMUokau+ciU1Q5PdC7/Dpb/tAAu
MNtD2s1Pvqb5sD0cFvpf5Sq1095kR1uXl5f7GMU4489KFD52+19MhbHdZH7q0ScQ
4/xD+Rq1plxmXx12FYNKQqiJWkJiPLCZiy7t1iAXSt3J9jVTcdi1Mt4AAYIguxCm
y/zyZLmHkSxMPdL0/UaT18BMDTofZxlQRwKgbypK0i4AyvbC60J2aSL0rzrKVa4b
pt53q1mAdu4z+YFZ/p1MwU8Zvrz8vz2nbQc31gxFycFF+EdWqjjqYkUghAiJF+qS
g91DZCa0Llnd9AmoywtT2whS3b1n4+suZF+hxFOQPrQ9V23x88b6hCKVUg3xgQrU
QwgoMRNTbPCZ8z5zlpp26klGkq19OIztbsQ42rvoKwjhdDKMigXpUiVXsDpfqmiZ
n02FIfYCfVQ9CuaE92cH4fTwc60DmMUZvrwL6y39uK39ZG9yGCSl+radwe86pF48
yhg6F8vd/RDkCNASuIYungAM0wqclMJeOhzSovRqtKkNpbPe71OTZSU32OFb7vNS
J7xoBVpl5CLvcAhdAxuBFFW0YDk27Iw90LPEuT9ORQAK6efuU0jhVNApfeTJbTwL
K2XlJcfIuTFwR0eauDLmSFzuV/sIrhoPIMCmH/oF+VwrhVi2SpTucj3hH/jR8gY7
7uVL2HLCCfTHv9E8gIrPbHqwC8YFHYlqM/z1mpYaZRq5XhN9TY6wS3LFJkijncAO
i0BXtYLWf1lG2jYphYft+3dNMkeXL0KehIuumW7G0a/Xz+7Til6SRAGtIQFTcHQb
dQBMRHldbU9rhXcRmtr2pmZdqbtiJa5moZ1lt/v84iM7Aq2J6iiMNIxNR8vojobM
0vlJTkkmy/AgewqLbvC7enTqBMYCeJTiYzZmHG1+9/r7DXAyrVtymQPhTY8CWczC
HHDssO1Cem9xSDLzSPCn2sBgadudLSYSntbDLk8cQXNfjc9q1m7G7BiaHppgAcmL
3yLlt9x3pXfjnxRfy6m0k9kDeAlewp0AyPbdyBPizwrdxn4mLp/gzOf20CxpiZld
WVWMJe94ZkFuCbYjE00caDh3G84rlfLkeNTx87WTNSnw4Y1cTlRrgL0nEvV1xNa/
7aka4x+F97pNSgQxU8Jc13Zqtl59SSlSrd0stTdLyJK1/RY7A6suixF4qLOtJOMd
AdZX2cQUZJV54fxT+U2364/UNbOQj3uGsiMR0hLI3JYUNm0rtbSy+4y3xRA0om2w
Vte3o21dSSm5p5FRmd3T1Bui1p6zbmpb84vRbT266vl8fvdc4OMOuh1G9dB8RovB
0L8BpnZMSwaYhQEF0RxzXfkQQVsTp9rhuz5YgJi/FUVRiIpHbD14GVAfaYij/fH6
2l2yvtzE5FE368rezfsGsOfbrUgu+BnF0+iOLIPF6rOMax0AcR1umWGHBOlo+oCN
nrjquTHPl3fYFs1lB6r6BJJ/9zZxgdaeCLMfc1GHL5E2H8c5BkdhfCAlKxvcBsQr
pvAPQcSr8sQcTLdaZVY4pZF20cHIH67YnRF7UTgfOch2llPYX4EdvkyqE4Y8jwHI
9FaGrctY8W4CV9KEjaYAZmhD/z9++3tiupLThXpeX1PZA1Hiq70GdbIJOAjBMXzy
SphVZNKFxSskENMcoZofMvPPr64oE8WnBOJD1w05D5aTzuBO3EFjQHt8RfmbcgMY
E6XCngyZNvaTiEDc7/XKLypMzbanmRlGUAHMCB1kczU7MZprbgNsQSOZ5y0E9Yiq
hLef/o3+hc6EqNSM0QrnASa8txCiZYztHIwXvSiyGiebz/iEEVFWGLVoAW6mtrmr
ntvfNjrDyT9UXp2vuIwUiZrv2eLsYnlgwFg9ZOLy4N/BXNyVpn9ilipxOELU8z5B
ClwlALpy86HvhADPyTQ7ymKDBDrZVD1KGUe0zv971o9whxmaoSuI8Ikw0qxKTqWQ
PpUDHCZx1ZgOxffw0iuN2EtYoClORr4p8azNXWWRQCnPUUVz1nN1CeqQ44W2pHog
mr9lCvqssFB6vKCr0E7eymJEDD3A03V+ASXQLM1kvRUIogXgM1fyjcVFVErDnwZv
OoFYO/zX/FiEMw6IGwfdr57vpwhb5BBw7gR5i6UiiVSMuQcSpHr34eUwI+XXWHAa
SEAui4+SvsgAK6oTGDI9X6tjxX1ESPnmgMhSdo5BRiINwyrq3RbOrVvCurwQ6Iqg
9r/5wq3pVHM5KKJmPqFpwyTlNHgGU/bxHeGySkEnCSRtc+JQ/7/B8wYg9JmTbY3B
SvpnjtWKueMTMpxCA1sERNE0FLeK1nmLeVsVWGqhcDbudiPZHKSQwwz2zUlSPnqr
WZxHYMRLUEjO4a06VGq41cPURiTHklFVb/a6tezkIgor/486CZ5u/mcSi+sZckD8
t2PF++jsZllZcQJXl/L+V6ZTYcg7nYGvkN8NAV22S/M2Dl7V7e6wZc5Q80QEr9DG
djWDvu7lRLAaze0viNZMZzUzAmdov16SvmC9RBs6JSFVRPBJEWL4ptevAnKXu0+l
x05i/aHOL9AVcrJaSCPmH/4sSwYdI8N5G33egIKwE3xUL0AfqqvLzkl5ME+YjSyE
wIOgzNXTcuWrL41gLjBgUaEb/Hwf8962WOmuhEyzKPcnYFm43G48/wMyenW2QTja
W6gTYokE0NRDJ+JimrdXkfI3fb6ZVxf+NaJ5zYjSEzgYc3k366Us/fLNZ+ZLHial
ctIF2ZnlXbIvcJl6sIOEAXVAdVapCB+GA+wnGA0aAA+zGGJrOP8F+eiSp3oaKLIB
GmvNUmOlk2i/mSTeUcAqd+r9vYzESaHyDqnLu9VMkKSxreFvNck7/BVvsuWOZYsR
XVgZenb4ZshXqindEr5JbfHkdfyo3k2LEt35l3KTrLvx2XTVIO7T7KIAN8hetisU
fxaJA3p9bI2jsk2sXUMspIslI2Hz1MRfQKUxsfKsgwMy3LIZxTqBU+ADmHiaTSAm
1w7rV+8r6CuXlvU4PkhU+sy+uE8a6cVipK1Pxn3r+G6bUqdD5Y/yjtRsPqUwMb8m
TMpOmlMbcl54i4KIAAZaM6juoDxDMtA1GdvG9Ilu4pCvT4/0CuRwSVM2tp2u+Ka8
WT2b/GXs+1QfzW987a/jevIDQecKqrJjFng5PrliK1kPGU8hg6kw3qE4lR3eRNfR
16bHOrBJ4nn2SgTpYbUuCsqI46vxi6iBgqcF0KDt0/ptMJ9vhIBWNs+f2+JD86a5
Uprw52PmIkGQRWW0gdvFZosXwAbRKPpV25YKAVyDfWL4AXsiyaMyi7cZg2H3DTr6
truGxIBwfC1ND8zalGa2xSTaF0K5sOQNxWcogS8enl6z1/giXx5Y6OJKmVboFACi
6egFNEfAfIFR/+76jtVRDm00M0kuv3hVXLqpxDpyXZf/5sj8Z8fj9c4fxTq3HNWs
h4El+I8zPnuPwCvdAaECXHdEXQXazPuPRAPQyiW1IXhLErSbgxl1AeFWEIFB1n1B
m0fbti4j9g2H6iUPD3R6PPQIRCbi+nv4G1IO7ftqNGMlUaghnz4AHayFvXdIGRsb
+FWmwPCGZFnx1pkNkydRYUw959dZWQeWsrjYrHEpQLfWheEvH8lj1Nom7hrdmA5A
NIi48oNu/oRE8prRToKlLK0izL+RE8kb07nIe+SY2ubrmhDU3P72itjeG1jxiAXq
DV0lNWSgqFjdCuDSpXLlw3c6RfZZL0X6M3Mb5yYJZH0vQuLf9p88FQoOl8VQQixx
/zchBkK8yipYTU9dl7K5xhzb9omPzJWD1ZpzW5j9vtm0YbKDOisZgUruN8mfrcqT
nMGyqjvrkQM9fb3SeblUWOha4E+AdwluTATUyq4DGzU0AQ/A5HETO4AejYaDrSME
Zj2yoAPszpXKBbP8AWz4HzTEpLVi1ZTvPmsyoq+PR6sCQftyCoJ7QntL5xnlrB46
5/4Gta3c5Rh3qdWnD7S5KYGFbUf+uSft7sUNQZXrdPkDEySVlyu48z0bAjC5l8U/
6SbmXLJhljc1EFcMAsxDitWQQCwsygW7afB2xzXk4zmEFuHWE3FMO40avhwUiaZx
WZEh0dQnlRRK2jI37Dogi49L0iM+8LKkwWujIameUbgZ56HU/6bOlZPkaAnRgUJN
lCKbSXOsidVh2yK9bMAf4scmCpXsB7M+rGAhFy0SCZ7usI4C5EGKkQCeqboLRZRK
OdK+FBJbQHXF8JjRalSRU8qS/qPJ0blK6oGNQ99ZHaL/zsxDXqpvABU84cRNTCjK
2FnyyQgGsV8F/5uBpd1DPZRE3r7yVoK20WV25zTcF3EdECkRRyruKLIECz3TRbvu
ULwMTiXSQ0YOcze5mKgMSaKzJa+Jg0p4DMQzPwwnYGyawyu7AlrW6goXZ0qeraXQ
z+noMR7m0eSFP+izyqGuiwpR1Xhtla98pKL1XKWiMqIMYI8vE7Cdj1NU1K+sHdFx
N5d4BK+lDknj0SQpJPLRzelw/l4REs7oXOSOqKX2deLXufXhVjm/aX4YdafqGe6l
5owidLZ9T5dZVkGakcutes9wXVIB8e6H7TjJO6SUagFTFCImTEfxcJikRXUHOfJe
Zomvx9NwoBjB54oEZvIh23z+is9v8TYjQ+z0YTliX/sMO+HlJO1wCCu2L9AtRAMU
iCTfSbBuJrZxwDPyvb/GS05YbwHPUkyS3hA6ITmku6Je0Oby5nl8xl5rB3bfx3jS
yJ9PNE3NLnyowVYJonAlh/fFcGqCpPJvupMrcJLh5r8SqKALriAW1dYbalYBo8Zg
DRtklrNKDJmjGqmj4JYJAN6aKj1kScza/5oy/T2xMPVzR1XgBPl76kIyrXDqiOiE
VgzHA5WnzINnXz1tGcReLxk3Y+jUahmkXY9ZQUVTRjbzx3fXfZh9yIqGc69YetPC
6qbJlZ/c7Npz8VnhZny1vgh3OXN7RTzbwMgjI59KC3zHBooyFGGteNiPmtCURIcJ
GFkqfnRfFZPhBs0jO5paVhCqDWXw0UMg6OnADVeYNJRlHQ50L5FC4o4tsTcolFw/
7LqqmHoGaN2yymEcELPf9kH/HGjplKAKKQgjnJH6EuJjG9Jzd4ggLC/gFC6MEEzs
bfEPp/hfNpIZ2L42DHDMY4VwiKdcshR8Hd9G0HBvBrtlQ3b7Chbw/DSwDomuCoRu
Jn5H0rGJ6YbM7xEuFy0UitCk166RpEgOjnwW2PQmKyyJ51iEd7O7kVUAmuDo3fco
T0egwJl7KfOu0wBsHvSQqF882n4s6LlfcgbcXcIfMD6848CcQr67sBT5sqwv8Rh/
Lol4MuYUkJM23VeY+jrnT/t23wN24l7lG7+ljxt8snnjS9/UwcNpkmYhcW+c/h2Q
TC6SJxfheuUqG/2vT0e5Z7PMtrTI62FupIKWfFkfXhRkkaAf+wKrFCkGMuOBLNUo
sd0LNBtGu4KWTuuNR0ijMwCRAs+BOgZh3eCNatR1FM7iWniuIp8zH+UfGb178Omc
xXYiihYDbLsFEZbz33n4UMm00N+CZDZtQoNOYbNXATYYdPWywMqmIluW9wn9JZ7r
w3TE8yO8iTnzS77V9h21O24zBDfKUv6D3rcYew5rpYmv3WZ9vyEc5avW4NP7pR+W
pKi4xegZwciw/Vv0W1DG1ZbOttATPvq1hoUAYP3mFdfaifJfkUKQeMmpWVbHF65I
g1/j9viTg4GSuLxd4Ll+C7NTpX3VJZVzSSNlzSefz6sRe3TelA9ULzQMbNKykRaB
cBjqNmVvGLjwliWUYJaQHcsFs7UjpWYwK4yzQ1tL3x0riCsy6YvQCXyjhtFFWp5Y
QRdMMfEMCBzNQvn2yjUUtRvWmD81daKLhmyDaK0fh7rEuQoe9MSHI9hxSPLgH8j9
+m0XnSKyYHMAyx+bIn+5cjX3Z93UA8bQKeZVASpqtG25+YnKsAiL+qBXB6i4tSIt
0smVW/qUsMpzITAyG0nP0syauM+1FQS9OdJMy8eW6OdJYzHEb1y2RsoEKd9+l5Y4
80OlqVQny+1/NTOJArz+JjzaGTktzCW7BPpqeiR8KAgiYgkz25szJO0KkiaHrfjs
r6BznlMreHiuV1JkKhedkrbqxwmOJRESTm2Je4Hx2x9/u0k5oHsZUlWFC3750q6n
qoD4DEwZvM8WNro8yWuKHKBCtcD+LvPxl1iTRxASgUv+1G+z56Olm6/BiJisCRf1
0o4EoS0HyJMEQjjPuUYpXVVjTf4KPHT9mWhA+Kfogo5VaQwhfzR8AYTbeGE/Wi3A
jfVhFRh2d+fIsuHhxsIg7Q2CpmjrwkWIjD346ir2q0fqBF5Ay8UTLul1epB+psY0
+But/igzs6F/cPcJ1gmbVTAceGGx5oQskKqAY7XQ6oCaW8FrOhse396k/qSq3bQN
a5xIM+vayFFXqIjBw3S25gs8N/+rWZcJrQNhfa4xuiFpERlFEOmR/CqUg4RFG8cd
4OXTbLvtOGEbgqbEf72yP0sQuBmX16iObi0OvrwLzFSKgWbqhrA9QNkz1lybRiNU
ViRIuxRYOIeaNb8NMkED9KMPXsdFqapxLmax2xJbbwFuU7Zu5D/WMhMifupJLDRU
18McOAgRkuV2aCHntVli0nN2wO8HkYw060CRR/yMofxr6zA9KHxiArhiYoQ77279
StLNcBWOOPl7yIsTnR7sahMqFK3LpsxgKOdNfEC32KabUpxXc0G5gP9Oi7evytYa
dHqc/hey3uDL3HxwGGLBrMJmGjGnTXWNg130ltU9z6y60rWHkORu4ZwMEREM4geU
Gh/Bjw7tiKd54eDiWu/gX7i0VmwbBzjnVrOxe3n6dZ1O5dIW+f/+4WiYN8zSO5Gn
qcEK52R8Tu3meyYxenDbK5H6paLFRKlyng2qC/ni600GyKwfdFC18L4h8McK+tkC
/yVa3swlRMtBakZc6nv5n/D671YtHolBaOGrhmjp2kmoMG4teITQTHv0YZPb/Tt/
DvS30F9OXnbLBU6/lgpZh+WQpjBDQNy+e4ipTmY43Rh88nZonSyIKGpMEBTVX9dp
DZYxcUr4FAiYO/QYUnkwKW+5q7EXzIQYn2okgs8KgKp3KnxKN8k0kIuPci/kdVvE
H3YiowGYVqn8k/0TFd61enKCQhGS7CM4NRIELwxN1ybED4mmmrG0QmFwz1tLTxO8
ywVIGNeZ1tniV6XKMBdZwPYhhwtN8sOemy2s+Nfpt3U3sbI5XqvvF+4ch4muQJ07
JLYkvcUJVigfAZmbWVhlPzhrs21eHspyudIbrFKhumtSvc1Sun2o5t6JKjmTIAzO
Vxg5Pe2JNrjRo/ewe5mRmhSGIEHUC0jQS/iuH3NykMs8r+8umbzuNhFT4Z7fP4qK
ujJAjF9jzJgYPH4n4wfwFrk18ypQT1lUDGu9otB85IciJiekZ2SJzjw9MDbr39fz
CSq/ssPFcthd9y/d5bzAE5TKwbAzA5c6bg3DgyqAtZXS1okk5eTDg61gryZn2mvM
TGxm+8/qhqwLR8ScP2HRzq2lAfD2T6K0WgKfgUXQ/ZPRpUVCTqeAzwCZeKylUyFu
dRyosFi4W2kDnVvD6c4VS8AKQDsS57lhuW9EKMuLWS+dxGQjeyBOGuAsNYWjl5Ac
7lRjT6Y8vnectZ2FjkDEEpnsh5ZWFkCtI4Hl4F8LP7lpie8Vsq05cBFpfcUX2GXX
YXrT9bAkuJOTwF8eLsQIZxdOcHednroV/D4Xmes4Sgc6eFPifQWVcKTd5qdIAsdY
Z74klreBqkZJWjagGi2JsGuUfbSAqS8MHiY5DOxfSOIB56E2W5xJLW8mEVkUJyu6
ds06q2hK3OcbdV6TVXkbRr/6I3MvWijb3C+Tug/2vhhqtzWYlzvjJoBPIIbhIb05
cLfAagfQP160Tvb9nh5sUftr8edjgVMW1yWdZiEmJja+uA7JlL8DjeN7tqmgWgih
fd0Ni5nXD0IR+tayusX5Uzqn85LUcG45oOKOkdcnmuN1iO3ddhfqalZx+Y64YzXC
1AHU92NdKRqaZX+Gh1SfCOb2q4yAtyw2XCx2su+IdIqclgXGKy1YgOYdRsnZmqV5
mARToz0rXV9e+39JF6G9XBFuSSffH81Yq/gzncfBsOVjQN6j6TVSCAWrzF3TS6sf
FZoyBa+hHOI0yHlcRfw++tBx2gMGQAWITKcacLzNMUmvPV7OHdWwnZIFhhiE3m3A
04UPBaOhRr9nUeuLO7dpOlfTydHFdbGXz+H3I8IYtaxQrXtDbzlSrh/eh4DOcJUf
2gHyFpdtsZTfwyKAgVfJeafYfl0EOYmK4fwj0GZD6zWJWJtF9U+arpx/j/fTV7Na
54W1edlRRkw+T+Y13iuy1uiMzXl2WR0mpECc6kfq/irdpxfIqwx9sSOn8OPhm3VN
sEXn3+BLPMiqmE8d891gE/r51AgAOibSgmkGxc7kWh0McIFiNqiHWu+CF5rKCWcf
lQySyPi5UqW9MEgjwvWTDafjsW96i31/9EtEuB3rb9d1dXBvGFkGv8hzqn1hiXuE
NXQTfX+oqhC6G+P7UnipZrHhi6povw21o05TG3X3ywtrPlV+UsIMyip77hy5oCE7
636vSZu+ADoVx5TGG7fwr/jL+PXlghuk9W6nm1/uIhgnNV2PLEDKL9/X4mUfVx09
gJIUQaIENr1nY13SD9Me6AFhWuYQ4f1TZYyrA2l0kwYnuIxbuz70WnI7409kuoPh
uh9oQzPi34sOdXPH4sf6lulbaqLB7zLnQ46w74Df6jiXFtakiR4nRLbSikifvqRn
SBihnJQ1ZdzUkPU1JbyMuinvgMUfsccR8Mfsg+cG8v4h32ICnq7mgtNAGcZeHnrC
5o8d6P3D9TXHnzZFg3OpQIow2gKzlkQTDMhCYInp13TpbjJ3O4bNiinLKW+W5YHD
gcF6VKPf8tkUgDYRU3wGIMfSxz6TmUAtGigziM/tiAbIKpJn+8pyOoGYnn1LOyHO
pJF2bl31BJA5Cs+XnBf1AcqDu0AawLYx85AZlqfzdwoOFSeTU5D4xpI/uLXVdVKz
qN98RwMu14yPTFdVj3g4HuB6YB4PGsBW5FkQwrSaoMN4PjoujGgtDe9z6s6SW19I
UUbc+zXTPwzuUyWcYyUvdJmskDhsgKrRCHs4eCik2wVSn27OBByyux6Us0yy45Wu
pZBtTXj4ANdKV6MOhKX2gmIp8IJ/yEXXPf8Rnh2Bse+7RhdnhkgHd+WGegsezuZW
fKM+CUdWq9xYGj/M10+3YfMvpvWv30EUQA8Xkp/EnpfNBh++fEWNPvnkpMJyt59B
HK2unZ5l4rYOoX9f1hBFO8N1G1jJ0Y6Yfidtj/lrV2tJm6ZzdHS22MF+4g7JDodn
FoWMLCEwYG5+dmy+/MvkAX88ApDihOxUop1sK9835sq83R9/0Qx4wn+plPVsQ9nQ
Z0NeqyKIHW4uMEPw1+RIqwkN2gnpPq2hy46nVT6DW2DoJTqVkguzIhJgoDW5Oq/B
HzDa2YRyxFA7tB64mLeXZrCYaYOFrqBzBz7rZ0gIKuK7ARdLNmdox0tAOC6BeKAg
y1x043gijq5B3yQOUWWkvKcmuFelZJK0X0mpVYxlFN4chvlwO2EzVaQrPiZndXAO
BqTtS8oky1qJmlRd0+LrHh5QA5atdrSKF+VbvJ07rnWcDbYn5ZFGs4qP5sNNQAO/
A1Fy4rXWnZPhydLh3VvE1p1Bw8T2t79K7QOpINvyDJcvfBR8D5RxAn9K/WxgNxql
9xaqGYqpx6IINTSosph3vm0yTCfUbjkGw5T5Lb4wtIgERR+Vcq+MsA/GyLmi2eMK
4B/Vd0Dxp4ZyxlGGHKLAbFLGWtPy5uRo3DUTk4bxMJXKJ+4Ad4N4wR88GdEp+pjo
a2GlnZVzGG/zW2+PmcOhD3XXnhc1uUCIiJD8tAyKnLiB9MVCMKINruXiWcEtoHyC
MoPDQgFNCqLSVfULKwNB5Sm6MqQ1v4x3+upSOUfEl9GZxvz7RzlpJcPZRrj9CXG4
3oBpPXcvvqbycntjlhmrOcoA0cRIJ524lD4AHsK3ZjUsE5574AiBE6UOOAjrdlX0
59azKWUyFd6aEh6j3fb4OGVhwNaPbcepHJmKhha3z5dn/DAuzLV/cRszm3AWZgIx
Z3nC++9cwpJ7rlT0GuoedmD24pQ7i9IOxPLl7Oec1hswdNbNpYJBBa5aE4l/5sHD
KYMQqa/+uWaIMpoWJP7EPcxFkjVdt1x+gYXR0boCvY2+oESjxia1CtOkW2GpCNK7
mvTmbp/cHStcuNZYYQSnXFI36hQaOjn59nn0DMpz5XFeqdH5mT74+TASsgwwPg0s
tVzJxAV2Oxf+dSXDJqEjHFBktbxkh6uIYM495RAHSw7QviealIj5u4dv7g7ew74Z
NNa5NF6dM7jj36LAcoQAQkU0D4pARgjrNQ5oTirkarto+ZKQgtfC4YGKdsjm9ihq
F7ATdYQ7Hj8fIpSAslDT55VFfg22HQn8Czq7f0pR6hfBPZUQBf5502NHSPjQvbG6
WLHJlp0j9Jg9Ja4WWGlwOOyKNrEs2Yu/8phQB+Yty3dLh0Nic11ZGdt+IqNFmVVf
Tc0i6eEXYq1R7vZ9pQ0mxEb9wC2snRFls1DqzfZv04tzBJbQxeg+uec1HPXjDaXh
NqS2ZKW9opLcOO2SavfArwaJcEPPef+0d0LkJVhIXVwYvxhvh9oHoVCTE8GBu8w/
RnERndJeBTjogMEkCrsLBBca/ZUi6YyNV/EOjEKh/gM1aZ3X0t3S8VJ905y9yurO
ANId6DGySWZ8Cxd4A2l2zRXUSU/XjuXlyf2QmVg14XKMR/ErVV6NsvBvUw6IStpX
JW4N6VBozMCoANNYA5PuRLX5B1kWB+Hotn7y7ks8CVMxKPdNo0pzp8mMK4HQfnqU
BkEPrEHn3gFH3YzltmsCGNZ6Nib7X0Vjyt3cQ5hdiqII2mNzKtEm2CkF3Rm++uYl
vUmbg7/YXIRhwgVoi+UQRynXp27bDJd8m+mt3tyWshwrN3mGysI81xVRPifSrMmf
5OKxyh75xxaInWg38Q0d9NqLhZ58eXZzxgxSHN+DgR0JYGLVzIrBLsFPJU7KWr8b
Ze8rKTDYrVDCH2xVm+7u9dzlnJZ3gP/qEfB9kae2vxNAoMb7mLJXHt2cSZGX5Waz
gkAjpCkGPcxSe+dE7RH7noPAW1QH/rXp6sBURSxbO3dPXCqiH/Hps8CErVzxyJ4L
9T2X3m26rr08xOeaDF+xxFFvoORb+lzfmJ1swWKyL23jok/jkj8tXmaBsTWTVg47
ISeKJzdJDKVnuGHmKqQw9qRh+otKBhFqyZPWfxCiomVNSf8pZRDHS7uo3BgEOZ/o
QbNAJYgIMBmgY8Z3qCRE/q74zaYCl3pW7rnXIXTsOB9shBOkyP/rmut3E6DXhG8h
QOQQnDUVElMi+GL1IB6Cq2++YKKDJZ+5u5+T0XHpJU33vs20/5o1XHmt75b6laCw
it9lNAKSwmo5iK96dIMl8GFRcpasfyGeihr2LeZRGrQgoPRS7H7Pp067xsIooNUn
GFa6Qsh+qry0OYgnbpFU4CXCPvwzW4z+WXJeQDIrNqEpnJq9evygC/SzsSJXspm9
h92j7S7QcM4NYb1OKAudZH3Ut9vlF6qHDYI/Y594UvPs0YHyxYvKuh7Q9dk27XNj
KPIWs6Z5ZkiuP0JZJoDMICP56AD1myaxcpXilYoCu0EB5qo5OAXlNxL6bAtt6IWt
FnIM0WXPCPoSEw/9PMJMpiGbp/5hqYiqmQELwHS74evaRcWzHuv6hOHNY7yDCY3C
N1zqP0UcxV3vMR9wKBTjbg3Nw8jGPrvf8jkdMWRAKLIo/ok72zuAQQzu4tdIB8ed
2+T3/66Z4JPXXHsLtFPJ6jOohtHf/7dhptPstugSMEWeXcA1mfwDAxH06IWyTFTa
HhYf6bEdiQ1cOfZnuLxMPSYy96N/lVTgDl3AUYdpUvkXUZS4ZcMvDMzamiYBC2Ka
NFgnUi70LKX6H/dZq6cLw5xBKuaueWQA0Ylqvrcu4i3hc+NdFWY1S2X4nl8NRr9N
1GBbufH/cyTXfloJ7h1gfsG+zTjynk/PI1YRCTWU03CHwml7fNkrCzw+FC0X7j0J
T9LX+P37X5bST6KNdIrpTGqFs4/uH6xogxFT/y9x4pOfcstUBnIedPRXtKj1YCIx
ccrSA6fQzBX/h7wFuQ27oJTp7jqnybZTyYi42vz5oxTQ7mW5s8AZPQhz8ba9dFvY
IcaJb/yKf2HCO9QJmkDJE4rPLXzXzGruoIyp0MqUDVenwhvzrzcH+UKjSMRNaDGu
BHGE2v6K/C8cr6+L1n9gvuZf852KkJfZfREFbJWRybB7F6yxdu5yelvTR8mNJlNr
LzWLMPBiYt2LRq607nZmcwpvbs/n8xBQwG+jslrQxwDOL8df2k3dfWawTFEJyLuC
QnlyTQL7QLJzxtjGGOh4LQ4kAxqiK8b/F4hWB4sTdp+bPgM1w7UUqjkcvpgrjrSH
k9XdLsrgE/tTBljqHgBIYvpRSrHwBDBGN2e/JV8M0sGzxsfJWpIflzIpHbEEGY6j
rjRX6UmiDiu6VnfHTNol2p/x05GSdBDWgckkw6lIJ46vo6ZV8cMwuM2KK1sUu2Ox
mGEo7Xun8KC8THNttMAPpOrifH7o0+/Ebak/G1uxtg/uwiXTZ2ozE+cFwmtq2b07
uzaOfxUu+Du4MVmANB4XPlsvtoEnClfDj6ZYG0h1WlXOsT+eo5+7wKAoSYWl+NiJ
ug6Bup/IoTilXat7pR+gqg9uu//Cwij6s6wu5oPA2goZEhvn+f45UWHYZtdqgrfM
C8NsGK3Aixvb1FtsqtYQE3MpD1CUGFhcZMwmz2hx3pfrACNtuXx7dExUoszFCfJN
Adko4BLdaugPaPcBp5MBH1devNJj1h9lfJlQQcpX7nKzcA5B+VSEileab76cCZAu
IMjpE0WvzeUW7FWRHVi1rApz1Vkvd33tXJ0J8Ev6TzMtGGSiEWUlKq9VXZqRYWLG
0Q+IJmEs2v8tdzKYc694IDPjzZqkaKf3DsIyPAjW28C4bJq1p79wdi49QjTZKew3
/1q2woG1db+ugw3mRXiVSZ8f4cLHkStGizMgcVhAAEudpaqunXQCyaKvRCyRc0ch
YgLcZas7tkNDY9YTRQTFG4sTxVjwQdDIT1MjhUqVDRnhQtG4DRJVQ37JcEV1W1iN
AgPgUgCs/DNkD550xP7/tQR9OcVGUNJziAPDMd8zae8wod1Yjqw8Ig1mOslrfcxb
/o5S8tp1i2wucBjka3ZhwcoWEGxktbTz/q7da9qtNFHbscC1wqm24LqVX9+yhRzr
IJX8SPAJt7QUi6+HgdicXFqvZE785WKX5dNcY8IkUFfcDvUrLsP31xI+xD1R8Rv1
o5WVWJ+holvrptSTx+F61EKgYYJVmOpEp7j/Fwz+t1VAtfTFy8acU4rIom1gU2uI
CpK1Gkrg28DY0o8OA6IIBLkC5wAqdzcI9oYSr7jVpDkuEFRDt0f0ejxTpiPZcfpp
kbjPvKvkiqR2t9I6uAJ8y5QtsLPcIuMQsOXd1SYh4t7YuMkYbHD+TaXPHoiO29Fk
y+rUi7DKLkOfFbVY3ZhFPNlGoZ9x+ttHB/Kj45teuk8WapPk77zXgySgoqVwzeAl
OyXOeGLhjxEFkHr4W7QQJQpE0ezK4OAFKClisvHvqPVfS9cmuOfOqjpJ0QOZ9S+m
A83EiIiTvUIn5//AxkZgj4rq/emEGHbdScqLQiKxM9u/AQXQBus+mDkmYP3xjxkL
yFM6gtIUrz0FnPwFGO0epFVBSGCWb6o3UzK1+O+sskp7ZQ/gezzKkh0DFqv5Jcht
UhTTYR2Du4ND3d76YKBGH6gUuQ2blzMGdT6E3Py6VPSZKfFdRCyR7GeBffCnWo59
8UM9yhKeP1KD++RMCOngnYcvdhoq8vLL0STP7McitfcFuPd3qKmBoT1AH8wtZo1x
yeTyV24WZaQBIi0HKtFARSoclM/XBCxFLMY85Q03SwW3oJHD5uEjRiW4O8d+kMo6
FRP1I3Rku37lrxlXjy97d6Vyc0CeQxLbk26Xk0J119phU+ci67X+fXUOa/Blgy6s
izR8kRrkJKkh9YXM/N2tCBgd6wZEu/xfK5Iq1TiDoovFTnMzB2xhRj5dfX21tfXo
zdFahwuaRuVX79gLMb4EJktvFa4IRX5iu/tM+3YSYSbbGPXmKj6aEg9D9hn8AvTl
W5c1f+XSCtlDnylUN63dYJ5IT7zsb3S4DCOfXOBOrGblV5Ipy/xWvguXQ42Kbdu1
Q4nXtACL+7kvKeCTWaA7M8HR3eDzSCoI/HdLraWJOP1jCEpHtBqGKUxwl0u7AeVx
B+FMLPN7K+9SOmqRnbL0qRfZBA0F1J6t24xgxNK2F5CWdxt2hYR0omMRUACoj0KY
HMLeiNdsAgfRadfxh7AOy9BECBX5/PN60XLj8AOdCXBoGNMku2EEABiTo6OKX1+s
SQNBTofvr8qW0mgNkBZ5DSGqHXco13KO8PMwkkoMGf/Sj9LlOBIDVDhMPItKlREZ
CsirPb0jWWolb5XkuWZGNyEmjkU1LdpkCuFmJwBfbI3aPROUMLeDLYindvtJBO4J
0B2waBP0QfwUAkQ7B8419LcO+eYUs/Y4fMxpKBJkvgR27gsW6gYnxyDNnVA2UVjp
QZlmfdDbYboILJgJLSxtCQ6R1GUaqBdtQmysC8DFUGLKBZNsA+AAVaYca/sJXwL5
kVFdIAN/gJlE7WjCIz1QWYK5mAFJtvN2VZHXYKQbV7QdRAqjePqKOI2PrLdJ9it2
TUlWXRbD7jsUPYq0l0p6/OPAs2PN7GKhh+6h++0r43x4B0xbbLCN1u6+8tvtKq33
XdI2+YahOduFw6jWUDCaJwKnJpt7mS7VUoCrhXhqZUkdZfSEouzjUZU5BUv0oL3d
E9BuMyt+vF4/rxQI7Yl+LZ9vFE9HNoMQE84Sn/SVbVoucEXv6ykpCm+v9Zr6U6ib
uYsKAJeq4rkkK9Pv9+74r7cr9o6hDthUWfq4m23fRYGV9IcXnQ30qX/I7cQIOEvj
qy2GZCjf+mxxqAdFZiGPgDsJMac1ePfGSjeiagjs580ZOrizrHy9dKSbXIR1nMfH
0LxIbEB6fybW0JFPusgACli7xdI8QE6kta3m8dHILgWrBAGR/mGXlEYCL9Bd662n
zniZn0v8ZYIC4nH++ZWl12AyMhxrThBJJw5RKMmZsTbWaT/ttjaxCO69qKvYptla
iGzMUuUdrizoUdxF6FpDLpPqUsNUcxUHair5o7c2/2eN30d/kLY5KxXijlKQRjhT
+MuI/vycwhosaAngtCL4e1SLFaVPqjzqDeSXk65BLqB2itgGapq8tpHyUpUSvUZh
TYkwuhsqKgStpdjgkdWLVRzHEFp4EzFPpjtYtMWkwYeDmc0QY/GMIAa1MBgyceoR
c6DFa+Blz+rXOZfBE8qCnnkcZwaPNA8peCwL8vyO/tLTLHguYJb7O8QDbFwmMxMI
W7tXA18emDCJ/aPEv/NVS4+YXtOC0mWATxOnHYBUZ/1sjlpRRZvEh8Hjpi/GMJQ1
Wno4Nq6J0yOaE2jV+GmxgSOvEGUn7u9GpQVHtBwrbY56WzYdRDMa4VR5CwZ96l+l
erDWI4gnDjwo9yQvXgV7QtvDbV7p3m9Bvv5YbcunWdDk/2N2ySH+J1pQgHC8DePg
nLGYbX3/SpzF+QaBNwljHjsm+JQfAI/TzGEzT5NRqkLMuwzoenJiLb/6BER0wCxk
Y32PPH/rqm4+q/VuzIsvOvA4Of6pHyxbYF2Nj2Jr3rUWyY17XGSp4mjRaL0qZA3M
nd58hEJaTb7BcBfezT4dfoy+1hy6LArKYlkTnoBZlKOX3EyKYhw2UnNWeB1m/E4l
Q0A67vj/4Ej0i3ebjivIT8UcI+CKcLHbWLSoFzYYJaq5Xy58hVYo/wMbgJLxq5Yx
kZSK9N67U3DwdGpA6bNFKWPoPatvgEcTBQndIBsDBTHvKXnZJmMH4QvEnelr4YR1
ELZdA9Wrjp96HW5lXiitgcbP97u4jRhc5QaSO3PzYzkbtYkEgZOhYp5U+e0J/ig7
IA66zhwzxm4FAZucV6NVNGpXpSdJ2f0+9+78zLY4JKMuS5x2zTLf3qQCzzZmbX6/
zeAEImekSswHcakLohiU/eR2+x90UmhXDg0nW5yz+m8ux5gzuVU6UylAqZZwpXdc
OYjCnGXg6T8KLXvT11zzQiS4jXM+XL93cf7A2tvk1zWEWIidGWJarqFf4FE326N2
P9J6YbGbPPU8fplILkhlYYKkl1Z5wssnZEtwBBVgD+EPAcN7777ciBkwegk0OHxb
WQI/xB86BVVsGZqinOESFd6t12zCtGW2pFSTRirWSJYhTJlHzBPB5ePf8L4V/x+l
LWgV8SZ3sW6Kj1UYyrVJ/grDJwsqse9kot93hUTdK/np9t91iJqZSxtHmPdNB657
IJhR7WFeOF0eNnQiBc/SzFs9g8Dc6mii8wJCUKkFhWMFMJ5u2rV5OAjpbl0slD/0
z2B+cidyJAXLePPmmFKhMaIkaaYyYqTLwFhI6VIY4o909k5z9ncR0eRteP3cSUJU
an1fFPv6fBQv72Zs2Ugar+1dDeTKfDyEi4n7G3sctnGx26doSK9A9Fc1XtCqy6lD
ZcmQRGPZPqDpx13apvPjAxCqOwOIMwg+roGAD4e5YgPCD+YgD5mvLwEgBbl7ol/X
dUM2wYQ7A7iOy+Y8RUBf5YEnPFTWDfYAaR7tavfN3Tb+DX9vbcXyus30s8YxWLOP
7fFIWvuCfSPE3ICpeFZ0qcomZKl0Ikedn6DKDLrmnGPDGYOC1kC8BD7ifcyCGCxw
64hOE93k02WPQtF78kMbqPlaXXogtypAKdlJzxvl2hxmIbHComO+qr4ntR0ip/xi
ys7Qi2/hbBNz19Mpal1M+FP5IKlRD9rxNuy4gUZgS5FvHlOV6gM6WY50rCR4AcDY
on2lkkD9LHqnH7GoU0fBNY7GExt2iL5n+0k4eUcSPahrZcvq1xKj5KhYrw6PP0Hl
/95tabMjpgVCVhKncRb535PQ6ZW5L9PWpDQl2Lm1HwSvvV+fGTQF4zmwd1z/WZZ+
9MO4NeI81tVnQBPzCYKWeR94CqQnr6s5350MIFggYIsGgpq0TlxwMxhgI4ZIQ+kv
0hJ7CFyeNIJI7c8syW9vunPo6YSZQH5geXzpCoffhaH2OOL9GgoUHW1rrvhBERcE
GDRlpu16NhMROgY0EDUOkhuo2LpLSRjT5eoMuQOlaHpW8uiKhoijGk+doebebyBC
YNGNe+umNVJYTYw3hevGxQAAOeu9+0x+U8rX54jfeeihplKUNjQFVl/3rmXtwuQu
hGMc+d0FdMKahRDZd8JvV+XZ1Pka9U44HJpKHHQdsAK2TPz7qqSCc/SMOu545FES
Hv5n+sL2Q0ubqZcLauf//atKEJTpDl6LZ3fIos7I/GlgIcsOj/XRodqgH3PmvOqM
KJq90s1Oihwd1M/6pk/mDpupANrhP7LQKyT1ggaiXrW2jnWxWmB60xvFYJ5iB/2W
wnI8OgLqULMNybOrT0NfRsY1YwJlWK6BtbF9YjuL4o2Zndphpf30Zfge8/ZsCIs6
iUMwTPhJ5U1HSM8kmzJBYBp84V1uoDDhfTHOuSdWDvxk1SqJG1AvlhhnHGx6vCDg
sF6eNPPcSDmE6gWBU03oiMWpHHFFWCW7iP0tTQAFKYRLrT3gMLeObLxoPoyeR/Zg
RRmTMofXcrbaaOaTkJMa/G0NAvdUxvW3SQ/55Ys5BXxf9Jm/I9h3a0j5+6iCSJ60
z/9ZGHn6kSPHstgk0Q8Td7RQiSaR4JHvFAwZR3dfFkx76S1LZNONuT9sU1PRw92A
sI2xxdSHNm6HcT62o5zk9iRmSMCsR9Qyz4vk4lhU1kVIoAhUvQK2nlbaibAWYblY
BlyWEsuzwquq1KYTh3dsbevvObJFTcZggmcFdT0yhsV5P45vg03R5aWVkWIokkpP
/A1w+XarxVE2qEPBliilHFAXFTktecrYVxWOStcxabLzr2WgbvL7woKDqCBsOYgG
96gXGap6F4ecHHS5+C1uL6YzNJH0K0Op+uCiEwlxbnM7Wk0O7l/BM5t6E9t+5ktV
XRhkrBnsKaKg2olegYMH3SfPOYxB9fd8d8htiGdwfjvb5AfXSXqGjxdhh8XiQNtq
DkuKmuGfEV8u7yD/yXhmohIPjLeT0BSa8l8fkfh6xmg5REIlobmaS+OkkCiRwe1w
eJIIfzC6A2foa5/d2BDxc9rIIAfjOpY9M60UMWF/Oi00CvuC8GtnuE4lTQ2R5++B
1UlhmLjW7hhsQ6rPU1jZ6YuwobU0YaZuDP8jDoHmwnEj0JpxDVe+5DulyGKim1Fa
/bsblx/Vzog4ZQsdwOQQLfYeF20UjuxacXf7R8cqg6P16cs3eK4kb7xhph1Zi1yr
V9U0KLePe0vuTlVd0UV9C9ghm7LiKENtGgAdj/gyZaV7gOLrtUI5vn3LX8mU5Z06
NR+PxZ+NhmochUYy50i8rhN/uVwstAGljhJJMY5qgJiK7bpXqEGrHHXFs0/T7tFt
dLvWV664KRU1D40XwCsMLt/Uwk47QVmRI7tD6qPJMFmEQxQuY4GKQGFWI/qvYKYR
EAci0DNy/v3dvv8gTPwhxUhdvu5jrUQHJrDhwZzaQxI+w8NMdPfnw3lqA0riyjNS
qGBYK+i1s6MIu7uZekWRpHQ95xfys0zDYaJYkMe8DeDzEa2zpnJPPnLmzHArGpNt
3B2KP+6Necop/bzcVc3hE7XJT++YIL7Bkou6E2W+3LfzDsw0IiXjg+jy+oa6fpDJ
IhDFrSVSwTmYgoqy0egQOC4AlePUwpVZomlDqWMerXRrZi5DcLNJ1mDht+5AJOj1
RSxEo8OW0FIPuIU0zrc99uWxFFbpqwDIssXNWLvA1NOuDSnw6BWKI50Ht/ltzTtd
nEo3mCH1Vgec50jqHX+wHxsvXUXkOYXAsfT4jECnUeadcGv8fuAWjqwZzvT6xGzu
fuOcbNAaL6hZykm+NEXTAFrYczGcKPhZLMvrkx8TVl2F53ieye3FuPcNBv4DNnNL
x8Mjieva4B+d/uTaHiQmhO7wVNf1X05Evqk7SCKr1ojJNY3gPQKoEnh4AHxHT1dv
ukAy9fDGoXKAgxlJ+/LCXXCvPy3YIjtJL8VSPCvPca03mS8t5z0AAfNrxB0wCzoC
L+C680QJRKBqXfPcJPANjMmowIqUmDyUFqjSCRF1lIA=
`protect end_protected
