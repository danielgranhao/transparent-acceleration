-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
R+WLuu4DA/P+PvvqlkJpKwUsJ0q5deedD2yufpBgJvaDNJztf784On36k+dciaJI
DF7plEu0QMAzmesay2MPzI1PDZcOyRsyNANxPn0H7uHSiU0Ex5Bo4kR7qxLHpaCL
A11NAJphuOiithhgPd20iH5PCOF0kyIsRifhB1eC9OK/mexkF7vDFQ==
--pragma protect end_key_block
--pragma protect digest_block
h/6A9HCJ9gEk3zj8zh1AIQUXsnE=
--pragma protect end_digest_block
--pragma protect data_block
2BTcsSqkI2V6CHy8ZzXCZnJ+X6z2nXPNuMSj3dv/fFutdC40qv/+Ami0JWtWeCBX
wFmUbdVoLxxgGdOLImltzQTZff17gLovv+afdMAjvb7XdPj/AE4f2vadGwm5+06V
3BVeRqgEpv/12W3LbUGPeBNlZVpUBz2bn/xR4By6nF4AtbzLPIRfFSOn5xVnzQ/n
eWsMi/OyXc7L8SNYtaHfaBRXv4I0wM6khkCxQveggbvyDFh7NCFrmmxZIXaguCrb
kw8Us9ho2dpNGXvqeFKU6LMdnMCZIzxo/CM7xx9uByhrahZrlYNa/aRaklAFl2C0
p0CAJ9sg2F/2bSB1dCcqz1ggcbZ+FOe+x0qfidzrnaWKMitpovAVe+b1pE6lxJp+
ZTLShdIBaPLF6ZAPmlB0Q/y0+mw0CjQrvb0F7Qu2OTpRWmHH0KxguMk7sWGwhboa
FBgpxwTK5PXHcm8MBVpcrf7YnciGru9T2l71i0EjLTBy30PWPDqi/yowSBZK4S6J
6bGAhwtLQrUDhexoAkLfxNbuFJoihO05thNyfzIyHJ+wySNTvbvAH75jVDpXn7lM
ewKDaghPO2gBVQb/ogICURTf7vVz1EQWHPH1Y6bbhNy12nGYIhzTHlESHeZq0kN9
HlaQ3JryHTieH+nviBdQJvhWBGSFUEi8lxDpqjvQKMOVdU3cc2Lq71SAsqw2M9/g
2vnuAuVddGQnqOcbqKwVBoIs9GYpxerKliSQ/YRxxdCyLftQHAc81Bw7oRrG7FA1
CZYeiddfYQCh0eX6PawnIiYO7z6ejIMyAU2VjIA6p71Lr9bGMD+oqq9ftEE25peh
9Ab+/pANrtck+zyC6a4ZfqGF2QB/uhT+2mK70B/7c0SaRXrXCqL97Q23WuV244Wx
tcmckJqpMP/UXO3yPu4SIfjfrpf48GFxsr+0K3cX7X3TtvxqFRbpJ1CNZy1yFxXV
+qrv0x4LvUcIzv5Ba58gmq6P6yAhEk54G8d2irkx4xPoLULG8YpC1LCz8DY4hbEk
DQaGLARa8SuE+PRxWxf78M7Fjkagn+d4xmf9UfqPAr19HuaIpb2OXumlomwYkcn1
kHKEjgu99oZisep0af0PcZNOE01zj11L6s0bkJXgV9lWad2R/X2h+wzOEhq/+P27
uG9Yx+F3FHw8aK+Rwr7AhuMnIzUi69AXrieYq1GH76nYh8n9dxSjbOI/19KuaY2F
H6q+KGBTU2YzO/MQqvtZM+i50rj/m0waozsytpVgK7/8ffveUwzMbS0+d0DNotp9
NZhhAZ+smDkZgxhQB0VoppbX96eUSE8P9PUOYZtsaN40CiQgksWVWhixwKgB6E2g
ADUROLYTvanKI4PwPa9FHS1FbnI/9ad6f9NjjsCzZnv4tpyYU0XprZR/Vd6J5DpY
RnhoYL1300NQ6FbqStIFAugTWy7s0ahOfJCpcL7ina78GyumQ3oHEXDCFUE2HSvT
UdBtKVv3YZIQ4W9mX44ZKsscoOqyeGGtkz3Jux4JZeksnVFmeTzvJHNiaJetAzCv
xaq6jjHO3eGkCU78T+S/75VfosChWlwDdVILevmksZ5TC7TxE+7tFeBiDNz/M5bR
5ZP9M1fqoOz4Ev0O7hmS0bTxrPTiV+uo39krCmp3YTlRNO0Z1182OgYPhv5IdwEV
3P5lgX/SPP/DxjgVQ4r61e9I/ABU4mNcuqrIHVrNSoedoTih7ALrv1WwdYwMIDRW
a3/DpY/ID1a2bJ57SUf1eqXBf54xeDimA8BbuuesCgldEmOalWceCU5X4L016Msc
oZWYAs7nAAwmCgwh2fiwJ0LFXLuBIv/lPvV1+WenbnnnDnt6txVWhEM7Fu8vLuNy
4aQLCg3gtASeIk9B1e6kuZIdA0tNePfaUP+jBWIZdSfXZT3DOMhs0fLboJJURSup
ZDC/B5e/45mcZvdc6L7DGCXXQiIJbSjdyRs6v7853U1keCpjk/th+DfUgllJTOEA
IeLQ3iJea6G6YjcLTB4iuqhHVhPkC9qjFFYYdw986dcxQ/b6Kn9LnSu1dAkNukEx
GuPC7vDIjjdFkjyfcxkPtNDVAtuq3iVvVrE03dFNFfGqf1sWVFKdQxV80kGlgPuQ
CroKH3fRy144w5Ryw7gznZSZ/nFItIiR5zfi+RgGJm0etUGc2VY9opZ7OG9EKLYC
PjJpGOXPy3hov2qB9Xm414Vz0UcKMrBHryDV0FHoYN64lXfCwWRKFtqeMh/UmW0i
3EDMswXQjC8maGla1i0HRDYqk4rJNmJ55zsqyvhNw7LwxlVK++DC3417y3sVfsj5
ssqkLzxdhjC1ObZRYm2g8MEQ8QFg300Q6fRnVzdU+fDgb2V/F6RW3hUb9+VBV3L8
bAd3GcJBWTwGm7FSQjkNGfKXUkrbNZFvsTYd7Qa/cXW02WxGjl6YDmGIcnhR22pH
gMwx8CQ5OXP6z+gH1tAI9jhkgzWQxnHQ1NL0rMvyom1dAPKzW8v4V1bWIdqzdCKA
78IeMWHWpyLNlkUwsILjsudahnycw5l7S59NquUt3+Xy59bDEWAG7Z1Iech93Oo0
mj5v4TE/x2l5Ur2mDzSiN/SzgZcIA2qLqqEOL7gq5Px7LECQNqZX9KYCwAkA+zyA
iZmpSE0iHfygW42T2gTBFjq53NeOHkfroFKKH7SHAjysLlCbwXT0u107fim9fWve
ANb/vTqxJr1pYD+kyEfs+5AOji0DsKwGnu7+ioAxCEfPwnRLlh8MyRPJPHlP3OGL
6yJECnIN0f9s4/r7fmIFQO9UZa4NWwo6NJYk2PUgRGEq8gCJSBN4WflBwOHa9UQ9
GH2Q5TZ71TVCZpKzheAzJ2k/FqyBuOMJh98OOKgTnllnrQPJm3pGlUuIGMrg8xBJ
Us9pvT448wOWeFYbefQP5ct/2R2sZdZmzliMvdevCHmZxZWnbP3lxS8yWxe/NbmI
sHqJqKLpPUNYpjZXAJ7kVc2kRwYOC7Mv8fDlXLShbt8XENNI2iY1eL+W6H4MBsns
AhBoiYHj6HrF14Y0iZidXZFZnSAztxnSK/QuODwFKPvxj9Bqws0j9SK5gmn9gxqb
8bIckJUH76ZYy71ieb4tWatFBCq5dToAhinZZERCB3VjhYYY8SnTPaLQejIp4+CD
a3O+qahqSXoMgBHlqjvHf6nQtrEB770eX+3jKD9fJYb2YJ0igu3e/UkxaVAin+/z
OftnF9RdfKzWD39is/2CWBtrkzy89dLMcKKCNfZs/N1u1KDOuQglqZGNcQ/mRjSO
5/uVGvP/zEJvOaBUJPDxVkucID85urV9lgcIwoL4G4sAICp9y2dAOO4qOem4b/jd
YurLZWuAfITa8Wnkp5chrCaJZsA2U3O4ynFBcEMMfbcL2N3iNiDQ26IzldAXVyeT
qVFrnoOsoxHIVLyawQRaMeNXKDYdiPeXqz79ufWxiRoDu8p+1nfsXAvv57feoTEI
9BA0bI4SRtczA2pp8VlUi/+zRQlUG07cDza7b4q40/RlVyYKogr5Yw2XzFmks+YI
pgbtaX7Zgi6civkn7DOpTH1Vkl7/7jzOwCE6WioblfzesvwZvGunmJHSe/bXeH7j
4RrMJOvS7b5Y1WTAkYB4j2ZeYlx/+WS1OMLmUe1FM+I2sDpDTXO8GKdbD4EXS/JY
Lcjh7HV6+iHwBBNHd2Zun0mcug/XrbFGfTn8tBIV9Tl00WYbhM550xlm30vMwB5a
4D7dJ8/uaguGPeUslVAwHtNdtBWEC2ZegE8i/27P0xGxXdsRAISsGeUktKnfnU0g
xLonhjyEhi5B/jOzDulOdZSOkEX7WjObt0eEZyKtzvqJLEk/uN/xyl1lHFdFlv5V
PMscd+/clbMrNSMuQE0vItTPd7H/2Jds1g9IPy3T5Q4qN8YkpdmFNwn+wDnIregW
C8IiirnoKFEV3akJmYWCisDBNYI4eio2+FPtjUn9IiqfUHwz+U6X8nrSv89+5l5U
vZEaF0B4NN7aXYXzSpNX4MT8EuE/8hpWEug7elxP/ZSq1WSF2oUGW/27OW2PaX4d
uZD92C1YPQ1K6cpRxhnsL9i+DLrgdguFpBblVB9J38vlj086+Iz/7ODTNRIIBLKr
ju9ZdxDLr7N9mQlMRPODZPydZ2K06jzlsDPWI6KqqJl6yxoTLFv24Db31YilAXrE
CcGHnKZC2iHnBcRnWYrnbB0t9LFi8Ofg4bSQ/3wCkmbxXhRhyIbXCkUmKPsvsAvy
ia590u/WtZ4WTCekT9GXR7XIZ3hfsGvPKmDUgvGw6AIXcDvtWmwx9tEG3xMmI8q/
t0r4+f4ge2/1Q8Mpua09yXbP9Dvg9XTKB0ySEnd5xXRDkOVcpFxRhk4y3gK1Agzc
qivDx7A/IVkQrOhn3nf66SLkC6J0CFoHKzW+wpzTH0vVe7S3zUnxL5GVPDLOd3DJ
BkYS+BZVIewjHp+0NhoDftNEvoiMhryxQliwAgC/pTVT3ZAiqUPhQTN2Zq4QNSds
5vIlAxTj0d8SolItSsU7xqZxUgkg07/itEBKLEEfsdwOWvNh59gsW+IYVusUvGJ7
UuOXRsYC8QeY1nAHq1AqLdpj1T/SR+duqKhAucuLXRMM24zH/8yf52Pquheej7ic
sdLvZ86P4wtJO+NA2qHYih7CxIDA3EqDv+gu99qDdUPbtYHAKM3ymRVXRQYY/RKj
qeeMudjNvMCa9sSBLaeAgwKRIfwH6zkcYKmsuzedilMuDJ+MDR/+vfHWISv2wYZs
W8INoWTjSXGqij6gFGe6zTtzL4O+Wgf06IRLuRp6D/yF7Hq8Fx9st31Y7/XyUFWi
ny/lNTk1J+0yLlyb7FbwLOuEgKqibJQnWYq0Q6crCZrisuU7Ab1ZG3atTYgXa0l+
m15kPQznujSU4U39LF6ijxhyG9/RpmhmBIhKy0/21brxrw7ToflEq/a0bd8P5BKi
ayj61LLNm8NlFaDqBzoB6n2/P5+mDZd/t0ntCc1STf3MjNe8SFmIG6WiEzNV5+/i
tYH3OGBZ67bqqaJrHUUE2uakuHByK+SrtqLa9uRD487EPzZTcvqWHWSjyBRbXoQv
MCb3jWbSQucoBY4OEnT5N3/gQGVatWnyTsE/KKTT4uYBE4bJTQSdb6Uh5nLEwNLd
z2al8oMTF1h9N6dtZX8WA8tJ54aoJ/cDyOUehXYUuA76QMklcY/Q0SX9XndG/ZgH
tqmvqWI8+Z6zxSkAxGw+YjkOmVNOP8uv2jmuIZ2QLgTRAQpfkDXDfVHnrjNmsnpH
yv8mD7sg8BBPkMtrN/JZuZHHfQnReYXt93Dyp8Zh2YoxGZtfHQaumuoAaTKmFPJO
3GCY0bGGzM3+Yk7v2VYw2DClo5kI0O0RT1tMsigx5Mu4Ni8eV7iipxwd6VPmBgsm
k6oEeqXeqVNNlwCoXXOcTQeTzXtinnUxp/cEOswlYqBOCxT1YjFPU5JNfHtjWYji
E78u3OJQH4SbNBH9AYa2uC8TgjPO/oByy5kIqCG3W394Ukuv7ziUK++74vTKjzY7
5HthSN01Mwvw8xZef/mqCksJmjrGXyDUNFQpUeZ6JfEJVCj9911xwqPgLcAnODJO
A7ASzVheoetEA+JrMYbeK2ih3IIniEa1/9n4xxAkvsRvpzLxLvgSpvaA7yQEeRTj
b7VNsiGhIZmOZPaCyFvV+V+s8HHOajoDq/eVbG+1f14df7IbgPLQmaYVoz8cYKbn
7HuLR7ycVUun0WsA6dOMaP6tg1uqWYyo7TkINAEUzs2Ilcj7+iV0PNWmA8lYi3hr
tjP16ZTrzzaGE6eDQDcEIbR3OW4Q+6Q0fjwnlbcHbpqNeJUztTQqVAAB0r/rpW4d
DhkRPUirG10jvv3ZT+WE1izIg96TFXpqFarWRnaCcWUeD5bohrYLW4V4JZaDzdxK
GoWV6NDZg9QEqLU+ynOuslOb8QLD1g1TpeAAOhLQ4ILd/5ODM5Cc1Yy45MVCXtBk
wfwMlvFom8qRySNVfsWeZ1E/jYtQreQJ0UFvkyayzhOOuv2IYrQOpsYkDtzzM7R7
KAN2BR0KAwCCY28eamoAcHb+X8ZQqEoqcI9vCLkvXUFh3OWjRfkAkNKY7vhygUZp
bcUGUzbELF7caeHP1TMXPBH+7fgV89TBJcubwzmtLVyfHCTwme6lSZcXTcMPvtRQ
DfkYl/4jXnzQaGl59NEWlLTnJbJxGlpa1OPD6x7fZWb6RuCrEACMq73mA28V5v+y
PbqwsMbpxGXhR5oX8ofrH+pqHRnZGDMWYflPCSI+uuE6Y1QsQRQgFEw3HWDOXMRV
/MORRqkU5T6We+wdAYoK/cHpJJaX9kTSkQj2J0mxkJxNTARt05OYtjcn0sXUZ6gP
eeluH5r4JFF1rmeONhE5YLeFQYqGO0OD2PX1V3QJHaFE7AUi7nXdQN8kh8SS0kso
4Ng8/E+KkrE+pzOoXqOrlvT53z59DqYVMwYTeOxtQZaVUXH2OqmPJmvj+hgH5dJ/
ous9DM2Zxt7PTp+ZQKxVc0fBGdjyjthmg0BYngzmRjnTO58A0ZE9COFveyJFrSE+
DvyYdbjZz3DsX+cFC3SQSP5boI9gw5vLF+OsdHnh1E6vt5+nwNMD2wqi8bkLs1nW
+5IYuvZC1ymfgCuVvCeuGfb4CL0qLhWVuNUZ1KvKz8dGrAr+OBYlI0wczDCftUmC
H+fLamXM9SCgDTjVR4QVSCp5s4mGK9QdmLF+TrrpWgmuJYO1OwpP8N9pzx9HCl0E
u8EeszJNt52WhLKDtrXL42OKd4LoYrQJySAQQqItQO1Htdu1NJbo5598sfmJLQ1n
feTJ/AXBaG0+2tkrTl7LsmTST+LrLgai5vMOMXydn3M+Y/xnwltA7fWNdHK8bRYl
xxiNQ+pF8s1iLyLeIOp6YZzr8Qul7SeTpnF4plNDxl7SFgjOXtms2NbppOAl6KdW
2Bp+lTXynhiUWDEFLn7Xp1/vxwwXruNbAbFkGoi4y+KtEow4E+0GgMCxLJ/pxt2v
UmR/psyXfREqvpnTfwj2G5fGhzXLkbqqz0nF6+bnEz9DTFxSyWxJ4yjLEDv9MAT+
mYO4xWXZLX0UnX35NzHHRKErQ8qU+Y6wjEruSoMcgiqMjV2FHdLYMfyoNYH7JVAt
t8Vj9lcnV1A8CW/zvWg+R7GqVWL1ZH8zWnNxWrJcejOyNzyd3oUcPO1GBsP4hyMM
H1y9Ly38Vnw5AFIrj/Cxbj5eYGEb+wE8jtMAWjrWhg2YaTBmOEMm/nYevRjioJ8L
sDRUfiiV2tflANA6lTA3B1TGtnqisRjlgpXaoi1pEecymCoPuTOfqldy6eFAlj55
nscs3uOXFArTIyIAy9XIJpeDveBh/a5M2ZDlFF/6zZhYce0TiYnzz4NjafaTMget
Y6+V1SyV3C+VBG8boca+WFOOqzv4d6L/8TOmRyCNN7NZRZFPrHHIh8LrU0eZ2DFg
328zq3pHRVOW1Bdd42kqb1ylSNMP5D1SbhgWJhb4w2cMIANHFcz0GzeiZNS7LZkb
38eYAfqYrEVlKEdGVSQB00TU91c6mIXDnBZUsZezS6QEQ9ulRG42g0wb3XLKhrAu
k5LBucGsdsyBeSv6qOubrNbDz5/q3QG+NNvT5EUR79TAevi+9qK3IzGuRwDQlX+D
+mQRsLdabEKzcd0cQe0u2WNL/bL5nS15VQXgghdhlb2dXRSSGnAvPJ0FWXeStcP5
pgEMOkrgdSUJAGXx01vMbs1eNN76s4IRg58PAs2UORFWG0eecYVjV2moHPasnoPq
GW/MkupqNkXy/Br0EhehxLVKJpZ89vE/MJ01P3Qe7oNp2jLv7c5tuSl4/3NFFmAR
Y4REcQGkIov8ccWlTslh7Yx6VYZELtwhFi9+2Nhmzipg/O4bnWMCC7ym6uDsaeEH
eNI6OYQvjp96/L2S3J8MOcqBqkfYAvaeJrc+9UShYqSbEP0/4BBAJaIUAfzBWJiu
H1YVLE6wg2ADQcGK34VsSaTZnU9/y9ZFHRYl5sWmfbBFPg9h1zPrDTczSprHTUBU
x73glCSHrGQmb80jRLBN3ACLW+JytgACAtFOWFQynnd2r3IGyqfzsIf6DEmT8uBx
Y4ztOkGowkunG2BIRVX4BjaQ2+ewP9qO3KPpyR/zWfT6wo4orVeuFOLFCTtFZDts
wTrwWytp/P68qSAEp4ziccR4djFLMsLAUJ/RUq7xwnZf7zSiEHRJf0JqncGVxmdt
FoLUJGo1peXXLQaNVYubUHduzL0tQHsv2JiVzHxiQs7fEiG/yP4RGSLDgvDyVk8M
uRU+91WiyoqoGCdned2MknG83yc8sz4pKsXWxZQUYrk=
--pragma protect end_data_block
--pragma protect digest_block
JjjFN43as2EAwwLrp5Nsxp/awFQ=
--pragma protect end_digest_block
--pragma protect end_protected
