-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
V39UdIdXhoc2hFoi7SAyrB7Lhbvx9cTGZfdO/b/8jKJ/eqj4q92gzElVvdMOJa17
8gARf82Col611qN0HNCLxiSqA7MT9R/8LPfyuwEFaTzYi5iYmb4oLFAhj7B7MbDL
cuSjqtVe5BUbaSyklaIxOqgnVyWIZP86qXCkJSwRTpJApA24L205OQ==
--pragma protect end_key_block
--pragma protect digest_block
zP27JQiCXYFyfpcpRYsajCqGUPQ=
--pragma protect end_digest_block
--pragma protect data_block
K8I0hVOFMsZ32Z4njSt4AaKrYmh8UdpyBh28/wQV1j7qRHKsScC7RILxQ6tsFGFv
lF5nM3PhYPYo1AhTS5Ab5I23Xrpdt7w6fP/YW61MoJfihqnPbTlkTkzEYv+amim+
1eZOHwYDI4cEyBAaoh0vjp6QUznjkxt+ygfMCDDR167o1an8cO90AnqItxKdpeh+
ZcJR2sg0lqpSu383GKP2R4ZxiMhLvDA0vPaf1EohAxe2uKPYonSLvcyOtE63cZNE
1p+hwKVuvY2JWN14Hn4eUZLARhcrVhzcWE7FF0t/aTAKmeeM0Z1qUCCPmGwpxus/
I7ix66xFZdL5nlCAkiBN30RZ3MwyXNwhS8wNBV7pA0L3cuA88xxDh1Zth3XFQBA8
KFtBkq9bP/wYntVKoOsLtI2Q6Nn2SnaEVxKNBPE5UPZ5xeaY1yCxVGW+N8eUBwkF
uZ31fVtRjHM4T4DB//klqtFvzfJ7WY+YV+iYIaOK+nn6IKKsgLrK0HRG+AakGiF4
WN6w6wWIPIqN0nK+dKfyaxxI57pyEJnWrckEA5pxfb1WB+ckddrG0ejNAf615HB2
uyt51b3cyobccMl1FRZbEcb9LItvquBtPPHNaWSDvFkpYyR/5qQuwiNN9mYFt0It
qQ3wVxZVB+uA9c7Dw3RF9DUq0P/w/f6TcsbIQswEZwEysb99k8gqgKvcVCLwiufI
iFSTCVI5o9NeANDU9VWPm8Q6PDEBJEHTuLWJJZtbx/buItPM7g6s0DuguGbughFN
nrQJ8sthSn3X8God8ryzVHpWoxiA78+/spfNjy3Udltio5NsJ+094ZuF0/fs5mBP
uqF+qeL64oEW95qoUgtQVag7aEG2cVD+o3XjRKdLqfrnfzWtG5LjthVcQoa4lT5Y
ZaYqpMojBtX8ECGcU4Wyga+p+tqCduLamdkj3ehDdnGQKvowNpQH+KfvylaDj4J5
vfw09FAUMT+IIebIA8KR9JBuFIhhIEDtuocllLZbXkLfBBEoHSeKvJIcWZZ4BFBH
klgjdEZnEPT4GfnjpCJHehYNkp2U+W1QrKLjY50W/dqnmTormLBYgaFj6a4v+foF
YSFiYUXplwh3woWTl41TQJLETY9D7pH34oVQ2CShQ+LI69SPI8YT1PHaBwcBQeKd
l8Os2GoJfeq554FrftH4RdrSBYjgFHfWi3c/k9uzFiwsM4ztKKXbjGwgIer471EP
mu1YrStGGw7hFuw2/8F7wHVTgh1RkYZd09GgFMAtjpB/w66EUUhtJ+zzDXd48YXb
AfLA2se/VtJTJJbUJe4Ccxzc6iRqe8n952w4BgJuuK3olPM8Vax/2y0gETnP+shn
hbbQIv1YUyuXJmYT0GHExp+40YbZACbGJzsbha6STGuXlME6xrW3gC7dDcUNuAUT
uTM6Zvrmed73tTzqGH0HcPKRZnYWoTvV1NyqRHO5jb7Ej/LifLAXQniFLo4E7PdG
y9XJ4TqygH4K9qBeaeHkp3Z2Tb+KpNzWSxwuCJqPGqsPc4kry5ZLlxVPerIHMBUb
4LbyrIHLQ4zxZaMpOKY2A+VN39wjxcLYJJH99Ga35RMM047qvnWy34ozOzKq8ykI
Hzu0cGj0JTje5augRk5a+1L1r/p83fYnp8sxjm0ENFKVVxyRAkcr2MnvSvxjUzDs
MccusOpjB6s2zODj4VPQiIZwCveeip5x9e4IwKEBmHOXfMDdx+//6kc9ae2Y8i7Z
ThgChHFafWSwgPvvrQKxBLq8Nju2HlR51pHCcy9hV5eMZXi9fD71U/CTdkMXCrin
lav6Ud2OWiV4mQBCB4/N3+WLz6kv151g3/+C3iv6cqSDzebdETIX3GqGgwX5Bwu+
N5dswD2TPAs0GSE3S8d7V7UPWGelFlSj8GJPcFdroXYbDOGyhmoYQQ2W7BoKtjax
biekJ4egJxuZWQ5iWMGcQkM4VasIKfEfNtB1cFa5Ounx9xDCnuvraK1bcPrlJ3ik
vSwlLMnIZWky+hX84SXByLGQFo049MiObXzS9tBTywVPRvonP0QmCaubbTEGlxuY
Ds66kYSyvrm651NiUMlAbDmpxyb8j9HVU5Sp1rtiU9ZylTftuOmBT9dJBmY56sQE
fbCCT8iFmqkJnrVRoE5r1fRErL6HhxhhLdydwpGvcaBMjVETXHIVQp7GxpPWafyd
EvsXZP65l3jCyuLvdTeWi2xbVBOcTA6jjhpPPg83fK5D2/9Hm1PTw89CLSjFwDtZ
8b6zaSMnnc6ZfFJYZ6n2GXxs59LAkN+hQgGo/bqj1Y1TTme5uDDk8PkbU6uKOkUA
72NtrOM4JbZT3sNsASgGCrmp2tgaHEq+8Ho04YE2fDc6QQSDWq0UdzzZaHe1FXex
rnDvq4SoynmIygT/q5TQRqhs8+D0V1cC6Hr8rAbE4bdIvpPZongMTEjRr7IGdc0P
F67coy/A6o+8yT1qHHvxvhWNWeyDxyCToHYrYzU9cPBHuOVhTyBh7HL5TElnEUUk
KueLa7q648xZCWocof1bj+NNZb2AYiEi+La5ppI9gSOTRYhQTLZhtrzQ1JA4J49C
4zEweZfr7F//ePzW87FqIZ/lY/WC94HaILXtikOkgKt+92GRuYUnFeBsl7RL0s1+
ozYuMwdn4JbE0clCFTCdlzgrHbG1CQDuLDD94jS4fFxR3xFBDtpO3F/TqLEoVaQs
wlFNkn69SdKWEEc/mDSVuqxi92/UnXYkrPKbBwvkGRHn5bpB+ajiqOveLj7m0j8I
ilxERIAdF0a0B3njUywcRYBNxTurfyl6UYAQIUCiyWOFFGW9miSqQA5e9Tlc5PhG
DQBarrelNAQad/tpEd7vgHWnSzI+THWC7puUsJoz3AIHuxYzOUTjmn+xU3pNm1Cc
0aieYfrIrjNelPgAa0D5tBgirm/Uy9rb5/7PcpliOTmj/rbEW5oLFQ4x+Kan3mab
/J/TbBvVJmQl8SEa90mxZtngq91mdvy6WVATSu/3+Qwf/qwxGAIuV8JjMjqkyuXb
5xVUkIASTK3SN/qTzArZSk6+6v8yq1NJwG4ZQ850PTUl9/Hg4oLYRw5D5bXyqyiF
zBqxBzpXKxHm6q5dwmMsPO1/7+5eYTK489UhChvxIcTuHURMtHGm1YGDCN60CjWV
xknDJpEwTvJe5SqlREohzzSsYfgNgmHL/WfnvFbwOO9qsrWa5YPhWwYkMvuJRDg7
64Cm/kY8wqLZKg7GIE6zRptuQiiPRUjVAvxNNqZrutKzC8SROg+mWI1Ypw4RHFxo
OIAerGXM1i001DyEU+IXWGPsmDEwfMa4rJMD5pYFs0GFvNF7AwCkLnaNqK4J0Rmn
3J01DT8lUxoa8a0Y/sxSw+bT8sQQM/J1WnXLTR8qL7Hxo2ILFMLg8VthKkkOuK0F
uaptoYiqx+Px8nkpodg3sPHq3QSTmLPXj/s8aVevDJr66kftLgDLuAusd3ACavRx
9Spq67nm2VQsqjGsHFhru726MYKqoP+rhGy0PIL6YrwoSSx62unvWnkgJGWWFIz9
WTgXyC3BHCpOkj9zlCCm1QNlnBJdnaPbDZACUzVKM/ce3O+bRAnBWpihefhneV3C
eklo8C97bDmuR6eNSwPpPlBsjxuLkaMqcBdKgIf0reQO8LT53QbnFcJiHxLo+6hs
+aQFnOd+oAuxg1lw1GZJmm4S/gwvdgwNCMcM/BugRhhtPxsXtQ2SiTpYrC27QCnz
DOX9RR2JPKKZCyQZBqS8fqPVDcW5/ky2VeyqP1+3Fvn+LXQ+HAtzqHLJ8sqQ2Gsw
vyqt6Stg/zhmuSazVn7HsTLhrWWjksPvxhybLvRUVDba0s6cQgmUg4Bi4NK0+lMs
0VPDExIo8FHioNLiFL2g7BMjnpoQWNH4dpZqYPZjPGuYEOd6xB3yL+bfS8dYRidQ
pGkSY3O8x7AHOLvptO6FhossXl0gqQWkgi9OCys/iRVblGPwKQBzbugSCgSQJL0f
3Th2k0Z5jlBJcuHU7pEBRehEHH0jVi67JQBIVBjkHTc5jGZfXPW/EkidWORlKq9h
kou/zAZLzZqqA4NPfij4oA+uiMDMrM4dlYcl66l2/RpsuOhUP4UwL8sTxNZeCNvT
Pa2gC5Mbz5dfkSraa6FQpP/NbyZiC/UNVn7uSDz78p2YxYLel+ur06MPV6k+m/QN
+VEGtjGAdRUvRO+wHYv8ugOnwEsHVHC3SVCjUxCOyp24pWpc1pLpjAIWPv3GJ/ig
2JvfOhjaHEeSs8bxibTydH7/U9fIB4iBPWLnkw8wRyjCOI7rE5gf4798EHWlnA7t
iNwFPJCVbLpBO7eXxGBp7cEZ1wgYgLfv7r8RYG9or0Usv5guEIl1p7E3tjj+d2x5
GANqElbXjmF10nAZbt3S2faX9Kr9svhlDZX05oZNelYEyJTrj+RgHEQzEDJWC5v6
W0I0RFoENtyNcwCIJ/C7QX4brI0/iNXNsllYErO3tvzOVBGL3RGQXycb+7/vdep6
N0WIcDxLfV1Jzt97+ascswV8x5N3R4/JFt8Q8rkEQr+6Zs5et/Y9tppsOGn3xWwn
ysl+UM4W6PhK2dAMkHCw2Nmm2L49GkGPYCJ9h/AVmBRrcLkrPD2KB4DphKzrFc6r
/9CIJSNrpd13I3Nm+Nff6na9d31Ux64aNHHuOSXAvTSoqIzB7+6vRsCR320NbBJJ
Av9zjW6j2Z77p00YQXWfXOPKmH4ualZS+14dr1r+7Ujj5niraBLsSvv1gsFVQJ9v
c3e9Zoo6TrcUU/ZmwgJct74DG0V5Fz/7y0jWMvLXFOCBUpK/9m5Swq5qoU3i07K2
epb6BjnnUObBHvw12E8uitiM2Xs5OB7YIFzIZ7+7CbrqsrxsfiOlY+MstsKSZVmp
AyyxqTWlzE1zbvF3MkNwiPYg055tVHBM+p/yOnkWzalqOFtzOjsxbUCh7ICEpYA6
vyip8fWIAm87PVus8bSnPyVr4kgqxmtmDwJ5O+9bw+jwlFlDspJwtk4MGdgrQvdL
aOFLeNpTyY5Hl4DUCLBzXe2PC4j08Nmh5crN+xjmxON39kyWwwSAq1dC+S2nODaA
y8lbt6b8fN/qH4m/FceAPdV01svQDmZsfo9nYQJPjdJBWPUJasws0krmfn9Bdyty
Wdu+6NO02/wk8AA+xZ3U5InfIPaF3+KPpOc6fWqB6580G6cv09h0CUER1Z3U2AVP
iwIEIhawQG/wqza2v3ywJiAeAyU77yP59HEHmlusxMnN3zEGER/5YOyXyApqjVcG
7yhycE46gpRnVUH5VFfjbYdOQ7FSvNHwrIFKBGyYS7DDPAwEpnGaBBWiPhSvmlAs
1ZCFezhgKG+oBTdTCgAlaXvEbEXgsDStpPgHJldJDDifvoWU1qxRINpF4qVp7R/l
GovmtREyTBkYd35h4TNqEifVWs1Lj7M3SjNvOAplB2JIXYA5sFhCzJI6DFc33oJb
YEgYLIjCJ/nfnYIvjAl0B0A+QxJHQffQ1u+kGRbmp4cQ5lRpfxUmsOv5oNF5RkBu
qDsFYioN1xwAxzF23A75Ytww3dgoF1c6jLMBlBxxiguNKCzoPtuCj0BTEzust7ea
UzQM03UR1NICCOKrpEDCzOdKgUTFGcdaZgDMm+DCXeffrbcxDFkGtnOODFuPnnJ9
lMJoVRS+vmil02ZMz4YbljuKA1+8uSm4l/Wf3ouWMI5561TqkaTOCihT60Ef56aX
JsjBWw3XVwwRiLX8M+p0e1uERUZFvmxw27gCmI1mBKgluT99Z1aek9amOl2fCHU8
H1m4Uh4mrM3NoNAMEGeQTjw8cmzdrWdzm7Wbe/MDq+hvc/ZinUnfMaitqMM/N+n5
D4JZd3pXBjmLa4qWwc0EQIN0lQvGHoKeIqgP9XyG2K+KDfjgQTp1Hcis8/aPIw8P
OBTu4jEpXrMWqGL04wlBR5HI4Xy8hzQiphcSV5kRQ0EkH2KliPygxadPiVEIKg2B
rxSpRrOOyIB4bI3iKx7d1nicOlhQ2FVHL06fInw/4On9hMmD43rV1sZDPxhT4epi
gfbKie/rQmPUorj9amQ2UQ+oLVC3H9IZu2bI9BDZS56mibV2xLqvPTl0THzentOn
hxwyxoR/WMLApJqLCvS8QDe8cr5gWkcPnapZSJoQViEMgZ6d5CwapKnGuayCPEh6
mGpD0rt+x5m537yhyVXpXkSbHUsG8zEdjnBtMXQ2XLrMIYaOz5Su3yhZGct5PYhw
PBTLgACTxF88SRMGtBZt/QQBsYBDYOsM/L10yKGeAnWgx/odl7FEV+oP3l/hskQ7
a1QH0gjIahLliD0Az4qOVlhSo0IfM9TGuh2/yUZg8lEpBK49aU2pwEJmaNbIVUvZ
TmMP49o7vO1lxt61mdDr/cpq7xwKyK4Bveyf14YoE2P28Of72EzpCgc2VhVkYVKl
ut2wgUh74pmLVEvlqSQgq6VvWlXsrrBE4gwVcWyzobWjF72NUkFCg1jFkFWpu6/y
cmb+YFJnPgX/aLh6Vu5bZg/HwHeaZlWJK1kMhoEWJqITQsmI/Hp/wNdb2Avg4muG
jQLVm5xgDdVcYaHriQ+8Xnd95Lj5jU+XR6XcWKVuPpw+PNMPBFSbvLUTGNJkNIHL
FZXEkOygcWLp8zqy2KKE7cjnGKZ17oPAw2klcwkNHnZAeLh2GouujeXm82x9mpox
H/SSBr2bUbyM+cYIvCy2OE3xq+fvxawpn2XmNVpsbktQiVPmbj9x6ISW8h2VVep/
7O/O//GcjMHO52p7BP3d9599vduZHDW4R3EgM/YIvun/iCjLzcBGXhhUHtHbdWKb
mViC6EQ+PGKtBp+Mu7rGdj0ULFW6JHlg2qXyFVUTshTNNXl0F/zVJIFO2x9JwUII
Hvxme6Y3//16GB9IhCzyBoCyjKV2JFrQ5D2aQV17omL8mOnCjYa+QfMhiec2bLbV
ph36xqjGf4bevGB/MW0HlqypCZEjsVxQbUqyhU8SdbO6mv7yCQrZGGaX8wgQu5Ys
6d8yUBaUyyeRWlvMnohEl2zpvak7vT93AyxifBuNOPleZ22Iq+UKiWLX8U8jUmgh
GKpnkU4qpmjYg69YEF44Jlzo2XF4x9C1wI5X6hTnyzcsgnR2V3h5gXSprEXEaclV
I3o+MlZXmz/PP/N25piK+oncYmwVnWP+apDOF12dPIVfEuRsqxXGDxEXvZty9RYw
kO/sGPENXfBwcxjuq73QsnSrI6RhU3NjdgQShVAuC7CF/jaJ2o85BpqQaW1fTeGb
kaMPvs9LZGuBflfbrjksxQXtAlGmQ8Xls5yQoFcKHBc40clxqQSLF0mj92my10ur
10T7SeJ9gswQcsKSmuw9YRB27sF7FlIfGgNRJAVgoa86iR5ykT3OZCuA1S88AwXI
U7p32Q9b5tH+Dfn/PwU4URLksH67qAPtt8/JxV2KcrtLLEL73mqd2GL/suBdufER
5Oe341cVf13IfGhav6w8U4sZHlu4S0KKAWelw03PQ4jQi2+hkdcySz2ROPZEvnCr
uKNU/tmctirqqoosilQwMzR8n9PyJxAP7v5ejEVEOdK0QvRbicZWYKhCM96WwJXa
q3zN9ABZ63uxyrUdi90oQCfo/sNitVxpHAWoTwW+NuY9bUcZLNAXraWrD0/hQ0ps
w2glHhxqTPt87O4soh3YSoJ2Mz7r/JqjPdwDqXEpPnKCbz5WvlIXH3lk1oSsDUz6
hIwx2ZJDpxuG5arJne3rY5amcLSInuBu9BEwc0QrJippqLVBFC9qbTYBWt4yJpsL
q2hMTes22nPZb1Jp2qi7e+23PBb+sytWDXHPnUdf61cBSXBf8vxWD99sb60LVtIj
YJpn2HVNy2PrYeVWsDsM733qmpxQ23ZlpNM9gq3ZCKzP9i52fMyRGvwKqzo8p38t
299euexmejmPXSZ+1ih6H+3xiJJU3ykZKnA9amlZNGOkKeUKKxDBEj+h2s0G2otB
yKlyHnWieO+L2uFaUyJ/2cd7zOiGt3xwn9wSQjBq8GpdSHz0C8gXowrwElQgMC6j
0oSBRhHWfKNzxw/Rc53MiuOQrUMa9II0bSxr/1mJPrinczukAHNzPTroEJFXaycC
j8axUjYMoqHY16qqHSLPS5uePNI8n5/S//U+IAU1dC289K9GjwaFZlR3DdHAWpCf
RdZ7v+0SW8XRWoUqfP54PrA/S+iJdoXEvUXO4I4d89fX79g+kv3oFhd0KsZij2sS
3BNcMUvSTQUNJogPFWjLnHAWkIcVlo9tVpeeUSBkKDJQ61ACijxV7TdQoYvQpo+c
cqnwdOmEUpJ5Dz5M1f8Y9x3PL4pLfVo3gkB4e5dbh1O2O+IAxJQ1MG8xaz1ESKV9
gGuTiRHu1hiMaw2JuogUgnDw3FVb7w+efXTgCv6GAv9yLs+mkXBSjfpZgeTQ+SiX
iPgGRn+Q+VGoGmlz93xf6OMvvkOk0T5FyZh6pg6+232k/nU8Zx8ELTk8bJ+YZ6I3
dzpIty21v+mVSnd5kAn5jHzndBO9EPViL2TGKx9g+nW/2yNl1/D5ERuyz5R4JIQi
VCviLw1K4ggW2JfqvqFejCiEKBl0aMA/kQI00ZUs3kzO84Ej5xbkbhhP+gVz64Vr
FkTsvI9tlNEPdOfkyJ+Q/jhG92A29wh6Ei92xmDTfhytQBVnBc0QfgCIoVcYi9eV
71RAGcUBFn/AllZB9xBzSsM/5RnUEO0OAGiiARXqjeNGEd68OFLA2vgSkyYgM5cy
mSAJzP9Qfk5/ioGOFNHx4dBOb4K59cZpxuvw/Rul0Ei2ZXlezd74joZY50uGC6Lh
8iqd5BjNv1lddBUlKR2HJayJuYswi7AaoDUkzN5NQauzewQIZgrrJHyLj+Dgz4rC
nKIs2GptD1SQSH40aCSdBAsrZ+DNG+k3hHgzNRjCLsVnYv38OTqupDgOzk+lPmVB
FXjdVkIqK0cqQ7QjjQWleoGkdTgE3tH3jw4tB/MUvIttN8nm8YWdouZd8umTIIlQ
0bD54Dj58qOKf2gfX8Dz2cE3447r/5qpiJoqjtkuIHEe1pazMQyhQy1M1E/ebVCa
61SQUkCyifBmNWJe97bEPE+klkQ4RxzlUu698QU15dSEVF0bBjYA16uvd3Y4/yu6
UwgUWKs7mtNOfwNsAS8WTKflix2fbVMYCHG2xqbcXr7ecrHXBsl3xf59cO6IJMdk
I6e42Sv3adgh0QMIVa51yye8ajfneeoNmKebcVu2RUDroZRhdmNUu5ExsPwCjvEr
sV0XpPkrn3BHLUqkS5nX1r5JkvlSevufpkfbehcnrge5OECqOL+1+kPd7eC97/Lv
KtEeMdTkJ7ZT4j4ALlKYELaNlhi9R2gQ53EvHEEXmiPNrH5YADThfNgNzC2zNt+D
uv6tzcw1NdiMovPLX2kRByqNcYGkbC1Pq4lLgn5uuvDais0AEvGXHK5h4BrDtvY5
iFUTVI7n97IBQ13COFBrq3ZM6ffZfFYvKqeRKQc3Q2sW3yWxPvHZFhp8gw63211m
LK9q22Enh2nN+kkvLnTasw==
--pragma protect end_data_block
--pragma protect digest_block
CqzUI6ydckIN+ObZWLJVLRZ5d5U=
--pragma protect end_digest_block
--pragma protect end_protected
