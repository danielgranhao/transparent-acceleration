// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
Y+A2ljltQbbe7ru7RQi/Htk2yhVnkm/kHFUH0+LJx4m3AuZ+UTJ82TbACHasyAE7y2EpiYLdO6p2
NHydsxWzOR+4iYd6HFmtmjtj/6VFt6iFU9dMCDLy+iop1aJS2/gufSZIW+pL1Libodos1+3HqBkz
gKizXlYmTpsP0csRfbS8/tPnvAWe3igwaOlw8ctvHtnbQrNOFvKa6JYuoy1UY+TviffB+wkpzZ2a
qfZ2NNvEK1fZMrBmomVbKz00mtgL9mUelvDK0gFzBVIGPeEdgsfAPHgKIp45bqW/vLOtNnIGEHMi
IIv1qDjQQeyO7D9fzuf4WeVZzeWoOeTF326llA==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 10384)
qa5nEe+nsVXDHZG2N6h/9bt5U4zo55PBomc5DhzNQUXhQL2KipL/Rfo19ZdRswYGYw3nG0LD9JqL
g9Dzqb47y0YDUP0Kqm3fLKhl6DSXDDdrzSEgrdHWf4GaMMgTZf95/re5SKjOayn73lprxtWZPi+l
BGc9vtyiSQYOuTMZDxgK4eMF8NYfunKeowHeIax51Q8ohnmT2vtAET3g8JuXYIYoZn4WNeshUA5P
sg1nwdHMtfAF9+folcDl+x027oxTypk9VJ6RGA2or8rOYNXoBxZwKnuJ6TKJH9+JmwNqLWavQ4VP
67itvNO5QqyCiRiz4zLfshhlPnVWmyOM6Z0F+EpSlMMbpC+4gcxCTzDFvxeouFZHNQiNrjD6LPWR
pB9IFe89wre5U9nZtqZvWYSnzxM0iwJAHvR0WmbnbHHpcXbxVOJBIZS/p3+tgYTTMPUMI81b0dng
xp9RG7DaPQYgyuPAAwMpuMEaNonKNzLj3/Y+emKLLdQvpk0LscUAwpjlbBOVqicWrt8D4F0EYoFX
eWp8X4DjWUgUepMQSu+dIWlkwlkHRaAFPy/Fw9X3czY39MKDlXnesjYz7m8OPBWlZHgLICoHylLH
cKafYSKiUYDW9vd5vD2Ig9/Y7RZPUSl7fJbgB65C/nLokxGgom0paZnfFIHR5Pvt96JyRaPFJW+7
XN79PEqJ7gmJHRe1a8awYN5sZmikkNmJ2L4HeC2KFnUg2Lp4ZO37FW/cQBUSRwVi4Be2SVwls/ZN
JgSrYkuivCCPfrrQuDrgthnL/0OL5D95wZbzZqmS+cMuhkDZKVIfzYZXRym2/m/RTTW7+ZL5YgUK
imd2XxWAlDzWeaQBqnvQ4nOfTkmBwC+fPG4Vx5UHclpR3nt+2fRa3k/pfkicpIL9UJ/GvUxldp0I
IpWnSfn4Pb0szULlJfR1UZGim1B38miEal5BeRwfESd9Yc8OZsQqvVcMTd9qcl2oCywlAOjgOzah
j/EwmVWpejKmrYuji4zbpUVRDGDVk5ToPsJ9+gZGFc7B6HapaahtUY9HtjRro6aOtGDWcBliK205
xPHEXEPTiInuRK2OowN2TA8e0Hvn0nVePbajvkTZMCjaro8ZWaXfE7Jpiba/jtd1c8072GavSDoC
KQC/unHJGKDeqc9Lk036Es2sjdBeGfmTY/4gKJFB35NaXWsCt/h+WJqDNAOHvjbrHOkCxMYC6caJ
RQRyY0mqoJyVYPmCzEWLxCeWX34DCXM19qhoPjOW0iNO+6NM+hTOJsK/WWtCmvzvEy0NJK+DiMqg
4b3vJNs9a6m0QfhW8a/GGt58bH0z/w+i++jJqfCX1g0q/GNZ5OPluf1iQLbnk2avwnyiMx3k+5LY
H4Q9CQ78vrxWS6As68tlCDi5fPaRt1/a0e1PB5vMqtTKEE+ktaAEFEsrsolz8aCxYMHTuoaJZGZf
6zx/qdTPNlvd7gKXJSr6A7w0NrQxfXtyAlle5bSuK+QrxI7OsIU1ac2fsJlaLonqJ+f63xj6RQR4
qLNPV9AriHzOy+IM4N7IscItTzHtwhP+6guI6CvJPSJmcoqM5de+HXCy0w8/8rBWzZ5ae6VNGxqu
vEsm2fyTzqZaYdJG2b66yXDY0lK8SzptbzWU/kmgjJcanygT9OJUZueQJWj7UZPvSR3OgH3EuhrN
d14TMwb1fETEala48HBSABtuInCq95oCzKacRp26X5Ehx39o0HWO/ZpC/McArG1IWVnBL/uAjH5p
YO/YeqZb5s3E8POajya9i5/ZN7qoehhn5i869aiOp2Gw272iBC1UbuHJqC6TZBzQ/hpNjnds40yN
exEfj8gH1A2H/Tlp1zxXBhpvu1JScw9H10yYwEWqNh78Qbwz1Qa/2EdZzEiunMPBoe8o4qYpHVeW
aGJ2g24toERF2WJbJ/2OHAenTgpIrTX0DwsJtMSCiYWP98bBFExeieJe9ocIchvpMmgIkp4XSIIq
00AJf2B0zgSNlZ3sL8dm1Gm98w4YuGUKmmMD6BxgeaSdIau3itLh7KkqPVt5fQlMxZC590Jzy6LX
23Mr/aNzTj7Cl6b2HPiekLEVjyPCmRuoBgTVqV2xTCuGLY+IbA1Vg1QqjAUJIWLnbCXEe9HfXPOf
a9nEBVsWQ7HBbv2kC58bNeupVGarhL6lvnqYugka7MKsmcqzWPrNrwGiJSNyabzDlY3j885toXXm
rboGIeCvFyR5hhmkp3HKo/fjqHmZvtK6STQWOE4olxq1FMyEiQmkGkJx70tjjv5TisG4mpfAhrVl
ciG+gxV0lQaCnmF7Xm0wrcO4TpEosDovTYBfIjoF3fbpKyYDGQwFusxa1rspsnpizeyUA9XkVhct
O8qYLvNwe9WoQrhYDzV9+gR6w++9sQlPPp8wIdBWtCW/i5nNVS57LQcZgVQilKS/Vt1kNWJgIxoq
BfU9ASH6tvcgUQrWBicuxinaekDTRliOKD7yB2+0SCun2HCoNxh+Dpsj/GIomQpMdSCebP8LWxY9
mSryl9AOBv6okzz9rfM3HLzWdORqnXg+5Wx/uBoMp4EusnLi4NIg2rjyL1NF2KUQNLzLnqzKEqH+
q7UX5sJRPLzN0JFLAfTOUGyGvyJA33rj6yITgqDN3ab+L/LTCkFSHTmldV1NllLfK771o8c7NJES
qTHNwCdkJTKBkX7vLsujO+lbFrfTivDHhI9PWJF0/7Gx8cdqi0vLeHDEWJtyw8zY4bpyP/p4Di6Y
R5l9mLt2UcxRVVAk/jKoEcR/JJ3FYBn5uF39ZTZKi8qQu9cMp9vPqrbgkCc+JpjZeC0LZ6/tkVID
HLv4ue+xHutt8cqM0ivyTbwa20qh/clpW7pbrQx+xGerkPyDVTERhRdxJJ34UskNSvOYX56CE2+Y
P4BBHyBzN3DhAB3rTJdPlC1NqFVPk2YwMoNj2hus8zk2eUcuoljwDX2t472D6jX7EiV/n5nu7PXV
eTBpvAYYrxnQ2uVBKzFacuw7VKlYIcqL4hscpC6wch0GQz9ZIM0CaFIuvibTOOSs5trvhAlxvlOO
1BKWVb4uVQEhADjEOwUEAwjNyJHI08A0rqTHXEo4ipnBivJp0RT+hapoKjBSaRUDPZRRGd5O1/Xd
L/9I5c3/4uF6MPITWJz5uxi9CXkisWnU0K3cGqf6toX/mUG8jpM66RSyCmBMdunuHC3cxDO2Co3V
Uj5Xqai0NQcTIbQ3J/N+peFno/WO1zz9JWyr7gBD1DaK3PrPnlycF5Of5BSmuD+gP3DxQR0Piuen
8B0I+bUTmDD9DtFVvNKcBFWfrVgm6aD1ywNBgD6kTjHkt+aCMQHc7m7rveUHh0K/jS7dI7L1j0L/
Bj78mIstx2LONFYEN+HwldI+caslQWPiYuibSgWKbjaZMp9TmCm552r0xn5+JT2X+UuGWRGg8PJM
KphdNQOmU0+jNvbHbEdNePguU2ahkqzb13VgVeYRXARu+9txeDE+wqtQ9fTiEK29Iun5e6CYXF0g
/bMBdk3gjdDXFRK9PPyWusqTFBe0bIPbyiEV7Uf6UPqko8G+rBHbd5bonrF4hNiJwlwfGa+awQ0g
Bf8nv++SCr5FYWu/eOwrbfmph2z8G9bHHGimC+73dqdFMG2oySXsJnc2/EaqCJpdPAatE5cwNOdb
5wQbHMYFlfkBVbLteSuqPXZ25excXt+Z6EUlD0lRwkVZ8V3r2LlEaq3EZ0zI3/vSM58LlcueB2zs
zyvpd16WC3x9gkjUN2EGr7IXrtW8DIIPsk7GS5j/3LZ5s2G1SUSK1PYvRWfs7XSl5xaGojtle2MD
cXObd6rKoxW1xXdM5Ky/xfo9QnWt1v1ExQ/3BgWVNDbns+yF3QdLU7EoiN5Dg6epu1Lucs5aScE7
HlZT43hHRaxvc6t/XnxnliM0Up+KGnbefbHZhX4bzmrv7h4y/lBJGEsA3mMoJpFbbdUCsRs8nj90
yYR1h4b44aPmRWVwEnk+y2Q9dejnNlQShMcXKYD9BzcOLxVJf3WXzOhs7a9qFPSLNfB4y0tC0r/h
kZZaa5TqJKa8hQ280bi7Vgtxz2WkY+qCk9bH4AsD36Cg1GgrpXAmH/TMhsCRFAVbrSqWDtyk/Su1
BYS8IktJACLJHq6MqHv6d7IYYnnFHXU4+PGYsvSM3DK4HxbN0OzORWdNZ8KX8LppBvtDwWP6SW7y
GotsvMpAtM4Y80Y8iZP/MtDOj1MwE0rJiDe65OPj/VURSk0QOqyurLY9CzjffqQJnj2T6gcJXszi
VGAtWS4Tf7wTFXKXRKNErnI+kgvY0dfVNVbyd54B2w2NWbGS6l5duYCOv6uO9wrMmSX9iNkpEswq
o7SQyE65TyvjTNw7Ja14KCUT8HNU8Quu//HPk2iznYZffc/XBHKmJCuSR4IVhcgk+5rygEwhPQhO
eFZ7wwxKI1IRfoQkdIJ74wy7pIzRF1rdkseQAO5YxOO/tUSoJ4C2dz/CRl/JetSxY63ZVjKsyvCW
6F7nP9Ash2QsLYtpVorhb8xL9CB4M+OORP8swjBuy25r2orY/jMLwEzGumV+HJ7AezIi0kurjlwa
UuFYqvTEnncTcEayLFQtXpja2j7BvJzno3nh1rAw06SGqjAVkHc4IrHgzFgipdYGvoLSO2CsShu3
XCjAl3LKTe4hFujJSGzJl9VgbTeg82rkS23H0uxLS4BjHyDLEBr7JrUSSzoXo6EFtxINTLkNGfqb
XY9zjNJ7+xL/Fl2btgIX5G4gG3HNM9FX29P+zS7OGr7UffTGzFCgvMQkKtOTpZL++nYm6GXM+E85
BgtI1hdaQ3fZL9zZw5gcZ7zjuqanOp3iyWRiXdL1EcTl9PSxnHI5mZtq2ICBr6mQewA2I9RJ7yjI
D99iSqDr283uk54YfKYvfFluPHIxEsQl31R1Gy41ZTtg3i05jbWdLWTCHlnrOaQbYppN+t+0ysUn
lBUwK53P69w+v3r5YD6q/EOouB/fgj4ymcSaGsPY8gl92+ImMC+mtfH+rV9w/o1vXt8DzPsMDTTQ
le52/8kdnJOVabnisN6auvadFDTVC+g9niXX69S+MK1WU/iibRYy0uOitFGC9+qzkXRr6IUyRWeo
ABbjIPd+sbt64V3ralFezZlZT1a0WOFNjJgqWbv8pb3tp290mrVub2htVB5G0CZT40B3qO/6ka9B
Cn4BDJ6etArRahfku2pb90RwLlRxwZBgo5pg7VZMDqX7OJoUb/f1eh5b6DQhjIjBhLiUEngmmanj
jLIe+2+DH0MYV3tWQzgrdjKyPtMGYuXExXxkPvjKa1esfpxIWiblVkKi+DuFIMN7rwicUpoqoZ/u
O4YgEHFIZhT+XFdnfDWlxGDGftzeDG6fxO38IOytj9NrSUMCcqAqsV4CRIPmc2XeI7crIJ+q2dBO
aHHzhQ9SsU382kLnqVgiD7laMaUwX2QB6UbFSyDQZCqmPZN8zaMd95Ia13TrL4p3D8kH/BHD3QJI
7bVwL8/dOonjSR9k7Jbzb3/BkrUtI+YtYt3El6lPCA98f//CWT+0xaCMgYoKxBV77TQ7xOle5ziI
P6T+o/jOVqWaLnzgPzrIrxdOIPk42wax8BjhmalWYjhGRF5eRoXDUlCTAmpPP/YUbdshFDnoFAQa
lSwWFBDOEywbYhy0E37rsN8hTDYOKTqgPIgeSY80ON7L8t/cGvqP/+dBM0Vmzah000lirODKb56+
fXaNLihvy0jzKDVhEsO7rnjyQIxYy+1AjcrRW3MeVScmZgfYtXFzkWcYwOi1YBLZ3+4nc4bNH15B
DifChPcrkMJn5L+dkSJcRuWF2leekl4Q0Gbk1AhWfSPSca/OPVAQIOxkBLjcKXEHakcyCYNQTml5
bVmfiHR4iI9u7+VK47CkOkUwX+5smXFHOUGOPVljcqishDX1bm+9cxPka/DATal36VolWG9Wmqe+
n0ceGweysW9ztPvsA6fqhLsjaSYuxPD4fD7Gj9NEPORzh9sb36rcwQ9B1gwCwAc06xpgyVpoBvqH
M2zhIYNE9WmLfbLsP+BwsjjYdv2Z0D5YHiNlBkOeh8NaxINJytAVo8Tw65vL01G8yr/MtaDk2O3Q
Wk5KKAbJZ/TlDJnU34nSirGLklvM4EDAb/w5YgleO22EltPRafh5tFZO+6oYT54VGh0AmKrUuFPL
PiTGNq/PnjIZuT2RpC+IMBUco9Gt8cGEbR2edykVkLDg+doVF+W+bM9YCxqEaEICJV7C1lThdhGt
m6LD2po5LANV+dEnPX32ZWe1R/IWpCwikzk6wqYb5wz2RzVtj9SeMKxeTd7X2tcE0FbqafTP6rL+
bSpALquYI0o3Da+P3ULQ+V24yYQ21yByLq72dTTnQM34Thzziqh73B23PcDzVP0r2yoGKaA46YGR
XdK7i+BqY7q3PxlsE5M6nQt9tBs4Z7wga3vpwgSNMdTiKV8YEt650raB/Fco7pZ005k6kwmai8Dm
kKBMIgfujSmn9U1dUxcSQ5P4XdANi9ty3mCW3r3dZn3GIfjDG4NCVwEmFh+Qudiwa9cpjSUGfn0w
gc/rPuEu2Z+JmPS5YQQHaxZaZlJ3qNf5ZiqqiK0D1d7dl8ArJzLaWfBsTHDZ0vSqIQVCSk4vs1Fj
9UsGeR0loOfGbWIdI25JcOz7PNzGiiKbgjTVaTI7fcdP9n1KvcqRgHBjKQvF9Fp5emgzrox9LMe+
dxTuPrkLHjlS0uUOi6EUJ0egzB/0fTt9ejoUaEFti25881YxgAd4H9L6WfOH5d+vPsXoZdxMk6hy
1Qz4zbL8pIvyTwoWKUR/Xz+VxqDuUC6paaHBdZnB0KUEiZ8Z6IrWQ2w5mz9sAD/dlhvWE/32V04l
y+agd/9ABJXYiQA64KEUiZ8ep8ERG0/ZUN3rjGenBZ53juuo3etEIoQXdFIIiwvYpqjvE/ZL1PHz
ATkqCXPOazZ1s9178DQ+lxemRxAcwA2ybmmRSeDXdzZcv9t9WxiRIBYZIvsdJJT0lr7wJlKk55ob
80BWaLw5fuToL/sQEtgv2J6b+fFG+c/7k/RlYVsfjq7bFWTircslkwckHMXtRo+lx/1mWIgrf80G
/w1TG4RG9K89/lKY3OsL23H5apKn3dydKx7GUI1uAPr78tP/0mul0briSdnPmSe3k3qYYg46GsFS
DThqRjx5dHFZ+ersWZYJFRJjQXRwzy8AmdzLWpjHdfm0M075M+QJ8sPs6/gUnACVq1OYMqkKW/yo
XzWS424aTLEQNhfw2fj6qrto7O3ADtxBuzsfOJCqDP+5OH6HVPT43meyGU1y6bGxDz37Noum16Xw
NMsrNnouCQkTSgBqxXfpwsq2UeuvgDSIRMZW71aXvdTwN8zN2J9iNI9cvOmQatvhxrUZ/eGmsGY/
el+tZpnWronRycVLVKdb3z/guRe/xJJKdqOnSAzqAYTX5zgcs0O+S5cXq9NXHcy4LKVKiZ6GHqpJ
I1kLEm09bWxbZd36jAAoqsRePrSh5wMlYE5um00UfHoUtYT04rm6fMLFF28fAly/yC/H4ZYP8qy4
1PL2OiR/hnxhTAWxAbUPvYXAgqQiQy9sdDkvuUTZr9PK+wGf4WjbfTOw078GvsqUovGuuVmHg+db
ZwHrpRHOQHOkjJ8o1gXwQj5PoeBT1v72rUf5DvBO1gvOPxO61zq41q3VWcLBCqF01nvXk4Mej4ZK
e5xRVTCbxZiDJGXXtVw/V0wICjKd4wotwdh8GYpLb8Ot9lkviI3YqyqHNaDYhJE3h87Nh3a8RhQx
5NPy5P7EjkbEi3weTmkMmN9bkESzfQMLPtELyd2ZfMNvWBLxuMXsukLNfopI+PpLMVIorxtIdZlh
Y5Cbx8E7RZe/F6Ake2N30hWFtqu56HTkGXT3kQrLJzNNgaqWcNEuDY3CyPg5yKhKc/LPzzXauaA1
fZ7DHW39I9XZzf0qHCHhP9ZbZBrmYBgk+pl2ZcNQxnfaxZSZ+C2qeRINteCmT3ieSa0xrIgMXrTg
2U2K13VS7Q3lqymxm+LCus6YtU1WeGKqUL1LPZaUBxAscNxg6RinikLwNrDU/W5XYmmN79U/0/o9
DcMueXYtBCEBLD62oXkmlmzcTX8UaolZN6HTaGUKK3i7WbX5sDaTSxLUVDxWuTF8uV2Rbsn20hmU
/zwKhcVMnWYZjAyGkkyDYlML9bGarBcaXgf4p9S4IK/cy72Sses2DZzV+ltwXz5wJ2SqI+ySJhBT
7kWVziH0B6yl+lWpMlJpA1bXHPfzytadu6nERP0Ewf9PiSQLp2lVI4b/LGMwZ+Em2dxCFCUeKXmu
CpdCSqOPP7AK3MlmrQD+odA5fltUvtQiU0KiA3Hd+yMHS6Xl/IJAmMZnM0TWA1+1ZUlBZb6kLhag
u594F9sEbnfZuwWbEoMCXSDqOTilj+nDul2xzP8MAF4ASUPJjIXxlU8n7C3WfDFvX0hVxNLcVtjj
DM7RlIDqrCqA1ZruugUJLu7XlDYrvN1FVqjzVQfniGFAshKzTlK8nacCkC9Xia1RQxwIP2AFLHFZ
UJOxtXt4MAH5idl6CFVoGSVuEBEhhVkE36NjxmF5VpbKrmsUz4D3oHFPcjf4Xd2Qd37FH/Wv5EdD
CpmYDZ4pzJUwAG1r5nh9smkyVGikdOslyU3+bOroy1hQ7nHIF7kP5ZO/eXmTSzpczGgERTu4kBHO
1GFdoI84nO2nL8S8UYVoxGGdrmGzwp8WO0GT4NXxIl6Qz7RYYpywjPTujnYiOxh/q1FOu7ZEfxuA
0YlZuW8NQFJLOZI1dw5f5xAMm6mKbmONgL6KQSIVcoT7irYS74rht5k0kkyD15bxS70LFgb3Ueed
maV0pQVZCNFebZEv0tUE5/VotU3H2urdRhYeqkaz9XYvztX6wLMpGjE17mz3s3BI1XPU4N9Y77rP
Zw9SKPbOZ9Tb5UAtHRBuG4VKRBgUfvH1/GslCJ1r/9V1RGERxcb/H7N7mj34JMLgcMr+b3+zXPvq
BWtIyqcdvW/bNTV0YarJiFFldq9hgnOuRZS5Uhn+SxX0+FoHoUFdur9Uz7y0gHjvoDOkGVymoRUH
zWaLRLJsp8/zPyWk1PPXiv00P5YqzBcjC7+115jIQ+eNo0nA//7JdkN2bdyGgI4UTj/Fa7v68XI4
3CdcU+9BvnMGpVbbOMUP5D03UjnjSBKkQqh83m4WdkiD5PoEGQkXqjvfNSbmazCeyKzLl727i/E3
z2F1dtZolMa4sY3JdISf+qUE878x/rpX1C5V3d6hA2JMHKe/faRf7KZYaKClTP3e4HmceV0UDBEH
mAezd2kAX8lTnv1COjNYd48+27zxUSEMvXHbhHtr5cUYHnl+UGLOGXuI4+ndbiMaTNHrGqWnLc20
kQZQ/iIY5M2aznvKH73whAP16kmImOIbMrSZREJt4KIcWh5NHJArIQ8ut0plQqZcY1dnZ+gB3maF
YwlbOQoNInxzC2Tfy3xJ46Ek8ypldFUtn/nZE6YtE/T2aISkr+NX/wCO/9Ly4Q+z1LlcWRfv/jyE
8s8ZzYanVKkniaQGgUsNbA71U3DONvNtzbZsKpaVk0LcdUbBSWUw0LuMWVrM4bzlpD3i2Xj3BFl8
xF8uwQZ1JT1vsRtFxde586+yBzTpxOSxSJW5jA0QR5dudeN/5jMTqYNW8LwmsRbmbv1x9bcTTWhJ
OE9JR/Mib77i1pzkZPZ3swgqBmUw9o9dSw7/pzpE54qyF5o6rUh56v+a2SI+l4wu7LH8sNmvkI5U
XZbVdDihaFR1IyDxy0VXXfCky6XtMO+98O4YYInIwEoOTAtZn40mjWEs++HEDYg0vEuouYgtVd91
5B6MAlj7mDStMMb2qrVAoDh/zdoHYCXFaS4OWxFJ5nbRliB4VGzt+l0zSLBA+9q1OxZxgxQNVWiQ
lBjna2VZSJxMWu0nH7ThIeJ8JGyb/ioSoCUgnhdWoc+69XNi5EcAs7QEXtCUukOwjTTssTuc1LXv
LcnkyFQmEhSoKgTkgHF+g9sl8eSynHEgS7QqkFxDOD6k6BiUO/xEqLVl3gI1llueg8Wx/kyDmh1o
qF+Psgvb9u6lhd3IAT6pCkk0Aub+gGbktITR7tEZ59OSB3qQiCDyxyJ2hhsLX0mvEX15fnvVOG9p
KRPHhYF5taX6Fq1Clnfq5HS/A+/hl1L/QR6YKKXuysQxPLUQnrSyO1TxOGqkOyltoichlxIZNv9V
pREy4uMV9SYNw6K1qmQjp1LWpNxki4q8nfLZ7Oq8ka1zdeeikl2wAPGA+6Uk/J0XKrWOxhNBlOr9
g3SV1PqR9JCmM7ksjc+tBq/QLcJpgrvzBkMxHDWHKE1VLOCP1SHIm8DiEIXzLuW/TtcwKreI43Ck
irDo49OvQ1V63vLswwBO7dkCfW2n0ZeFBRKh03eCjw8WKXxYUnVY8ARTQevS7viNuAlpC7URRYr4
DXDkCj+p5dHx16s5q9bzT9KX3FumcBtAcCnMC47ZS7lBpQK0w6kykNrPSfsNjrHyqo6nSKXd3YQ8
CcrFnwm26+h2aDSnMfhRAfzdIbI8sG8aTv7fEd+MobWjhVSJlEQp/ywpM6BX6ybxko9jmSstLu8X
4hDhCTNx3IDiIJg3Q0mp0S+MQrT3fCuvHCUCXXpm+t1/EECtTwjsZzZ6RafR3BDjuatQzvE716B2
7lCsoo+EFCqm6nOtgzeQB0trBAb0yu20c9d1v7LX6s01YN1PGEz1XKBCTHxQJo6zhUW+GHvThLJS
Wb/ze/XuC6LXX+jJsLJEFEJQOm+5mrTiwvuVLRp1p8m7nAhbASs6ZEFAv0XaIbu/rPLdIrxp/Di+
3yzzZkUb73DGY1gTIKiI9gLm8k+rEh8eNca1fitfnreicsyFt4DPNGyKJiYSpklxJbKYk2z9j74p
GmOLGSZ6nrjyhmh8Ufob+aWGT+xNVLBn3Q35X+xDAV+Ib7j8GqMgVSPK8ifqbLSB/hUvNfhiowzS
xkWdmeEHf9EPNna2c/H801K+FHY1O9DKIo0a3KcE0KSweoX/7t3jT+BQ/j+INcdluEa4DMcVOti5
o16SJn3XNjWMwm/9XRak2+Id6kPq8zSCPfAbTVSDVtj5mpb4kXeysJ3octnY6qQeYNn8vAE5it6D
2irF4y10q3/7ezuq2S8bTw9Hl1Wz2Cmb0GWjDTCyL1WoANUhY4sxR/ikA4EJGDJ22Q5+h+FrdOHu
AgtekG1zvh9Cg+uXkTOL3ded9DWpbF/qJ02OPlYmNodQccdkSFF3SdszT4lNcFj5F6ZFHpG96jZV
+hw4i9QKui+th/b+12GbzZLuo5Pws8Wn9XORVFc7cJuXAsktKOg0e8JrAx2UrYtD4CtF7VYNDFOm
TAx9OxzMOWHs+Zp5bocv5YNt2VFa9HlPft1vLMp6/duM4MR259CW5zQ5lF76ZDmDVw7I0zcCL5B7
a4QcWXmNl00i/dbLJXOxd/DTGBLfNMiTvDkR5MILlnaGTeTmdna1a5Ga2x0zdsmpaYWHyGJor+h/
gXGP7fknt4cFGjnksUgnw0kt1lPTExnUN+f2NMhqow1v7s+wkpMzfjOopmypvT3AXueZASy4BpjK
/Y6epnMv5OWR1cSmR1uwnz0tP/WDL2IWZqh/YG8agCZwnBx+8F/vDVpTmdx2SmJmDWtsgGC9O3Dm
XJMuBFe6RwV6cOtzXufW0JzM6eEpe9rPkhnwszmf/G4xjtDfx1Ep7Sqw/Ft71+GCN7PSjUO7i7jY
OT7MBKtFQoTRG6LiDTCJ3h2xdQF0Z3mJn4pvdNdWrRYvM/iGvSIiQ7ae1EFyeZdxkLbbItQHieeD
aa6WnwMpm3AVvaHnqVRRyDA42fZF4IWrUDCPMa1gZmxRTechzIkhjy0WXryzEQermdMaZbqNJkDB
FAjL/as7HsuKo6LppbXc2mjsm7VscMTZjhyc2JW+PP5cmWWBVGTwb04S+7IkrtrOjT2Fn28ZhMU8
JrnWBdvpcsvXrPhdJAXwhYlpfNAH9pyw0Af2ef7y1hrgQLIFrfrsbxhD/wkRYZP/oQvVztlVAfg5
MVcKG/EwnX5ds66CI16GWKI3gUf8+lTlcuvH7zYYTYLafy3mhI9C1N6TcAiIcIRo8AOKrCsoZrCY
r9rYkSl6BpBK9DDj4FcVten8i09PF+VUddIZlO+Jq43SZ7WhgnWCjxLlaImQBjRK5jw1x78rNHAG
lVn4quLJnGytZzn+qKYp+ujEHghagdPLREKat0k8ohQA+LMTkvcIC1VHF0/dogrreJ7QELLr5Ezf
3lUwMkhiu6iBqOxdPkDys0yadGdPaq2w4DM2bSm83nIyognvYcT+lqtNhe9V5tEPrR+TUqFFggEK
uUwp8tPVEz1NgZKpUkhQ63QPxWC/XpGC7IXtpkejl6jL6V/iSsZWsIUJma3NNaZyOBuCCxanbI45
cG3elI+T52a6aJA/9BtP0NkmPRtHvteMS/LJp3UGoSWsD9fbLJ/6wC2WmuYrFYwdHTPG+7QfREGC
WvUG2J+f+a510Ed2Pk9Mq1enytMAAnOCZt0+QfGhBydxKkndFJ3OmUu0QdhojBjUKn7Dn6xWX6Uo
7J15qapsE7mmYJsFcGNOJX6DdATsiej2X6ttuQ7DqwBmSf1aWbUaIVKqk4pykEV0w9hWLBG3++8h
eaOSwdSHtoYUntOHpBA2cNEx8djm+467YJ2jdCCiJ+GarhFOubvdzEkmZaYY7S4D/Sabl68q2WqW
ONfWN1h3bVCMtlhw2w/4W/CHgJ526snln/Y4bS8P7eZCLxXL1giv0F8qqZpCX8w28Ev8NRBi26Bo
TgYNwlaNs3pT+kfk4/eEAJBHl44ymSABTwvthFDgPCpuj7YqK/pBgffkalUis64DuQ9OBtqK4jEs
ZY53N5Isgd5OqKkGMl/tZQTpLJwsaGTwEu2QvA4yUXp93xI/DJ3O4pXXFdips72XSwQ7INhxxcFU
1czxnBAr6U+622xH1Kb45TFqnpun7IXnKgdMxRtQsvUYPh2sqYYp14adV3L3+pxQ6V9GSvdreUiE
xeMglpDrAxNBDmyBqqGtUcfD9jgPT8e9TvFFfna7r2oJeo8uInJ/RCLoIHZb1484ptypnvtE3jWv
/dxZQZCWJLeLscQhHpVFtHP+hS49oZjEJtU3dEUuFRSyw34gvcn6T72gNW5VvebIgu3REAkOf1cD
wRqljxZJe0pZorhMQkj0KyDm1Jhc8hSFd4llpgxOlKTeIo6aNjW6hxiG+zkkTv/nUOl6nX+OhAEA
rqkq0r+RJtgB+CoVtSZE2zG78V7aAKlQeDEFrYtmZiw3kK0PGugiDoN/1hh3vQcPfNqvxzfvGGYA
BvYuPuXSKRfTS8kSBnyy2uh3kjzIEF1i9Xzhtz2HcUBZGNYZCEMMmoh5mXP88mv0OExIRZbsnbJ+
lDrhzxMe0ya8qz10ScWdSvPYKPzQaswoSrKGjQf0BWLpR3erABC3y4ym5v0cAC/JLcym2V6rUp6w
KRCVez0BCUEYJD9tP7e84ChnTF9bwEIRg1mgoZqKKylewSaGybfNWT7YiHIBZb4razW7svnugpch
cIN3dTOH9fOvtiOnjU3rZ923EWtKoB9sNG385paKNUAc+QyMRGfOnK4prNxl9Rsjh1ZloM+uGdF1
hD7645ZyfM++Zus04hN7pG6vEO/QkPYmaQ+QOlTeB2Cj/tn22TGiTCpszxzzuMV46l3HBhawUh6U
PmTiXOlM5au5iRzwAQdtcnTzppQlf9omChrB5g+G1GEEldOCf3QKOLvGjf0pkFCZznGzY9fCYOKt
dsrTNnd3IpT//0vGs5JZwMSMKQKW/zJLBmrT7iTcZHb8xOUm8U2Xf2dDHoY68fQFamb+6jlRaiE6
nBFT6de9unJerw==
`pragma protect end_protected
