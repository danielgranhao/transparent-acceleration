-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
W1ds5rOActpKjU0MnPy0N59hLWHebwDewMjV01nAUxr29nuLQKfCx7lqSEUnXESY
0LReSCR1o5w/fH0fDv8DlAv3dy7VzL07/0A/vwMe44DP9CAvy1xkS+G/s10Uux7n
Xl4CX7TRSMVnb8RADWkKVhD0s9O+Ze3uBSlmTv1feNU+aqgGhtP+Ww==
--pragma protect end_key_block
--pragma protect digest_block
7B+VDBul4ZHzGcjngQiUHtgEO1s=
--pragma protect end_digest_block
--pragma protect data_block
RHK3YVDaypAhRZFaLpPwcqK3vKwnjWfAMt2rJUIBTVN9askYJeUcu9fb3h8m0mt7
SKau6NuLgo4BleFejKRS1aVDqjpBCxQ9paTBpv6zDNaTt0A89xtJRkuuo4cTPDNG
GH0Pm70vnST0LagDpLsE/TlI73eaW5ZwNtXhokInBKYchKpdenpShNzF2admLbn+
PBp+6MaqpOjXUkN2nlzVk5RZVGOpiMH3TVJ7YaY2SMlwMzTm7+OClfRYOpqTJ4Sz
O91wJvroLdxT9Czr4PUg3UcTWFTxRIDQXiO/h+poMJ0Umtn8ZDyE9HYaCo2S6oDY
ZpSk3Lu7X6lINUwq/ixOpsw6jMn2KhptEok8aoU/GMhiXTI77KIHlFmBpMMdq0eb
yzUfJf5e7YQ98t8bjHWHoUBN/3di0dRmql625UBkI+GWqs2bpRe/Q6LtaU08MeQa
BBJ4E9Dcz+MnvI7vxlrHvN1haRZajCEybQ6ruWklvBbhWiHnp2/XVBVE/5VG8vSB
cPkwrr9fxXtc68XyIoFhfIqeUY23EkThYqu4EoOdpb+s4By2ZqtvGMPBJlPAMAe3
7G6hEY0dbMZ4f6BFUCcsTsnOwyc9PyqUtEDW3f+sl359KPuylEE2z9IvkbbHQ+Pc
GE+ISdxKoAoYisS8DXIKmmsho/5e/blG+ae83Fm8S3B7wD3zfuKxpjqVjXhTMnoJ
U1UOYtp3o25H2Cbp+3oFd5EXnV/iSa3rYQI4VH4VCOQ8KdJPwq0LiF0gA/wojLSj
FqfwfxFtYQKAUpaY4ULYu7CKX8OR8u0yIffDpYNfQjtM+CsN8NdMftjPaHGU7txR
TJfPEMqmBQYESHl/+86BCLG7CfCeUactR3J73Gatzptm6MReTX+GzSWppjY6NjqD
2dx8+z1mJfs3oiHMfioqRDJRLcUEiHZlH7+GvYrnvtaAdZmMGck12haWeAL2qwDi
XB+38r3fKaTiPXuBSLOvjqE5UeXM59FJDSd3RqfE7yTMtiiDVdV0Yjy3ZhIPefTz
W+f677v09u5hR1Ay3i/QZN+/2kB46wd7iJzAa9SZvStapb2VBhCsl1re0IfBrJ/I
xmscVkmVye2anDHkAvQT5CH3TuT4M8iOwv03M95nZK/gVXuWC1CCN1roPUgS5+oK
oE5X5I/x/USjYrTPIJbAj/D41H7EeSdTRX5jbV4xycdfCMd68d6Y6yvB7AxFb2uq
/+3BE3LVSXF7qWR6G1ebRLDabydrufDTiH16OcijgX5S/xskm1lLzGlrvLE4Fihm
dgf9+DZYXf6mWKClQ0eb+EPtTun9+8XZzGQxgunwaSVJ3dmQXQV6fJ4/EatzAEbg
dJnBWc+KrC5Myim4y6rd2gSfXEKKVtyVG5gRthhRCV0yxDl1J/rtI/DLNenG25yD
CPxgHCOgf+oVui44+76AD+yx4k7UDg3y1JOyaiszO7LIsH9OSlHdJq5VhmBeGTK7
3nlXlTfE2aYdR/IvAHhhnnFt4uR+QQPuIPuUWbXSBGv26l56dm9PE9DWlahyPcVS
23pJF0VrZsW4+syKWMd0YOVBxb4YWClxj3/qhaNfn4K3FAfH15USgVrV61qW925q
0QfgpRhZdaAIOKZQJGXRckPJttX8uug1I92tOi2743unWuIef0nN1eSZACHL21mX
SuOGsd7bNmSTVY1Xv4iREgRthZx3zQfvRjFLkqvQwumpaZHqXZ6S+u8FgxFArcKE
CxDqXh0RjmrPzgRRLU3TC2ZxlIXiGYQ+a2Gmn/PBFMCXpLE5JhDV7G6oR87MeBRp
wMveWOrNqImmAgWefgE2uFb01f/Ys6CuBWlw5U4HNizJ38NP9L9t7q4YUupn6Zam
zyICkR++D0xHOHSlvZ2at/aMDInWc4UbKaq+csZPqyU0t22qQtQIVBhfl29IJc2m
qP1IUoxeqv677TjXdfq++yAL47Vw68Gh6pUuRIifLO9bt13kVr+6O/5shh2hxrP4
61hvP2l2GuSanJMaZrbHF55foSnqaXnn58WSJoUOWDwPSBM7VooblLVN7EQStBAV
1BNAKmjolhJ6OESwDZwfATN0DPOo5yl8i1IJZyBlmqNOT5tTQT+o0YIi/0ntj7Sp
neZVDHDduouIz5QLPxpnRXqk8qqFSHSAhPmpxeLsJSOm6KYRjTWIB4QRcfDJCH5i
0zzLkxslZ3tOOzUdzhRaeCUZkRCZUX3wozaLPkldjkyxqeQ93A2YxkrqFVzXEeCq
vR+1MkF7tGp4+egHcHwI8ZDBA7H6SqFZvQ9qpT/IuCIV91l1Sbl4wsliF/DlKSoY
IdmkuEQtIJOmK2IOl8F/F3cmm1CScZyJzUETZetFfsK0Fv/AziLo1vXsxNChXyK6
RDWtfdJW4OKDYcdu4EiOBNCU5BDJPPO3y2lqYsdnt/mSJMxf0X83uqZeqI9NL5sE
1yJ/qGK4th0AyLa9qik0j6IPE8+LF3OhoDW0Ot4b8FkO1T3Iqi048/LuiuzS33ry
o6uw2dpC2N1CqGJuHV+5s2PzUsYj6Vpsw/Nzc/KERjDS3xpmCCEKByJ1rjF7n06C
ZAEHeTKUQmraql01V7Zyj59eUToIxRXM43QyW8ufo4NtUa5tiH3IxtTbKAFssthE
gmL0Nq0LB44FJtk72PqHn7rmFrKRZWvhEn4jp6r/6k4xqdHSJ9ZW8JTbYH4gHRF2
kv8n80eWRbpoQYTvp9Vcx/pZGqplAl7mBK5Z0x5FH9DTspgq77D1oVTRffTm36WM
cYJOmDtLRZzWzJlT6bFNQ770Ec0DIvNmXNIbfX3iseP3ZNBc8C+55YbWIeEDBmh6
wS4Fa/lXlpCuHegMaULeTnPQfFbSbeEQSUD9YGAnwzvpt4x+3Hsk7yShW2AgB5pj
xylNBhmOkHtmU3oAjxdYcY3do7ivEVAUYLMQhoYm5qVkn0GsnoM6eo569a/UNlbJ
/T8rtjxSqg/rJEBERGrf0cix+TafvbIGbX7cmzpj+Mjn2B1oRsbf/oEk7Ah9JKm9
pI3DjbqWYoPtJmAbun90Z5UTcrYlixoMonk7djgZjCZSxaJy5xXK69r2dArZGJXr
KQKxuGfDz5rSiCQj2qpQCTZQmLP7W1xukZXG7KSM8m2pUo2WxQR0Wma2Fp3KQxTo
hRhnmPvwftSPYYidM7Kz+vY/0n6Bl0eUUdIxjj6nh2bS9oFgYEM3oVH44vAlpHuh
qRGKC1ZZ3SfvpKMvlUEcjYR0N/Tl1D0UTKR3x1+wO3QM+uhbSFSSM1u84SC+Jl0X
RxFAvdkFMyyHqY+kvVXDirojyu12cIadu2wxJVmIJliBo6kuwAU6JRTFLj9Kz06e
UQos3wfxvvbCXAuUsuZZnLVmJzTvPQNyaRRZoy38MJHAYG9QLBUvzCy/Abfb9Pp4
8RiancgfJpf14V5/QuGEXjUGjaX7RQaKa9qxOL/JnNPKy+XSQckqi49NOL1/xVNG
+4mj43vIOY9h8Dv7iq/eFGV0uIaNn8I1Kfqfp43bHdxXMhsRJDtaBvO3Z/2HYlpc
YQeGn4jEF6e/os+A4gG2KEkL7CLdfdY18brKGQiWxMYNmg4no4GI6gsp/iM6UHkF
KpbGwqJ/bk0iq71mOgvqxJokYAkmWdPwTY1jN94ZetKhqdP5cxxIObFTS+lSda1U
l23uLzrSxdG3QsEfDVxezHCPsEF5aalJbOwKhqO6T5fMPH900cNd+k3bgx4obLNX
tDBri49YdxFDm4j7XiSKL6q3oUDiCBrZtLIgSfRgwIetfPqutdRyYCrg89quP1J5
foXeZE0RRBOlTBxkDj0GROV+Xyh+WHk8LNcACCj6e6/Nu3eR4I1gFz7VFcgOETGc
/GCzwdOSn/op0L/ES4UMaaZ9RmItRfqwckZZJ2oZOtB5/YB1qsCrd3Oy70uhhHZm
4ySjstAwdnjjxXF5LC0Do4IkNvzzFxHBCZROBJnjbAHByVUhanVeCE/soeod+EC9
kDqFpog4qTaDoCvvlRSl/TK6YWFcLjp3orPOPQwykAETGEGC0+Vr1S8Z39kElLyT
GDN+KHRrMrjR6yR5khygIM5m/qvbfnK8TrkxfLixfF8cW8dFwk862jrIkYSOzcbk
jm6r+PooghkKV8USstCKaGTz2HjnEEwgaOAhZ30b1NK4bOgD0mrKxU5D19stiUMt
iTwfqCRfX2vl6/PgojyaFATZLtGJ+5czpXbXbTzx81RSiU3uW7rmBHBXZYZYGxok
hdQz+Y9APrer/ZtvYLKtJjJfm7mvtPeR5FHoeAHvKt9CncLtNuGv/V/hCuVq2RFD
m2chWciDEDj0GTvJLXSs9b6hEPpxEWeGOKPmEpNQ7xLOHNdVVHK8aKGvqG4+Zjy8
I7seceIhP3rdPvSdewyGXVlyG5ii7QWygophR6nxkdzTAa4josIJZZ2dUht8q+YE
WRiSNrpPoyL6zJfxN7gNFbk9nVZl7XK88UgqTdC3ubL24Duyk8IMM2NEKphRpjOy
8HyV7SEPseYFzTpFz049PaSfttSaOl6aXj/f8MAhByAqlhnC1Jn9xhis6oFTEXWh
Etb5cWF9RNVM7r9WtSiLK4uREm/N6iMZ78r17D09QI4J2oJT0pkuEY2fb+Tx6tRm
OBSw0F0+5pBuGQ3VPv1R+G7iWnWqz/SkN6T0D0ZKsn68271knafgpkfnwy0xn9xy
gvK3px1Y0Cyd9NXKrst5mNcB8gYGXEe0X2mBCTjat9Fz4yyMPFVPGjiFAiWjpoQM
RB38pS2Tx94QsM5bB+fEHHUR1jNntuGwh0I9Bqoc0l8wOGYs2L+hnORFWEYSsIjF
GZohgK++wXAOywdRO7LjEr+4qyyT+2WW3X2V2s5nWdhMuWxrd9OntBc7fl8GAOcq
dOk3/XOHFx+aBwIgQSXWO0xgDTQmvOz124TmLfRRuD6I09EkhGW+i/Rr6tOs1Gbj
bjnF7m4ZnQ2Sr2eTsnofDA+YI9EjGFoYU/t+wmtiJZJqGGbWgkDZfrpwIsRkDNYS
uGdUjWu3UCJO3uGGIKiyH+4Cxflkvl7B0MrvbRvrSV5NlEzIBAXz9X2MdmcKA9Cj
ifG6w+WBTqKJYisoQvQ6XVkhnqnkJv0fFPJf8fZkxvj29s5RncqUXlvG6vn2b5Ze
LILMFNXk0MbXB7l9xV8FWM2cHxwA0eunabxv/7xQaB77/CkeJ0QlHbmYDz2Z4Eqx
cL/B394+CWYHLsgDEtYABhnJCWeX+9v240Zd9to4fNevt/TScp/BjXvpkNZrp/XQ
eC3PzAJvfUBVoOXok2+u2U6CUKQnBDdkDYjhivajc/C8imRBbacuUMef1tufnmu9
/0pN4OEa7Kf8HhlN8KKsbBu3wmIxIFS9bmQ1zieFngGXkuzYTJAixJNH7VPkVWEZ
1Z2CDBNVYp6i3uBQAvl7R6ipMVQduI2BnhGPcNRA9caqX17mYwpL/5ObSFADR8ly
Ml+9AYEEBNajeQBVB/6p/mqk2v58BrnOAJpxqAuKfCfq3EG1C44dLNd3YGQflBCT
WA+NtoNP65bgtxIWVzRkPViKDz8zHSXY1DSa6EiP5uHOx6damzQzPYgBWPeW9zZo
gburKZV41YIlAZjC6wf+iK8zXPkenM+r7iPDj0jwDM0pmqbA2WWlUXeQYns61kX4
G4NFPKOzv4hBjpmMzNJrL9L2JmkKzAduCa8Nqy8nFL2hM6874cyFM88Gk+M3j3vg
q5GtJhaljmW1h8fD7BImvA7ZTlqAIKdPvqGk4n3JHV6kOXH0crBUqK07Bz6a1VXG
QTUUdEWrwYwf4UvtKKSfn8h8KLKUnRnvbcr8Fp7JTsiZ/+TNzlREAEHT/KfFlXK7
IRw7T83zNTaUi2ozaczcN7tzdedwVZmgyG6m7WOLw4lQ5VrQsLaOFLOxug/LavN3
Qp9FWBti7CiRVebgwAoczsc3N1SzL5ak8KuxQ7QCSIdzxxlPF0HBPqsWnzi7lTZ3
1yeu+QUDqMnZ3hIP3jgvn/3eJ+uMflWPnFvtezF4JtW8f/2s+A2jx5DXc2l4+BxD
j7WYiADP/Aq3fF1jyllJs82MY53BG9vzs6ecTQUz5wGXEqYmlw+2Zr+1RMn0V+vV
szb6bDcQA6W0ZwbUM6rB/4EjsVsAqZyJD8bm5BMhUcPClqAW6/W0pna+F3MFXRPr
QhLrUYFueIzZ1vScfwTc6CQHEuvcX4rcqaVqJC5dU+X+iM1iGXir2UobWnjT6NTe
CF4U1Lc3QRd43OEOvBWk8A6LhWEhHJ+YKQr3gzNBfJNhWKSD2bOpwoEJQRZ/YV9Q
DSQzYDrZSnRqtK9pDmR3imFVIX5kA0e+QKVANrjl6tLL5c8nOpJwxJbWzbSw8kh9
5UJ+RoU5g3cTpVYt8G2x3lcyr0rnAPjp4z1Jbs+cCg8jTjh/C4Sdfv53T1W6Art5
kRusqM6Mmrj5Quac/WIuknpiVi81dgQTRNVyn6YPjKqd9f2ve5gKT+/KVEfXR04l
HTuswjpH+wUZmZmPvh+yq10daYI8rF1yizsukRumuXzkfOlqcmDrY4t3fxdaMstr
1F0BtA0jColG+VXIkbi7JABnFeCrKux0pskbeHKp4QaxogoZdNfCWyqHiUjgh+Zw
HJxqXGscy4anuyZfMsK806/i+aPCQXyUVdjs+PobOd6TZFBtFhno8xfzltOraN2D
xg6BE5bGPNoKxVTuDJmbHPP6Nw3J6jdDeZUxgvRu6dTlC81aLP7j7pIliMlI4nh8
PFnUJ7PUJlVgvKeFo0jc5EcX0DfwBH4U2zhRV9ffBe2O9z+yhGckTfvpNqGnSHmT
/TQ+dSHZ1RTmDPZKLDzFPyvDI8wUzrK1h2Z1Y54tteY+5I0khTb1Ff8cCPXWDVHA
BNHACa7EXJzGxgYx5Tnjey3zTYR6wOwb0JxBVgG0cqUpOXGiVdj5sVgFT6DpNFvr
1uuQymKG121lhrgXPibSzSmcq6cmfJZbBkGyo/oTU4M0Wlxz/8lOrbY5Ycmsbf/+
Da58ZfG5V4oa6TDyb/3O6p7/+QuwTgv4nvPbn/SFkzRZEo69UecGjp+6XcAb1vEK
VP2rXYXQYrKVvrYBK15O2wrAYcG1UEh3hA4XJYpLXO+1D4JdabEWOWG9HAPKqLIS
+KXu+m2n8WLq27F3qQGn5ZL8GUjATMYKA6J4uS0skZhM6qRSZEnYaHNNLtVBQIFe
Gu223ffxikEPr0ZV0AO22BYnBUsMw8aK+jD8IMIhW/hHa9/60DfJsE6p94ycQKCY
6Y9eNO8HKfuX8FgXXOq/fvUoQTAJNxnkO1/qvnVma1cVYTqAB7QA/CExZ5N05Nds
jVpCycTlT8HYairiQetwNEGiTosnawPmKgwmdFzL0FLBvHIMcKMkBP41xM/t2zyG
srfB69SsydjNIbLXumDtpIES/H56CRsZ00gyGT9cz+9mwV2eWnOtonUU3v2sJw0r
n/bQUqdyN3PhZH98u8joM2xTYop7dHgDLojDceBxP5kllkKIMwnoV9+rH6YF7XLK
96txcQiv8nxmV2BhClFkY7LWAXDQGxsw1n70gYVlinNEolgcQmMVermGIlRefs3V
8vyguOUYAcCHXJUVEF70mssgHWsmGJs5Jrf1OvSLHYbjsVFJDaGZobAum2OzNTxM
8y1a8FQEhzkbqFuPx1OdSbMqvkM+viwU8eFChCCwERkzt8HWQp7BoeC5yva7MFcc
AqwrbfX34IcKHu7Q9yjBwU2THQow6/7Wdu1D563tP5dS/HI/5sgUKJrQjBEsUJKN
/CU+mYce3VMJyvTltu3Qhlc7890f6zrfhNjtBU0hnYFF30qHisIgcVYvzuI6fWrD
ljY/wxxq9cgtTxWEZv0DJMzcPirtU9us+r7gD0+/mYYPMBwF3uxWBFKQB1WE39X3
U/soW7GfhlnaqeX/ADTWZO8wqQxUTmxGN3Mg4iRNfKvJ9b2W/GSLI3qJuS+QBdcO
44Fe3floCvoO2dTdrENnqwGhaSOzuAD1sw832Q6btIyGpvjVq0aQmRAlc+Exba23
XTrSSdhWdbrE+3sYi2LU6P/uNoJURj0B7EDFf1f1uYMNz7sZBIkAdAetAjZRIQRr
zIAEtGVewXoV3XKG7W9bGNvREuMttMW1suqBgXdSe/D0Sp/AaICAzNZKUjXXwKTU
gMt0sflJdoJAS+Jm6uLgbMjPepGBa1EIcIBgdSOoKPSKYruIK/K/GLBEHmwCs94v
U6TRzJ9qi0aGV+Qco4H30nnrvlvwIU1/NpyQMQdHXBCqjofnF9y9A+Sdj0ukepcG
XjGRPx9HrFNk/oUTzC/16u2IT96RxGxlh0uJUN4zpmVRshNzNi9FiXasO/GTJcvZ
/pAFyND66M3/Hj9NJCN+4Pn5l7rTdrSRuSItfoVOeEwAYHOy0KToesQCwAvYADRh
LYKz4trvDZg0XXJ0ImS1K4GH5+8KJCFb7+hkdYkl8DkCMSzJH/Q0n2SlmylezqRp
EauzRxailWmmdR8Wqq7iSJrL0jtPz/cuxVfWdADd0k82LD8O57KEaSttq+pEeB0C
NHFj5jTmOHWyX+gFbne7jU0/bMmQWDswaDBFyK0J6m8K/weSAhY6b2O+dDWL7xKk
X16T0vaSJmMM1cVsiriOJ4CJAkjeJwCjUzNEtYVGf88lSnPhWVayV6mN7sdvZZ6U
NDWvY1XRTcY1UrYsBRwSEzbP3q3bg03hlnAh9HRzZIkAbVHG702lg5ccPEUqGwzO
SDPU78Xy9Mtik8GJHM/7BYaosYY7SFJjQEznNzL7HvfRSkGZY5mZ8mXoPenHg6Qb
yzUim4CXREViTbJIYtBBLnOM+GTU/ENsqwIRkr/NVR9MDJC1x9YR0b5/hE9CGR+e
TH3wsdwDfURws+i4Arc9AKXReoILJwue480NBgbT8B8QEUrC+vhqp13pmQec1w7N
+tXfPQry7tIwX0ZNC1cON38fVjjhRzzFAyJgJY4ybZOtCHVr97Oxo5SlbKgvNK/B
lvwiE/zfP/iFqCUg9QT3z3G3O4SbtCqvPMIsT9swwEVv2o492CZs/Vj7ZcvofQ91
76mbqNVVFEVqfK7+qkSK0bOQyNg82yIvxkiEqH8OlfayUhh7yCrTjPG05BvIzvPg
4ZbYa+pXWcdAmvGAZ/hW4MOKPsRAohRZbSHM8rveVUfkmXh8WR6M/xiApJhlav8K
C6UYKgLc3G2lfn7+Lkzu3zcVar9Vk97gM3HyKQHwXUr3C1ZMlox+gnamlFMGc/Iy
DsqFbdSo3ZakdMc7QxuinsVcIXaMTT8eMG0N5AcbbGu+dgIntNUw9+036HXbTg8u
ykUskZ+ZLarAnibu4mZ0CHfr4dLYgMMuS04eC8bu18kc0xs9Kr/YaPU/jkZpqwQ8
mpwb5vwWroKnlPf5gFYehys5JFPD8TVfMbxGog+Sxf1eNaXBLvim0ja5KgLo6X9n
d/p8VqH4KHckQnvu/uBDse5ZSslkkCfKUKYCTBxGtGirL/TpGaKV/EPfjXN2/6hb
zGkNqqfmKfOEHl3BQu3Lmo5PBs/CRUt7rf+aEok2A0fyCcmu9QH8Ce9MKbYvdrjP
MAy7vDT41pXViQ2rWNdOc+uyroeQ2/sCnQJHJ1Uhon9hwnGQYkVq3Fn1Va+KdwXr
O0ZYmdIpSm8txnanfVKUcwcKkde8vb3S1l5N0uSQAJWTjkTICN5JQP70Q3a61ovQ
dy0K9DT2LyrhsXvZRFb6PcoxeD8P2k83JLdxXsS3Q5MeWHL74IlSbauAvvee2RWd
7IBz5mKe5XZBJ2UZmYJot7Z2uBUcU9FljR18Ahqfmj4y0B1kpKshHr4S6t6xajj1
WYyxpaTfNmXuTs7i/lCUnmxxCUAvnjtcBx5tfT+yKmtzywzbnhoVp/W/APqk7Pcv
mpU/ywmZkFpmTfxWxWFupzIU21TBhL9COZ6wos0Fi1DOZvpizbdu/h/PXX6hLnXM
knXuU+qcMFa5TtLb3qqWFD8b3ogeCvkTUv7edwiMV7EcED+r0JoOJcPArhBN7zC2
Cx3fAk/hHgMizsC3W8S+A4N5DT3cxTA0rpAbnd6ClM15/itTR6po3JDW9qvIDbvX
kNpgIYiOJQX/PtvsX4nIRGtZgUlf7jU1AqeYGo2kMVSo1qny1rX/oNyeJnMR0Tcb
LnCv56FMyUHrv+olymt+ugA2ozROwP4eGiCvMvAphJ7SE6eIyNxa0OXmVqZ1cIcI
fMfJV/XQmvF6WK3CGq9GsMnhL1+cJG3PWBqsyClOW0S41X3Nf6luMIxS1BRNuZ9S
7ETZ1zAY6gUnZhO+WJ6jv3nRJpcTcgEJrZwv+mxwUizw8SAyZ4e3vuQcbn8P0vsU
xSUeiS4U0+pDY72wlsaCLmfk7eFcegLHitkpY7NkRxuzBEIR8jRXkFju8rjZEk7V
6FFaogajOzpu3bOK6kwmDeO1TewUypaJoEmnN1q6Vez5xraRtoeu82a9EIz5ftSa
wD7QSxWpaPzFf9oEyLs146S7xQ38nIJWboBH3wk2N9sC+/RrrsrmnS43EcY/WaGM
coWRTDuUqI/NhF8fcZpa/griuZkCfFC9U8ZWGsrTjTkzUSeZR0gpvH9bwRM8TbMe
+dVsjY7/EwaMMIVvj/AfcbEQm0JPUBllSGZyl99wfuANfao+hNvUUBBCx+odcY7d
eoLHtby7XEYpub2cImJ+aJGrcr4HRjqgqSHdGr2B4K4Uxyqzo5l660mvC3lhmA0p
dw9HS/2scD5u4old6O5in7iaYRUrP99wQp1BJzQpIEkP+z7MOhNYyzObk6WIDQ0Y
uz3QcQXDKVOOaMYbzbFLBRRUaxcEIv+rk+zYxdNvoykyxP227p6Yg2B/U5WPK4ou
lulxfcwda5Y6BNGINcBRBft1ihDESeVXwKC0lrvs3nMzeHaBqnHfucJSqCbUO8l4
lUIyEgQ9rqfIcKg603++W5vB0sxATi2ipGMzKEWSmN4bXNxAHx6wes7pry94l5OJ
Y4fxCZT2HwuzA4e+XJdB1jCVVgNmlq8Hub7IP/ciMLEBQaBxMhsE8pharwxOLrIC
GnwGSX85xnuKUXT6qbOT/Cwpv4RII/07ZvqgbD7xqm4sXosHCPxrseIfGGvkzZH+
DJIBt5Plae80YdyWmLinVlYj7pVSJrUg7Bq0r3+NMxX/rKIpWPLr09FmFs5z7iHS
51TR3FDa0cYV9RaY84uHnwHH7wBsWl43G+3rKlE+UL0q0xwhdGj+IPM2o/2iwlJP
NZITnxWfC0mgAeftOPK/2epfZgHKK6WJFBjtTJ0FmXSxJs8ZteOTRBP+5XTDhxh7
rSvtN14jkRGDQcIzZiGOBneqloFcqE2v9WEejkY/p4r2IhHo+fJDgPHV3wkOtdCx
gEdQpkDIl+GfOqpFFNMh8ACJ+AbUfyOP6knfs6mx/DUQSL/HJ9SVnW3cvGbplUs7
OosGiRDdJKJj4R1tT4E+JpNuq04NkEy4mM6MkM8SKS32o1Jw+Zemdo7kLbz7drme
25ryGmooJfhaNgbaLPEu090CoyabTwAimDbMus1/+aFs9YbDJQ5dP1vP1H1fh/Ph
GmLFJJnlWCGw0zwJUbYqgcAojAX8hqfSMhaakm4cEACeWWwhhipVEk4wseuTkGWj
CkKh5OzL9LLmCXprHkwIQVYIybMFuv6PywQCaxOp2JZmCGWowmp8GVe2trdW9AoA
bEyG87wvZg0W60e48keyK8gSdwV2CHp0j3w/unTnit9+ymfZSHhMCucAjs4H3NP+
0ByKOtD58iAocjdkU6mYMkm3TJg236HGrc6K5vhcG5NmJYZmUWHSxPAXfSfDdatH
bFfIl7dCEYQnYtBhlO8RN2v1KdEytqTbVFyl2OpXDX6/ayVHdiDEURRfdd4zhZ3Q
E6waDmrfYnfQNppm1W1ETkboShaxDpV/Dh+TclPRJOazm3xhlLgI2r7OIz4yElyx
//3RYK4lazGw84yQAGT0QiNBrn4qmApanxtp7aQDm7Yj9VrPJgvWT762chPNfJSB
94bioH+LEA+hpwSaznRV7xiIdr1QlkNKpQ1qK5hZ4HvzqLv5Ng6mder00mJMaUWK
PV3PR8x73MPUmwcB4Osaxhv9kt45mF4/S3VLUcUMiEG1UjczdR+2iuMcAl3HTJ0z
Ox6cR+94rsyq4Ibu2aylKTuqV0PT8EUGmflb7ZZXPg/gkI3fmgZemxqZ8whBG3dS
wYBMaBw3e2J3xhYfRIv9QzBXMfZasZvehy700SHHUyhn1SHFqxMhdKboJdGYFzew
hSAYVafoZVPopxHd//mByX7tWK/PEZOx/BUQw0dYMcAquy84qwg1f6a9EF8mqKeS
ggZ01XlxSblHrSc888EbCDzFGRTCnzKBHsKb05VMuKFYiyLHE4Mu7MUmnnY+wb3g
qeFiWMCGlwuhD5UKd2ES5clzwTUcktC+bTmHxxabXj61y2yRBnQ0VWEmPsVH/XiY
iaJ+0FF4NQ3Rme4VOr+xPpAz63desQPHa6jna/q2o3hC//aCuE5RCiwOsOO/c3qL
YjM5YB6K0+9GBhFSRxM2FhviMMWm8G9OQyKeTOxlPtiXo8BLIua1bLVIlQDeZ1Z5
wCF9jDuOZmq/36m0YSg+PUgjQhbP+IwXjO4mxhqtEpTgBvLp20xETtiaNOtcn61u
PVkRqAxO/sqHowTtQtyl0JQbyHza3ilUR7FVOJscJOtq7NfxMciQOrN/P4zaxTBT
CKoSLhOkGtsOPVyzuBUFWEtSPvNLYkbQyfSo4ZMQTagmPHS5/G6gNHZDyIabUZqi
EAPVu9uU1fcNQvTfBBRl/MyLGLNxlhrRQpW2GGb5D4mwfcdsyPov2mG9FyxwrztE
L2eA8urXmdoss83h7Ltmsrq6bcU3f1RmCA5HXfsqX2tVlDgDwZLm1LQ7EJsSSjjj
c73hAoxLMHxrCDy4sjsh+Q5R08oDTfyxdLiV4RM80WgpTYstaMtjRiRpryNTYNmE
c/k9ZRElgaVPveeuydI90b19hB53+MHcD9n7fsZL2xxB9NvXKKJif3pGLAF++puO
UXMB2yBUGjzRfXEt0a9A/f+cVPHjYpM3BjozEMNZ8dWdofzqwrLWTzA7CcYOZ7B4
OmjQBGHOPKIoPnd6CHE9WXK2pAcO+DL+JgDn0/HP6h3cOWp8+13lCUEkL/MbNGaQ
Kg5Dz+yEWAy31Im0ld81OdJPYlp4ICr78ch7S01rI5471YZB9UU+nhjjRgE244Ia
dt+OvGjuysePvRv2kMtArHxVT0Aueukr59aXRuIcs5N4k/xxqguWbzy4mPViV265
YmcC3u8c97A57VwRZITHQWzhrg9E/JbEa0O3rL0STVzngQcCYxRjg/QaIlVLprHP
JWIy9/sp+mqSKwtQiZ3x/knweEZXKU0vBTVe5jH8TS53j9cpEyNj6VvTwzA/gEv4
2WdYwA/PFGpQ/XGpE9kYA34ehpJIUXIMaIOa93/oNM1A4DbBsZygBcz/ZSeLtrwO
1xlGgsyDOf3qqk7y7+See/NbIqFwd/UaFI2piSnCVM0st8QUPPJbzFYXBzUo86GA
9BAlnaYpFFI2Xeci3Gvecli+TaRZDAJp56NZA7QhP9adrOvZ6F3Z8CUkVz8pxrLg
UYzHK0Eos5QUp3UZTU/nTsmP5JhhgvjyVk49u3OvjQvC/dsld+wXqv+LS4/Za9gm
ph8INaMfjg+R3iyowHR/GX96KDhTcXal6403BbjeXVlonhR8k0Hb2RfqB2jQUzOX
R4puwYIJ5C/Q9n49EsXP0BFD2033LHAcjiaIZ3VgGsZEKVARocGpMsrw5W6O3IDn
3ZVC8/GopZUogSOOYBIxFsYIxP47B/b3ffqAiwrsWU126mQh6DyNTmFnWtJOPfxv
yh7SbSrJJf9RYkI3GkuQUxoJjyoCoWyBq7Wv1lx0ADRB3hHPC0hXs+J9MBkMBilJ
Wrlk8Rk5dgeoG6ebf8KfMGELIMzK5kfZEPsByROORPsQn8lNx5BHwJPF5j1uOw+X
nzPRNytB34e9I4/EVgbz1XjfSC/pCvgoUw5jZs+MhQBKIaBuC4Fn6i7tHjDfbs51
h5UTmUHkAqAK+8HCjE2WqVbvZthHAqITiRK7OabnGFPTf7zzlC4/hQVOSAGe73IT
h65ubCYxXqUPmEIwEqv+f3e2crJfj5L5YB76X17shdGsf/ArayMPVRAtHG6FvAdk
5nFFjJVt1y37dxC7LNNS/htQSUpLUv1fPt14OMS48kocNZxbPaSr8WxGbWtFRez7
/q49QnRg/V2TBls6J3xjY9OpCC/7qbSM85MYlKRHC2hU8fG4wU5rmE5NUZJNhl+r
iNKyTbRbr/YlteTRrnNunLogLBo9ITe7dP0KLsuCDAUeHQhWoVm0E+udK+fOjFW6
ZRUM10b6VSRO13faMRHXx10ZpRPRYmKX+c/Ty4EgFAjnEFq/JROX7p27IVoh+D69
kxLNDuRj5YoN5LSyQFFjB52X7xbqJ9ltIp1JrjlpwK6y39/WSKLOO1HniX78j54g
AdDpiPqRcMpNvvA/pGf5ur+W6OaydS+ZsHX8NBCF5nszF1k0O4zObRHbj7V+36s6
lvUuclwWM+vfIcu+0Rh239BpKDScGoI7WXELp6uF8S4NcyFR5xVTzZ5XLwD1PHIv
qG/eg8oqzB10hQqoC3/WLez42hWUhcnIPXXGOvBz0u8lUa3xZGd1BEgD6MjtDZdO
C/u9WweGRJ8gFZ0Woile6VcA5pr/WZRWbGe0A+ZGfsM2yszhQTm6+OEcYWNGxt+t
KE8pSz2Y8lZeinDDA8XAS0xfRKtz1vfQ5FWmiZcs5OWQJMU32WSaLhX/liyCQ/r+
dXxiU0B8GZGJU0nsIG3NnQ7rt6JVrpXJxA4vlrIeMQYfzwFcJ3DDyCgwrI1/F3B3
VQRHOx/MdZjaSHIfAUKbxgLmhZ/Z7378qPLbcJ/XjZ+zgEgRv3EI2OJXOFvxOtr9
YNDF0wHWZPPzTZ8ibTFxf1V+5hqYoEazo+Om8QPwJAGqKLj1BWgpZp2UKWhWhv28
1hetfWxl6GHhx+YPN+zPZqGQjLlNkKQ4yeu2tbuFErohUCjlVA2FV6b8nHvOBc27
cKd4gJwenUr+0EIMjXNoCNtsGPYXFUQ6peBoPkDJ45oNggvnXveMYrEsk1y25NeG
kemT0b5rqMNkG+v5zP5J557VJ+pRTdjxAMOCdkmoILaorClIUYq0Jxo9sPIUerTe
3qJmRKfYnqhSlm7aLAzwhCInmRjK7mA+swnV+7Y89E6NaiRjg+g1+jUIAT0uY1rS
SznSTHOOFt2uKRyP5Y+sllqD29eeil1L3B01lQFCYbTshkesIuOSQTsToWeJFdOn
RsjzWrHYjiff6ixlBG5chXHK+kf54JHqe2QBJw5kYBgxq6DeKeugiDfRhaV03iV+
ZNc0JQHjcYAwKURfz8Y3/9FJ2jxCUqpSfgM9XFD2b1bmT55IpCmUKgm5WPxics7x
mTr6hhUY7U7/ztLdjGM6jcfId3qlFWnejm5CcgdBptzb7xxuu+zduSCzD5U6PvvY
iDaGu8JZg6wvF8K/ETrfZ6eOx5O9iXuJmpsSATD6+fRqxpzzI2Gs5k5ymVwa4Hhi
A4toYxgytdD28eXpXs+OFZhB20L9dNEUyscLuOqORdGWsPpf53NR37LwySl3lnTE
/D3RRwj8bCIFtkLR1FiQz6ZDkaZ+97XIrIp4eSNTmAh/ldjhQbux7BiKZWTyk4bA
xjvWwVeHl/c0nuVHNqRnhuq8td92OmClaAHLqioCr40hgQvsJIBJxW972qgMl1fP
BAPKnc9Uk8YzJThPHOWweQZdsfEb7GaSm37YdqR8QuCxWiAooN9naYTb3ToNh5+x
i2MZ8IlN5hUnnW0huk+vJHssyUYTaBksZVp2jRpmHFnjgtEChl1iFpllIHMxJLwJ
/olLOWq09sOQdWsnlHqnfXZt2Cs95FocCMFq4NZKA2Vu0tpStSYAg94yu6VBh3Ot
yZvTbs1DmKIFTpEiiTa7L+BQlbdPY5P2QWdo7DG/bhDMAR+ZaoTTn1qFHqEyE2G0
vS+X2fKkunW+/cMQwpyO7ykG03GyN1ZChQPCoLU1kuXHTYYnXw3NjioW5tc3fdjH
GlmcoqbkxjzZanUVn9kwAVovcn7pEwWkKIitsw1Bo7XUo1tVaFwHLg4xc7ErA4U9
6WJf5f7/yj7R1OPGULTUQMqUWDBQhx5SsEkc2PMp4nov6f2voBAeVZNGTpebhQd1
aYSbe9lwJyJ+2cizNcSzKaA7vQyNibD62hOJ8HHinOm7rqpPUPm4Ko9PGMejgjNi
CmoMy6q4bcWZb3nT2I6ACA3ROYaouf2XL8+PO/PccKEgKLfOynpUhJxAppHQrYaf
MPgg8E6x+dP58TlN3dzhCIErXTGPdnOK0bfN20nKvQER2ns654H/Mtrp3Rp2LHOx
4YAVRZMset0kJkgwu/iOjvwEpo72nHfVHgFW/S+vkZz6aMY5UXXajuBLMZlVUrhp
aIXWjo80GnOAgxjAVC+PCDTGf1ZBoqAvnyTrlQcPrsJHvmPsx9jnbFwxr1PiMVIY
vSjh/xB3/pUKofAF6kb4xKkZK3tWjyei1pCtw+SstDsQdrH9DJtlZ0lSt7f8MFXW
9Ser86O0HQjYJH3bEaohqGixS/R8paom2auRgr73XOFTKa+uzKNR74ZEHfwvfwPL
CuFdZhRGppvZBxLaxTuEHWrYHdFmEmm7j3dm19RCv2/fyRPrzC8e8Wl/+OEJdZS4
k5u/mqZnKZA1EaWkU7XXk6MRDj1lRRoTPvIOE84FP2NlWPQJ+tsvai89fX1tti1P
Q7PJV6ujmWw3QhI9mK910oDOeRRBTLafirCzek+7RKOEfiJQggv72fI1oAAAZ1Du
xDn2ElRd3ATmHYexvumCNgRL9gADP88bvPcwFVVG3Bc++bsBF1sWQNj+OQLDuyEt
ee1igOKLynUrJcnAjihvh1A7gRwrcXSJ3olwkxicFcgBIH2nFgIDxcLEPL2lA6u/
ZSIeakdkndC9BGi7lq5KB6cZ4b6H7I30xsvNct8pDi0xjn1DVVtbkJwwXxnZOpqf
CtZNvKqD5Q3u3jJ7LTIpU85jgDTDYQI3qq8KtIAvy6i1kx24KudRYjg8MsuCEabR
ejzY7BzIk5tKQAd3S+AFHMaQFD+WHf0NASph5eba7pL9GRPpUpLxuklrgtbb63Mm
9CbZJcK3OH0GSyUBcAhO1fDpg9dCSia/u0rYdpy3VxRtMzworyeEjrlAwh2ZLN7f
53rYKava7i43ZX/404VG2/A/XzaAPr4zmWW2LVz5jq4g9K/G8gSntoJPYwsTNHsi
e6Qdu7mvvcDZcg7c7o9++3gg2SZ/WjTktFWwCPErIY9H51OKuU7w3kPz1YuzDiFs
BL+s+wd7iBdR47U49m1gVX2m2uFrTI+i1a3Z22tc6gbde/xzXeCXg0IwOCVpFrez
TLwouexfrO2EPksmvZM1pqxKS3OVJN86QZ7tKnU2sqBSTthBWJiOVZFfOkG94fRm
+yBIXShEPG/B0eZffbEgsH2q6caPxrQJP4YrpUflLs8Lg+9Xs7IPFJf1KYAZWDAP
fb7rIlTSOGdNlAuf/rOk67wJ/2waKlmjfUgDgdMfPJLvaX6Ry3H0zSJOYm+J8VTN
8Cm7l8bCjv72ZTr0xzIjb7s8jHjq20QrTOoSSP2WDUgKoz130apEet/+L6ZhfAus
SOBW7EiTyloxVENP/yl8jssNqHcmQ00bOBDOW8KqGsmNAfBTjEhjkGclC6ScICBV
wPHKDydkAdyjAbTPkozw6ao0y5Ys2q0CRS75ZLTtUyjQKr8WPOR1/FasG5IKNT3N
ws3JTgUiNgvSXNNTZcL2I5sUBIGRPJdPe4VodnGt3xbXDFoDNWv3GDxY4SEo6yK7
V3qZuk+GUYYfnSh7x+PGhB+wRNNrzv7T1FX76ZtRsKMLd8iM+tfyPsXT4pXXfC2i
Y6Q6Ygz9JKHGPLMuvpcioa4PdRIM1LHYZhwJENliBzIbmCE74orItRSDu3M1OA3E
L+5bBKZFNbxS5HCpbOta9yWnvTZdpJveRiJt3xPZQ2AQKwZbTjjMG6qcPPgIhZDX
+J5t/9arNo28bQvUujT656AxvkKQL8021jpQzSSjt+DV0WypXvOCrWmQjA6Y/mqm
KBrYcNdiKVkhs0vIFwMfAZVugbPPqZlI3yAEAbULOXKSce7+aYDpbAfTTgJg3BBW
K0QVl7lltdUufGdkemNuRRkPjTivnteh1Zoecl3z2Zr5mYWbCbeMbSQtHSQiXA8S
dExe6OQGaq0cjDjCgE6szHsjXhQuT7AuFx+itRmqpAhBzlnBuzVCMar7FsZbTpQW
gkqzSHBQo4f+L8Yad7QyRX5IblRjYmEx4IdXXOnIZC+BuhvsbPKkGJijGefVKk9D
iX4t8Ehdwz6Givzdfc4hPgqZAxBnHNIJM4We04YBbFwHqr2Ngw5LU6yTZ/QAZThX
0p8sqJLke5Po2Qi/meP284rpHzIFCGf28kByeS1+mIOHIYUZ0EFadvtCv2pCkbfa
NGHb1M8unJYrFLtl+PsJwuFE7F7Ysr1wdsdbuDoLjvyNsj85iI0s6qIf1XQpC6Lr
8BHN6jGQn/aYSqkgo+z5jOM6chjABqp4aOzlAVP0r2N3HQ8MSOBDbyTiQFRmpHjU
RUuqNMxlYWWETYghyhESTD6GVUlKMyNGQ5JFS32hdWuzFQtIl0XMz0c1mb4aXrO/
gQkF4Q67k28/A+fZHCMbmKS5U1tgKS4LjG337RiviqThSSECJu/TgXGYJfwd63Cy
ctiH4AeuQSpnvmBkD6POUR4JlkpLPdLoIJQ5BjtLAe1OR2FP5PimCDUKXIVMkUzk
4nLAbd1rgWCwumvHdqfUZpOCr48rDZjlb28uDaV95tVmxn0kpxK6sqzfuyUjucUO
KDkYnU7ja6d6tJo5614iO3K0+zrdsHkZqTarYwecZRGUYgK9zj20sdY4l9OFiZ1L
Pd7i5mk1YyhJ88yV7TyoiMjLstcBUTdbrfgziUo5SBtuzz/m0BQfQO5VdfpgLj8O
mqydmLnIx9pj0yna0Nata2CuzmqyoyTYIiNQkgUvEuemHOd2e8d9mqqsUthowMUW
Cs4yP3LothqT6YAXC+jylBFyUQSeh2dgirP2iaRquCYsMKt8TUCfmbS/jGpz5hj6
E/DdGz47f7T88UtAtTogdpoL5NIvRqZx1HICFEptZvMnZYK/twH2bxjXP3EyMwLA
CdgV1uMqIJD9hxDXa5E7u4q1NQcJmrqGDCorera+KGN1hgzyRGm3DVZoAYlGF53t
fkaO/RkNqJW/ZMuBCS+qVNSWC4BRnNz5nclNT8nINS4cn5al5cK3mGN0+ntS3XYm
/nctQR1xyWvYsrZWCJbgzr/HfTj+zXY09A8csQys1AegxBYao++0zWIPpn1C6GYj
0ikWhSBfarpk9jKd+YcSj0tEEy7UTxhDtKP0xZ8PbUrfvmk58jq5Qe4xQcYTtzQs
yDJ7K0VCEJL+3ABc8qG9eahfylU2bfTWtZ4NL3wNmeXdyIl430JuScBinaJL8fT8
Ws8IfuTeF7jutaUPiHv5BnrZsvZZw1voac31wRYli6cXysT5Ng4lw2UFWAM4ptK1
RRYcuJDeaA/xg2YnU2P7X/GiTjebdo+NkigqcL2C5DhP7Dng+TUPkQBU0r8HqjtA
hV6+hpyIELnHbl/uJ9n9+mh/Yrd3673wHzzlCFsdreBJ/wKjj0hQtuQ91eC0BHRv
ZQAbfDP89HPq18LKpxymVlElvLUBPYzHXjS1BWPCBY5VzXrXrVxyz7gd4QrrPN/9
XgPio+eL6JhBYy9Vji2Gg3WFrhMl81YiYQ7llFnEqNc/ds9yfQHdbXP9aOT8dVRb
nRQlRfRls9jd85PM8eYE6T/hZ7d0UHLty7Z56SeNnh2HmOiyoN5n20ZupX+CXZlQ
1ftsXqXJR6kMLfHEcAELkPwSr93sJaTHsR6GumYDcS1Qw15IpCwTZn1cgsyzar88
JMUfIagOPQclaJJnzSA/iz/Of4BGLZD1hC0xbZ/mj5Ef1k5kOHOMSvs+g+sbx+ZU
oFi/BHwhZHYNb5RMQiPwv7xA+AMhjCAjuzamCczbkVtarIlDYVqBDYI66lOZ6Jhp
d7zivWU0ScTcsqwUFfNezELQ6yMc//SKdY+oC0mUQ2BoJJ42axh7CjS6aPm7vkc6
Nvx/heCOVPclDj8NXALDO3C84CerGYljI7odnN29jDDumlxskt7dlLGbQbEpFYHI
uf6b5JnLiN5YuO7o5Du3qzTz8eGlqFOgqhYld8i4WnuEk+/wJAow0eg5/d1ja7Xv
u9RgofBv9XpKViKZycfGkME1HL0FHdtuY4voDSfKmgY+90M/x9wMehJ6O7LTc4Bx
OHD4oKO+zNt/yBbEri3rrPc4NO5hScUmxnD5INZre4HinRWzV03YIuof0sWUDMwJ
GtHuGdOrR36/IvoenZ4jNnChjukLma+kGVX8MBowz2yTXbipbYwwjHPJ0jJd5G90
dNYkRrHGc5vvCdzH/SsKkmasE2isjZqJC/ej6LDejLnWhaydNLiov4A5t8a34hh2
YtcW0XPBF10QsgC61JzJRySbDsy2AUcO8A28UBD5B04v0BJDAKAPuzsHLx9p2X79
Hy3sGY+wg6lCHytQ5OnjkE1TN6BMMdZq8lA5XG+HOFeZ0+ra4+ZwpsU4+eaHbWNg
SALc0jF4+Rrow85AqaTKgOdMUQJ86dpQceegf7gQq077ebv2hpTIu8y7lIAttv9n
6aefpTso+6dbJdt/ckD2bdrCHsX0cQzAv+slYwOo8o1bjrouMnxsaYNmAsh/OXac
nzoIq0CTWf0VNTGe+BTEgav50fARSftwJO93vRZY5bPs9arB/n4RMkq1CPoMC6jN
l/yKCCKnyYrPBOrMEQ5reZG+4t0Mvtvh+bQN5WNX2GccY4nkIs+QWU2XnGrFL/k0
kG6448PYxUjv9z+QWsMe7aqXW/qKVfK3KS33tWVqTYKlfp5p6H/LivAUgIcUkn/J
27xw8zV7y6pPn1SO8IxbJPz/eDnMqV73KZlQFdthP2UgIdKqBTrd6r+ocmRARGuS
/hYmWlE8wcSmb9DUvWLHC6QvBthFMkQyxdCQSt04+3EcAKJISt4rIlhgpE6Kl3S9
l+1PThOQ7bAO8vznnbiwRH5zh05946DNrdc/8gvx6CqVFXEy2QXR6xS7oSJfVQKO
ywuQ6sFo/JeTzvlyzrP4ujomeCtsoaQRXVALW/jTl5Oc7HYGcuNKV2JZikF3A6Ym
uV7cbDCdTZk6nXy65oBsgYQLvwQTgd/0gVBPNqOlyYLOsrpL1ZBWMe/EMXWKGc9D
h9MAKFifRSCBkmLF3FxtlWH/W8/q4DRlN1I0KTZ3km4HqO6bJJgthaVisyv75LdY
1pQpL5NuJoiny6uqhTW6iP8G2Cxhy2BmLo6e5bUpX1KaIVsJX6RridObapJCwCvE
rkFhEeS4a8nw38+OWCIAUVT5/77IkQ3jzZTb3RF559StAQ1y0Mo7LbeGRbwghj9N
gOrCuGFUUUVTLjVouezte62l+p8m4kWjLieQ1C7GikZN8jTMiBMk8IInNWBFwtJF
oQryepzq7qTV5Ndd6+9sOK3cwbdbs/hmTzZ5NoRssItJgab8dlYgrErGylg20ogJ
8G/RiIGlPUd6U1lrS76MnJI5T6hcTstDW6iqy33BORTkJmnc7R4/TYvTlJKHBfDW
l7WSs0A9kZjJSzAARPiXwmaZRHzQn0GewaCCFbAw44F5uCdEZAv7FvU4ZQjSU9uo
Z7XPL+pHKM74YXMjpjaG9M2DGhbaMWSLD04betYHke4GiVdwsPXJKTENpsA8U+Gy
w1BT3+0URrJfv6lWZYHfQUpBRPRkYjZcRrLCOdRQ2Qiis8gNtqqxFuK0wrqNerc9
Ql+qmRMzziy6Cnm74ugg1WeIHp2Rxf2NWh42sMV4F0VZpuH31/eghaYgB771Z6kF
wmSrDSAlEmxGmMMis2I2zqCuJDzDv4Osqf7i72BjDsmjn1eHjO0BVZ+qXW7JRD+8
RxD81UXgp2SihQzauDp6kvJKOabeFRWQJ3DvVoJTzYCqRflFjY6KunKbYPXDowMi
nL9sKRTHQamu0tw/2+OaRY5v4hOEQ2aMSz63le7IHjiLxtf1SOt2jGNuHGGdVWXV
1BSQIVy1MXnvU4PwgXq1FOSw71NebZ7F/YazLVk/MOT+fESdu6PG0M4S+28yUPwT
Gi4sBQ5vmyn6t1DOv2AdJZ5M8dsh9YB2xrdeztUampVZKgzwq7neZ481nBKcCcYP
xSKiFCnYN4HCEEH135ydapnr8djV43GOCVTjXyRMoH8iS9gJrpog7YoR/WOH2VXS
jkZkDByeBP3+cLO/Stvaig2O+rVapl8n/uknlzTkzzZlQL3dbu5h9FbjezgpLKaL
Bwfr+JkI+B4XPDxWNoKPSu0A3Ish0LPM/8HE0bwx8aEs+zhMtDp8PhdzAo8aQr7v
c2K43bGDdg7Lwe1yE1GAfrjZqGGqifKVm+9KaKk30cUqaq4fEzX/wAmXnQAtXd7t
IAdvutA+RZ558BuPilAkUvYfn0GvN3Yvo5p+5npWFWDOV6dEOm0qxy1/UmWiniHk
zAuNGUFU7qHogh+gLMgNSuVwSuHjecXEp73CpXSJcmzbpiNSel55SpPdve0K13d+
5mf/eIuCXcww8SSpuVe5pvqLEKtrTtm0gD/wuF5CG6Lu3sYeZptZdBuiduZ5yaTw
Qax6YzcvPK9d+/SThC858UzIpNwaXpl8OQI1fmRbjelkPgQcjkbucgkSuZdTJQCA
iAzpoOLegp0O5JXzXR/m0LvNM8xeDcJbmPpNWPEhROBd1ZjB4iK1jgtWM7CMR/wJ
UifzRIAT6FDZ9WncdL2o1sCpnr8UgOfV1sDlPtgxXG3pTNiabKkai4NP76rLu9cX
WOniElV78wwRQqqmCzdE1wmSqyS0O7T7jB/5YOGmP129prSo1RSRz6djTRj3JrkE
heVA8B0rvpAhSEJ05eA0k6J0ZWl9GUAI9Ce5htTRoeBNPeANdEIiVq36kD7QDviu
nA/Muv2bhIvlAflEIyg8u1v7cyZu/ei7N0b0h9s+puIG/APgj8QN/w8liPZjvnYt
H6KICvWIDHUE8FurLtBvJdXeQUlatNp4Ad6MsErqpO35DcwtcjnQYc8oghZR4EJ2
tpGlaDEtJ2pYxTQOPHSydQ5jd7PHjI+HfeaTk5Mj1gzStG5eZ1tymu7EnDagkgxf
YvIs5b7uNs34gw7IN0StqnYpqBLWAz3WFIE1rtVc3EaWuINoKfEREe27jK3bEgWF
1hJhowhkJYCvlkN8UNnyvcWp4d9bwV+RosAJDs9bbrTC/zGfVkdwmQHYtKoCWv47
R+Jv4ZqSdS8Obv9mX9V2uSrpnI16hsNeGnB4aa5HsHkR6jvnVq1ODMVCIr0KKBEt
Lt1YBE8RF9YWswhRBdWWcEKvdtceV1Yx3N1+/3lzx4/rovpPk2xesDkuqDQDHSh4
WYgNyhtUq+lSRnMSZrDr8jfOr0pTmi75xEffs0VF6sth9neF22dqqABYUQgRziOA
fccPoih/3sWx7lAeTgF53LYZxRon3Kgie+zBQur54GOwHciC6mv6iYcG9g7/xqzC
azhdQVWCN91w9UA2JQa1hbU1dfN3D4MHTw3ZZa8lk9ePp5R3LzFEg9BbIBYI6rqV
COanyIVe4hgZd+v80yUH941/zeqVSXXuo9IXTe4A/FRs3bT2VF6DNDAaPug03J0B
44IFO5c/heCUf0DiIIoOslgUTako0oqXj4C8/x+qoKQ0DjLQkXYeTVAojYyDTE8Z
jkxQ2xDennwcWYKuduLaIYz/BxXJjx0o2cC10YsGpIiCawQyYH83Ty2Xeeqw4ZFQ
uVsisSJ0RWAYMdsfZERviNLJ7UvcLHTbasxt+JyDhgpYJYK/I8h1TF2V/5lmLNiU
how/jz23h7mPXcJYZ2INpjZf7VUOSqMgvWMtfHoroO51qXuugCIHAz00rcF5s6D2
IJpsyyYBNwE5FQ/+ZL93S1Jxi4wx4CzdsnObY0VbQNFAKp/F2EAvzR+Jc9FgDf+g
7m1mdupfzFx+w/bBCg6ZyV+SJKcmjMmKD8CWLH7jtFd7EkhA5/g+43hA2Ulmikex
LcKOkfTVjZYyR7heLmVBxpc4YM39pAzR8J0EPEVvHY79QeMXC9ATCWzpGgvwIH1v
HF6EZyYtQy9HoqimLhMNF6QxnYdA+3/dg2QxNiAbg4yLYE386JnnogPWl8oM+F9b
cztKnL/OMZePxUbv2MI38f96lYxUc77/cJZHaNxnKUC0A4vGZ4/Asvhx8vgX6JVL
njfzEkT03hCjyPy+GSR649zCv08jWbYkrDxnv48fAIuj0aOojIbl2StnV35at6y3
1rhq01uQKMMDnE+VXJ6kZTLb27cmhKT7UyXlGFGS5Sw/JslBCKSlKoXN9wlchSSR
W9wlPOj23+HtMgji61ymXJNXVznBjBTGb7kVSq9uPr4UXWAdp/FwZNfooJSxFjmO
mT6FQ0Tp0QYDmstCGh2zKC/L7RJKnWljabgADuoWaPR+zqnOWu7ududW6ngjXHGa
hNHn1mbt5qFDQX6Stltqu5ZIyEig24qWitoYMZ3ADRrxtI0k86kcZ1u8Cmin/c2m
ngfeIiU41kupOJkr5dpxPThDV9Tl2FOvYkFEW5Wio5k1vSLc91McyRT8ULd1Pf0c
U2aihnGmQR7+e7KGAlTkA0qwczHwjaY2PngMEVXH6fPDnVNe7FTN5/JAMeCchRbv
2gg8WTJPOJ7E3ZG/Gmq9pwY9t9PB5tVyY2YOv0r7sOawmYUziIiWUFjziyCG5Pdr
l+/OagAo1y5yo+zK5+kj7O+hQ1np5WzRJ/GtjkznAPZDS3Vd44VKAI2XVcg70k3c
YTjcQZeyMmbI77NS8EX9FSYqH+4sb5awNpE8gu2sUBsrglWF2Os5NEppUYa/1RQm
Ra5COKkrh/APXvoGI8LYpc+ubH1pfdoPsn0N5LE3pAeQYu5ruHzsaid+PpUO1Mk7
hP2L/dAbN0aRNa02gU5favscMo2qJ5/Hxx5oLD9P96DVIKXQwJoyniwvKwz/gbhc
jnHfO+V40cpgKxjZCbEkS+1+SLt4MrQT45B69SJfiMDY7JIgSJ3EVaEDb2fPB59w
GC8NhmL7vup9xYFE2nVhpBZBUFHpvtn5dlXiteBmg9f0SWWLnnDLsU/+0Zr2Ai5E
YSTE9Gt0N6cQavFHm3IZ+/15NSTDureMT3CKL2T7ljurfgfK8GiSU28Dlsze27Y9
WAeBAlP1sS1DjSNC3Fos10MNX0KN2ovM/zWnhaxWZ0IoaGsDgIvC6gi9oEUJPk0h
k38GlLE1WJoCA80gpsWaTPvoAGrn84TfmUDVkGBWDCRxrbg8ZtRClTxxb3L7agX4
hrDkCCtM/CAn1yyexJ8vb4yu84hjhqmR9GDbzeBmNOJBL6PTpTJQcjr9d2FOpkSY
TIpsECjvllpj4wHObHnqTt1jqRKWshBAJzgjeQqAlogP9eJkVENPP8xHWk9PXHrt
R9nmTGjhh2E8rTfO3KL5ww3T1GSreVLLXKLBCeQGplk/VUBc3ZBO8QiM7DhPyocj
gzDFncW+JorJo4epgl73zh6YbhmQ/x4gdWt7f0ZvWTQpgjQ5niAYL/YwMqHk8IE6
Fpki8mNO2TXufsHOD+Uyu/d1TAK9BF5ph+OKwjSaq3zbfupIjT+lUVQUS4BY/NA/
cTau8wOo6+zKZzrirIbOD34tu1rvl1j2wq51Hmtdy5diXaqSXyKsi+YVgtNbbaUR
43lfi2cPvcDKx44wCzNa833ql/gMEdEfYzRX5O4wVdH2vnXMTx/CPc/Uva+myTv/
+WiRjLgMDKGiHs6t7U9KXJ4UFrXmGRS7bbIKSZDJQFFaY38APpGhN/AKlgGnX7Z8
CG2BXlXWzguObVxaL0aO1lETiNOpqdFHpn0EV4Gd8CdKRX6ZZagoXfB7Ls0l/P3I
wU0vaO2VWBlbJD9tbbKyWtji9zNXymu/hIetJtqlT1oU4vOUOtqxMuardgoSxqV0
uxUZZIwnwiuBP0ivm1uRh5EyZHXvur9c8M0PQRGCUC9/twv1tlCUcQZMduJmiT6T
ms3EiArZ0gHhLlJmjciyje/EP/3JEPWqQWH58C88qp4Eioc6zDlAW9/V6t+CAHdz
3gBVmJajwUzCgvk2j4cqVeI/2ySCn5C2Eroqh7p83M6uekEUZhQUrvEB0EOTDJDF
9NVAS+s46sa5q2Sl820XST47bDwT/KdQTHK1kbVw6kGogkQScD2BaoPTzf7CqFER
pA0gPRbUTIc+9h99l+TbuYRHyzv9jASbqXeLLzmy9lJ7eohnuORo89/zt/2W25i7
A+F7rpclWIfiQS+ZPjQsY6jlMgaJc53EhvFV6HOlW/4ENHdaa0J/YEnoT4bg1paY
119OIPj+/AV/cCEPtzE0FbHpB/VhBym5UMro2dwqZ2XHBPX+0NCp7tut3mxEA2i+
MxBn2J2a4c9zlf0egbYjbMSEw32/rlGX4FTI//KcmHYa3ERKmTwFW+oWWdF0xV/7
4lFtk+j29EY7TcDsZIsbixGvf2wlCuGbnM1CEGoWV4HziaAJiZneCPDtgKXRAtbX
jCz7DlF9Lyq3Trc4lpT7jBKoqTopguEAnWI1DWu60GPZSbUxq8UIDvRKEJXE2n0v
j8/oUHLYlQkjBIUtTiTivguU0Xt8TTRUdvHVwPpvFqqew00+ygDvmRdWg7gAY15u
/jz2iMzp9LPQBLmeBtuNyWsUPkTRmIPBDhDnccWEB0ka1zfSD7LkuAwx+iTC+Xf6
DLoXPZG/fQ4ttKgWbTAI2ogIKehCf1DIOdkWvEjrvVsXkR5eMktjOGrzwBuYNyX+
5bctvL0KRg7yiYfUT2y2eRYIH6IbpxpVOTtU9L0A9lNWXhSUb8Ndac2dGFF+598w
ThOwD38zNop1rb4lYLDiqB21iu5fqMjBIuRJixGAKhmdbKDDtPyB2+wkeJXXWIq0
KogIHyeTLQfNqQZ5bBvTaXoY6gOKyq6xyhgvHgIGjD/Ygpd4jGT+qhAii2fnxKz3
ilsTZMEXl1BMiSJb0Wb4ZkA9K3qaXoJmb50PgsuNGjNo55j2DLH61vkaY96n+jmv
GMqsSyQuDaQ4DYceVHa3YQ2tC3mJgZ1oIdVIcGiBZXyCVRd06rTE+oAb+2+vpN4h
mfdUAdZvjmwFDFoEwav8i8dI4/As1KZQ3YAC+s3sEOX4AIoQKcECnpjKrAP+XI03
KpYI5QO8j3xngT8LVehd2FeumBGsLalDjzXgCbbJbiSLS4c5p/BhkCFxm/iEAxzw
JK7fdnTl/nhEpL/kHwa6Hd7qqxMRtEp/BZ8iEPUvi7I03vkXIsnsaTYjAbTMTZn3
cxgymeoG5kkxss4hm8BupzfnJcpemN1CaA0KNErziLdFiSp0tOk/8jjiu4omY759
eCRzECS0hyRBaPV4d2IsvFdHCNOU8pLmM0yHHlyHfce+c5XUU3uNcyzZgpnwNUVq
sj4kwoBinbSw9GD0j1H8V3idEoN9m1iuW+2/64DkGYgARIMJlwYbST6jjFNqETHz
t0ObqMn+IVRZfTNPDH1u9OLS/zRST746sm2Ud2S+OnM/bB0jnvnwHj2CSLjUYLxd
WQXmqMbJkF3CidXoJjyFqwqraA9MJ9H1+YWuMaufzRbzP1ri+fdj/J9Yg6nxOT18
r9/5x0FCAKe1I2p49CrJCk4XN8K1TefkZf4z/LAiP3WEjrj62qEWMson3nQogRYo
CVgOWza/HutpkiiUKnQH7JwSYmjssWtpWJMQ+M5h79jcF9RKqwFRz0dK1GMVd+m4
Ch5f7NN/gsZFIcywBQwhqDFUpMGG09sqxVxC+3VucwUUZjZJ8zUaJVz1hXIwbMfB
dEDkFr8s9y5gtG32x9/s2nKn6RqyqwNrFlBdQAyKNNpMaaJslRZSo+5nX/vW1nec
yaBD0TZSb/cM/mN5/gZAeXxSlshBu6XIFFz4y0MArvcUDH8QJSbl3YqW1/xpGTdx
VK7gU/lR4sx9Kklo+QY/2mmkqYlYAo4kTdkm5ZC4KXQUNPgLrcROdjwpLD4jaYcY
eEtTvw+azjE9mQj+AO4Mk5fQYL8fd+5qihaESgCuoiudFNnR52gYcNKJak8CVC5A
cmX+GVMB3BvvrXZbeqPZXaBPLhgvwFB8XqOQcnySBS30umLNIZzZ3lR4y31UyjUY
nb4M3VkXwRPfXyaR2oVrAWOJdbXzAg1wKE69OZS0rFrqDyPeIeuo9UFJA8jFa4DI
3Bkb8sJlJWNUoTzzbrqagCIq+Ctj/CDBcfrv6eq1QhnVJYR2NypGlirHqypEi9eb
Za1Fd+ShhZmawYBlEh6OtlJovhdUDm8tH+fmFxItrHdwz/zeC6KR9tN3wH/c3SN2
08rVHMHG0PeNB3R2cfuVGYA6rYutf8wUI3nNwftCaeLsSLSezHKjFw4N+7LMMXc4
078Ou8+Ji3NAoArFUwzhDeIO7viCd0rNXuQ0/VsIyL/Jcm/3GbF3ipqQmdJ/Ijq0
6O+8kDUhhrWeuVIn2Ho29DfskfTj7+poO51pl+IPtZjhPClv9pDmssQLv97ZafHU
EOXYRdcDbfM4vZojq+HQ8+UVsmzWLfSIE+fafelmUr3FPstU5kDTbvjzHOsMtgmw
F6ZmRTw4hrj3etPOfa/qYqe0sQO0aedhPGMJsu04u5MKHEIBZ/82Sclb3xhUOEnM
/s+E3JBDyzg/BYsMQ6Flk5KgfCz1vvqMaX6IkVAoOLrADNKR0r86iq1k4F0WV2Az
8pvir7jLMkgHV4SGXKbnRIF1UP+Bx0vg6YqpaWzvw104puFoj0t6paijmMtu8FWA
3M4Zk/l09GeLTkmNmfpu5o8n+fBuwgmw5N/X9PHHwvqQnmIFVLzqUp2052ZBAE0j
SNfVBYjlSdGhwvqV8VFvNbwVuOjCCaj9UBnGCl+Fiw/IUmnjbGBvqbrlJaImuWkj
U7GshrI1PtexilCfBlC+ogDVsjeN7TIVMzMxLoPtK84GBtVLh9+LiPUf5rGWosEv
z9w553+gsF9GIgJxHiguyFKigXwsn7HW/ON0pQjhwEow+wfPQGYhSnDsbzBwA3qa
NlXP0dhLihEh2T6X7Av7y++TqGSB9hHXicnSO/gscbu2U6UCVIoAQIaqFitUTbPw
abbOST2/7GYlxLN0eZYmiwiGsQd3RV6sbcXTlS4jHgWZZDaRLepnKByIApgwtDRQ
P6+7T9bLZUMl5kj+4KgTTZ0Twm1RpngNLCZjUvNIDf3fZJxN1uEnQJRJLxtx9ylO
8M5Mo7agCSPeIcmxx5C15j8ajISGGflnHvtkXEx5r4LX2fcm3UNCKZltSXJjyhIP
EDtQLbFRqZr//3ROwL9Ri/0t269L8663UuiciKYwUf5Es7aiVCq4B+7pKFdxwK6t
vuR1rcJrrpB93gU2mGSS41WQu/y0hifQ8C1y9wk0ZlNW3RiAIQiziktfOoKTbp6M
hUV0AwlmpZpZv96dhePDKsOD+Zk8feGTwleP2YqXdarQEuApA78qvFPdeg+Y2lW3
pV+U7dUQZDrswJtmRAPM0ZMur5aOIqzrP3hL2H1W/zhIKIPdjhQVgGtlmBlLHhRq
gTTQjrV/QWDvrzWmERMgUFAHFkqUs5jOlsDQoXA9BWfbCa5DguqMBMkQoU4hABfA
M8otSpEwVJwkVOMpAlkp1f1tS50HWpRfLyfn/drpluGcp8OJh05klSgt+qYyvyyN
PTK/0xBLrXbrnuTCe3cNtaaM4ueRyQpJ/du/Q/EBeYIHhg+irKFSVXn90g3+16nO
8M2gkcZFYyRvhlEEQABAUOwjSfHCVuTSF/9a5gXkiUTgLIw2n+KmmLVCZWzL3piK
ahJsiGuPGnMBloxc1rwWC8ZhUi5RW+WfZbeVoD1FaSGC5cKugXQ5xqLStEFCAiaz
sPwE1NTfQKoEVlJnrl0qc7LYV9SSA9sxp1kTsSd++WY5NfV9ZRJCNqFJXyQ4toAn
PHiEZDJ5ksSJ58fyKdChBvoV/0P0Cd+keyEGVz+3DnxMZKoBfXoGCf2zU/r453CQ
d9YncSJiwOJcoFsMGs1fMs2q414v0/51WQpl4/hbDfW8EP0KZKDMkY0ZCEVLtKIL
GHdiA6rguRCnEDJO3y7DYfR9cn1+1PZOZW0x94lrF8jbP+pLQpr3l2te4WR0lBpn
7GNdkuzVG6+gD6BvZtYr3WB/eJN11HpmuHA8+9kfBC1YxFGiMryEtQC6nWXRrhnc
FUMIMS6Xxm1dmP4zW08sIVbOCji/2fh0tadDAZ4VcsDnj92IhGnrZ3d1nQQTEat8
0xk8gvRbTdTTRi4rkE9EbpVvW2Z6wbR161bHohffWsUxV89G2kptTgl+Nt1T0Tya
9D0zpgX1TQCin9DKSycfbpNZeo05MAvae2wlvHgwETXo5a37fyK1j2WBkA9QilD/
3uMre8JfGvGv/dMQq82EQ9gF3+H6EcNpciWfw07q0Y/p+VjmAscCilSsqZ1o3HJc
a8QIiRX7vv59IMw+jdsEIP6x5vZ8LAJCieKJY7McOmwlICV157wgMObEuyWNrSn8
idYqL7rAoVRuSnFKzV7Ykv1dlor6tu+vP0sfmjwdQ7mT499lYvjYQG+xb5wml7t+
UIMs7kuievOlSXaCA4H+Z0exp023/0pXpQMjJIiS0Lkv1oWNOQlbGQhXJvGWScyw
GG306MPzfYeci4X3yfd0eFQ9D+b1bZpp5enRAyM8Ei0/FdKeWNrOfRQk6x5XsVge
IQzMmzPhBlr73fCWIfmRoIv2TWbRsr7xEtvcclcMu91l/aamVCUueaxN6yyfvCik
x+e30E0e5YrsPQ0M+LYsfEuNABhrKgte6o3ZbZXlxsG3LLd+orzjDSjcghgQb8+t
yBq8onoOg1YdG67vyD/DqeeCFT/IAVuaTRSqMywC55gXk8gKYLwzsxeL+aK+7gMr
xIjRtzpTK8aRpN9Kyx+IOYt8V5DhVa/VQTmPI8wfQ/Yae2RaICLbnMmmx6pw/0oG
rcvalJe2InnTj7YmucPg1z64ObwdXmYD+P5a1AZaAhYN5/A2VC8jSqpTvMrQBS07
pAAGws8oV1gwZ8I6yvA45KHzA8MKqkDie2M8jPdosnbaampti1Go9oUDlQBF1jtE
fed96xDZtj/1NgX3p0vVmA53WRl2ZzVLh/P8HIM3yyRNvWg2p1FW1x3e0adrkBYy
qHrS5oEaIGGstfGwPeTqQmdUE61yAN/zREey7tIsVaAL2/K75oD7ICz8I2OE/AhJ
6Kj5arPM2Uvxc10LVhXrl0wK0mK8wapc2yMZ+EgkvZR27qcLkVGbp8sgBDMdziFx
QaXJCWAe3lR8Re0yPC50R9mDcnPnnE8rn/8UMDXdwKcyBuXg9+Zkpj4Bq4XUkp5I
AaH80FB1ylx7XxjTLzaKyWthUj4l/KppOW0ZgKLagJYQli+7+PnretOM+YduwOua
ba7v1OLAG36sEkCZHWEXA2RSo5Hz675cLSXz3Az8Sc+7pSbeM7ominWP3I4epzxg
zeNPc386lm8qRoOdtaOv81ZjD3GTpU7HPMxJR4j77yBGgNxGoJuW4810ZuAT+aAo
+CbiJbUr9xeYOq8auiyXvxAT2nIsL3myQi5bGdZYN1R/6QNjrSWBxJBN7ydijt8e
9CdOHyhOAX7IRKrwCVToX3iX7fKXiQSQ8+daOWvMgKxNEtXytAN13yxrcjaxaXhi
WaPSSallLT/hDDO0sFsdjZUQhW+UlCyN9EqHUMmr2/hp0vLH19+7278cwLeYkHHX
ulpay/DqFHA1vT/hU0m6/eRFrKJkkwYCLLlwZE7xZ9NZC0FzMwPIhKScAFOCzsHJ
+KzKddIAIEglf7Pq1aA4u1n4TdFtX4WFsZTGpQba60QntfVXNJfEEfHGqN+hdIno
n7fsutNVSO0I34FFPZxy98FcoG25Et9TQZ8AreT9+wO6S72bc1d1FyB7o0y3XpxS
1RSuWo4k4FaKlIy6USTo73zipmjlsTWMZ3ST/UmhO3kxUjZ8wOeED7hKlegEzIZD
O1liIPJ1eMn6qtLGf6IJjgelIGOAyyCc2d0z0prv0mSnWfc9Yx+2RrlkS7kpV9we
B+j17IPenIjzQj8pR2Vr3dfshS0jN3oXyIHa8TWRuX4NMyWkUr6JALO0rCbF5tra
2qYrNHgjPFG5ge5blwn6FJ+AIZEQcuwUNzTDC0dA1enQGImMBksgIDycOfApOizq
1Vhsoz6PuS8LUXPWNkBR7stsVSp9ma/Lo2qUDXO3emiFeMp2OqSbbTfUHJ7rp4SO
WSNwxA6rYGD+xEM/U56Csy+MTmCormNenB4S91BuMbg8HkkkHRmbNw6xF2DXOD/u
S7MPDcIn35lTdBJFMoS+JN+OqNUBY1dC5WqjnHRbX/ZSNi4iOdW5txTIW+FR30Pg
ZK+HwDLfyLOjPDqsqb79jpAvGU4ZwCe6KFWJDGZIXQXvVFiIHnaiI9A1azxYt3W0
GXp+TpyrivLCvteYjJYsNYt026zJEOzXicKMiZDf0XtiZ6kUtYuMGHT27g6UuVpz
19w9qyKjDwQsH52DqzKHgkamo3Llj+EqTQuCOtg4bu6JL5kZObkCEJXVeMFnvjA+
laLRW37ILCnjzs7YHUn9HvS2Wl/V4uvlfNBVXo4RSQlUNFZHiMtm0PN1gelOAGRF
G8QKWN6x54Rd8rdkFOELvEjPv6SiYdZO4n3MDERSy56gHc7JmK1/azY5DMVgUsLr
sgTqWaal6iBIID5n1cKEDdLSnAjfNFtmoDUFZsnGX7VquHKI54GFXxuD4grAXmU0
ELFVbuZs0ZoTRxFK7WN4KoUIL5vC+ieJ2Nse8r93HKcnLBCiSdmiSDqMfuQtnDoA
3Xk48XA+YImaIRx0BsmHPNr4lvAAkoJMI1bP8h+on4rCoi1cgF7p3b9lsmRaES6U
4lTjSt05lKKG1RdUJlcNaFKwKoEyVsthqaackzXAEI+z2aHMZYcR7NY+fw609TJW
DakrH8wJw3kC+iqIcsEi6rHdbg//UYvCMP5CHISX70JrCUTzythIOUQaZwGwDT3I
uOEKJg+eXh/Hd/NscQWYNQBEtVO2nJzaOAfPDLF5Iipi1pT0yIllLnu3MQUqbXm2
FjUPcbuxnTnwumsAUw4Yxn1SIy21i4D8Lzk7sPj1uptavGlKAKfULDJiu+F9WPg9
lNnOjCtA4KvHv9o1Jo448JCengr0TzCkKPxHsjGYhlxc240kOheatsWWFJVr0Np3
kpQuwjp44n0FwYf842EUKiK7rUJcZZ5XjpgXn5eap2pQx+tDU1i16wOCfDRUD0++
w4dnBuFfWYkfMCVp7anHTZiizvf2te8x4QoawnGj6ppdOdykzDhNFO10o6oYZ52Z
r/Tsgpl018lCRROcCbYPPLVpZ+qrgiK49PE9t9HgAdoFKPmEkO+ZpCW4MFqOcTwU
gAX5OuYsa/pyKn3jm5NznBvfy1UMuhUVf7jR1BFi8heg0uRLb/bXfxewA//VjlSI
vu9/wTsiSLX6isbx9dlE3+F7YjbnW1zL53p3L1GXi94lobYeWbVeqh1PlD8giA3H
q7qOYwx4QLOz6uGvKJ0ISrFnk/uCgReR49k0YJQC2gYPCfUcvDj1a4Zg0Tr71eak
XvWtsKqzootJfnGI2u3Em/kuUpTQKVA/RjJJMjMKdglibXq2E+aAEOTqIDqMtQXE
Ba8J4YCy5qXArxH68cxztyO7jRBavPVywn0bzTf8iQgpUwhY4P9mDQ8sbt7J1IBS
yGWLcNdAR5T9ZksyhFEN9uvvXF7P+SWv8p/khO87rBHxBFk8gV9gkCGJEalVW9Fv
q1T62+kH1NrufR7Wl4oKME61uzE43mrFpSKUWRHhepIGMGXlzXeWjycNJDWpVye/
9IfjE5+VWbXqYyd/O/s+8juIa29ZYjRkgRDorGKs74Cie3Zke2MOkeZXdEPX7+0x
bpowyQYFRtB2SJQ6A/4MBwPphlPnTNqppLSi+YObAsi3Ua7C1W173j///hfSAb9J
7khosVWkESEpkqTOAfGMG/cih+y86/f4ghXMEciOligvBZVU8oih/USNFQ48GqRj
IornhaNifKWBMbdWUg/H6Vejlm7SpFlsbELHVh8xbidss5wojxbFp4woGuJGk4f6
Zf3JbZyLvIOwNEt+a1LVpnCKCfCxQMjjmdyPtfCsxo6a1LXf2DA0mjc0fAK+pCzf
zgmYiesciQ5DUufT3vHGubYQ+U23pVFN8EqNzcGRewpAj+8R2vI6jNb1CYJvyKwS
2li9xBlXmMH9cdWgTqBMy67XmMqS58SUQaVjypBPXPokHz1iwzPAAAkh8tPa6vBU
ozvA4MIsk/srzHGD8Lcb9TeMuCtIcosKeTyicRNzd/4Bn10lyBlPWEnucf6V3DMf
MDS4T0lMr947WQ/3StgInAbu89proEpSQBKHaJsKSdJXl/MZSJRV+wxfjr3lMbVE
Mj8++ZndnvHpaXx0+XeJzBatWssCHlSoAIrPsYVM0wFUyaGem0ljpLfodRNa9ZwK
ruobeFJK7J/viQSVee9ZKkrsP0O9rPMcs9BS8rizEIDus5vIGp3xI/alvlkf6hye
8B+iHs+Jphn2qxVxK3JfZneMbLMlZh+2xjFfuusPDjledQuBBt44BR1Iu1hmx75U
CCddeniVKrn6WeSoeeoLyUse0rlwTbd887SRbw7Zdng6gcdH25sAnamnH738pir4
t50G0UaCRVEFo+FE2rjbvnTNBe4TRUJ943o2WNlyKdoH0fmFI7UvZbdvAc7KDwvm
WFVf3lSpizCSUvJR40aw86grPmIC9k4d2+tHPhi5bxDBMx/QXdccOtEEPYqIsiCG
/m5RyTM+FYnyTBOoz/5FDhIvEsx/Aw8khAYHx3KxCjSTJq4JP0xZi3fz0EER+ziX
jBlzjE63xhzEoDR5BfRtejXWyl2CxWkZZpawusUx+tPxGjq2KIuVkw5EZvgMWwU6
rV/ThPHK0FGQt2/PQg3jdTCECM989lXDRgjf5cgDioaiGxvyWsjNYP3K4aqzQ33h
k/yb2YAUFWqYKzRNH5IokYMqYtHTjTKjRSOvg2gFR9dVoBD3Bkk8/CSeLVxAIFJY
fmOm7qQx1tjY/HLDkQeI95inSFoTc2m7H5C4RsJa1gEbxnIx88L+CEafgGwbK7u0
PwZwO0vtLYH76BQVJONgbosKOjyxG8kO9H7963C4UmjCcceHlFZGWJopgEjWsQxj
MBEW0XACWa5D8vUPLfeC+boow8AEv07Sbatw7NHJ+CznmmwlREuh732P9xuos/kO
2EAaUZvB3vEtHVd5xP/mNY/gwj35wbQC8oX6WcWmvkNRcKtP6srhibAjccITHO9+
aedCPiQlMsPfSqH2AwFFDHbXfK/MQuQrt387HM11/7qXomq9IFHAJQLcAQHJIllZ
cTO4BJVSRQW2YOczNtqnA2wFrC3lZK9Z62k4T8M8BksXF4UioAeZGqfbaD9sTvUf
G/gJnUjoEEKPOOsI473yS84hBa5WyoCG/fh1kp2+ChN2GbRCg3x5mPEJSUJcba1Q
3HNn2ORubPRjogTbOlYRgrvkDmKlgHkhRjERBdr7VbD0S2vXCaqirrgFqNBJD/Tu
AnNLOWte25+UKoYyojA61jsVzYuZDHYbnwuizGO8qOJz4f2Cmg7Udx16ooVL3AMA
F5+Uf+yBy5mjV+xUTuda41SEEmzCmDu5TLfXLnCJTYwJpRC6Dzv48wwLI0+jO3Ms
tAxrhKwQLyswIAq3GRyLm3R0ti4RhTc5+9N49t9VNABdkieSv+04AWB0uIyLRwGy
rV7fYbQBNrR/cGKbEiNko0tRVCLy6k7LP4rfGz+CsmO2SVgFB6uIr2lmZn3zKblw
zUab9OCAtEsienjrghRde3RLkS4Hhnwm4vOO5hB6rh7onUW4AfVt3KbY5rpMZ8gS
1d6gM+PzvmxbRcIHx/CFwbUuUmyrknLLXvuvgrvRLzeMqOfbzKVVH4gt7mhbjHYQ
d223TG3XQZZVPoZRMgk4BBJpWJUArytlcJJZYV3PejPzIPAnP3n8KDdhkpPWWISl
+EINKXSyz/H7nbbSS2vzS8vc9BAL171OnaFriXtMsKQ5zHjuFS99gKs6ExKDfowJ
gLzR+piuiYe3tmycUBBtmi9fG/3ycwP6BlVhAhzOwmvTD2jUgqWP8vyVdrQiNm5e
PWf2AKSq73HHekV8Zj1ccN4jojOa4hcMkk/BUL8UhFbNsU8iz6WEEnethQXSxJuG
oWrT71EDcJwQoYVrt4pGHtIRn378h1ywMXl9N3dbUL9n9emLgWD6K3UMhPMR4dtK
f0NKt8t5bVElA2QGAY8luhLJns4GyrY6DkDM4/CK0OKTae7KG5pC2bgLh4sYFeyJ
kuj3nmDlPWvfJPf5C6gYdcCDE/lnr2Mu1aGqC8k60ULZ3f8pUPxhpkLALNi/Xlrn
7vuTSushqBo8paM+zDltda+SCq7PqkdiXEgKfJpNLbF1gJkHmsqI9TKQ+6vcPBHz
vu8X2KGI7UmxA/lGiRDaf0t5G7vGlILOoL1Aj6Ub+uIcVtkcer458xENg/4abkC6
/Ctt7xoGH/LAyDw4ULmEnuZAct42w5kRX6Em04kfe9ND5iubrE7Wa594iy1mg0J9
NKkvnPFmKsLnThGNJO/p05mbCArKo2vjltXA7HLKX7AcqIsSAD5l85hke9VnT8qh
9baa07Zi6wVs9o0rdikWGcO7EC9V+qWwRYQ7vpVK4iTMydOvkud3//FQ9gGe7DLZ
IB2UjgsO7MSxOPcQih7y2mMEt3RlmN0lAuhomJ24B3gkUeJ1YFAnSs0Y81WilIKB
C6rOMTkJyu5CN8aRMg/TZKjkQPS/E4nBqJbMLehl7p2qW3YD11c3XjYU51G6IzNZ
j5hhSTNZrdRiih32KiZXAwnuUK7kbyliq81y6aOLDKhNB8IHPxYzF7D6rb4jGgtK
nOMhMQ/d+0E3qKKkkI3JmrOjka91y9q+LjgEUS4L1shDUvgFEQX1GdUsVQRJpt9I
ezwkmf8J0vv2xQiVB7rH/3Aq2oV1WJhyWzkPWHxikeo+ORY5rSMO7GfBjxqOUNUA
AngxXY7bXj9WdvEEO4gspE2s/tMt2Ge5rCZwgbSbXlCxJAGG3T5AvAAYFuXd6OmB
++njef5jDX8mEmA8yAxcLjLxY1tkbMBDp2WmXULf9GnTz/3V3wYKpUiR/xNr8nxF
ZVgn/VJe/7Y+82IQCHkVodN3Q/BPWf+I4aKiC+W+tUDjtZNSyaJ9xPLOIUmFoqt1
ZvbxcxCJytPUsrKPhvb0LWSm4Q+s1zPylN8hvez0sbsQblpya8VPmCOCKdyDvFCc
2PredOdHEU/9eweZdftS8eDMTKCAwF38jYJLG/pxzc07ExuJc3oxN/D7UoeBEbo9
IyY99q01fZMuWFPxSJrudWjrCjTMjF+woRSTzw4dlaPxwQaDdBaSbA0uH0voOm37
Y64KUydo96CHMSxIWzBxx9jcASDHOO7AP0NpP4RG6yol9tPZX9FlM30rpOz1dN4Z
H3Y3VqT0A6/2wSXknM0Um3UI00mb4csQroYfqZzgPUtK8lVxO1dYzUx63O72hrdx
U7yotx12upVx/Cqpdmp1Lg+pMVrgo7b3J6ANG5klKiIfULVmrI3J3neGFlCMt+8t
KSchM9NmdmKvZA0Cm4E0qYY3CU94vYMJjRp8UoJ3xTJQOQeQH6Xuv/qPYa3+TEXr
4LIMhAZLiv1VDRm0ZZS8Xm3HSm5QkH0kRe4iy3AeId7gcsl2EeTHFpfjBJriIuyB
4HMId3PYJMF2cxbVpjOu2xP9nN/ImBz6BlXrX4h63OxQYzE67IDIXxnsZAgqmwBP
Lf4s00dI8fRW3iZ41viWBkgWZAamMOX9lm/TDPCvaib1Hj3o/dYOo2OwGYd7iZy/
VfnVddM+fY0wRqVkKSQJGVAfKLeUEyLP7UQILSj2RdVx90G/YuZ7Aa0t7lJVzzZ5
9zi6lrX/CTUo+M2r+F4jB+pX3L9ErMc3/ZRxteDffpXGLzOo+jzW15+B5ChdYcAY
Fr3Q2DgBv1VQw3FqsD+V0UlhOyjkhJ+TbSX265uLJ4o+klXgr65NKOMIWaj10Njx
vGxI6oA937uY/SjcXM/z0MERwDKj30bHf2JdSC3vmZlTVT7BkI86xpUFGP52dZoI
nt38FVX2APbNIAG0NYhvF7yWwq0Xsl+ZHDJ7/oODHQ8ipcGvcsSXzox5gYXaeID1
IMdGDta6VpKeS5eB3+MrdPiv58Hvb/6rGkqRa6QgFbi7wmGzPDMTXstIRvcA/WR7
K2ULjnjyPp8+NmO5yjXQcK8Qj02vOHHZcboShbQ6bQYhz4dmd93kpgRaT4bThITg
PEO4aqfAVVzeHUEQzWfTWAkjPi6HPTBEr59dMsmFm4/JRaJQlhAYkpQalzeQM+X9
ehspJEiMXnUnuP1OXKfqHYeHxAHJ2H6kBHv6dfzNDTavchmSjuXISSI2kljZGLBB
vb9+a1uUxXHWybGiu/Ef4GAykos30687cePFywcDTpT8eMxzwUMm6Vkv2ZsI4oOQ
3IG30KNt2vDL7m6QgmCVgGp4lHYtOYeoJVHF48rOSCQNCToOsQRgHh9OQSAktNCl
imPv8VzPqe9hsol00GVvM0RMVboCz1ua/32lXx+JziHF8ogtc/i8ygcS75IKqfxG
vTGXRQ49uaTCpTdAlXns3+nbJ7DxqezU2e+N/8Lchwsv6mTB1B/AW9JzEIYlYDMg
a0ZuV++0JjeXp9WcxczfmKSO2hRupBpNp7mCOrCQhg9iTIVaYHOqSZc9vLtr6d/w
ef/peFKWJaJy7Dv98v/avROq2ylKcUKq0BK8jN4HWaHOCrp50b5lrTQlXQ6FmMQG
r4uu8st+Ym5eRNDUB2jZ2zZdUVnltXJVm5nq1vztNyZGNHxjvveQtdg0b5eAu7mK
IbLAa8YGDY7bIT136ydGQUJB1zI611J70phSLV4P6daYsp2ijzouGkZf73qSz4LC
kEC2FlOMd5ARVqtHVq4riFtbufpgMUQgBhkfcgpGIBMPO4lz8wedXC1pLCG0XHvH
P0WRoNoavokluOGnG8Lq2yF9AB4KbRLy07y67pGK775Pr+iMOPKX7m3QWG/CyZc9
5p0O69+PI1TdjIobKW98wLUxoxNoUJ5CqGZr5ZRXLgccfzlpwg1VGKXvKNniTL+p
IPXbnNZvrwhL66eTTy31W8Y7/W5BTKj2JW1VoxwUCqGg/Ebeg06AnuJF1+mCrUtE
6dTkXj/1jSt2xnc0KmEXKXf0uZ/Od98RH+oX0x0892u0v7OyYCjRg4WAWx0g3Lbl
/EGRBGiRZ57WOwtp3So6vaObYHy0g/UGxfeb2X6RJ4IDtOCGV/ZSFUh8AHeAmBV8
nRmp36RoXXJyOMBruXXA8TM6UD5OV+zuCQZjSQWpHlu1KzEAu3TqQ3nJv1bAP7CY
ZUJzaUGZmHlADjziL34MmYlgjsoeJUXZHB/mcEjcC7bHSRxrGSxcxtX3jM4hUHYL
eNms5I/juh5V9xBTUI7SJy7rsoIppD6gn+N3cqV1+MR1cBBZMBYMVUaIhjSIBWLn
aXX1PgZITeMWe87TDY6UT8CnM7Ft4p9tewXe9kFPZmcUsbgRXHy9y6bPfb67YZ6K
pRKce8FlYRu9hTnPYAjFUa+SjXaFRn7x4Kf+LPD+lGVZLK4ENdiQ6UWRkgQ/Fqld
/FKN8tWeAd7BJ/eMdehipb5orr3qrMnUyjNzaeBjhtY8RBLmV6fBzBadJK2ik1QZ
795x3m8a4VL9Df1Ex6YuKaZtRw9IgU21ertiJ/R+6QI1+ck0Him9g0r5ovgHlJcy
8ZzTGQ8fADNdfba72zdW1afvQWg09QS5pc8OJPvHhFWP6bNPPdhEYkfr/k0Zr240
uN59eH7DW1QyaZ7ol5JxyBpBj2+b0nL+X/5aBeS/S+7E8HLz8pF+J0zy4cemJjK4
2c2Vvo+jeo/HasBG6cQX7wPEL8/Yy6rU0IJxZwG9NNCHfNx/hUXZyAJrTNOTSche
ckUAIkmtQv6N8jUHV4ckZlrE+5MiDvYeo/NQedRoWJ74WsTOK+P3ovqTJGco+oaC
Ms/B/vzyDXrfgRp+B3Q9OIUyj7OE/6ZtypunTBHBT88lggrdxpDNLqmXW2ZTp2N9
AcxSIx5q25reeYOJtFrkBzSBZkYAHXWxlkyWBBxSQiFl+WKJNmJstOaFuJ0LOjhY
0vGKdE7eHjckgybLqjrH1DkpyZQSzM7f6UUwqsLnHe0d9/duQhPhCtoRofuua7JE
aC+aoFT8Dqs3oRW2bC4TVC+WpoQnf4QkmbdhnsbzeYTasIlLzB+3/62S0O+IL5iv
BRKYhRQS9TLjTqBj0thlvnoWODRM3QLs1fsonVE6szR/KdUB6/u2edNu2Lq+HZq/
B6B3XEs9ZLTJssIqWqAAiibDZWuiAE4RXuYGSRn4kAnqy/9TOQKglsyu49hhtCm9
/B8TbgLg4vTwtAMVyDz+5Isy7kb5VR76zcJHXA5gO1+BFTxFlnIgx4chOXuViq67
VMvd+hFkiCjcih4bY5JqJnQU4dJr1pRJWS57voaWxQakH/lWYI7nZ1aJNFOoEN6z
XGfs17GsZfRb+RUgk4Mq8hA0km26N2VtFA+S093uV7dc6M64xYDoIRvpfk3ZmJsG
1rUcZFYkrXPwqSglzM6Mhc/lEjbCzHpvao6RGkrn01gZWW5LCF6oeikjqBWr5Nw5
SUNW77JEngngNf7me83xU9q/IxIfJS0mdBciW3wt9fXdsmcMoArnYArWgmEg9MZE
M0+mfRK0QBEy1bsKk8zANVu9aLHeFktajolH3txUe94Ohu9sBiPAefepXj0xZmxp
nc35YXLOa5FS034+CoKf2SnCWEWbmsd1YBtN5aCjFvux9ftCDIEBPZ9cz+TzftMi
GJeE2mWm3JiC2/5G7em5kUOjQuc+UgKOwLiJiu1iE70AQw6X6mAC84ayMHxrxWak
nYp/5dHQ5A9Lc1KxMiUt7yyAaUMPcAwNhjRl0ENevrr6ppAgEM4AESJWbYG8jwp6
f+Jcof73xoN4c6rOpW0J8pOUeQ0L6yVHuR+Bapdmitvd0AuwvXUgS0pHosfmRDU1
z1Hesga22ZIHljNHY2QJqgQuUQUJETErKe84pb3kIOwOrxuxTDeZ/7dlbsXzzmGh
LrXkdxTzVj3hYl7w1FlRH6e4WEcRYfQEnjo2Y2pUPONjIybohU0aLDFtFwD9wECb
XKD/0UaKpuGQvamwC5Ow9ShonpV5+U9vLLbBQNbE7Rilds1f7LVWpv7TM7Tj7H6w
k4Pt3KiHcJxXGHjfiop6isAk8u1Y/e40c6F9nATl5U9S/fTAhphwtz71dLxmpFZx
DpiriFxyoe7tEGtD+4XiPWtpr+GelvwhJ6tNecgTHOpSV3mIbFtWDC8YYMwPCP8k
IRx1NZU2jw4kKfRgz36PMCquggLLnqxb6sydZ0Mff7drZoM5TxxphgtIQCfh0H+i
l4z3B1Fr2PWZvnYUEWx/SmQhALJfJGz5VIfsU91vF8hp0wmrlvmoYp15ZG3xIlMV
/YpprdGoGwH4Z70R/uW3qwE4hdRNMUP9jW887U1VWhDoySkumJyMZL7TWgUtbBh+
sHW6IzwaS6NvRw5YHbQWES6IkrtbZiHmy4i8yNgpOCGFBYhSQq0skZ7lqjjcNg4b
T/4PVcaootzVY9d1EN9MKo88CnEgURIYfS+lfP+debdFkLeePbJ1uMdNoNi3Cpz8
/aHk3Qd0FbvYd87t1W/bahbmZla3TXtkLB6sucxpavMQfzoMQWN+/q2Gd/B1rEog
LWKQjAIojONWakeX37hZ4wXmrMbFsHM85b5+MyV926Wyh7wyVdGoK3dvLVGBCnx8
olLK5Q/vgX8grWUijmh/aeacNZ9Ha6MUXMqdTUVM2W5qYhMw68ebuFSy84of+4sw
+7rKM/Q13ExG627JUdpj27f6NDy8oJJ8eeOHIMPqHibB7i+MrFDlykvblg0D6nXD
o2cotTLfZy38EMG2RIM+jK4uTBouhD1Z3UaWyRdETigD2jPWp5ycHb4L1OASjPGz
lZgh/CsrZQOVK7cWQCT1WqydaISuOArHx3Eyk3lN2EYlpvO1ge8DadHVQ0OmAu7q
Yf1mHFPrsc5BoX4iTWfiAP9Y19OQdIq9YqRsY0gCMOw9UEGw3bFMrsqL50MTrrgZ
I/DAnackQFxR9EU5fMpuJvWzqh3Wsslbo/65aQBaeDgFzlt6t/A3Llof4+OvFoCa
BFz3u3H8pixAVjX6eIKLupN3JZU1R387CG2epYEwmiFoyM7VBInka3JcM10dDVlY
P0ShJpuC2+vdgoDtWihhmUGyCIPQQZyH+KR9nb3ttrR8hdmMW4POnfjHf2FrCTIF
21ArQI8M1vz5KcyGBGfnc7vYD1HlgJ3xsWSGOvpchb66w9bmvd3vGLPbRH5/C08z
ZgObzx+h5g/I8GBbPM4YE4dx1Fz0Q4/wMTRj1jBLqe2D5Up/hNx+HhOzZusHblL/
FRx9nw2lXxHAuRFjHrnxlT93qwvaftyfyqzLQq4RLOTwctBzVT6y3xq5QAE1j28P
69VBh9W/OAuwg9VRbFM3pQL+cugTnCnZiotgnV1QijIEwBioqivsMGWdXAMjmsjZ
j6bMu9EtIovi6uSW9wAyH34o+W2A9/BwUiksdKFGUzM6TSXH8d63V2I/TIMvUHzE
lf62OzRF+Tp2LBgoEFROuClemnhSp3zc63etSp8xrslDDXFpk8Sl2Jd2v1n7vCeE
om1rLY/iu9jsOWCqra7S5rjHtCxqP/N1vwdCBybjuK9Db84ZpqPsmz/dCoyDDlJY
W5qvI5HfTy465045EdM7TY9futH/m/eYn58Z/QffWErlFjasi+kaYphhT5YU7UGh
Owvitq7n7AYsT3Un1Mms4r3mWQC9WYx1RSlSgaQSRpBXco0BBfCiO+g41fiQAkAn
y8QGXp7mGJ+4uT8aGnLtFRZnOb5pnpqScq57CVv0sPP5M55o8sS1bmWxRGRwv7u4
bbgJ165NvORgsIg8AGezj8Zn9L7B45oGL1BamkmhwcxDfs0Uq3rbeJzlRppXY9t+
mFz+7Re4uZEuYxEtd8LWJ/1pVT7C4A4H6NQFJ8dGCwjn4Mtp+zC6hFesPkySb8Hm
OYpPJtth+zpG0BNzxwSd72ckvTwq/J4A9ISgMP18EhTnl3tNQ84UNshDLtjxXq9/
Znz9p9DxtXjRMKcNT/pUVNSqVwBV4sQV4h2UufAjEBVBkQlsbWE3OgkUjujDRYRp
XDULLBCM0ceuKDjqxx4rfO3m52mfORJvy+6xUXwayc03tdTDO26lU19l68DcOwW0
Enh49XsfgluDoAKYfRcXhiusBRt7WwsZm+5NfDaxbcbllhei5b9IDuTIHzD/2Fsb
eZbwff5A4npNVMm/8jOgkaTewfPdbgRQepdAtn/rWodzl5+Cpj8TswSdXOPs+POc
39rZi4tzEjKHI4gxwmjHOcKoLwePIxOf8jazkuZ+6ti6t3Cb/LvRCVxv0E62huV5
y+ygkrzadoSJkWhJhv0lY3OKytO6/fzq9HsFUlvLnLf0zqXZ4MGCMkAENWWIdzU/
5s5dlKs2ADlq1MzmKbstqy+hcgrcuHBJiy5bR7ylm7iqKBnv1ehxQh+vaZfRlfUV
mZ4aVONJZLnXyslO5fOmYIOvggamOsUyKbmsjFAMRPo2/imMKHRg6vsva1xxYjCF
rwE6lszKmomtO2bhUkCgsa31QhdtDHdq1j9gwsYK9N2ILIXeVT0XQIiiu4VaaZ6E
oQP2Cl6PoxwMkbmViI0FiUtqG/o1ZZdItUG7+VlFsFColKWYzbcGkAtnIhvE5kdm
28JEGOvwj5WgysrctcSGPHI7aluj5QVRhEqlAs+XKDAXgHlYtZmPGSVt12zCGBmG
A/Msui07r4ZiR0rqJILTBVKiM1MYRhunlnwAGs9ADwbNuwusxJnuTjDmvvan9eHk
TThIPjEYNh0xCOl4+Jqnw/htD+Wj95g8n+GT95hoIJR0FWJviQlMcvTLsTyUjH6+
bQDXjN+efadAR81dIKhiNdK8PdW90pKe7CIZOVSY+8TqxmcZyejZdudMKx5ZQleE
QhUscS5eUP9xWMTuYl3U8ueQw9ha6Cjjlg/KXplHvu2Lo108FhsqZztEEt50ORst
Ne6tnmKae+F9EPrIKdYak4ZpKYbqTCvPQUnHuEn+0VCUi6JUMChZCQJcj8jxpyfM
V6c3E/GNeYYIfqXYWaS4TzzZOKLT2QE+CpeNhGW7znWUPFO4ELGnwCbdr39at9PL
qwdH1/wTToQ7IulH86nEZN37l0zJ5IT0BZo7zicyQuGHeCwrHwOFwZw3i+v/sla9
+qUZyshOXYzd+BKMOkgj8nXCb8nqMMFbJiT2Wv/XyvfIfGBAUi8zXj/My783XGro
KJBkkcD8/EI9iNJyRNGnKKlxfrOsxlsDMjLWKeE2YVFAOaa8qLl4ZPYU4GEizqTk
uJw0fQxLSHMuEVVnT89GEcVJn5QuoSOGc9wDgi1NN/MqADZkOY9+GyEQ8uYZBswz
fxHGBNdDxBVl8drTJUZIito1RUeuUFV5AlIp7c9JUKUktnEerErumHe5wFAKVCrY
Fo1v5Ms7OGEG/91+Hl7L2Vs3/Kdqc41mf/yxShRcQ8tqIMf4OfVTnIP6jKU3D5G/
z0AjXkCZL0sm/ol+Lo3Zb9elkePJ4oauw3soRV55bl66QckzKg+dYptmr5wL+lZn
kL0kXMi0BF/tOZcCR1vnO177wl6lfgIhjsRvRCNvCyvTxN6vxOSEpElDJo4ZrwL4
OJ+RcpUkEVg3XI5MY90Qc10qLDeEcFpidQqqyK2wlqIm98D+zB4aCLOKPPxhdlDi
HGK053Sm3tQuT3JMdAeJdJ2K7/J1S48t6bhBQICaY8VrdsDtUhH6LYSy05Okuqsv
XVo/1HyfC+vNwyQkHOUjGIp3sEFECQqByvGnimIi7Pkg7JAI/J/uOnMxwjk1NJeP
D40I98eMhRl20OWqZRQSTaa1HGg1wjwENe4y7yTE58SnBKfmvOydZvDFSbPvD64i
YP4iiQs4YB7eIk0CYCLa4LqrgR68N6mdz1G1KmFHCj1iaS1tJ+MJXAtfn7zpwjxu
8RmK6Z/nOxO6VOMBB1P1ekJ7Q21+oNZvRqRaZAbF+BUSnbWWe9hblgcyybJRQL0N
SwqqT7Ow16RvePxkrSmeFXbeoyj1WxdBsJInYW5vbw9Re/OjlrYg+AOExNta2Xsb
bQTQHeJ7XUy9Cwsov7+inryquaRdHVTZakDCrgHIp2P5WnD9THsOqguHaWdIlSBI
CAk2493o9p4uTQHbBSk6ShLNRvFsEeaE7+ewYDrMwA1LxLJ0y8zzPiGVXDXdLEDc
kORrQUlM8wzdn7S0eFy51Luex1gV+xcxaOUtkm6Bb1SKBcnLoDQB0P4diiJ8sYOj
nP6trbPrPMYRyk/twFVyfalULhxH2xcx9IuM2a7lCVmIUEgTNXfbPJq3Sv/LXvr9
mNws+N3x/qg9+J1G8cOLonEhr68eb5aDoSzx3glLNK+Qe2bfDGIn9gxEitCatsVc
UOzRI+A2kwPuJ9gJ2eyh4oBaJwkUBOnnI8OUQzU+P9JiuqhGC66wxbZdgw7nS1o6
DLhqWCTiL66l6huEjDsY0518nGt8eGLH4QsU9c+FBc3NASEkJvJCE4YPuR6HNWkQ
Jptjt9tpB3hHy/qliNJgPZOa18nSm8RY474ZGSwKBJCI5lqVBF5RBU67vBzHNkfl
g0QCP+1YJCfN4J+kSTXwaTiDgK3heb0Vhnz5b1gRe22BGEkHmlSkVuYgW4l6/quC
NTsOyPfLeCS56GzoK2xy/YUiw/klXYgdoC+ceV9cArqGUa2CJ0FBuz09z7ThFUO9
9fhwT0Eg8mb1voX2F5nDNcsAMrQfyBkMbXs5swTh1Ru6pA530g4tsOGpPt6BI+88
8QSpud+VPQFaKdoyVXTcSmnu3EsktMMtA+0sjsT8sz/uYoOis5++e3JVCCk+00KS
KyXo+d7hB6jdT3viuIHzlR3f02oVIZ2+KDJQyI5XfCK00W4w70Vs2ABKYcYEFiNR
KhQLZ+QyW1aEvj5IFzeTCpX/qedRUO0ZZ6S6uu9wQPBrtTHyuGgJRUfoccSqJ7Ef
mCVtH0ZBYIo76s1YUkaGzMVM3qfUBnpADlGI+Nmz2tWX88+0yXavymZWKN3ERWO0
sKeLnW42jQAYAmkXkVvckZX3kp55rM/Ul+oSoZPqo8Gm9sB/WMH0n074WJBE0p3K
nW0OQ+VRU0vdOePyt7ZEs6OUGF/Q+i5zULRQ1jxowPXV3CZ/c9njxn22lW5BNjb8
st02PuNJNtEE8j3b/ZXmQehOicbMZZBn1K3uiu5q6HICb6urTRU9MfL+bv2pD/Tj
VnUS9zrY34nYeXNM3KxM7dh5YHmkZo3OejALgNAa8fOndbFbhv3/9i0F45tT7eXe
b31WpO4fsva4pWoui9wqrMuEzQWBxEHwZBRGnMerEZ87GF0JIpPMyLw5GXu7aS9f
OikGv1ZaqqN/tUplSwbF5dt2Hj+GqpeMAf6qqVhLyoJ+prrlz7Q9QD5QSOdi536s
40QSw2BNlJ6ROFVGjnFUn1DAI4JSiDbEZgtUWBrgB5s/lepsK6pqsnYssB7Ai1E8
pGxFEpRF+nU2IJPbjhIFS2N2uJLueSvhHZjxFxs3HrIKxLEFVkayhSiDCS8Yf9Tg
mDFnllcFMq+OjPVUDOvX8Xs80GXkm177vutR7IfT2POxC/7eK3Qw1kmFDJE5ye0c
A2kJLkdOmWobHA75BKhsmWUQECgJ9NgBrt5YmAr/K4ly7DIhQmWrcZsLR2zskxR4
lqXnLf71qcTvIBOvTIIGJ5pjdsXMhe1fDQGYAeXHpc+K9peu68wuIUWRLXxG4Bh3
dlOI+iwwD337wA4UVo9QGebdXeWNIXWM1omO7WW+w2BruD0BL4eTK1tiZjzzdfe8
I7AJcElRzpuEPYchhg4mT6TrueayDbEzwt/qP57NbDbNiPWsEtqyE7VSG1+AoXQw
mHEtQIoB+zB0/E/KgOVFpQ0+LJ0OeDtgfCi7/y+/qcl3zKZt5OqCKfVDWi9RC4Ra
3NkaSftnE5u9tsRqKRz/C2d0BCwN5iy5tFUmkQ+NWfPtdse5lCmzj92wSVRfRO9i
GeNegCjNDxYjmAUDVyP6rao4Q8DaozGElHKjde0rPOPrHsSqKPumXpLYcbdT55cb
NzPluAdqhcYVHrB51gzH95j9WtZS/DKnO3F/276t0bkxZCS6tMJSIULK4NmoNqiM
gEPmAKR0kl4ho43LALc1YlWVGv3dKhjP8ur1xkpi+6lis/hNOTPzgu+bS0/zAoyD
niGU0RhvsJqEbkI61BScc+jUpWgqfYFQK/0kTHbIvDeqp/riyxzr/+q44Pj/nxSE
a5WDor9DfcNbie8L6pbdqhUU4SaJHtSDKocO0BW9xgGcPoK2Ash93NErq3fol/7N
hGplNYHByzDg7s+gLP0UsZ/rGgfItZTtMI6Ate5ccScjBTl6NmbIcTb2JJvqMx8m
Vgh0ftDRvP7mG76/UiNEUULi0blAkwWMxbt0gR1zofGK95XOnlTt+7WXTxHna5Vy
de7z6bweCt/FB3u7fjh83iKisw4K8koGwmF1fiF5xJCMkCtutrzl9yikQrWNp/j7
qBxCWLvUOjwTrlOXZhJgPLppy+3bY6fwh/bovixbp1EFW5jUt8A+dE8wXkdblYU2
qDrWuQxufQcm2RpIcffxS4iRMG4zKLvXntMFMZo/JHBC0fVUpPH78k8mwLR3O2NH
+Y7Xf1bo6reUs6eG5kSGFdzjXaVPnbODW8CynxgKFMZ+u9e3h54ASO8NSZ+TYQTz
ly/94SdCYvMWoe7V11D2B8wldD5XHKfDqS73N5wkcEprQPI9W5yY/lVDtSScJnIU
nRlN4f71TAgyhge1DfiOygbXFRudLZopMqtqo82qbm9fFdj7k0vcdpzhIscN6NW7
vsthacX9u03u1U2PyAcF3cn8gGazzngVxcU1pwC7a3cUzRKmbOosBmc/Qn69ABzb
OEu6Ps9V+4I7N22sndHbNNEMpi83uUmcgX04a7oSzMfjcNLVd/xmCVKYW3wn7GN/
tbRuF8VOOp6AmBxpydDIPAJFYOhoUaG6g2jsxT4OG/DiY8X9nZ4/agj4vl2EebDL
/UjG+F4Z4Jkvbpo842DYyIdr7y0c493/dCWWNfsAF06PsCPNA06ieX0lsuP9b1W7
mDLsWbkC2cOmHXj5jZumFViUf+uRuGvH6xMXQv9D+ZsBCQLZzYbgNCNbMUQcYk9S
C9odu/CSUa7aCCch/2mFeSccSANT7mBZ/1K6u4RpMVFvp9CnF2wXp/dd5uJeX+wY
GgQQVTyCl8du7fc8p0XmhH1fmYU+LLXgY/WsuWQqUp/XU/mucSvUB+TkSDW1zHfH
ShoHyBF+st9Mu1H3cL4CSC6rAo88IOJKrN9sol9YtlVPh2hKRP5nhy1Jvo02/xDP
GzCM6DcbrQS+xKC5d3QcYf8hjsc8b7FULtGsDEvxRCffah+trpBlQ1sx22Th0hzI
YLHBwawbjrzfVgG5cfjMjyRT1eloUDa7NrK+WFHzI8XQvaf3F+RJZAHUvBKSGtec
gPIjWGEdkUr/ov4pn8WPAZOMZYbBiXgx7Tz713Gwb8U=
--pragma protect end_data_block
--pragma protect digest_block
efhYYiTG0QAAWD5wJOszcvA504k=
--pragma protect end_digest_block
--pragma protect end_protected
