-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
n2m8c51C8gjLJ1mmXUYPY5lByxOxJumpq+/A9ZFyROQ7UdV/+GBFY1+lghFY808I
Rr1Nzr7S0uSRz6Aw/eMdydkRJ9RxEU6f8cnWp5neMQiclMMw5R9r3J76QZIMGn2q
rdKw1JK4lX5X8RWT7MQiYAr4LCWVv0fBBp5JH2PRffk=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5664)
`protect data_block
z7CuK+N0+dp487jtJnQOFo9ybrA6WKOZM8PX7a+Ikwsr/264/FU6ooXC2zBtMByc
4eb4TYbkW+wBqlV86mAREC8V4EyAtxO9LqKhYeNaQ8zkB47v+fhBIAm9fIdURvau
PPBs84y8IZe+7OsXkVFAQXesD0KSRbLVPFgfDMl9hMqoJxVTA09qQh2+39Po5OTu
olt4uLKnxsWvclT/yTsafvjA/powoZZx5HA5TDSVPMlQ5/IfgfPN3Ksxr3/J/mLc
Vk/g+7gzpSOyQiC4fITazFM1B0vKY/vOEGDQjhKCeuPU1uErD2V5ZFlWGESp+eyb
3ygAkvGvWAI6M3Pyand/byCfCuUqYbqGY8BZa1zbgvcAKExn3jCIuyV2cUv/tXl1
Jpp/K5iK8fhFDbdt07WxgxJUwkfhblw4TkfFkwfvyWoUWQJOKYSUxFYQce6cu3rS
4plL5PR69ig4VXQP25i/gFaPjpBngdXxRpNTPNMIAd90tPK7VqYNKnbANLLkJsoA
u2i+H4JvXl8iLW9oNNyEscEin8MVjpI0s5F9Jk50pKZmhFesUmxXc2BMsp37y2qV
IBrHct8+UM84R/6YtDVDtJe5fAFtCRZEnlB49Ro4r7wbilMJ3EMiEbLjAYhbQMNU
/IoY73jFSJPcpvqb1BGQr5Y7vBr6Sp/aehSoPiKwiG9j63UYSRPdPomv6cDtnkqY
g7HpcoCpfy9UEj7WAzhnQdwWJ/BfY1FXlaiM25tMJSkNkPp3hht8MAV+34FwKfob
l1gHDzZN8K3cL/3x6q7o6w5ScI7l10rWb3RV8ZZd59+/D6gGotRGrOLdFYeJzqWt
H1zWT3nXR5T6EZ0ROqWw2l0YLIyFE+JXu8eHo85SqXgYjwwl46t4ha2fv7Jv1fRT
jz/J/3QyXfSDFF4KvBF3eWrJJ+X5Z3OoPnf8Xb//kV/Mwc1W7hQmrgT5IkcOm9bv
7/zZUx+ILz5tZwOPXhFU4dqgHmWdSErEUOhByrI+zRoXJES7AAE3Aiw3Nd1Jy7O0
1uCy3Mtcm4KmwDtgZGloNrE5U5SULOXyh56MPzxHWsFX7Jmj1zAiShEwWRkbXfKG
vM4svUOB9p/i/H8sVC103GouGPI7o2ZsE56mWSxouSulxaQ7vUi/5zhgfoL8YYZw
wBSvOopufaB4KahBrVSnA96PgUW3EEyTl57OX+iDWBUynRl0dXuTv2L+gQrdbaax
u92o6kcfVtLh7Kdkb/4mFPQLyG4/+n+HG3WsnKdh2c1vYRx1+xSNTPnhCg5JA3oO
n7dnhCyH4dD7u6Rbhr20UL0+giTocWmmV13TPDb7kzhki+XAQaBd5PK5SsOcqYFd
RG/IwIAOtDEx8NBZhbjvq6J7Gn4/eTgbpiNTcQa1FrHlZlGDPY6INFXFAk1A+mbb
g8fN4aALq8dZk8XPBOmQUrY+s7zQyfkvsahXpGBXXnt+rMCfTm6oUNtoX8+2N3bv
5UPpkNF+D3aOLrXJBvBMT7VtzWve2oZBWhltYmANNG78gqg0e9qxZMhWrnE136yZ
TYEGKrVYXwUoJ2SO7NqIs3Q4UALIx0nvb40M420DTbPIIeikB7yXBenIZrCb2y0o
dvYz52yz2Wu+rFgak1NsczaeHEwqthXlfUh5iv4yeaNT0hEuQzHqlv/Ca8qsV8x8
mDTdVo3/lwG9qvGsF4gIy+vfeRIV3Hhe3AZQ+oy9dvNWjYJz71NIEu6TPs850Q0y
u5bbjJg0ohMsDFnnBQRqwBFZrsEqU/PxFARbw6VSZeTKnkloXX+I0SVVazOi1FFH
qVJOdJvijoMvEIY+6EFzh7rH/GE91wMUNHPdN5e+LDYWqgwiX3j6wQGR3x+KiABv
u/96zw1UGgt6rE3LXKerJw1awiFuGUAeTXfApHfaLgtMf8Q3OadLqdupKSrIFesj
aYWr9M5OLFwKx7F4mnD7fgOMIFaPVqsRdr3RyNgQU+2z2mPfrEzKzn1cvLjBHxY2
8QX6Ps1FlAmZL8d7p4yF5RqlxFGy2mbg44RFDc+04uC7Ul6JitbH+Rb0509TkhOr
mAJtlRmosoGv0XWvCza/yGfjmj08esz7ChdROfM7E5txyYS59r5HGNGfWMOD2VVw
wNFP+iNd21M91Tx2BMYe2HxZuXe241wfgT9PCB04bdwAxR3HS+I595iC0z+Ju03E
f4Q5SgoN28DNknZr3Rfa/nxvanqdNSVexlgtBUklSxdcF+G9lehPbdK3tIxlRobu
khjArgqzEpysDVJRWqyD+M3+/NRxT6UC7XvhxdldkGiaJCJr4NccGrJB6cyaa0gw
NeKt4PCG/NP/vvD+PKEe+XGp43wlwoN9PuVTxq/lg3bM1E8Nl2636MJV3HifYHcE
AruZfRcShKQGjCiSEePu4ho4T4zI3aDzCXuhLpArMyio3lIH7JWsgOfPiw+F6DfM
guwM6c4n98TkfVyTRpxkrB0qj5ypjjXQuG9gfuJFG/gdG3PSKKFaQpwmrN3MxB/9
2lQMaNBbni3CgBKmiUZQTiD/gQ7gkBwR1ibxcn5LuDwRU+Ub4Nm5ld0yE0tTIkBc
E/cVzqD+xKHB/QwIheSM2CUOD+fj3j/eJjkKMf5rPTaKkV0J7CGJvxZz3Ejwcuxq
npCnwIovTo7UYZmWudFEe4wfChYghnvB3rvNjyushVssHPM2oGmC7xQiQEXHINGG
NHZ4WYiGMZwTMHWQT938q6ZtA24v5G+EOQH9q9GmiaaZiZaC+XXRDUd3ObUR4OEx
tSBCnFNEvrRkS4WFJfMSRyB9M2YQDi2n18CUzV5crVlC6CFL1HfdGPCqAmCQlvgk
znAngOOlUpmMT0z9WbmhdQeX+i8OQ8mSRuEWmlFwrnYczR5ycMfn6z+1M1+/lgFO
XsATDSdDBaWml0T3TM6RNtlV5hz/O6L52c/WmbjornCGaO5KD4+JQKYOr/lJcaGx
Vl+kjrLkCtamX9w++sDy3rrb1EwxlTs1Ir9Dlvl8sYeo1BX1c0FxMQ3dk7jzvkPE
clBWqN5rFa5ZwCp6KfhJmFGd5jVFNg0mNP9rwG5SGP113qAdr9u7T538Shb35oxF
vX2XQz9OQYk/1+RFSBzmL6u2o/ioZyCCXo43IHjV4I347qG+InO/KUCQHa8Yfnaa
mi6sXokTEhAnhaPYgzl3MQEMZl9BK9nrK6yGA8vzCRoZ/eo6UKfzzw9EOqvOPXdl
XrgBiWhVE/JUsOQyUSdlRXgQy6ladiZHYGCd66C8ff3eQ/NfQqBcHz+UHHz7Yu+I
zEW9MXQVKq72rzqrJpFc5xbYEkHe4KbXhdoOyLxy1o9aHUUvvppM6wKSHGvz8QMG
VnpMv3e0K9r+QlJ6TU6RRc/dFyLwsgHyYgDXsAp0Eg1dxO9AYYSyQy+/1/tpyP16
iKU5jWNglAGu5VsKhEvQ0/164+5RASY/4Qrmh/1eq4tDB6DwBJfyxx9uX+BCppky
1+Bu8QxrsaUPozcrqOBTyuLiDF0/HdpcoaQjpeI4RMzraVEzcdy62LZvM2VslsfP
z6E7yNU/SQmCGRxX7X9MDl1aY6VmeAFQdgDI95vKcdBj79nDRE1TIMva015f/CTj
CqMB9UUlDxEgr2dP2rroVNFVZ3/M26BAl5AuhvCKQON4QAC71SKHGa4V0shv5L1/
0bNWQ2NsFJxGVo/L8dhaRSKH/2Y9Wne/cmy8UOr0eXqBt29UKcEPZxOx+d+IYBm5
vMlT5MfMHul341pLGydMpYc4LqbJL/4iC+T2WMpTo1kabPqMkevb1TPTxetckQGL
LK0hO0v2P6j7x3VCniVhk7qmQ03G47u5HG7gFJyoXKvHzZmZxlGXfbhQIiw37f/P
bgsFqANzVyy9bfSErV+u8xzIpLjbk5Za3ibPxTgnzSEHB8gMfHOUTrFkVUCPmU7H
vcke4miUelZaH4Ze4IqBuQZBNx4fGhC505W1CXk9tJ+WLiU3/aV69qg/yLjQogDs
I7BZryl2II70aUlxQDbtXT7ZcHsIIFrlut9YTD0Svwg+4cKix5FjiLxixu9zPe8h
OrhKfOAaqVNOOcaxw7FppBw5KcnIl28URmJVnoNf/2NEllr+QqE9Frg9Aoj1F4UV
uker4hgz0iSI6In6f6p/7p8h9Hbp+GkHZdJrS/qLqUt2/DqIpmsI5qr6xg5hVVhM
f9qX3ElxNgTo7kd11oTuAmQlCOL2zZLJLtcjdoBPdz58+47LZAK8oLtsdmmZrjGj
X0oiaFwsMsIZ71UgZ6I4XS55ZLHNAKuJ/7o+DjLZCHZJlf+E3aIzAPg/YsJlr+ay
ZU1iENt8UzaE2F8zcYQ7a+Cxnk7+UU0NxaFCy6wa3ZG4TquxkRl5OqaEEMM9n5oX
zrF8lf8TlmaA1sep2Yj7tQEgtNzF39nKa8+Q4V4loauBoEDrMf3EpPOEoVN+WMjk
sG1v2GaGj4Im+iRE7eOsCy9whyKoPf1TmuBIUreD5C22MIiKBF7wZFJ+IjE9QeCp
ekmEJq1XTWWXZYw3QFGc1+f/CxRBL31Z/neu7RM5adeXyxyROrKszRU9qr42oX1r
JWhmYNLOXVPr6kQbKEaKy8vS3TnATSE7oAaxXPihz4nOi9KoVeUpr6m6ycBKBwAL
LTBh9uDMyVRcS0/TXgkbGz7PNf/qh/961hg41KRXbKM0uETM+MYJx8Jm0htI7pud
A4c2e5RlqrQGW8xyuPHwhPpIS+vfdY5r460O6Y6FkVhG55l/J5iqVIB2TN0cZyyo
z2rVjq192F24FisBcvhRTauqZ8ZOFds3CmEjJ9B85MrPuTb/ic3a5YM00ge97q+I
dfnuGjtQqA6YwPXZ9L4rI5nuPabQlWCRcifwVp/u2ruzx2IFPXh5qwctlerPYrjm
Np7uqsuhP6bJDjLEoOmpREDU8Ntx/xNbftNfuIEIUrqHvh5vvNyrSOdULAhssii1
D3E/KvF1PeB8K/PQ46rDLfGuXrtH0O1SnFlgID96vRN6u1nsEbqDHK5vOB2XTP81
Mi1ZaraOBarwjLL99k4XfQPCGwhZwtwdKXLRmpPGuuhRCd0+c/9CD0p4ookTj3MP
vi5HTErO0CCZer6n4ICtac+N9fcMuLPpsPXusrI6NXrzowiVTVBoxYRfIT1YwdUF
LvCAVKD0b3xpzxYYKSbxk6L8/zekIQvgbhmMaE0NlDFe6Fg4SQK3YIpaiYIRe2LO
dfrd85ofmt2eumgWalsNwTcpxnwbnZKTfJFJBvNYJh3I1vcuri5nECLr4JROk3Xq
rXM64EoeG61w9O9YSKoj3YvOTPq68OJArL5KrchdDzsetUXbPqla7tlBNjkHJgWB
rYfDT0Ttws2wUyx01sqwnQLrIe0+s3LSu2rz6JU6oQD+1/9xHsgYmx3veVVdvNq8
NfHukcQWw7VljJo3rwQJ2kIoGKUpi18Ch/VZSAj4WxBjBPx5QdZ8mtiiHJGiGDuC
BF60TDH4XRS219FogxT6u792Kc+T9IV7B2lzugtGiEpBND7ytkDlA01l62IWeDmp
Gd4GCnXPBjAWW6C93RlMoSBDEfbtaaFJ70pCiFsdWHmjuIVKG2IjSD/jIjV2udMy
CIKXWfgftV22VuvDE3SiVvK25HwxCBt4xIuahRQBjADDzlw/o0c3h+VWM3VuqxYz
tm8372/bx0lcQyHby08lgbjigzAUm47srR/zezHToNep1qmrE7vIkJrlnhiOgkGJ
SyZycnbxF7gYkcqTksRqTaiE9jXIfUKJhliAbXOEAUdUCjfGJhfA/TeiDuZEfml2
KhurzAn3rPtsjMZCAOt1IjfetwNS/CMb+xEHngHFTQjvimxz4H/Fb5J6ECexBIqg
gJ1WQ5hZUGfIBwHOVuPOcrsbq8QfCo7KfGSNumd8M1difDQx+z/73qatSdB/ft+H
fFzmgUJFQzNjFR9J0qrz0FVAG0rGv50yUWMlLnkaweDb2CvVMm9tQ909i504Px4y
4yxImPDHdXfsgO7Ii8ryV38kKKJzrOBUK1gHDS0DVKqS47b2Hor2yn1KAq/xN3yP
IRpPzmUFjqTQ3JOld28A8HIPEFAsBOJubwCqU3VE4mPzULNlzYLTnJIO6of0Coez
zfxY8rzaxTFVi6OWUHJdNaCV1XLdaDymfCXDQxh2CP9aP3bUw69ao/t1z5/m3d17
FYn4KBGmOjp9v7V2rdEp3NCjaBrBW5jNuEtaPUKByYic6+QXPfOObRI6PeVi75sR
3YWymjlFG1SeWNWEFCNzk0od6z3EbqFScIBmccOkzyBPjnGbjIU+Lu6jQ2TYnOOX
jG3LkKzLaAEBGTqPFu8aTVgGwJY/WBZgLaIbNfpF4otSiFMK9/nXuK49jWLFEO4g
rOwYm4M72ZHofXmdSLfn6rfhqs3Z95Ihsa4RADudfoa+/G6+GtkD1PK3NT3mO8B5
SToT0tbEd9FIw7LQhJtMJAqX6J50R2d/NoUEKtomT3/ljbePBJpl0vsQVIUJ9T25
NNrjL3zYDJTA2NauzCjJ+n9+1k13VVPkoavGaKYgip0biqzT9+ykUaYkqi4XLFK/
/ycl3SBYUb5OU2riZoqNtM4bEdxdZOa462mnZSlXKnvDn/HGrjIatQ3xdygI8HjF
1Gpa9/Bzsmdpshd6IZiwIWpLbANkqOFVGqhBVP7LJ/XKT5U88Bn8TnYF5Q8/Pwq3
0869XlYFrXN041+McS4gVnKoT8iq6H3nz9KoAO5B1O0x9XA+lOFFWSAJC7TbpDCX
Zz7pgQeMi2YnFp4BvGouLlQEJvgPRA1wbJKhG1+U0SVZTdC1NMEJiq6yCpgb4JJd
CepiHnyjhiS8cKsRbY7XDQNtctZ0OuU26w7YuRPuR7XZRyZMnUa+qJjxOV4XsT/w
OQQLtWY/Jrd+rZ7GpFhOZqckSSJlKWhp21SSlK2azaOS5lToWu+OWEKdVUyFV213
XjxBj2TljTbIGDMfisfRYrSAYuHwEJLnNWlGt1CT8ofHVKjOwQtam6NzyhfBPe5f
u5KW8l2lNq2yK9nvNikBOBPHyl/qQVayZBuBiRl0jmOhB5HlnxDZvpP/RZa3JgL1
L5Bx0KrSxJ7k/FFuQJllRKHMEJ3APdLakJ6PMWyeMTKl03RFlSJwqVeUkFPohLUs
N2HSH6LR/4Qp+c/q4zmlPOgHEwma/0UgihpCX3ApcJQG31jGUXdOtcye2DNfZ08+
agpHVsWiLmEKkS76ZhvUQdv80d3iHW2LYnd34rFdcEvga5Hl8ffit3d55mnPErGv
ACqQGAttNd5PPKNZacp/snQVM4U9hgXECp2Zfvu5EZ1pvlYJMBSkE47a4KTD9XrE
I8fLJzY841Wn3cXXW8OSA7sCcJSYy2k/9ppwGrEnoaXeByGB2/5FaPsTLiDTgEmH
xuh0FdcznrP7OYA7iulJgcHr/QoLcnSJ5oJt1yeu48xsX8FVK9HcK2qu6iH2WwjV
JEeHA3e2f6kJBtSTqa5dCaTYqGHqvKH5eUHGGWXEWuAp5IU5M40f6Zn2H5QpRUaM
Pw6kG7zwbGpvqtrmT9NMIbqnAgqEmu9C+tmlBnQmOhPQ298SbZdKeb74HElFnA7X
`protect end_protected
