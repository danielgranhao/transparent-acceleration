-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Dh8GWtIMSoBncQ/7K3zwUv1wbv7k21l+WNJqWlHgbUFK6uVB/lpYxCJnOsyiWu9w
SQRLRGoMnZxb4roZA+vHQ8Z58LJXN4fv6ZPvS4Gf/cbL9c/BQ5KWez5FS5z5nL66
yftnslrVu3xnXjcoyZhc1b6y35HGVESzHo8f2QDc+H32Y7w/tdRj2w==
--pragma protect end_key_block
--pragma protect digest_block
BQmYy3daOUojOd3MYRGSNUIDcpY=
--pragma protect end_digest_block
--pragma protect data_block
pLc9IoH630i+WhFWtyit1Ud6yf3yUtMEHzhanfSWYoTo8hhyrJjG9BnTSX3Iael9
Fj8011gbIKYEOhusGgrPokUVldWQLD2NCH3AszOtyl5f1xd7gAajO82mdgKUi6Ar
+EvWJMnAu9oLPltPgHfRa9potqGjtgjslt7OkeM57BKxkYgWRRRXwFBSXNkA1ez8
7UGPwLQN0Wi18aCSPMBZGoAJ+4gZ+mDYe+Wov+jsNSimscLFU6lmMjEU2BZCOV7r
0/2WNOFXXkemxxYz2MFPM4zbtnQqcFhxg2pIletSpZWJOdTZcJiCzK5eW2UXROW+
STS4yRRO4LpsED1VhU08KyIV/6QoZUx9yJJM8gZrXLB9IkilQ44KJ1/A8iN2llvi
lqbMqB/X0H3vU6hYjUP0MxXveOhctcSFXi3X4JHREpjez3IFHZSQ40dgjjBPhUc1
pyXG4BpM+kb03jJeJbJGnlY/lIjl4wWsj5Fo1HTzceFbyjx5hJ8bcAHHZjS3b1wW
D4/lbDYTo/EZllGPGJy37387eFHOG9I9zoKMd0JMLgjdRsZLmYrY6j71XJiS0C1/
0ARFTwgiGuZpQkEinlbRQsdncrx1+Jrq+ziaWB14euwKOEAxTezZF7Spm6/GOP0h
Xh/jP9BCE+CR0mMaW/fG4GLbJ6cZGJyPWSpQKDJR0n+oBKVsIbT8rVgRjeLcDlJe
flA9eE2azMgTJENvH2JpppeZoAAb5mWZX1lNYWvW5pOeRQWWY5T5vmaf2IT1CTSB
AR24nHFOyrVsg4fz7PH/obN7+NJMQ0aBAjCcKLMAEWZC5QxHPeY7SIjwOCJcyCcy
H1yfKDprxqXH1pbtb2pWYyBvt9zWU1y5wa/fqIIouB68omgioUZfgBqt0RwsDrbl
XEBtDjyQcq9fMOpR9kvQ7bcUvZh/YlKYVqEX47Fl3rMFzAt7IaXl31U/1Zq+1guh
LGWqeQwg6GmD7vHzp3SyvgKirNC/7zv2NV2vc9+dLndDy78DidYNowttJ6ijMiWU
cGV4SKWxTusnmhjssM/wOFrvy6GVk54t52+zgf3YW4pSFAm6mnt0/+9anxDDaz8Y
j/Qj7LQPxmhR0/tTmverAMJ501YAbYz3FAmHvLyvnQbQBpTWg1etBxaTPwXQi0SZ
EZbDdu+fOr2syHCFIEjuTJaYfCkVcFjf5dcymdxeMPzrHGlDjsv33HHN75jTDUOI
Kdctz5YlUEb536bh52gh4Af8+f9pJs7CG0ubcza6ecCTo3Io1hLhjg1tYdKUFus7
RbNA0OH4pCdVFpoR3YQ4G5jULfZ9NJWoroUkAssPVHnkKOfxsuJUIxFjm8QiYOX8
PZ6bkx/9KnC/jiuR3bikXp6rk0KdWt3C7iZQUqWvmutsctr+tTMhmGwLqYiIpFOe
Vn0KGoDlLU4k23fnjB3H247ct3jgcRWiFtvFNhNqFwXa1RghmviDj0ZzWJLTGByX
02EjmkLSlvjOKuryGE18VOm6xR9FrC7AJc3t6KOW3d7S6bh+U0y6HilpGUElIO8J
I8J+AYQVExOL/1D3/mNfTSqxvwqUntCGALAJmjWEOhNxLBw9gdQn4c22e9IhNhq6
OOaUDDrjV0MzYiY06+PZInXsrRxXljwCGYNabGMQj0SbcGj+UAW3zWmIC66tRiEu
18Q9gGb/I/gliwiuNexmr4s98RD7kw0RGh+HonBoCbZs4M2r/8WWU+WiV8Lojwmq
woLa01Mf8qa/bxmmAYReqWooobZsdh1xdyCcxRaWhYOwwLwza9E71232+QUNLbXi
oU7N4N7U1yApkSBC/dSqsLfV9125wPE7GxexnKO18oFP+xBg/I37zOGnKjaPkyFZ
gBLikWZMmrpYsEvwg/wfJRN9gKuxglpi6oZTYckBwBclWWKA7OmziDWesJzn6FHx
sKFQMgBKKeW35E7r2Q4clPdHuM2UjiL2qSUES0h3AVo2IN7SHg1WDYE156MDtGrC
iIqGx0o0lMHX1lVZ92Ry3R4IWSiX9+BYpkQnCCnE/YdrIHk2Ej5bsHA6aUsFt7o/
n5BaF0q7CSHfzB2QeprlgeJONNzLXpI390NTXEDa5zBHC4pPwwMyaBt4cXPRAhPN
BHYO85swQwzBygC+0orS1TIiVQkwLixGOuuFTKCCLh5CUNndF+fg8Z7eaddnrd3Y
gFqPUQhje42UyjJf1cNf4QWwBtsV28Bgycoj4gzv6CzY/20uie2ESzWY2TBL/Bj9
YIUxklE+NRHOGnnkVYQ+3vIay7N40a1/oIFvCS6QGC0iJ/Kdx8516dBU++lyMu6m
ouA0iAgQ7Q7JQTYB30sxTTwOnRj/eBtkvPni3+W8cQTEsKEosuxPulMQDHodlSSH
93Ze+NRj/Gt2gfu8UciAN101Q1ljBK6awhhdCfrTO5PRB9/dgWdYVihJ10zbvi20
x6sCqjGJOJ43rETp+GjIiXYkseODbxDgbtFaYsYNOt7w2h6VC/7eojD8PKtRYthU
H4Oxx0oabYuCgIG/KghD8tCc8oBUnWovT5Hz7QYnk/DBlcFx3lvpaXDzSGx2I4jW
rVyVQfSpR4Wnf36EcQWcXDwwEaSjGt5NLg7Su8VvL8esXTgeG4D7PVBrAWFM2Cun
6vmldnalqyG8/oCzEiPUOgbrAmxJtZY1UjzfUnDB8sMCh02AdNIfuRKFAkdyTV1U
WNQl3dG4n9cWHbFHvbdYtUGZk9DZe5wt+c/e5PYAjOrLDuqE6ItVK5m4p+u0ibfV
hRZ8cakGdUXtiUQoNd1dCBZ69A4LdM1z5Va/r6zEkUJldi8pillNSypX9pmxJ7zH
PHiH6Mls2D24+B5M/oGnpxN3BwXQHjz5+M50S7225rOLf/ngpRatLkQSXmBfeDs6
/xhQ9tajFmtcfnHq+5UjxLeIGcJNSO1eAs1CCPaXb6RgsgPXnmMT6wZz08Hiz1a7
vJJKItcL2H0o/waOx2YuyOBLeXopVk9BQ1XpVMHBzHkP1Kg7qx5uVENQfsyMecaH
6OlJ9USj+flU9nqCIPEWMxJxkcQF9YAwHYIgy7k5rTuem+wMglurzN9KFNmFxWq3
WBgiDviyARA0OXnDagwGl0/QKRaevACbmQl/OMycFoFGkNPrL2Uk1MxfJT3zs7oG
vsqum/tQs+Xq0S1mNribYQuCEQQ3kGRMd05VvG0peDeLeGlTqAlSvlBwAPGcMNvK
3PRVCk05C4ngmdK1l7NfVkQsSayuFB1hOK1cWsl+auL8i6w5HvMH1x8hP6ZXs7Cr
QOpDvFMrbeOhKs/of7TWrF+3PAccfs2xhc0mtREWi/DwJ/JzYSJYxXha0h1sr2bP
OHZQjTbjtyMPdYfVMDHBy1XGerKIbFPqS1B868QODbtBLTAwWcycfpEf7wkOQvwF
xIvEuftmQ63g1Z/EufrKqTtJF/Y/bdPePumYggAML7sRJ7Ypea5LcAA24qxpkvlj
N2Nd/xbwIZ4E2Q0I3gsqdePAo1LDTcVJVHzKetYBibFpjCtlB85luOl50M+lbrII
vHhyfr2kQGhgcQjCFAPsewaedztbpr4MXd+lnwHFowAkm5ECDh6NcGqopgDXWzPJ
zlOxAgvYNiHYbObPnUXRPF+7h4pzKnY+nkMlzFMSkggkDzlVSOcb9pGX6UoTPh27
HNzpazTDBFZo3WWafkU6+jZObIb759qB/Z+QJzF1by80iWa+ZXm0uoz/BXxURKTO
7A6mKnO1FfGihP+bG8GwB2nDxxMsqod+Z8wG1lS26lDaTWPZEtTa0xTl9t80EQQ+
Plmlg5ArEPiZoKxaDXZEEGWsN7Mkz/KCw+30y3onNo3tJaNxrtEk5Eorj19VxMi9
Jq0aSXEmqolD1nRIbxl/lFUA07C99rAZ81sZc3+fcE51UdY1C+7Ut5vWVC583+4r
bDY41Nz0BJN3IN2SHj1OMR1hzL5Pl2Znj0WAHUOxEzcJCs/o3S/ICeWvQXHhTYjf
EkvoMvMV5RKRLPr+/QvsD+iPC84ghJL+agdukq6Cn5CCv7ZcAdGNNs+tUq4/SRhF
i1xfC5ut5R7o7uDqOQRZcVUbpDLIQaYQ0GGFyyHdFASWtkoJb24ULZhRJssGlsiz
uYb87IPu9R3F3jRaClyJ1pwrBEVoEqpOQyPE6o96rDu4Dm9lQkhcyFQIIxo3svil
hN7JjxdIhOMwsKGr9rOGzDAZpwuYTC0Hj8rz360BXabZPYJN/gzAnnYAnYwwyZgx
uTe/UNyLOO+Zc8+fRIHm8DTPKMFg6ipW2WS8tcs+GRxn+DN0zbWfqWncEcpChrru
d4Wy7/C/SsoB4DVsQdoFE2+fKCueo0wuQO4DIv+j3tyBsdEmNzaB4nhTw44m6fhP
LnxhBp5eyV0FS/3UxeQpngZGRUz5tiO+1jWA2N11BS/4e+BEd6ehtn70OiQox3Hz
SzqoM+w9PnMi5Nn9axbsvZrzcgNpYk0sIUeKJ5nLogUDmrDIWQ9oJoKUVtB3C6RO
ZORQ0VFGKcNjwn9LTtKJFbI9v9Kxs8ks+fY9F7GUd12xmgJ0NVJk7iuq13vjhkSQ
wBNvWfHxKyMy7w4aJ12FXU50WWXSk9MRTSMq8vC4mtr09FdjbHDIZE/IVXKbt0Pr
Pf+G1Nm1m/gP/uUE8yGQ5tu0bUYIwccE4TOXKKflGOcIQ1Wm4vXE/VCu0lswXRsw
1cViVBujXCeJQkqRK8tAS7GGMnev+T2EWhTgjT7Q4iUUpXPCg4d2uLfH+qExBvdu
gnl67gos7/vVuTcmXC4x4Ol5D32XY6EuQNyOPCh1OkEeWTE/7bI28PiwW74dTJ4p
ciS31dAEDmv38pVwQO63mtf5c2dOGIilFIF4jEYM5Xd7Ghhhhnwv++itRFFOGsFf
kLdb6ACYFP4wQ3XgXhxl9bdGJcoakY7ZCdh4ib+r6GXKg3Aij3I+60/GVDv8/O4d
+HilT5tZknkhGLrTgV4bSEPbyvJkg7T4s4llJnuaUu1IFxBtV1k20ixyIcj+JN9W
e/heMj+LpTWWhK24Bs6XMcHDUM7YiIBMwOM7pSO6erVL6d/sKU3L1vKpeL0K5Tns
4AISlVarnJqIADebmS9Ys94WoFvq3r2ZXeMfNYcnm6H1zc+arSbPR9w33P1Kzi8K
umkJ2Kt3xR2GXLL1RU+ibDSvoM7T20cPou7PnzvtoNa0Tcyb3EEaRbVxZlCNniln
oyilePQyCWWYZzeqPfGaQe8VOgb3/VovOrhp1aMQw3JuQ9e6PTLyrNjTzTCDEJgK
lSwfK57OzSiz2VwL1RepQvjPT7vV/T2QIonMqRGb1LYX0kqgw6K6aOqnc1jLmXct
EIW32fQ0DifswjB3ZwBiTx6f7G4hSdoXlWtPdUzk7uGDQDk/3kNRsm+pbMB6VpTk
qd0HS8M1fU0gHFK224vpV96Up7amwFP4lKxovQX74BwXsy8h0Kup4wHaFOGYwL3B
NxPnQ09CX7IpIvynM0oMvG8HBehsh+EbTMY2rCDnZLdKnLK0UbAS9PTYuyrJ1tMv
pzIQAMnGdDhTEV+2/uuhVC6RFL3pRG7lbkm82VzvcCmMKrFzV1nZURbYaSVvim0M
Xyl8107urVBVyjxKqzPlfImKH/yoDZtASphhXRuQ72UQOAaOZKjEFK/93a6W7lwX
OjVUFq28pfijqJ8X6icJKS4dZ0E7EtV63uspmNSbexL77Dg2qPXTtwJvv6jT8kfo
16Lorl3NnUfJqm7/NsrGINkiUjaLgciHGax/B9Tcv+9Jc9H66gTBxR/7AOyO58+v
Ow13PeVpdvS5YqJyn9TdIs9SIQyIS7hzvTiH0yu7E/k1iOh6MJqNZFelQoWuAe3w
5Gki12RLfA+PqZhPdocWL7GhYNyEJFuweOwQfD09rniTtrvW0Wl2GmBEvy4uP/SI
vMLAdwNaTEDqyuvU+qpOVESTwRhGMzIiMukrCQ+yshS/h+GN2xb7GWD9DCDY1zzR
e9hJuYu0Ml6a8yR8NWIx/cUgok3ySPzP/xgDqcRuCKyDXDk96HYJrxSrthrb8jUn
xFlUVq5e+rrSBvceTIhV/UPyG+4VkFmha0KIYl3TUJsoLZFCwpzW5VjN/HPJO3zo
1bXEmGetllr2zSIb5XxFC0KqyaDKs1SgBeziHqcTW/XmGOViY4UlQHMPWLZmeft1
CU7dpl596Db9ZPPalbhVME3yopVQnjzF5yVf+ZygFAs416Jxk1xkElUr2g67+0tl
kW5ErbCbej5Y3af+oLjoPSz4u5KKWrswTD9lZK1YWVVpqFYDaRHO99KRtIZLE7Nh
TrWXI7ThCLwuu0HeYpF+xoSW1jfG4pR/fnb+dhiut3WFEshvuVzOGUch/yW7PK8S
vdFRwY4Jnx9iCUnH6CkTstvCuAJA7v6Ed/NiHulvRAqyxO5xtY+0s7MF1ekf4NMi
BldRJfYMOXrP7kuA5P9Q7lUbv/vM/dFHEHjkdqNkem0RBY+OsrsccuQPCUAhz0H5
CB4ppLwAQI8VsH6WYLgbc/VHxNW0vqIT+mKZ27FCp3wnVO8fEAvXjs2gn0v5x8hn
Fq4mDjuI6fBtW9i7GBMVhvPUEv2XWWoBDLgBHm3Ek98zUyJdwvNeIZDPCId/tXn6
6QUv5eVqwLSY4c0IqtZDiJAipB8gnjANTq3GRfC/FLUFbP3xL1NvblIOiUMWpwkq
q42KlfoseDYksbtYD0lI6++tFa9XTizQgLdH9zzQfZOgTgOh4inTB4X96P6XkaKO
oHDVZpv0gG1Ou+VqQcMP1rmmjkyNs4QNh6E58VD0+6eKH2J5caej/TERqPrAiFru
CY6/VdMAfGXRc+UTMKXRd03G6q6rMmMBUuhw8oSc3nl9f3dYa575MHOaIxdColeV
4sWDP8kVCYBTpWKo5whsP6vrqIKO+vNDiZcuxvWlK1UvykwdoPx0m3WfxI3qhcWd
oyAq1xXuuSmYuOIs6IrvuLjaInM2QMo+3SXlRlCE2hMM8ukevsvpEYhZO84h1Kyv
x0IXihGn9xIpGgYAURGR8e2WLHkf3RWy709AeddNoRHi7tWBrZie83pPXY8RJaTb
YfN8+GGC8WhjW67iqPdWWyJaRwFTGj4SHawJg2BsWVjioSWpx+qqeOnju2QSwarh
oklAiOTH/TFWKmfhjNnGwgYfi1FrrrthvzxLhTaevCbz+H2HW8QxR6Czfh8E2Zfl
vOLxBzVDtsjYEuIcBUa4jFncidvFl2LlFXAgwFIEzj3ubmnKTabTnwgV6D7D8Cv1
vZ611JVNlwEIvxYbW2TEuw==
--pragma protect end_data_block
--pragma protect digest_block
Q+1lOIwu0ihk1xEwLEf2/aW3y0U=
--pragma protect end_digest_block
--pragma protect end_protected
