-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
kIPqhxdAADGrIC/V8kMJNTdpmyeQD/wTgoIQP9BGm76WwrgPMTqzXK7kieceAbsb
+R2twO3txIPcD0IkkaUYWczzZuSVuVuPDIYdytLB0btxhJ1HqijR4T+yKtmmUiKF
szShzm0wXsoV4Tgj4/6ChYX7UlK48VIartKu46UlFlI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 21424)
`protect data_block
lPEjuXjAjdtzBFp5NQycsHTkWrmHyvbC2dhBveROblYYBIHTX0rZI5bCZaG1R/nT
xqsY6n/XNap08HT1uzH4LjxyzS6QAPS2XJa3VFwBD3r+wmpzDfjh2mIki7EtF94O
L3kdn5YqS1pPhHxR3arIFLcUG7PofTbdQ4hSYlBjgFBAVorR6VaqfbJwYiEw5P/O
T1GNK6o2EOIgiM32nPKgoUd6cJBBM0DCikfVyeuJEukTzOY/nc6AE8Ht+3oIe5Lp
sqIDkBl9OGpot9MhKoQi3j9SrF1YYYUbDqmaix3xIjhC5aMNFA2uOtn7LmvSTW+1
KieK/DdJEnX8OfLUFX9G2n8b2X988CQndmr+5PJ+eWUNkLswlmkdq2sGxdVKz+LQ
jKAGeGTA7vDxxeVi65qm8i7nbWvOp6YknwVzG2FVcoemjv17Nk61r2OAwlgx3fQQ
V+osn0Emuq7lNfG8sX8NTieoGO1Mm+C4XiVVVD7PHWuXYPc/0tQADLhhza5fq0Tt
iXAUH+5xsyvmLp8LyXXBvOBqip/zsJ00l+GPil+8mbl4w5nzdCWA3ZdD3XJ97v0Z
AsE1SvviQR2147icnieQ8ku9WQ4b8qM/z8WL7amY/HGlKqGi13hbXs0U/Ofzq9L/
T8A6flS/GrIEvfexP8/CXe17MRuzUdaChtytAe+DQYcsJ7YPQ3ywFmtn213htoyY
c84gb4zvVmXd5TmUkC9vCyri+ovNI9wdRNr+xUTQ3omvEANsEl6bzShJfLm96h9j
DaR8AXPzuKDs+Rsn0FP9fkKbBhOR/bEOGMHuPfHqmjQZeyfYPwDsOACPO++ixXYL
b5qojKxKgwnXNrkYUe0rYWXBkhBklZ5rUl1tDfTcfs8bsktAaKBOUa2yyC5l6V57
+q37c/z3SyVHNPybIQfhbAtdlUWDBI+93ynTILUqTzfRlcJgMoyvNaAXOVvvFcpt
PRX/Na1RIOho4SZO1thtV8LkKVJSpbLY54RmwU/1DZCtB3JwjFJhjuLY+f8T9XdW
ZFcQiGhOLuzhZUF6QVdXZmpwcxR0QDvCPZ8V/srgpQXrUzL48UB6ggaTRhQt5M49
3edyU9is/xflElzAoXNh5JankjVjQIfwOrmgYZtCRt9C/EyMEXz2/44dZAeFlo3i
ox4Kep4/jLLb5EhfnpCAPrtpW0hqiJ7W/nByYI67z/TBKUBoXCq76xvpJ9xW7Wpl
XThEMrWE3oyQltYmXE3j0Jj3Fk9jkjtmxZhVU0AiTJeeN7GzU/C+nQjZ9xFN53r7
/sjS8lHRjOZp/ojE6QL8s7e7gjsq9OX+ic7kL/VrTWpGDYNq8d1w1T8eTPXE6Bxr
H015/bLpmveuG90O84s5hOrfg7qHQjvrD9WqRt6nst+PWmF58GrQ87Icc/sqzzo0
1j8gWWT+Eiwug+ueiQce1TKVuGfnor/WtPr48/EvhmCvrj4GQ7j4fblwdKSHtIao
vmbmf6K4vbWZKaUidOe1miXO+Buzgp1tnUJx6YrvcszIdaEyhCVyQixF3Xa4v425
H4VzhiKdP7ImKf4LhIu4zAOsclNs3rZAdQMBe1yMAoyIWQcqFphJN0M41aY8qlnK
KT2IViZrVp1vK8TDpb4ocXTYzdAi2Lxlm0sBG3+/CJlGZv0ubGmSUdNXRBgSbqE7
c93mDNGzLuW78OqwImDeXPf4OcANeXkC/dNeA42jOnqhh8BDSaKu/FDGqDX5xQCW
wOfCKeQmmC6f9qi4B68SM+5fWG1ax9LX/Xeyf8DJ8bABunONZ/1sbdjB8s/GSYPr
ex1WnCOjhqmOFfvFg+EEYTjWSELk1BJMjZDA83KFXSJO2T1WBd0KNVPyaEMBTtRv
1H0BjYIVuiD3y3N02bcTVHpzIyQl2Joprrbwx9vNplOaEBeaoOroc6JIG4/KlNUf
WKyTVcD29dQv3AFtsfZvNKcYEoGDcZJrEfqbUSiQ6pGbT+4W0Ap8miN4UdFbvJ7C
nYsYn39q8OEOS1RoLzxHxGOEyn0ZlwiojJIrapOX8m7tR1dWKkBeMZjhH1diygvj
j0sWzOuUi3t9sCz6+091sZbRlTKIspjMcOJ3HthucfGIA8SEMfPclBzh0vu2CpPk
aB9BhwaHrtCqHiv4pKhTJGHNhffpMonkATWBcJYeY0XSpGPlEStK04AilYRaNfAw
Xsv865rIzR9EZ5uVUcjEYlc6DZJvRB41eCkBqCynTrSJLP7kQbUmB9oaCZmTp4LR
eqNTNTHNr36QpJOBvGK+9isUlrRJAZQumh0pJZ+FgpiksqrmAWGcIDeN1NJ3GoGL
yjWxFJCV1J2KON5aa0nfoyfyAc8qqS6jI0fXcP8iBSZ8LMTCzU0UZiDL+5i+Js6C
4wA3F3UkzDx+AeLl9MuJjvRsLshvk1WrkYld6fUEma4+Ut/jiZVsQtGVj4NNkJVm
pNU7oXVswF7hkP6AocNzJh6zibSyD9TzbRGPf0GDNoGWJ+Yk64WeH7al3v1yRqdg
1HMzEfqiRDtEVDFTUXzipEWtZ0L+9je5A7unfyFuJeiRcLr1JSwC8ysfGVAk6+zV
YfThN+67hX7BAm6xfXsBaZjm5zI7NuSYmxO49n2rhz9q3imaJn1EIoWY+E6n2sij
ErTK5qektp8Wxxc7Ml+W1Nd/xIF5sebSLuH3fGITuWR3t0cQhaCycKmkWkIU4F2s
lQjbhCn4F/e3TdIiZqzyGn5xAjevZoPTWGaqp8o3J/NX/vMP6rG1Ozf1zknW4DAF
pfrYGtJFjYx7VZaeUtFQ6Tth2uhq+u463gseoczSlbHm+JBmz1M5+MneDazL2+3T
HBWaDfcbvfsQRAOEVsT6ehgpwYS/SNx/J/2FqVaY7/RGDy+/B511w21pn+wX7Py8
P1KLNI7sWIqHat0RX10A86Ei+Lzqt+vUaV8kCeD+Q/wQ+c8Iul/2znqq4YKhEJCh
WJL+L045bElFsPzByHurcJHUw0LsPzjKZRvXuhDi75/Zt+nzeOE+EotvUotB4k62
SAECwDC5uGwhqVC8J+pMcaPdzAEJgnyHudXqtfWtP7/dDMfB3vZ+bH2YKZ5qXQcK
0VO89+AaiKgtTg9hQVoK/KTCUtJ/ifoLu+keFunEidnhY52nuWvr9Yo2DEh3sAIj
yDDWO2uNNAZPRiT6IVVV85wpkdK/qx87PwmFxVmtCbXMW6V7pJnzzqwMwf7ZMf6J
m29MHgmSZLRh/a5kAxGem+sAoPwC3Qa0q2MaBzc6nloMLZ1Klr6Avyf72NlCtTg5
LI0QVGNbsLV7tplqQm3VXdutDyyv0TmdSZmF/htHaCEeGihYx2B8d4s8wQr1a3XK
PsT4GV3beXm6TwE0EcZFSAdhRzJSEddeJsn6Cp134n50jJBBXMSkI6gfACU6qOlE
H2zDwzHyN/EhkCop2981bw8KnLefzYP/MptzmUhGb7TOIYkQpR07XOY0GSOwxMfT
xEVoPn1qWNR+zQgY5VCpusRjO0YQv2Xnxjqf9PkFYUqc1Hnk66xZ14DXSS0N92dm
a5hSF2YEo3gKl+Thl8O4NU9vfWoUu0IlgGRopDxuyPzbHIZITqq6p2opcNbNtUiN
s/ASF3KUk2riU4gJstmqENK0xkj5vczjP1kyORp1kGvL6Fp/zNTKMjebtqVN7SmK
8G+wjv30u63FRZCy90tvvhHLkoeeg6TGEonmj85OcobZPfxLMNq/FaMQ3TuoeHkO
aNGrVae4jobezf04icGrV5I+dECnClv9uyKmNz5xJs+Qe3LTJ7rYhsF2+wWfhXT2
RzF/PEyYWBlzK3U01m38u2PRE98crC/OHB3FaYbVvjH5cFRQ+885wQAzia3q3coU
LC2KYoO2JW1OlvXyxoaFFpA+rNLC7zXA4t/BSpQKy1f3yIvIA+Vh3mbyTN2scyB+
W6GUZVynRlJL1KgOfWcqicVx4/0RmwTGcxJ3ZqB82OKs8yfKqloIsbHgaCOtobIF
xFd2MrSDRQyWFRtM+YIfd7Ns9M2zRXZcM0MdUjLOLd8bmRB2hzQO3EM1yiI8xJ4l
MuqXRV3PBeTIUhccmKOF/mSiW2Kc1+ipN0vuftT9GHrLaPb9ULrXqLrQG02qqhO9
m7F2RvnDqYstApQ05MDS2rjBJTYxYevTz7eP0QocJePw+cTv9Jj8Q3L7yn33LwQm
CzyHfOhnnOZ8rxNdIU50NcWlq2NcdPbqXpmi1efixiDKksyxeIdtJD6Dwcadh2l4
YBGOV/xt1wU0m5H8tj8vkXGMoBj7hCq0N/Ifuiaw8Ejt1qGcJlBNH5+nPH0QRv+Y
fqPwKLdY859lyYiMADOfOnE5WXTfIdrCFSoCeFKkNXIu2QEICtdqGW8ca/tjrZXU
0rD3jfipkOohABHezRY+sYh3DHNSADsUAaqVxX765mGewUI4DpIMuQKBfw2E/7iV
vPFTdgNMHejE6MoYs50welHFhBmQMSSTqTFkfztugZUELuqdoekBccn7H22M9Wci
rMG6ZjRBkCgTRi0DEvUiMj0sQfU31MsuBLDDJ8NFRi/pmLo3BZZ4ZwKuvEfdk2rr
ZTemLa0aYquHu94+ezNU7CL82bGLMJorJXSGy+qaxW76eZmZur7GXMbucwz71HAn
F5lIeUyGR1EMtQlHUHQeIB3xby3hjpTgROhF8/x2U45UbO11TLDiBRpZb1W1kpiX
s4JYMso604yWv3zx6VaNS9n/TbBxJ8wPNKw1f1ZMLHHh8DnO9kaZu+9Kbn3x1+L3
SQdFru9jmIYOfE6582hc1ywVvYNJ8TSuO3tEBz0mCt4/lHbDBMp2vChP3WS2yHjr
/I4trdBVfwmL0Qt5Y0OUXn4STnW84LCRG+mq9gFV73SNSEKEQzA414BNJG5IvkEa
ampdhoLcNmjxbeYsp2k42+HYj85D0E4aViBJJLdiwdpSsBiErNrb6nFSicdQ6N1K
tPWqn4LttVZBDXQd/sy2dT7tHwHKOxqCDEFFWClg9Zuqr230At5XNEX2H0J5sYm0
7NwFjUfriRDXHx/xJQYiltlYXzkhmcjqCgcflBgpeFq3SyU0eHmygJNS4l7q+uLo
p7n/W3RpAmEtwMPSr4gZFFhpPk4RZ4pJJqzy5eMoEUg9AuTfo6H3JjVfKhuU9lnh
CSrzegDNThTvV7ZLXwhnqADW9Y+8ipOYZxWLHt3rcadSmsC+aLpacwd7OnTjoF4D
oDuNxc1j3Z8JbhTbqHPM7G/GPPsM93ypCGi2CRN4HBCxRDgy6F74NiAcZzxbjukJ
0e82i+syi1cSjjKOYz/BZwO+k3iI5DfAIfTnR0lccHSEZoJ6v4T2QGXy3oYHfeDr
kpF5QBZOKGPwtShGDXIArTNr9RhuaETLDwMG1GfhIBa/PIuExiVT//5lS7LQwJeG
wB3X9Arm6uE6cucvjzUuKss8aKNE/Oa4f6ToQ4o/Z7oUt/GRHb9Ui/NGIWajHuGh
nuf0tp0wG0trJcEwFapWrU4d8YQxNa9DQisNWDAN5C6lmHVHQPiwKovSteajbLZB
zoJ0trBWCMqQIJUrW46KjPN60qP3R7rGTMg3ZwoTHJUe6YT1zK3l2PKZvFsWCxmO
knPnLieYsCqWy8yODol91BEyqiWvvav0TFH29NP7hyjwVFDCXx5HnIjbHPDDmWiH
pvKKN/NXgnh3FKlDsbI5cqas4vEgZlOOJD5FTi673GG7x86jPqoielTOcCwY+mbz
01Edly543uP+LX/2wCGKmR5FsN4GfTEd+Ikpe0ZVMmOs6x0PJ0Uuk3XVkuCec8Dd
ItBAZoMxjEmsoXFgCm9+Ni10fXN3SQQwgbMhvbBYillvnhjSr39+AMR10hyrMRUD
ESaoM/L8hpYD7tLFukiSw+OOkNZSn0Eo29XmS+E5y0Kh170ZxLpkYJ6GJNGzbaMX
jMJ6KA+QbiLse6RBVkGUEnG26aZv4ApXW+5T2z0Z2JkKXmZQHs5Xq6HihgWqJIl/
/Ud2my4EBt4tYiogpMvMlizJwHxLTQnP9j6VJqdcIyply7MzjKuKHnLhdb6XhQOF
1eJjc1TIGShAl0xHjwDfBnht4wlRESveRJk+3AB2B70lwyd8jucfqmqTNOa+jzGs
ArB8DOfGlK+BzOFr9faPcY8SIkKWMH2I+fAN6v3yIQi+DWpsOYGMXXTx0zNLc+r7
ulYiK3BjzcOShiju836bPpdmunI1yF1w9tTu+e8YvlwTfYLkryst+yEvZjSYVRAk
vj+1sH1WpYkUy4Om0Zqwj18YC1AcYgmP6LJGLcb5N3M5EUxbb1K9EHFcvoVxhiqS
SMQq4fb1JptSTKgYZgC0e3DZb+r3XzMLPdbU+rLt4fLXcuPaX/10SOcyTcoxe8Ov
Em2+8GsOYcfWsQw0D70FZhlfE3zDjpW7flyFRNQsw3n9mfir/pYyr8EjorPQWb/y
EUN47386V3ScYskiQRq2lUL4A0s7umKlfCCP2zfOqUKXfMlLntmztql1szTMQANC
TWdqZm6CeYAbzYYgIPH7T4txhUT/QhHqq0glYfCYvvKbGj8LZq5DgTjJEcabve1W
Oc6lsNdRzagXlQo0GYwwOBh0dcqKT+uvFHq9XMHOucJaFtLIaffFfnbLxgpyrO/f
qzGWkJ5yeaezSp02G0trsbehj2fC7cEi7iBZLQ6uBcd/gLC2LrrKGey277B3k6sj
4RXMVuamScN+tDamlCBUEFbfzVzFnSvbOzrfQYJwOuIb/XYHiy4E7B1DARttEgeq
rUcBoHPbRFk/Xzh4VaSs+mpptPCySldjPZadY2v0PJRb35cXXuf134mn5EjzysMv
VokuBDrqz5JnnNkdnMorU76rSfBE/N5WaN2pkbU6wcRzBOeGFE+GYsiYmhJtB/K8
3B6OjAdn2n8BRw79wKA9EbDn4zdBFtlPKA9gYqz4o9ITuJUrMS0X+sPJiPacvXqf
5lMgUzBBkme4teABrUlMJK7oPTUH+ghrVWYM1YzPX/VCWj3CeFcoI//rD/EMYxjw
NuMxGk8qr8/pLVZO0/sm24CMnvrLXByorHAiNalk4eCgh1ICKKw15pQJo4jkVJBh
uPIYOpZbiU32ROAL6i2N4a0L5AWLEJ2uPMEGD7YY4nWI3CilN0Pnc/7dna0IF7+b
J5/rXNelBQzgYr4Ik2GxgxzvAq9LldQW80bm6bRZwrTfJjblwEDyQkZ07LEzQ2Du
Kb7JgVLzyAor0wRb4PvePY9990tOKuryKEeAyfOMg9al1gAmwAG4TCVXWKPiJ9Cf
6lcSKmCic1PY1sUwuQbiCGXz4TwJUxoUuBu7wmi8Ah38/GWdlit8Y38CdP7swNy+
8HsAYyz5Dxh4YwcANAi5l1xl7KF4YUZHnfke56oHW24CjTBRdcMZAPxW3o75EA0D
7BfjfqL1pQjXW825R22qhZ990+xi5L6Y1CYPMm0Lm9ZoJsu15pPl7oUHenKoz11M
Exb9Yl0g1RnsoqG571tXhvvCYs26QnWqyF8yr17KMlsBuokwuioc/axnDWdJUlF+
LMd74jW3js+HdCNZAbUYRl1tp6y/ubT8Ih9I6q33Q71sF1Oa6mp2Z7n5/6pg8sYS
OFiq/bRl18vfCQIQkn3ChM6fPglqyWAPUysTppJQKslMPvaqrfWndii1h//mYEUi
JhK2b14RR3hVAvQbNp1tm1RU2GnQriditgsoQ8i2ZVNZJPaB9AF8yE00DtacwV/3
43YFtmvOMROiy7oTEVTfWO7S/hnd+SDP2RycNduzQi7dW07+zwYLIw2K6d9rdQfI
7hs7TMwp7v84IbAyloHRJEPFhDDB+5LytPGtpluxWKQxL/jyHLef72QCMcN915j+
Cuj/X60uL7XSXdRaz9fjc6U2tU0JflV8ozGpYMBO3VkZ10u1Qp5dt+zgdSGbvjnV
XMRUeOefTCTIJ357BcidJAjXRhcLiA9LpDUPRf6YoCdIrHa2B7BfIMKDfTn4gSSB
tCEmrXI82QZN58tk1+jNMh4keO4D/rlhdItOYkq/J7SNqtFsy6WjukB73VLVjVhe
DWgwXcNyEApq//ILTMHmndjMp42pN9zEbNY5WVfTFXIcywB+P5L/kgeuisf6BHhr
wuQnreizUS+fZh7u1w3JJbe9Ssc0KoyCbmN+O919CeahYfTDUNmZQfsRVwBzoKKx
itOjgVoupzb36Qw4VcRemBnxq6X9YEpKZyODHPN9fK+vxuhXDMG6u/hDcQj+jUgC
DRDgFMw8Mz4zsT0iecgXWsofZ5qXJCDjY8W8+AAT8bg6eXt1qvCk2QszRWSvkUZH
748M3quRG1V4EIN0JNZRDV274VDZJQCv3r6RUh0Ych8uisNdUc+cBRLOUicRCZu9
sRSeU60THG7U+gqo8AmKT89ZNyaOlH/yVvx3Yf/k8pURAJrvVW2GuVUnacYlOa63
oRmm4pERsSPs3AoPxTP/xn7cN+P7fT8SPCSyERrxf99fW9PuYef/M8Jn1UwzmjXV
/tE8lLxO4Cz2MqxZNdvpEeD0Cj5s0eVrfZMjUewUrBQQpC5cADZ979bg1N3z6gGw
st+s4M5VS34/2upaUuwUGp69Jdqx7LbmhOIZfqY8xO+EHrbPpmNFOHTo0eP2tSjy
5FPkj0k5f+rlCgQkLM8XF9lRM4YG2ghfKRnaYFMypgyIjyZX8muk0QjvkMOAhuIC
37T5OtpCtMjWGhbVcJ7Gv+rJsjvxtzm4RCKb786V4wO/adCWTsLvg7859mi/iKtd
m2xuByN8ZTMojEmWDblcJmSnrOCoHy2M8OkprNhqKvkkIe11/xSn/+3DkJQFApJH
J+FDUayQgLm3PKuP9idzIUbdutewEUH1JwaUwQAdDbB0pkQd77r+g0WguZGLjPkO
gnWVe9Y6IyhdoSpw6P8HwWfoCujAlOrzKy5gr55Vt24tPVsnh89dtcznKSbPijQY
pmqz6GXiuHZEkVVWa90/1/ZVgKz5EMkK66hlAYnud1+9Jqt9cNrsC4OuN8oRgIVn
cGCKXTNCD21FfRdcv21CCh+ivUYZAzGagZDjpZucmAZ5qKTcmpHL33wSHD8MkJ4k
JezbqRa6Ma8vluq2tcoSS8BVi6SYuuwRhqv0gSGaqHQ3VmF9SufgwZkWvekG0lfs
rtfuk1REFIwN762O5UGru6UFp65cXULxbUlLr7XJIO0dmQWu6t1+ZmlazoqqgK1w
ZTBljNKhCGfwDTTP6tu4gY1K+9h2aLYWSqn3fWSGE9KWRFa4xXLYyFmKnkPJnIAR
yg+UpkcWqbeCJopT49ilaaDPKCplcaazsmPmoOpWcsIuycBoCqX1rmcb0TWzSHhp
nYfJrcJS+AIrCxGUYiAbYhJE5UG2XwCAuVby/PhCQ/htVY41De359GL8MCZgoYNb
s8lkJzSbnz3B0W6aEySEoKU3QM9CrGsmlGRDnog4sJ6b854gQc7Xr+5IO3pFd4Zx
EV8WTuBTPZbJhX3yvek0oLx01cKuKUC2ESgCrQK7dL3TQjUEA7rA6rGXwp22B2JS
ZWXxa7+OOj641tVfQvD4rUO8+eXUTkkM7ZJPyHbthFq4svzig2aXG8tCFZ/JPtzM
MTtWtOuAlvAvcvxHoJlMINIoIAaEKS1QcAcJZQfT4/r4znnHQ1mDAMXAyS3o6oxm
JLEC57d7ka/5DGdo1YS+3ksWxs+qlrCyeWyYECoXYFpi9Hl2zFZHiIOsk9iMDa7n
igP1IbPtPefhHDUL2NwYPyW31OYVGBVDqtwk0i/QsYy+o819WmJROj0kt7ph+rGG
IUdTyjRLwYwsK8mQjxj03K+Onw+h912kXI2ehUrIPPoMJCnxz6sDXznVs2Z9VUzR
ZzDArEai/9CpaFK0bBDSQjeh1vlGtpCSZopvOZ1YZdqCCPlYqJn0mcw80NLXfdOa
/FfZFwc5wYpfVagFvtyqP4uO7Udc9LD6bghSB+rn1LOagqAUHzbfyttLxR45fj1y
LRunpIgHc8iCMizgirlrvBWkRq6F93gNm2KK5an/1PFEgqMz5LmIa2O4Cyw/sb3R
2V6SEhLww4eW0/VO/YPjemNSSrpbn1cOPtCzX5Xla7A5IF8/yVuLmPB0X+KBupAm
Axcqfdnvs8y0aoUDpggne011yEYwSzoJgTLVqERwEvgRc4uSd32WkHq4po7qB/uj
HrwxKahFG2NQmBwzcLGIaKsm2M3p3XpYPR26J865PR+jCZ0KR+qN+8UFd0rU22fl
Ge5VLyg7OJgEfRRI5MciqObc3B/f/a28wnUcQSrChhG0BbFsO7th5iWYqNVakxnA
pQqmumdOceALhrgQi7iL4OpAWz2N92FS3AWS5Vc6kmQ8ilD0q49Vr7ZlGN/ENIJb
ZuVsAtSr8/pneHSm3Y4bGZAqS7TBp4OQhRu7E4bZr1VOzX94M1OWUQEEfkstNCoI
iDfUHY5+d8RTx7j/NqlUaEVcsjamsyxZa535GkvE0xUKTooT9NnagwimigwO3AaN
dsHo+IbV+qs+pxxkX7h2RCP8OZGFJ5oBLEFVhrpArxw4L4nw6/johBtRK5ilvmJ9
MJSQbw8FhKbpWUpzOoO7XxVekjjS/lAtGNtFWvnwQcEghlYTGhqgn3x0WTNpKwog
HfIhZ80skm9NzkoyoMCkkhEMbmVqDwJb0P4RXkxPfaVvFsveLL2lftN+6F4e9U3h
b5U47ncFYdxKMM54PpuASUNEKrw0RgzWBTsGqZbun3OMKB0qp1Pi853FmUvI//cB
i+KOO4fgp3/Sbva9oqT8jXcl7ONm9NFHp8T6wWaXxm5UsQICHbs7M853dq1WT+I6
ODOETOyok50gWHea4ppSgbQBulA25Und4REe0QGbA3BtKTzF7UbGXr5o6apouSnn
VsgyYiyWzr5RnLtB28bp61OOhIeuXjSpyna04y2wLoXxg1SMGbGebAvme+jQJ9f4
BhAOusxMf5uTgOML4hchxSKX3a3DeqUmEArCvLOvu8QMjMleZNp5DzOorAAdxtwV
WcqgvJ/ts+g9arbtmDejZORhagyffwWSL3kvOAOL/yrU7xHGnz6daBD9b8eHgGBM
giCTMGmr2bMHgH75djJ6Skkyqog5F9tEQlHqOI36lfxRvyWS8Gk56uUIeyFt3U+F
37VoXsIp+7oaQRDrp7v0BqBUk79VKPpitEmgjlRk7qtdHKWxM9iBEAsZ8owfVotM
/Q+A0o629hJ6bgAeBvt2Aj3VziSp7dI+l4e+SNfJtPInRq5cHT6QoNiKbBI+IQPr
Tk7xLjo4EwP2y6qRKyX9WVDvNG6+mDw3nhjQjFbR38YEFTe8PSPAerwzwbFMPPkn
TyxTL3LAwFnXRfmQcFqmoEMajWrq3N3P1SrbHfo2Z56c0TE+QQnT69+l1kSAy5fF
fBI8wZbsJVgMTRcA4PUwLdsgXab1A6O4N6B93abED1spWUQCN7zQ1+YVMTVHMzQA
DdPNwwwhVxMkUDNUNNhrVQrq4AfQ+YvQWgkzMz25xwaSeM+3qDoetepRtpDPSkjg
82odIpOJTZrEuI1EhPd8g84rvtYhbBmd8CnZaj47/cmzz6cWXgc+LxP/MBqaL6LS
6yXbjyNNVLDyjjBP4KW5zr898sWcYq16KB9eoI41T8Api54auoEjESosR7GB0ien
ouHZu538gG2+14Y6k9FtOh3OE3dHXf+KyyyWTxVg5O0lAvPnHBMNoSktDzcmOOtV
Y7cm58RT8Z7t1y984nteErkCmU7mLF2DbIFIMB9YXh3L8TjrkTqWCJol9NEDxIR8
kb/ZBaraymazk8fMa/+vPBSKiEr4L3AtClGDl9Dqnfv2xEzbSSlHlxZBEm4SrzS7
/Z2oTuVBs3rqmUgbiHkQVXjJP0f3XRf6jekxSoBGxrHRT/Y0BePfRzvBSZf7Hkzg
yQriyyjx1cTOqk5fx0VUgVKA7SmSxdDuSWaFXll5nF6OYU2jR67XMGwVWpLxb4H1
w4Cw79tjtMokMrHFdgwyREtfCf7UllPHhD2Bdalvz7T2gU83i9qoVdjRJVYZXU42
HPFoay5Bgv/+EcW/B3/S3HKXlqd8nCuq+HgmO94ZS/PseiLaLc0OYy8RDPYTg6xK
mnV0ZI0dw/NgUf99UKoh9gSBcHTNLBGThnZ8EFDHlROoUsr2mJWavwKXtojAdEu6
E3wxKxNoB/DjO7D524Tv+Q4JWdMKrF0k+pWq1fC+8+kSFcwtWm7OQKMCSlfK2w3l
Yxm4gYl5VNK1DysA0reTPDYK6mHmGNRwIZJcaQAGnYgq/PWOqwHwLDRFruwYQNQB
kBDfS5AFFM1gipakS1TR9wcecC1V/G/Ek6YHgqnsBTbuikEal9fRZNnmwVjNZm69
UQoI1glhbd0DylQPJQhbx9z8kh3mCD4FfJqq35CCnWPxMc8gRS7L7VdIbPn8Vsis
sx7PoetS5UgxLLKQJuY23zafPWYj1D4V/AlZrAf/SPGThwEzmOMLwX+PXakxuQT8
uZSBzrrMWae4bhNyiPHSAj4RraLVOaeLmocLkcy4viaq5YIyb9pbvO450LVQHLAT
UMgfggmpKuX1Wp2SQIvjzLCPUkJT1kCU22m72Sz9HAvMYfreIfaiM44Cmu1YvuJT
5Rit5DVq81NshicvBU5sZxubyE4p0e9S7F5nYJNmRxb6sMC63vv8FhTT7f9PoKX8
oQS8S41CJnX9UMky8KlTh2yAwquNn5aYYke+Evucs1mhY6hfzYAOatDMk7Nu2hY/
rUtioapJ17/Ky2tLEddqnQ57wE8jdx8feKHlDOmP7ywzhCsrNrkHdvORf68ln91t
27+qhqIiut3PafGu9o71golbznybX0ec5fE9T3wtA+e0mXKZtuKV9/xMW0KQNgP5
DFmVJJqNj0nQuA2v21dIGpP7mpfVWEvshCgzhej25zg2ceZQDEvTXGglVLsrPm8a
jjwqSayK1JJS3CG3XUykVme6K1C/j2XRKdfMLIO/h6EBXgLHYjsKTJ54ockqxtIV
CBW4LdOYX3J7QIZifYQ80qmJAeGBc+WBxoJ0V0XS71Ibs7z6ojrzuCIlqsxUPBxw
zO4Qw9TqGnDeiX214TJfBzIOJv8such+wIgOq+lWZUbtktXwB+w2ju0kyez/2Tdn
6x/Qeu/sCaa6hT7Am0eruynLTCCRgF4M8W2UtLmSDjWFxhVzKgMzYfiRBqYVrHzI
0ATQYsrDOJuGHqj6LNB4Bil9aYtbo6gnvmUjHozZBeIZT6ZLluwBN+GF98uAxzgp
fI+X+GQRc7Aoq/59oDDDCRoe1yHD5Eg7xgnpjoEv02oChtcaBWn4UgVCXS9QZGJ3
G5zsKSDL1OpnZSmpWAwFdnx7ah58X1cdOVMhOYaVkca5TyBYbgrjOlGsnih5rsB1
VTmwfV3SezNF9a7pk1xECdtev9ZX7Q1jxkkD15a0tKGbxKxEupAFiy4gU5ubSoY2
ldkiqY/YVV8DonChfQ7pg80qjKkwIIpfnetBsLZmjFPya3dgzMsMduG+9pWSH/84
5Jl3vVWF+AjHm6u5RJzJpJ3ksLhh/vuRug8LQDNZPWTQSOp70zcmGYZLtMGatE5L
70GkG7vhhdA1NIuTciDMgWcmogNOpMYBm/QbHA2iUcYhKILItg/BkAqiwVSYoIHk
H4v3bCLHe0hYPBH7dnvgsRhl5HxFkUaLkflltpmjV+BHUpHKedfP1NdixismC4av
xMAV9+An7KXUTqqf+kBHq5ysMv2glCAI0DHfECTKatKHY96pWXwSkbS/bsCEJbTz
tIpsk6uWAfoaNlNcUEqRie3nigqTkmdlIctLK/rFCwwLgwvj0gqd7NCbRpdf850M
wPH7gJX/jX9ky5l7MQfddinJXMghhRJrE1oxvqmfF6yFpNE8NeWkcsM45BtPB7CY
XZKtQp512G24AHvVoxZVc7fJpJYgmpb+wNtFzFQk+zgKlgCJ7241BH33zDdkfegu
vG+eaQS5+cBywOMMCiuD6vqkT+hhOORdeHP5EtPLqN8RmY/axmpBNAs50wWZGGJf
8e1f9d1FKCK1+O1F8BK5l5dFBoT1Dw++4odHWloPlb66LiVSfD4a3PZQS5xwxlQ7
1eWrdvXSDKPycNBET2DPzDSlmYC8kqpWms/xcjPRS6m8wH+KVZ6jvwG0OMdVuARF
RMeNpV36SLszkt6Esv9gMxerG/apHK3p/ewPq1P6oAKlDjaEBVWCs/AaRSM8h3EI
YNfhx+doMZGsCFEIK91UXK2QPkkB4zrVQh7aEn9PV1RP4qKac1Hbw4N3jP00BfQe
DRQZaDAa8TE0L1btIiMBahY7h6hZcZ0EA29WdB5XNEGSCUMSuw7dT8kMJoQbf6nj
E7f7tb7K/+Xkmq4PeyBmJf5AL9XPeDNNXl5VSrZuZSGWYCmAytNHMonniIDAmBRo
apG5VoPx2oN/vgq3zoym1f2NXDAudXNY5uHZsPeik2RrkZRi2aiOlJijEv6c1lZv
phv9iVGXhS7P42bxt2o0sUJg5ZX4z7K3DL1E/IumV67OTzk30fUsmnDtoGG8+bnM
b5VbIR4NLO1aq5OGyV0JTAZj3lnoU9gwMjTnjiF6P75EgLhV/fEM8vOG3wk6W+7O
zJWYOBWqqQi70Xy2ChILdp1Et/8Az6uEia9pRG6E/ZOmNs53FFe1egsUhjGTZ3yZ
aAnvkbpx5dCoSG7Hb0Vetk7Jf3gLdje9hTYzjMsk4RjbUt8u7K4ChoEDUsawNM3h
Yg95yJgzrfDcfpAxBXtQxj4UOpe7cC666fHcakGU0w6EXWcM2NZqJ6ynZeQXRTwJ
pr4mqs6IHFwcHLRCncgxtktOqFbZg56CeJtt0aEvco44ptpLMf2lWkc38tfdlQIW
UQruBIYX5RY0dB3/D2WE2dt9totBWjX5dhlIJoo1ho3zWH9h6QqD0DFCZUAaDBkZ
abwpGqHy198qsKlt6eGxYBA88AKI5wB1+JKv8zQEs/V0XNBEjjGfvbeVe1GjAfd1
UK7DFxbBh+zfnmzUh0of2MnD3IRjjKyU64Y6rGzfWeEWm6ihxVQD37LR5aenByIq
MZpOwAhLwLGw1RvwA18/jdNdBpcCkMavx+S7+Avx1SMjgpa0Bz4T5q1euuVnkF51
CoTwgskjB0KnNdAoW95xDhPKAeAxJEPl3/qjpsCUZwCgnP8MAFs27H4gpu0G+TjW
OlkbxEaTx5WPBwtjOrres4g+ZyZQF+F3Qwf5qcIm4k0mNB8dqq5M3ju530lczpBd
nzisrrLPKIwH1Ynh25dPEa4Sd3wrL2WTIn963iOo4NN6IOXr1bASz4QGS3bBoE1p
W2y6+j/vqjaVswEa9HeDjU0RN2THCf4qAWprzPj7709WfacLCGolftYoKzQSh4AL
dzARVJW1tMsVExPFUG1/m7ABOPF7eukRyIKwC07yH6D7Jiijzjmtv028CtvrwywR
SrvQed37eY3aaoXs8nX9MamZ/TZ9Kbi8bZb5TNkk0B+r4kLJmqc97pGCpXqn5/bE
rba7qMaA18Ngzim+iod+e7coA8BcrPkXwB6K4wuRV3TAPhkCqN45JLgq0a9qrYEc
f+F7J9l8+F3LYsHFFC0Q+WOi+UASGjXaHWF0Wy586esIvaZM7zsq6zP3sWFE0IcS
KgY6sIepFaIuBWTIIsl4eAftmf5vYHmbPFaMdA/nr7RdWa83QCT0Z2XJ9xL+1tYN
m7/CXOo7LuNDo5nz20YxppwFl344Pk3MRNUO6bYBhfhjPsuPKNJMrY4IVR3CS6mz
ltlkVZTFjajF9mpi6hR6NQJ1QyRtY1TSE25EVEVC6+5SMGUFwyp2RVNKkEUAWbKY
aq1VbwoZIHMd1HACJDBg942I7A5sRK93M3NIZJb2daaUK3DcS7HqKgksp31v9Tu2
E+713YHUw4QA8vaEuFLCH8UG1vsknkSdI+YTFTKA05sEihT2wPeN0q2ty66sPHEC
SX7tLy6+B/0iVpoYWtgm1mCfpa6EsRVbaa3lqeyj9jdJlFwQTqyPsZbJTTyNmtL6
2/NRb2Gsb9iBW+E5IjG7IixEbgPeLZu/8tc6TxJ753Dc5vv6gnjZTXGbjXAiVnix
ZWvIJmScJiTb48TH8VEOHbJhRhdwezN+oiVLavUXNwMxWoP/N19ctKccEaqfmRfP
kaWXz+xTISnffvE3CUUFgU8OTBZEoGLSvkIL+EkCQFbuZoxFz5zvOy51mdjXaGm5
/5aJ1TeLn9ovzGl6pfUJerSGHqCS+mCscdg5Kj0z7V0+REt/f6m7pS/MtEjTu2vX
/FqVvcegaKVHyaPq4+Vcb6YLxRInGvsnURbhlDrNS3IU0vwOPAd7Vcysb80Fyxbn
lWR+k4MshL9YkCsUPqkOqXMqU820ArQT7ehzoVa3536ksa0jV8O5wtne6IqMbbln
NU3ld/lTWSU026i3Qt7dMVvpfHC6AAJbT57/IThzJMHCnwFsO+syae/AoPrCn++P
tR9W3U1GQimwIF/t/0aBJigVqVpRk2+JzoJEqYVfm9w5Qfkled+3ZKvLXNihsbtQ
7nPdkgMiFnBn+uqb3bh7FzyvTIqJqpoDsXIkvzomwy8hB8ll3WvdY2BwfrRTkTVZ
lkGeSpPkenZxg3pdCS4XFTsl5ia02kolrR93/5lMlG1JOgb4J319mM3eZblKzkKQ
beUMTU4P2bSel4t8nnfu52N0Tx6bqFHzXFesFs4dA9zgnuXPvoLli9ZenX725tPP
DmqkgW8qdmb1u2ni2p4d8i4R7mX1yloGtkjDbXyRwdGEKQrc5XwNj+QdbitHIPS/
B7Bh/Mu/pG9UWNZ0qcGXq+sy+k3nQ+9TCLw+ijpGPNsXXP4yv0JnggTxoC/MjPRp
9YLs6S0zjQWlFYla83DXFY9mEmBOumnZ+P9L4oBX/af3hNDuIZJAd+ASCDGpFDWB
rdJebohQQsAShGtAR80GmpIRI9Xs0VnYgLoPBoNC9ihYkJyxQ4bUWu/IE/FIm0rd
gno+PfbkY4R3yMSZkHpHfYY+3Vtz6vl7yha4iDIR0j/dbWnMC2uP/Bwl471iWlL9
RsOqzjYPaDusPQOrGamHnZ916Dl2oJw87K4rBD6j9vmMS/G6dPn70/yBs3RXrP8E
MYGkBGi6uBEq3tAMA01PnfgPm/KSGdajB3l3rmJsQDgCz7SdbXsllXsVUSK11j/Y
mAxymdRaoixtJ65BW+nSmqchaOBt4Dq4hRrF7a6RAe7eck/IZeo4O9ybHdLsYrZx
dbXf3bmW2cQCp+naukTd4UEG++PQIoajmNT7UICFX/daDNqhXnbpuG0J+DpZPC/X
pJClaP1bV9o/sxQv29lRSndMUI0dmm+2fUZjUDswbgfzOnvHel8WbpGtBqW/YvAj
beJewIedsCCvbO06U24FPMADVg14FRn1CpMxt7eIReFHcEiD7vJ902YqZWvIoReq
C4i7NfBUufN70ohVej4L+EOZlxXMUkqW+LJP2NECWaUqzMtSeWijf70w3RL4l4OC
Lu0RBIrab3GFGOtyDFMVQri7gsdejfzzUs76yjH/moXkAcSCR5+6wK6sYXtqdYFF
xBrGYVXNePNUy7UO64BMfboHR70P5dlR/glwfrx5wvPX9f0+BRWCmTqc0SSrDDuK
80NnUixnPYjLdo0U3ctkpOZT5nKXTMpzEv0fHKLL0L1X/ALszprNbk+yG5Je6wPS
BhizR2xuF2KRKW3DLfCmOxMjr8JGrRb+dFYK50+L+ljW5od/saoiNnyXDFJXfgl8
G1yt9p6WMVrMyzhIn+/pT7khsMVwTJ7xTP8MmNQj79xf/9dwUeZRASpx8ILamatv
shuN3qRLlVxi2v1TfpMbnZlds/EdXfCeCpsEtfUCBd6qgUDpiWBllVbVdkENQnRs
/XwNV2+YeQl9kgzC7YaRdsxP5pwQ3CY8YBknuePM6Wq2a1XqPaAvbh34eYr+vHiP
w1eRsF6hxdssVDZcC8DIIpFc8Iu8tHlhg/R+yjBf8NnlFDnMop+YzZYHLzHjoDne
wVMUFOvuJhl9twOdiHmxXub7TQSKYYbhIuqcHiTPIucwC3QEbnvC+8rn+xDYdv8F
Os16zCl775ouGu9Hg1tYMzzIqUFGCLn9z1xKwoXS3IZGmOapZ1dIA5JlmINv4QTR
6pC7AP3ysuAkCRV5+GEf22fXxmPjXUacVroNuM7w8gctLmbnkeVCP5OWkaz0yrxL
Z+uD1XkFHPGglTrySah7niy9xUIz9ZJWSMJBf5yN5w0ww9gEXs9UJfs0gFysVZ4v
Sg2aIA3c6SoSrwWjYIWhp60k/UKmRXYdO9IDP7qqUf6rYrPGe2rIWOMT18dZskeV
zPlgd/Fd6wPhp6vz6tBmj+uwm5/1sCpnt1V4IXC7oImbp2a2UO0ePmUvx9I8eSk8
ocdQ9c6SPD8eC5QGXxaRfdm8VPgPSJ6QVSwkIzoxFRMkjdXfRx0BIl8FGKfbd7Kt
Oe15evd4EUO/yWXThNhWzJ5eN1+PRpGR0WyXN/tXOH9OTF0F6bxmPcL+ovdXOd7X
EI747dRl6O27GugkkHaHOcVVmmGuOfllf0wpORij11Xsib9lnMtPZnC25klUfF6k
1xOHzZPihHP82G4YmPvbcjWpMULRT+BGCAMDnHY355Y+DIFt9zrDANStJpA3CUF4
fxKueSIkoyGGQ32FLWxUbLeoygNn1VvV6j4v03SgKvlVpbkB64ANWAkpI5U4KF7x
7Hu612rpPYQxBoP2vMl5Eq2MnFplQ+roiBGsa14iffibvugt7yF37rex9qNN/qtS
4/fWBihg+DipJQzZNJboyoLTNn3ZNMk8cLzJUZEdye3gIiczx64ig+Xrm6987fi7
JB1jH3qvzr/ebc9FxGRUOXXaUJLvoehIjtIdPJkWM9e7P0BiADxthUVxH4MoNQ0o
+xncrewHCTtcpwiOHv8GijSvIvNpMXvZdOLC+OW4mYwPaycAPfAKAtavoRF82V2P
/dG0K+agexkz+tRoAsjXFphk9t3ipJvjGkOBLdU4AxlPgs3BAY8JpsBvsK+ai6Yn
5DijIgO1mSX5b+CxdQq4HQCqXhOFtiaJF5pUPYy5/XICo2UrYodG5zU7XY8sazlV
aneIEGKDJxOQzxvuB/Z97vIfBsGg/KL/OX+c4AMgKvcuao1NT29dtENB9a6mb4WO
9B5vMAf/cni1POEQvlQ4+IlY30cvqiNo8U4/KxiyIlOy11ANYjK6GfyNy88dXa1n
4NNbLTO5YcLYIC2wU3mJ+FjCRyqEMVUn8cWLj9A9+vGNE5rf/kddkuqUTRQAai94
z6THCR3gpAycS2NL3cIHQuOWnarhjMmWnCM7xFhug/lhQ0UUMTrSMVszL+hGcguf
JPy8zUWJeZI+7Bh6QsoN6qp4zms52WJ94pGiM5/R3Spys1Nt497Nuii38eZBbav8
dT058PjmmmcMo4hQ1A0BsMsBrYzrd139tPGB8te6mevueFhkgrOm7VxiXvx9uozf
wkHlx41+NgX8+OkXgDLwcpc5qC9+NovZNKSXNxP5soOg56a0bSGtAK9+ql1cnBdF
IUb9bvqrYNm9L4BkdwjBrvar2kTODsOCDVlM1a7d5GTKHO2fWMM16kt/MnCS04xF
+DvW78Ivf65PdInCmr2sGEQYfbUVuNnkKQT6GfC/08wqsnhn9wIY3ODzx/F2yYZd
9svn2WcaTOBRpYJaMk0u4XRhwM7IsLz60sXJBnV9brQFpVom5XT2X6IuM5qNbB8g
ILyL0t/XGHSM92Pw2OUi+KgfmJZ3k1GBIQR8w6xfQfjwdV+3j4oElg9cs/+Y3dsj
ScV8+H22mnF9jZewZE8mlqWu60Ht+POL2xui9zfX/gqhltUvNN90H6tNACt58Sr0
9EGBs5YJYyHXBSV5qfdWt8Dka2Q8CrwHz5wRnlTn3WZOq7mZhTRIOpc+M3NDrRzk
7LMMH+MKmf6e/IHTOx6O7fBVPC78JX3B+DyfozziL400ihXsyynI9225MTJr9nbN
02RpEAq38oxlSNGicXGfCI1pB8euCqCGboY/W0rRbOqdcX3PJ7TLeNb/23lqP1cb
x+VT+iWSF1nw4dLpo0UZTqVq37gNZ8dEzviRWgaqXPgLkTatvRXpFZe2iBMmUNeZ
jyFIY1L2HeOOtQdl0vLG41OC4VQ6unISIebSPWJ++5zJw1XR8qMXA1ZmKgtu1xio
ickuzvfYWGJoyIJj2gYVoizo/G0r5EeReJL0Ks65EqfE6ffwxSuqcewX/X5JIHw1
pcGyxmvzEIHt+bLRrLSwJHFJG55nMuZThZa/SK0pvctByyl5OYgJnvRLCQl+WDwI
S8q6XPR0VeAQdifUhWxVdr7+XSkPNlpl4PHzbu4satM5avlL2R5xkHX/uCkj4QkJ
S1nU/1X+EAb1VAe4/j/BV3m4ehOofilw/YHatd5n8w1NVCGtRuccrXtHaa3ZOFOI
jyjaKsmucc5AfEhbcmKCB2kfN+is62CeNPMJtFDRL7nESk3woSC0QS9dFlSQG0BT
TYpV7D8YgMUG5rBuVVV9M8NbR5RsOW7ovHfpViW3IzEx5a4Th/ONke7nj0yd7005
9UDDu2Wi4chEUAw+xPTJp5sg2YOvV9T9QMU1uvJX0mCCtvBBC5iEJPzbzDM4THSe
Qws2/Aed6sbcXvr5hZx9xX0WI+qculFuwB7x/21yQBApX9+ELcZ2+eeZ03oxJ6jd
WXPhBZqmWYJT58gd9oboKnBzqZ0E50htHLYn6zXZQFh+NBn1KcX5hl+KRAa0rbk4
IJYM297OkycAF1COmVCntveVO06nrJmJb0kypYGa4IjC77K915gpifWIEXPXF4mo
SqYg3QKW6Rcz7KJnEEgqXpc1ct7ncLwXTXeYgTSN6/LDxMeUyi6YuBEuJOna5E0h
JFYj1VW9+4yKZVz1n3QdmGB3Wvaq/hsWpcX/QvlhRI4esPAP9Z/tWoflkN+l2IK8
OLQZ9+/+4JMSd30dbAC7csFCZzb5z7tUHiDeyp4HodgaEtMXOvur+JfFeRq5vdR4
PP8OcSfq5egNZz57q3Kej7kOTybZ0HAH9dMmipzJaNmAId2YeOMUc4ZeFbMC+0sA
FvBMOVf7XTZdTkDUx7apmswW9BfWvG5bDrEr2MyubldGcsK9yopbF4QY8l4TavMY
Mjww0D+28rtKjG1wAmbzFu+KdlbneIRD9RRTWFaLy4YXt3YZy6o3IQCmXpJwcudw
Mnw6HEu4eEt/6NQ4AYjVpuiwVj4MpauYcBZ4feb5LQ2OEG9P9I5rDVA0bdaqm5RS
VEZHqbz2atNaagQCeCfiQgvfcMfgFzzmx+hYLXUVvXEQMw0elLuUX5XUtxD/0q4C
DLIwZgaQH3ygECikUL/tKRcYtV/6WGOnqS3JtrNfLWzGV6KkXjqydmLyJn+dh30A
D8KZyqxKGzMh+DjFLvi5Mk2bhmTE+BGVTZhONLYbs6pA9NCDf0iZswj3U0C0PsGF
hUkbjb92tIXXhgH5uoAFOcTAbSWW0MyQZvHtEY8ABZ6X0GZuAOxiLxFjhNRsjszz
Z6u0/ellfQQLkxi5u4N39+TtiTp9JIiofF4O2MJsjrtq9belBH+QmySS7+LoIT9/
L2X8QL/7f1TSDYccPH1aNijBLeLxGRwQSFwWIVLYIWw3jQHRGRIUz5yJOKfHW7PU
j66BRF6AIXqKmKQweUh+eWLMtXfgDK+dbgruKHcuqiLeHMBDjj+5Opigqzbe4ovH
/zHPSHnqdZPW88njUy2Zu/fM1YxYMw1utIBGPEclx3O4qQLoMWin7grr9CgKDJ/1
EVBw2SvGVBxg3AbrjYZro2/QbRxTqN4hIE2j4SHbFwomD+MpgzITysDdfu+qEU5W
69goXpVKcuwy8I0c3/CBMAqfqfKDp85iEoZhCJz8k8MbrF71eT3thIEx9fMYavf6
5XPMXppCGt0yX66//OGGrtmvufSoU7FNRsiyGG/mXfyDWZTCYOxXNwtKZKJGTv1b
gr7G5b2n8vW0oSs+AoZ4VyZujJcVCGPSRfwJ92qsvVp4ELRWk2zKLSJdIWq7xRC0
Rm3A9PcwytPM7ynS8z5Gvtv7pnPNX5JuKlgglTEUWoWhlhfDqT5JxMkLOBRnWG72
HuAL/u1e8W+RCoBgAfO/raKykuxJAQWPrEKq6tItEnaWhFeNFBH2w/uEF+xn29tl
ZW/t2jxN+Ehok1eVTEHQmE6z1foN9c+Dj4S2ACXrjogtqWQrZ/vtoC4znx5sTzhu
3umgzD9+cwly2Cyb/Gk018f9tYPUhJfHfW/NvzDQ4Od3hJP75PVrQfwmBsbrcatu
UF2YB3r/F3nonuU2JspnaaipUG3BwlpBbQ2PAOuq4LwoVerRFyYbLBohgbqaiFLo
uQxrEV0uuz0mJYL4dMwQqwX/K8i2b4Ps9Q2/AWG96jcrAA5Ox5aaUO83VgtPLNuS
ZSTl7eUkkVdaC+2PUWrSAoWUVfBDeaLibGwPfhUbQBS1jIewFJeFQqq/kX40R2B/
LkIabJiGmq5HFA/vvKYoSdy3IVCdO2OhoSJFBEr+2mxq9aI+ds14YyVObQHH3EO7
FMAA3ssfVeiUZbjLoZDVzCiAnPAxC60i+gS+LA2z09JwrjxrPIXWIiYDON7eUuY4
Df178Sp/4svq+N6EOOKNgMyHzB/QP1M4Pc4un9REcGvr5pxJMSLBVzhya3E0Lfq5
ju/uf87mPsIkKBKr4QWSxhOGbNexiWisW4pkpwv1JYi4b1x368sn3V0vLGajPs6l
Zs6aj3f5NQcKbSAU125i2hTECFtx5xMINRK6pS7xsnq+zjShfc47hNfnV90j5dgx
LaRbnbtjpWsS2SttugNQ6rt/EJTbgMCTX5AreOHABuzYgFdkhL8YhT1kdTOCjAPU
AJMEfsjmGw5T70Cn+inhSqThYHz+TvPd6uYAzjdNCdnGCHnrgJnfKqvOSboOMfHz
kGnwG6/Tk5Qufk2oZvBn5qoyT4LwfSWVrH7QysOx41LIZawKpy6rQIq99AEbTkAv
uKnU4XNITOZELQRpIapxJquderxDGXv4ww5ag0ATs01L7KEUJdvlp8Kpho9jMan5
7wSv28UeE+jgF7ek6CuG+gIutt1oBfMu9tLbykEvyTdu7WOsfo3t0hRX0CZhfQ4a
Zd20wupvEMA2ho5+DzUDzYSPGIuS8vG8JY9lEGDSLk3tpsHAvNhpMoVXZsmEhYHV
Mob/SaMAXTck51VmPG7wZBGsdVksGLY76oDPWWTlsnxSUnBNuvCPNcpn8wc/Zchd
Rpc5enwjsw0sEZeg135gpCBg1ANLddPNce/H9edrwxpDYAVJ2qtKISSMqCkvxTMh
IYkn/7QOZsTJ5eQTkJPPDFR8B1GBYBoakJ2fHO8HZTFl/0uQw4xoaXObpb4QbWrw
tUrxA4BPRYw2BIfBj94NZH/lU44Npx4z6HX4b5OKu6XAVY4zf+HiErD7JR5BjbAs
PIvOl+XfyJ/udbsU3+R3tkJpc72Hfog00FGzw3oNYwZsNl5udZBkdtwZsWHlJv/C
d+nWXLVPjGogMhBU3VqLn0aILC+2OQoYvfG/03hawEFTrN3Xq+ngAkKROosvhV73
967J78x1z3q1Iuj2XWDGqgoEkh9M49RXy3OK/O82HOWKU2j2bZQs2OHcROQgmUzV
Jjc4RCxfhgnn3mT6SNBOieI8K+b5H5zP7Gs2u2l2Gb1dCvQXwn/bP3MhmjJc6jx2
CWHo1erhraV30DnHDrWFymzF/ghiyALEJ3s/1luO8acblm66tFOo6OcC8FzD8c3j
lVlk5JVhtd9m034gEAwXRinmERaHp5gypnYgd59zLb4J7kIDEoQ6JONrPq3+ar7S
tM7VP4bNNq2chj85YjZUdIWUOHfpsLUVckBv3jnbvx2TTCgetBmBNxqBcf+kwcl4
L2HMg37h2AdqXiR9uc24Q2l7cn3q6VpTNg0xIuNSpvxe5WUv0IpdKzpAOpDrPL13
WWPa8tyNIaO4szFM6FRtE2wE1zHN2b9s1MVuZr7M2kG9COpTo2HnDJIUEJoiI/qF
4C0bQuVz/QzsrGn3cj6lMv4q0GoWQGt/OmE60zyfWpNpa98DNvUv2S4EcgYf+MI6
CSSk0mzQ+IBl0uINQ/jDqAoECotsFU0hFwNeBcQ2sNOxXOUqjWqrDgBBU9qPVyuy
3o1YhXouEku8mcwHkwMTF7AmWHclk5JRZSF5RWTSiN6XCv6PGJq/hfb7fqSJaiAJ
2ZWiGf1x9KqZ1DvHTw0nHFLL0fjGT+bbp1xXyVL20Yqf2QWN8yxFZuWCj8vH5xnE
IU62MKfBNup0K5FfZk/B+oeZisbon51oSWpl2Re/6A7bLcJK1WvhPGW5Udh/MKzT
5c17x+wrZKFxXPdhx25SZiZ8eAKXTx+2arUx/w369kBKFr9us5sO6K7kXnqfa0VI
VxERf+/gQ4jNSd9uG1EiQ4y9+znleTFDxCQFUpzw1Nq4mphO6RqFVX4t43CIFrDq
lXZu8U0+fedYn4c8RhGFp9Q4/TARkcVxqQoiQ97r/r/g1iTKjPO3nHZwsuWzV1Bj
UjlnbT0T6ILV6E1c9oCUrTzLrxSVqrNkQJTgywkSfldwUrgnuPTn6lJs7Lk9+6Ct
Lt+jw+0ChhKiQCoQJ1Gthqh3mH1gdDa09CElfYD87/9sIR/9OaVwoAhxuxvErJEx
F11TKwmx25ipc8uW51TRAOsENPk5QeiBPFsMlu5TbC4pDmrD8uGuVGQkVtd6MJWm
xBRpNDsGfsp7tJ8U/zHEuyKMvqO71SLNuMtELPSPta/t4sAXmBvyj8MhoUvkpL7B
iUuvagZfDbyQ/yVVD58B+X0UwvTGYEirvkiZwuokzWdYXmDzBnGasy4y1XBKoR9M
D25sPNGmNiG39MKLj+IxxCJl8Aa0Y3v4oXono+I1U3e2qJ/sXUDI89e/lKi8qict
/dk6xxLJ0/9BEfPOXkccB7KcydlpD08hG2j66QVSlN9oC4Ai7ybUCx7zDSQVVteI
vsz7JmBw43Sm3nmF+gw74npwHBmua/dyKlElq4XHMeWG3fCb6RunyTP2HcNE2l4P
cLEPsq+LxXrVyqH3hqT3RCHd4itzpNYIBudWNbsiusf0dYpHmgHrGrOmGB97wpwz
eONeJXEKq/S3mZb0ssxbrP36EJf3+Q/28afw/cKcUfiEtlV9r4EK2LxzKFKi2amw
2W1pa1Q35ZgK3HXVzh+OukfUZTSUZuIcXg7n+MjgIzJZEYfyTvzjJj9itym4ycfg
+0G3eV8M5gASVPZhnyKq8phkss43pnhlkzQmg36QNZ3ApT1OmYp89geW3dwcXuXj
ov0qZixMLKAEeyHnX5OSn/Ql72ns/cMAa0JZeoKWiCnpKfyJjYnFurpIiGB+zM8E
WhZ6vFNGAk7XjwmqgYXPy5YtREC5QUCO51xFT+lUsMBJ2ycldYuCCk0E5d04xd8A
HYaJmRteZm1TQonFboJLg7pj0wj07svO/Z3yW8G3q44hELk7RTzVWP7XCwf5sAZ2
VRkezuKq+q1eefQaLWYomYGL/z5DHOawW1JKDDPYdASZe3YOJznTDk2sW3UgLMbg
+qz9EmCwM/4p9oS0ZAKIuGytTBZBsHooGud7jpRvWceuQqU3bPzYyWEF36ORY5BG
NxJE9D3Zz3M6Pfbn+4OUZ6I9wGoQCOXhUG5dq32EcfIY7OUolRRxjKuVVLhgJJjC
b4Cw7/zcuTgEKjFGgGELyUOX8OUM72Xo0bAF7MVBLDUNDtA6QMWiSCh038m44pHe
fnFV+W7NX3GMtdtAww+sRXXhx/h1m+OgXZEnGZ78yZUz41WCm49cEU1xpVfQO7hp
6VKxLbc3KNpTr7YsGtrQS1ztPJXb4ze5n6OS2/ELsgHSxdb5vlsC8RIyA/hWvesi
YqTY2rZTUxW5oO4x0VmeGSVXk3eDmsroOm2pVKyV86kyKiraIgPkEVPgDW7asNxQ
eeA8mXjWs2qTXUIEArvw0Y/My/tW7eWyYTJyMm0/Tdlh3r1F42o3KnAkpi6QFd5H
okAnxqx2tl1FfR+sGLwfCyXR+XblFtHMREHdZ5Ww1rPPTHERylAwlgMvyqCHouNI
bUs7DBQovVT22sEX6oHBednwQn9brReznR8GhwYZ7s+hV/LXq+fWTQksJciaf9Gc
m0XlgYdHdqG6hx4yJwcWnbzP/v/JZ8vRLCuzvAwUVJy96cDy8y0aKWYSLs1ogG64
frisIP7lYSeHjrUmK0F14u15N9rmGBVCrmh/gQseiUQolEU4O+WtSsvDxONQ1sS1
SnHGEoRuBowxOUVH7e3aoQP3J4mvqPDceZf2wwAVCQTH2z8n8MH985cfp1ncNDxz
bFnjdSNcsUJ0qhPo+qXVIwgxFFUkQsBsYvJP5Xulx/V/0gP+rwJ7hVoNGFkYmEAi
9xuleUdlTy12bQ0kaw5NODX1ZmHtvYfDcIItB0MLz6AXj2TG6RMpb/Pmm6cWBaBN
YQhmVT7dWh/4Fpwuz8WonDy89G5Esa2AEUMwfEoTHzPqVkD0LInJqxwNugJ8w/Vv
3Df4570os3b5vFjKW1nrVWmCMqB0FxnDIAv9eFIcmzYtC89V2IUA+9EdCJ3cJGqC
pwh4Jcdqeo3t4Zyd4eMmgp04WhrdS/OIWSecpwhL0nt5rGkxcBMLtNryYy03By79
sMaA7w3i2rh/aiHSZGTtoQB33ndULkxDpNBezOtTdNbiIN83ayds56fLg/3mE+Jz
OfMYOf2ntfA4AogDuQ1tC5zFD3korJOuQhq5N9XB0J1xfa3dnw2FepHTGj3238jO
Gwxyy3W12CwwWBNpzp7I8rpZ6V/DfwsrZucY5rOgDvymn6ar9/kKUpSbeUKp8oRC
NzYR46Dgdq1veiZ7bRCx2KGwpBDcS6xjBcZsISDc50hHJ1FzlcOqemIgLTsCjG97
C3kB3LLkcaHbsboPjzB8oqYIiC11s/0URWcRdAd3Q2kWBcGLG+ZtLdSN/ecPXHsW
kodtX1inmoiU2vG7gPi7JQ8+EC0SP/YZ2gsr0ym9E1N3KJYCuOptWLr6TptlOZWi
M7LaMNfQPViG20fSdswhByCGvm1xX32Aw36jOhPAS9JZFTROnQFXNr24Lj4UMjG6
hkTsfQniOe7UbPflU411xvPQb060uPBa3vrA4YAuT6R2vDzfYSucUE2FaoXv0Hk9
9Fm4Tr5tIuoJwbxcP1szdUqQ+JscvMdRBkX5Qd4rev92HeoMWj65JF/Gcwt2Lj0F
DPUeBfeUjdUjZO2+MFT+oLQFHByNSPsYidJPYrZ62bPGHaOyHbo8SWpGEb66Ih0w
mTkJvfHjKWsK2wD7iqdDheyT9t1+wNtzDp2iocy5CcUzNk/OdAk6+kZi/yD+0TPi
JefArY++2QH8OzGpKuZSUQcf85sTQJpBioWKQ5JG78P2imeBgbCHNhcgSEPxYLXY
hp2lP3ztAejsBpxBdnWGjLY4hD/U1pcw6K5c/4vZlC+xffu5vaJg1z1eTJfVnNKV
oAWZTskooagKQGHX6mIz3tvF/lwYXAUvEUDcMGyn+adyOXLXk3V1162qSwHrefoe
WmtqFEMEwCBv7ZFG35hOU2KAa64dLQAkpDhul+co9Dp2CcXjd/m3T8y1TrLO2j1U
tMUMelYykzawooEEQIA3ZvFyAb1Stfue8rpxUpGwHWWj7zEFt80jW314MVtq1499
qqT6mT8qW5QSxf006ipIzwuPTdggGOQ+tUPwuj3Gj7jsray35AAu4xieohjlXnjc
cw+8eqofoi8Lu/Ert4xpK65cTEjJ0Y6lKfN4OlXLKFYWb9zEytyArHTr3cLn4YDK
ftr8LJDj97sMyInEsj9xuUUNv/VDHTh90A0WC17yGLkoT4Qkwe2Z0uxqWM7GaBNT
N1y1AFsyNlE4M1eTy85otobdEr6UIVeVp/H+DEqgELekSDmq0mk/LJR0WEK+LZ7A
YOJ9jTCGscNPq5ehDuYfyhYfSV8ubIwLPpoqMJZGzCVwGowIOwdPNAxnJRoMhFTO
x1KJ3ySyEMax19J+LVzoC/8/CBFZ9Z64js3NYy3Z4lewI8iaFCuitMLImeCWVKP3
92KcJyb8iflBtWaV6vpMDA+FPv52+RqPFy9zTTD9CcbITziCTepY2gcy8IBvhdUT
X4S8buJ6MI11+s2kicEzarzhd8KjTcLMl6c+BB5nYg3tOErMIV4r9CRGDRNlEovX
iAN5oYsAsuBKDU51piE5ZYMkvUTSE4dTkQglBX/W14MhhupUKaJId5w5coOzPL/E
uNz5COx9/FVN0Pzp4HOOFWmqt83rhnZAwjIvJXmXFoiKpz9w5t9FUktaJogTrFH7
ma4Pc7vLLgMjIETHrk05Nc69sFzJo7EfeN+CtLXoPsUOn8aS1yQ39ZDWFvN9Eiln
/OBUAKTJCbQFIOpDwWhl6uauFmBSTXkBbBhsP/o2F9pXh5w2+zsDg6xT7u8PHrWM
ZW/uEmitRRIWFn3sYB7X5nID/DQ5DNjtN+TxXFRNuUywOKwjxIZSyXcmLedeHfMc
g6kjyZkyrFin+Ojosg4kb1L5XUqytw4OpzjqUq4nGIe+QgiTba7v+K0t0Jt+WF2e
APhFtY/EYV2tjBSXzN51qNNIjJwEwsAQQVSFBuxkRoQ1yrwQY8uFoteHw4YZshKo
ki9wKWP7DCTHCmi2ea5cfQ==
`protect end_protected
