-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
iMWBqJdZOwZSipwGzuU4LSDegEQvVowwqQY8YsrglHVD/dBYyxEIN1o+5LDcXRqV
eB57E3Tl1fbTm9Eq4PK7TaNtKdbsQ+vP3Tyxf3aQbejEZii7EfCt5HI/iWND3saY
kOGz+Ui45hohdnGDkozvewZpMCX1xBAANKoeFazgDLY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 10679)

`protect DATA_BLOCK
VJqhWlv/QTDkmHjz/sC0F+ePScF8xMzopLch3p9sk8R0eXoEM+zD+iHKNuPJhzrU
39Eww6PyS8+OTGaNX+fPNH5byIRSjWpW7TbFA/Xl15cw+MBHZhCw4cPmB+0EcnzZ
vf7Gd9tXeYp8ivxosm5BXDskL//tLFNboUJ7rIr+84qnpELHEcOmKi52CaPjnS/A
oe8Kyt4kA5wLFaO9sEqoHTfETZa1bM40++evPIqpzhAZ3Wi98hrmDn7JJN2UykHN
g2UM0XpD1mXPJ60d9m9LagW/70aDD7MBePohWrC3KbyTlCTE5ryYthC8xQjpaRg8
ki8168oIx41oy7AlV7xLO07uu2m7BdubcD/QwKjS/t1GhRbgIPpZqFub6c7E8mwf
m2PTbmQuYDIQKKlLHMlTTIXrL1V0obsIdHh0xiQ0EWYcf/Y2NOJX/Z06ClSTuNDK
Pitl9QiByICAvzdS7Fo98hgg+nZFh+XMQ5udbMD4eW5mZQkzi16CDvlWYXbdnFgq
7bbrAPZOPii3VEVmVCecXtRxmQFwywMdW552Hvtz5L8gPnxyeIfWEiX58UBbCMqF
3OfB3/Deqo2gqqxhR8zKf2Vidv+58/jJR5h4hX8ZQZBV+xyRXmll+WkL7RJvEN+R
5QI2W0R5qi7l41Plblmp2mgG/uiL7uoVkk4E/ln8gV/DxrB6hwKcD3MvZpSNNMdo
+9TsNYkCflW35Qf6okSTz4NGRim8BY0+9K9LFwt1L90YQVxmAV/WqK1hZ81WYPlA
xbKAeKvFodIKRqr5umqq1Mr8EO3XvDNyeku4RtbEqrtnqBP+xrKeLQ3HRbQtTuK0
JVrJ0Bi/qdQWOTMIl9gw7GkqOCjFrFRYT/RFaGjTPCxDspCTD7dxLQ8YJ7REIVuJ
YVygCi1e1UHL2nGdO0l1jbSZRhNAXCZS9mSSkbSdj80j8vECSD9PlXv9Mef2xygA
5AQKYcW8vB/Uj4lAMDTJv+qucYmdy6Uq+oz8/TH09Q1CxFt2NjbMfCMz4kKj07vO
ZnCTmA+d5caHQi+GvmlKwuo8phTM6DKKCBOShOEVCb06Jf8/2UOvROoaF/7FrjC9
73n5dT9jwJ04wwH24TwC5oNPNSuFFdkVahWe3WCBvXX+3ujbC+XqzCusOwZqhwvL
7rIEIzqg0gBRONsiGsFwJT8Oe87RY/rRFXP7g3/v6NYDCNg/niilrClw+MQJ2gud
4fF1g5RTxQ5rxnfAE7MyvML58NcTyLj4pQYUH4MizsCrx+i1i3T1CnGTH7PyeXQZ
0ao1FOrD1+0LFU688NdM2+fRAf1OZTJFO5G/qtTH3ifyxgukqRUxYnFxPdfvwCxk
6CgaVwsvYyLvsdleILWKTYZ2AG/28soEbdev8/bASr8NEJSnj56OhfVOg51s3HJV
m9v4aZH1Vj6UmDtJ7lgWiTC8NfYVVXHz05MkL1cO60bQMJfq8Bp4iw9vrhkpQ//S
um8v2wSlU6qSU+bun5CT0FuAlQTvPJZFnYcvRGpbyDu0zbdlF24lAecbbdx/OUj2
m7y07k1Fdd/U2Iyic+6rkYav2Q8cut4TcIfW2pwRgBbH7JXH/nJzRUxoeYNNwKv9
KXZVaxQ9YVXgBurWGz1lxaDNEziXzdPftRlx5DMYs/QNfocpBaq5iaFerrGIK5xN
ZZaNnOFibW5PK4WavNzPmjVpY0kUBpsxSa3ZJI6RoEUheHnXVKJhSueWoAJQE/pn
yALbSM2gi6x5T5G+XaYiYYm6JS16aP5Aez0G2CeoA2Z4XGVVBt638uA/gwZ/5qBe
K8e4xtSnayn06KIn6QaX09O7b1LJhpftuQ1YYNFFWzXvlmC0lpR7r1n98rK3s5AZ
K+9+uMxl3D4ZkWeogYIHSz2lrDxiTdRjYfTTJOp31yz0AwvpqfZ6/FvKeKpEj/ov
W+5KZnWaUGUW64/+oILHDPVWgRacveb1JMlEpoxTL9BAEzSMKfAYQ04tMUZ9FouU
+0Hw06AP6odS2zQsQxDLCw+5nZt+QlQuHin/lNhqw9CUNCm7Qdc08mfDEYQ9QMoA
qthtUpRW4+TIeEa4Wxa5Z2+93IE7tKsZqS20nGX5XIJOYD/VX27UZwWRNb3Sx3bs
nPkSbFFkRfCEq81DhiX6ELXPPONmZ1qAgBY4//f9tqgZ3qnPbmlDssoyc/QZfUVS
aLG/Hpu3HwIBQr6nQm5OoE5rvQyhwR2d/HsvbiLfRKMIt1NBPyCCw+XjNvEiw1jp
qokmMpQU3Z3nQmAUQECnlfUJM2BTjz4n+imaWDz8H5g3gEhDedryBz0Id8PpOamZ
GGUtecpQZZdAQpXdEzrHQvmMY5b+UPmrXXmDR5VbRZUiUtflEpE9ELDDf39kx7p9
+Kw39onDp4sD9zGajxAB03Pf+ueQgxaGrtB8zCLERAByxyiJcWRs7Gsl/ix/3oj3
suMdNlqYLGmyE1NdhUplYPDFyoLPZjYCIx0RQNnm1cojj616i/+2XmqyZF1DnsoS
UthRT2xSc5QnB0bIN89nq2BWCetvuqkxOq/JQqIx9VO43b4ud/7cXkg9Lbgxg8Hk
uGjppA19SYw7znCHpwVPRAXlqoNFcv725XNzeIuwU7gVc4vHrnoVWQIKkQN7JbWe
zf6Nc4NWD3NC4qowNkMVE4xXuvSRcEVbzqFPZ/a/s9iTHCSajFr/raNVveZjKWHJ
3iGodZZU1ukENk9vKL32rVwcZLmmYw9A9PVTt/Z1R2/iH6omT06P1GcSKYqaNIp7
szZMupcsHZHpgyYcIEdvv8z4/VBQtFYSl9mkoczEv+y17WLB5Gh97n8u+sXcWkUQ
lTC1EKi0NcdzLWYyTtAVI/Qb1AKgZCi4Rn71dY0bCdhq2TaVMcDKexGYdlK1OZm+
qIlUqhtmakrsfDBCcKM1aGu7E8Swy5gYy5LU2XKZf9UJqiRhYFporitaCJyPgqpK
kg1d5nk8A3dqDEP8xQpNZ+2syukjFE4P+WPbjHrs2/ZgvAuqYawszYJ2itApytv3
sbdHnNZAqOoualD6ghzazregOPSdqGTXEL089Ix2Xdwqdc5wlFpoA9B1a25fTK8c
VkgnwRe73CeGemZeIk1KOikbqUldRX0SiBiLK3UtjYlK81lhWctvxRy2dmJw7vlz
lMc5ROalFtqOlXzsBbhlJ7ncc7UlcH+/HvilPDhM5DkyO8+vF/jKoXQVIHJd7C1W
TwIrB++402pfJeFFMN50jsF3Pd/LR+FmzwioOVMRZULX2Sc3PlIm2i36ZlJ4a3UY
NQSljHO46EdXnPxeucwR56Q+1YOFt4trZcqe0X9dqVcZgvkkrVoaG0XSCjG4QL53
YJZyshgS/XuBCe5zJiL6Ff14lb1n4rg0q7XxZcywB+Cy4v+9WHwV2V0fXZ9e+8RE
JDEhoEzdJIUIXdjSAX07tcsmI9pFECEfWiQQhA7OSyujJ9sXx1rQ7qG54NtrmQwC
gV5JpLGN7i5mhozYbp1d1XGNMtAddjy6dctETRO9epuSkCiTTcru8bPVBCMCo0by
wRDtEFAZVKGMSwZz73zCGp95sl9j2YLePNdivSAhWHojkgR6WaDZRpQkaPWFQimd
1CWYLWZG2oa6I31aNekr8UrV89oqAEDT+WkfS4HaZu0PMyrYxDJqAWoc81NF7FNW
nBuyeVpcBPe/ZYdOWpzAOzWNjFe3MCHEL41DqUeebqRWnrfLwjY7hLC9E6cg5XC+
1AlOh9m5BAgi7NnMqE4TW/Ej5Vk0yT6Nd6q0BHzqQq+8nzMWXvDqjkDTcualHDGq
RbG/zHwp9jFs1gz6uKaqZej8hB1YwRK4NiD+eBJPy8WpGmKF8NeATG9VUhfoQE90
sVFPl5x0OHJfeupBbqdz+RFMBvcVt0wYnfcWVS4g0f6qrtT3/ti+KvOtq5e3/71m
33+8eH46k5f9HSZ+QEaMNBzz0g9nhck+iwsrZtzAy0w4q9kc8Z+jiigbZfdIGs9u
o1SEazOPSu0V3cJEjg2X1Dp8t4CEx6CI4uLenn2TINNnrbv+bwY1Hb5DE/RpQJN7
Grbge/pykxeEMGNXlR0SMMNBA7MIAh9aQA+vYwkQPbLiqYef7dqrle6TsbGhiSiv
z++lLzRl+RfDYKvcgqDrOYOxpNxgxbPFsX0A4f7uejz8FSH5GYTtOehrDvwjkkMp
yAUTGaci97/Ev535NZ64jAkiiSMimninYWNo1xzmKuC1tqYSEN+8z3cus0m+awmS
yQuenl3tteJkugTOxs8lI/UVWHCTrnSdfM39pofRtqHys1n9jzXlAdB/8ZQbUqT6
GlzNRuHYoxQsu19Sb5n+HqeOxmDAHwMjnRAd6oCu4fpbhbB5gLJh3yqOQykG3oIb
gtuMWuXPQFaMc9CNjjjgsHPlijflVxd7qNDS9LDC7AMG/MT8xf3N1oWXadaufD29
CckUWdlaZmeJ18XXcz9OzIfdcD6R+jtn5CcuxVejbZtNfTyGUdVXS/ZWTxvHVkZz
E54BM9UKKyk9i7VT/tQAInsmIb7+TpvW3OZMR2w5z6Py4W1jSNSsWHnoK9JRJKkU
9CE82Pna8mKgYHGJ2nMroMIEPj2se8/HlAcKCYurJVDtnbqhIPVV8MgIst06zyOx
DIPCVo2YkbJtZCoZFa1fK6ZHqjX91pq7DiyYMXqrCFFCD6IZMYgFA5GMqT3PE+Ec
pRNeEznm4c/bLz0Aivn/r74t4E3H7G5+5ggR/nYjqDmlC6yA8/0aIVrDkF0gU+LM
U6JY86WFJ3nPS32g0kt/PCcHhL05GATplrv1HICN6j7Kz4SmkYc5zX0NktK0slSS
Nrr13XIkXEsWT3JrRX6OUgFQJiFRpq+Neo0epxMj7kyiiDjsTvH6td33A6SM6QCk
ZG+dKlDRLOMqpTcRxB/hPC1INy0yRAYQzrtbZk4thUxaPMFJP087Fx9VQqTkc9Rw
jEwM77hTbSj/S2FuHo/g0BYYq6lDnfq2OmAZHjwFnHt7FtGGtmdB+iAzmowqjWag
MakkHqYcust0QbcUWf6bDQhYfir2WztebPZK/TU+woh6XQOVyMBUzK1QfphLjWrp
8laxb3fwv4DyN3BcmxblKpvPfKT1Cf5lmM96ffLEsBkd9iNhk4+4R9oG8AF9Vm9H
0WPsSn6A01b0I0lw5I60aXocdBqtMZljyrMj6c3mfQLZ65iuCwiZxo9Qz1cGQxW7
nQEdXXEvUbdHA3JTsU9RciR5XmnRbBkuIFoe5Yi2G8c+cR5OFczQAngtd9QU80R6
Y+7n7QD0m+kULF7dgVlGvyy7NSbEIqYYTssWIwl9IUKAxXi4ErL/6rPifTMD2yfb
JtubE5Ibj9ko8qkUK+Yv8pljtZH04i8Wj7XfrADpPuuUWCaKWI/uFxOhsrkc8U5G
+y7D+XYq7aIteKUct9LSMG2QmPyGnlPc31NLDBxaKYuJ2KPCzNjk2qzebu98zj9t
1LeMy8UU2BGzZYx55kgWkXAMclaXKTR3NAFORAXJYsCDeDSr9ESsM1dW3APqidw0
RYZJPRLKv94kOLLzDw6Hxj1PujumT+ZRtM5rCW9FvNPB3QLxoSpGbmJm4PUKDcb3
bzGJfcZDNKTwUyGKxBRvSVnZ+bENvHhrO3hsBaooXRM/RNghEwBRImZj/cm6K4AF
GV7qn5fnQV9J6sX8zojzNdZxF7yM0EJ60mykOOPrzU6SP+Wpzbo0HTWlAQMJWUv0
Q/Ob4cozkfsZcYt2D4jAe1RkTBFWmwRdGHSmbkEL4Al0+tNCX1xB5Sf/XCw5+l7k
iHmJEHGwZOCZqWGZOOUxcNg93n5FZoV3lJ8FTShVRcUMRUlWY+71NHBESCPlPvu6
uJos6rL3OHQSuKgeEzox5vXyyiwG4UKi9kS5AHFOVKcmsYoe1FtLIRc7eB8/3fXP
KZnbmZvGJHUQ6Aq1kHTqcGdan+NvAJcFYCLul0nH7JA8LxJSoEljzB+jg7HNb8xg
Cp3w0YsD7rZK7N1pE/BJ3+3TQdNOo/Ty+V0oeXj3oLEeYzhfTzp0fQOlPjIYS5Pu
aAlNPCy5SAPHdO5WMcx/mOoktWEW7tr3nPvUa6z0EfzXxs19fwudwmqOJ1E4ugOI
IFmXI4mnsSxhpJ9NLkR4syGABMmRx4Uk7Fn8a6Ox6cQsf2DJ53xhCDesaaTm5J4v
gI/GiXPCtqAthCnnc5v4/yQFTkInMNX0eNgwhNUCzT9WoV7nXDnZJfRr+54GwzXl
tyE0twHCLohz0OMiTEM9fKXpqn/o3uUmjdkh6QwY80oudlIg9d0paBOXD+S6g0Rh
PIUPNcC0LpIsVmsDZG9hii/q3E1X0yn4PFzJuMb7VSM5O5kLXhB8PHj+viKtjaPn
oacnZ81kWYyHhiR+SaA6TUwlj2laT6QDBvGLpI0JD6H5sABLVor1VO2krGsaS6oO
wcFAQ0nTgY5ucqIH8tcI9MUkS+sSD9A27+pVBTT1nXf+SExHNjvPUb+VZAhxdzEY
pwowIEDZcXS5pRWp1L6NZf+6Px817yT1Z4BWzUGPPgQNhB0CUOpAsaYmJuDEBE1R
fbo91zmH7VOwICg0D3ndQUKEFslanad4SHQwybtmKDfAad08koxGgcuiKqK6qtdS
6bB1/qBNY0VfpD18QuJKccDX3oqlVhcWnF59wvcw15k7B6U+5xFE/0fJPAkNT9Wy
YzEIg3w9HHU/guGcvoydFcOnlMcwy0Jwd0vKv6K5XLDgonscL40bWsRnClTZDJ+j
MMsZoZ/S/NW4xj4AI5MEjZMf1vRF9l2zT2rLlxCRI1hHvHzDxpI4MQDT2De1T758
SYMTFMR5EIMAJrI1k/iNim+8DO8ESy3jvlQ2hM0oLEj7nZPD0p7weaRk1ZwUtKxN
jYvCzVYzPClaoVhN5VarW0xjqpVkfEQBXe8L24KlUYtKoH+63p53PeLIthMXnwfe
oWf07RkCivIn0VuHl4Ys7OZb4FSGgEtc1a3QfO2n16UrWcnRLwNB0wXBiNrAsfif
u6X654MtWxBMpUmoRvyYAcdFWF2r94UdaobO/LqJ+xy5oxuZZZkk4nFjJ6fQqlnC
SfRcVnN6vUgxpx1PbE5CQf+YmrYncMfzZfk8Jy5zxA8X+GJf0VZmCy5YR+JvDLEj
A3JRw3VamMNet7zuDuKJdRP3Trjt0U/zcQ0oNUDLIU0YE9mmGTEOyAsoUJGxtrxt
dCx77LzjHMC4wfKZdRh5p9AN2VGvluR8Ht+qTuzHb0PCPJx//yBIsnBniLREVYM8
+Rvp2kINlFQYyLwHzoL8bn1gEHH7ZIYrfCMV7sJzcxh8TDAF0dILvE9SDRznRLWZ
ZOm1kRgaDhgxSop+6uHscktlTJU7pqojVE2BgkFcchKXcDg5E4kmI8KEwvhmPSdM
iwRg67VjcoM3w0C41rZpYxzLEYA/SWQVSSyba+FG16nzo4G9/1wAV1l5TBsbitcP
LT9o+sgkB2mubzkEgsahm3Y2nLzoeBcobeAtmSOUDXy3Vlnir1MsNgZybn+s7Fvm
x0Wudswc4lgHAIvuaLsn7deywQ+iujcmjJv7xRvpz5rpdTICSvBoTi4d3JgHxU1v
Ga/PBcGgnkzUAK0Ivy/P8Euc3Vb8vOb3bYqQr+jKbbfNoeIFPVRtVzKqdi90HgTp
gpNMf7TvzuZmSZzkMNoIGr2wMKrm/LX3s80ma3FB/PuuW8OMDmGdM+gNFKNw76SU
ks42feL5uOwevbCEze02+gGgvruMDRtIZqTmDuJ9V2LGAozto10b1s6ICRzSfwkc
yWCFQiTm2c5JfllxV3MBFYENjA2xZlMU5Y/kug/NoLsNzak/BL/ryGOc5B0EBco+
Ptaqkv1bkYdIFxRyVs4JXdtCl1/CJNc73rju/DbaYuhQexXGUiP+4GeGOjuOZH9I
SKoS38teqW0YhuH8rXVy+x/RHDmBfnHJGQLl+NlUKJSr4f2qpH0GGXW/5gQaigrD
K/Y55VBEZcasMfFvA7k1O0kVJ8Ygt9CkXXGSc8L/bfs+q5I4gyVgq837UmUOcBkG
EdwqXOITHnmEcgqpkPWNadEPsSWfSHe0OKVMIhvmmyqmOACOnbUsWlcf79bxXelX
CiMLiotk8J7g0BJyCDMETxzGiIUuhe4D3M1fQdUXWiYc/VZtbI+R6T92fp+JabUi
LsoianNOpwmFOjWGXHNVl3cQqdi5PebyvQ93myQQgIKmEoJ1EvJq4DGgOEpnEAI3
On5x4WhrHx95JzIFkPGuYmnBwCElcIudRbJuyiEgm/+If155Hz4heE4qVHSFyJol
P376V6UsithH8kn+Y968BzNBKhKvBslIuES6CDVLiKYMt+ibHXRwN/K9JeNRnFvD
VBCo6W5GjgtwcgjAK23VAO6bdzZZ1UEc21worEN4/I9vpLB1gW7+ASjWUi9cDwbU
yBYEpJREz8QRi9vL3VStvxXgJW6WIG2VqjlHU4e25t/4QX4iRpLRP0CLh7dAFy5Z
q9qG7Jgky4PCD0dt9o5oqVFeizpBAC5/7OLpErILrk7QRC0VBfGoFgqIn6EmZCm2
1Iz/tSbpd5rM3nOBzcSDWLliqar7uIwHVjuY1pNe2KretHyuyDFnN28Ku5tncYVT
9dVC5xTEwYMu20JVmcHAMUD/WUfGQ4a/obkC4n9HOe6O4V8U9wqwc+8kbGDYZ6IP
NQcv1kmiJyl1PP54VMsTpamv1vqtb6BDCa8VUAfkIc9MCcl9OSzDv5QLvW19mLCg
18POsQvpAlN5UC8IBJxVHS39vQbNnSWXUNwoOTJjIc+CbsbhzAA+8dEiRYx6kxve
4brVqo0gCzD809+xtmGsBVmZMSc3J4+4ExhxdlKdyTiAVQ/V8xY6TGc7NNTLUk8P
8a0YT4jWOyqjQAeRgC8WF69UaWM0zsuwju0R+LG3aPSIXMuBbJhY5+oHojs0KZeL
WDiRmFZeflC/KDQuUigymZtlfXTviEURTTHmCehwKXOAdmbGmenxan50sozOt+wf
t8Llf+iWK+sAcgRBGHrre1mqxJxT8mRD60w4y0q3K3JAX5AtnB3Mph+qvLucP5B7
UlrVbuK6mPU3BzH10YvhTHfh2FEaHEhq8Ld6+SWvzkKnWM/U/Gy2H/SOi4FEa645
mz1qa5D9WJ8HQrvfl6DBVIIhRkDLz2wgNHZ84G5D77Gn45Ytnxx8/AYrWSYVRbhh
pMo1W1rxA32DMIwp/35GE7HYnu6xpefY0cndIBnNQr2ez9Mgns32bU7ggcn7YY5R
TWrv050V7A7HWw4TscLxcnZc8FEpIm5M/bATI8vj0RwskCsUpd4S9bFoQMide3T0
bL+Dj4fn3grw6PE6EGakYtYCs0MJJv6nxdPGn1yW7SlCP363CCibhvAnjV1NLBwW
0HCLBhFJ3MT6lm5SDtZ5pTiaCd/CiXQxsZl4ySSUO8Oxa/Qy/Kp9vS2xa0qOmD7Q
Y1r1R65tW1yaV7cLUyc+w2sI4j7+I7g9oXmaTKkDbZewakgNLxZkBeBBhxriKpjL
sCTjvrXZiuM7qR17whSH84m1Fev3R5671MKxLjvmI6qP+FyNY9vETgNWwQWmbv5O
1drm5mOUS9VVvgsAkaq+wSTimUIa0CT/fDIZv5wYPoXzGb6FDsRw38D91G2lV0mL
BdaLSBz9cs7o3J2Fb1IdePqGtGev7LILv+tWEucBgWT+WRre57dh1ZFvsKbJHo4V
OG02aNx3fuPVGee9wXVZSsak46OpuJl0PDGKmigrdfz4p6K8FuKW0Ylmc58GZRgc
/eRVKc7li3bVAmMxPPDDTURYUCFFIqSw5vjRTCieOjWFqDk9JO8dpdrc9Gt8sA/B
moNOyp4vSCYLXtwC9Q/t1bFZlxuvN6xcTMOIgPZV5K1JkA6orKs1qges1jUxIuO5
PjKwBB6P690F1oE81tSgrGxzfpUXv83CbUE/hOS/gzNxT44H922VB8Bm2wKSmEPO
nOjFXMaCOAHQgHFv2AUeX4zuMt8/kFDi9EoUua4RWXFQxft+ZLkqBsnyP/vLDUEr
fvDLkffZPp7PuoYgUE4TcG8/MSFcdGG0V+f+rE0IzjbxkLoyo+1t95llwvnb/Ptk
hOTChxVl1l+D8R0uG+2AjwQVJlBUPC3vM60ixrK4B2Nr0rTRsXBcicCXDiJ6RD95
ge13b9N94a+2fhaGkX+skU9xLuhYzhOqbfFWX0Q7I8795OE74Vl5K/dwVLFLiWPl
uXRrPMkuALSV2Fug21echlXTlHwgA+7QhksrHVC3oawWLNO95hSj4MvvtLVlEVcc
m/PWyxNdVQ/8PU2M7ItYHQeDyHDB5mp5ul280p5t0mvGr2snvomtV7y1wXsMFBJ3
r7YUOYfA7RibRFzcNToaJ0aQsidnP2TMx4oCrNJ84CrOvaylW70dHTHTP1gkcRYq
YFF05Ghx9VbfsdhLUUbAmUjkPXQJNMsHyHH+jGMvlVG/xQHNd1HQfbm1PlrHdBq+
jA/E8PEvNhEyZpv87jqmmvqEmDA2+bMwX1zPEEi/PqnaPmk3z2bUJqSPhiHiH4RF
WDhc07vnEUDf939g+a2UgQUJ5hLU68OMgoaA6JPuYIRVQ0/FtOXZ4KAwXAjdj1ea
G7U9jFeauyfcpup+5+fBQ+jhNfrmfaivWvpkCIMB+Ze7Oih9+x8k6KKD1XFlkzgP
7kz5YvXxNkmoPevsepFajFKcwU9eg5dIKHe2/5rQyAACRVHr9InWQ6pV32WWdzgL
B7DZds2ii72w1uHfSdfz7K5xk1/MQr9ea+7YehYqkzZa3inRMV9yCziQzGq3t2ww
XDFAzuK28DnhKEBIZAQOgfRdHfRUeWgPGX3q3TbxnJ6Xk7L3E76DLGM9hvbftj9J
gF9EX2GQ6GkKllXK1eR3S/VZqz40UlOsPm5fpKCflGwHMaLCW/RYkea8tbnKYD2Q
eNaknjsaHYq9fKxO22ptzyPmo72l8ANpG5agqbAFbwHUmGa+yLS1hAuHkGSdNx4o
z6OdTBLVPLlUzQT0wRYYN2NdMWalbBneMOup8hnvlqZQ38B3pX1vIC3lUgJB1WsB
aeHSk1SkuKCAjU0m3ReqSG9BiN0vnKb/Kx5Hn10AswGNFRLVFiR3q37oMCcGN4Yn
ExSpuRVLbeXsWUdHilEKcP/kmP1a9VM+fOCd2YPyAWJWgFIYEL+bHN9eAYX/9jX3
smaaGa8TJRD0IlmERq/sQOGzE8Qe/uSXV+giGqDwFcWhenCdZV0fbSWloKnr/Cpj
QdYJns8ApjYvx4juBnZd2ykJEs+dlXAJpdKlkXMMQOwtFEiQK0CBU4Q3w5wPP7Jg
7wckEGsDP6/fF7/DTNKYzt0Oof0q5t4FeLHpe8957dgkfY1Fs/3cmh+6Lfo0B3aU
6NtrMxeR306aISkGcUmv7yCkNaIu7sHVNhnHLL6a+x3yjuyWZ62T4bxS09lf6blK
gHg8cAKtdhuet6wq899wE6pwYI99nMOqyNp4To8KpB8xILTUc7k35X8XSZuf17bL
fHkQ7C7Q26cFnjQqEbAPYXwTBsvurMLBxUhIYYFERaNLCTLLsbjgDnTx6OYXwF6u
ugfhjizEIorPVXz9Jsy+HLhIM5oI4rV61W4s29i2XYrk6NZ0lebW7hDmdTSTw2qA
thJ7w4QEnU6v8wxVXqTPf1sZlJ1VVCY1/10tLsG3yN/ZLnpJvtEVRcym8qG9nOX+
XecY4Jgw6TOzmQDKUrf2oHtGKoQ8rz7qO8g75a2oX+/uV+RXUibMYwyiDTud84/B
OcoITn0VNVtn9WiPxquj3nH9rz5okMu8sTsomRrETHC3eH8fizDtt5TAzyiizJsd
Xo/urln4TI4m/+ddg6EURMFWF8OCxrup9B+Nfiui5/0pnFEVE03OYaQtDJbh+cXD
jAvzq2ybQtasny81TtJB9gk6WQ6iRklMLRb7IG60D/WHgKzGYCwEicZnddrMmYfa
7tpapamimu2PqLNsVSO2AWN/QlCptLBZHalJBXBSeTLFb/44yXjJEzye1na8BkYD
6VWrHHKG/mABVgdQdqSjT+FpaC4JXjtjPbjj/RDKKcSnhjDkl6CB87KnVTxh4dvg
JAxlSxitC2Q5Q7mjwEdSKOOaGwU4SKLKmSbyjjeh9mItBE9EPvw0GfUQfBY+QTgw
iq8XiNJjrfSv7LZqnit1X69HaEAmChPdDLhyrEABvBMIgEPd5L1UMnUzhmoE6erW
prZjwr3zf0bRUvnA+zuM4XGPl7gAxQ6lxHj4jzoyqC/pyGhCXAbJ6K5tzPqjBRna
Rcv++6BN5mOowv0fc7crkehU6FPK76ZVm78vaBAJtxwb2yq4ukd4gYA9gDm6AtWU
KpD41oAUevMpOzJI9CSfyua6CvFnYCDMNWzW9C4wzstObmYpvHDg0rrH0tYD/8G3
P1gWPJH1h7XOpw9P2qgRS+JBDs2asOYrRCqPrpTdJ9pRpMWIfJhEzaFHyJZKlCYB
ftz90mrQFm0K3HCN8/5AR0hlNBaP/XLxaNE9NGeqPExPfqGZ6zXnm5Cbw8YlUm8P
kWqqcq75Sfwxf048CMZ557GpU6Tz2n8QmHbGbuPLBxVGLqppgBFH4hOofy6Z7pEp
/kAt5FlutlYEW9F8bqBzkY1XWMjDlkh6mRqdS+Yo7kbjPMCEzDorKhmN6Q4AuQ27
uXZtaLuAwgqMAem3l6saNswHKVSRXTqZSviYEa2h8bceS0EHGIY7gcChGP/ruxc9
kzf+eQv40JkpXhVfWC5bvObKFFIpmUGBMNdYDfttujxtgN18MIVZYfDxooihACuS
F/R0d/pmIBos1qTocPlPz7QDpcQqMN1uW7zQIrVBZRettpSSK+sxh3Lx3mCGapZI
dQIJGe3OEGN8hyMsFhYP2l+Yx3cxD3638iP4uvOkrk+cnUT457UeyEZZFmws7WVq
MBhPOnDsQ88GJZghhKSBgQnOM54ZntzrV9RnLV5/po896k58XRaY8DzeU/vRWdWk
LolicVbc9FK0Tz1WtLCoa/zcnqv0Up+vj/N4Vwe3ZgaehTyqPi26Rr05M3Zrlt5c
uKSfj9WJvlL/DjcWQtJAsmrtZ0qGEiR5nUnptNYLa5WVJSpVqfwaKbS7CsVfCcaV
M7X80yCxqKuPe79jSSzj285D/h5qXBDxzcj/GJhM7A+ZMjn41OfzzoPktQA3BdLF
Io7KCm9fimbRSDMBofSaXjYT7OtF65eNV/uZmzHdTtXv2Y5lQXxNKnA2/dMKJJKG
+ufBiiVVbw46JP7hoAXRRE6pHVxPsTSL7zTivmo4d8Js52/X09uv1ZDpQwJm4BUc
QNDC0TehBO5CJLwCBLBy0SCVh67ZctTPfnOF5MuxFJvKKGCoIeh5aU1HZ/cU022t
IzNmQFtWp864b2eXKEpHZvV4LxLq4DvNRQoQA2gTqfRlvijDBRY/qqmJqQY88hAX
Jc1d0Iy3dP8ePasnAe7kggoOnA75CGyIvy1Yq64qhuoLOaw+iwsOvS0EzBpkEr6E
SoPHOHRKyHwcsvfMTxvgp8ibP9O9qAx4uReGWByHE4iiYTuQxzdtWM42A5xrTEoR
pS49Z83eJ4O1bDl3LXGWZpPVDZUnb+u1NnAqN5+tbz3MuCgE1OrIL7Nefcpjbs3Z
pmePcNqYp3A7fuK/NRWepAiSpHKJWpH5/RhUwHoQ/+/3dwIEXb0yJbi/x9pTlzfA
6BCl7G5eTUIL4bLS0a4PfSwC3h1+Qt6PHkSRXOnUn/E2fJDesv3C2quXx9sCxC0c
4bc1//YS6NASstRn15kGQk2E9w91M4F1aIBsuCbelkrcjn3WYuMp1G41IykIKEVv
TcvM0kdOH2LWWxiHSs1v0XMZi2XBwFzHGIeNp7WUbudCL/rXO7AhbMMTApRloZbF
s42J9wXwyjysVWvdh1q7umi5iUKIU/Cm4FfsKOhD2iYBF7gzNQR18Y0WbdiOw2Nf
GmR7uvt8Sai9i33jpnR8WYyGhGqIwXBzSq6P3xAXccQMnF1SlyMbSdas2nuIEX1E
EHDndyafsGNvPVCjH5WmFMSFvJ4FBTW3Va13s8eNnjevUKGqtUu+cwNKrj13rosz
NTGmLrZV1Iq6fnFDsHxQulbi2TldUyqQsInDd1h0BhiSTIOah/TdeSRFIvNYET4Y
G3Uskb3cTsAzZQ+25sFKnp0ikxZOHt8eE1JX3rHbkbi+CGMogx0LSd/v/xR+rVjr
Hm3ELdfomQ/Fy6RepYou/IbBTmTroCB5RuWlp9xUR/G6ArsevibUaCvoumCRjJuP
P5CRZuf0KC3JdLnPNq7/9BqgrMRpD3ejBd3h0khM1Rx7V4eWKq8TcpHEbuuMQ6VR
`protect END_PROTECTED