-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
XT7y3guz5gvHh0l9KkxyW56H305wGbej2KEQpjyrx3A4fWEvqFcRXmP7AHPSKsVW+55qFCVr/ImC
h9vnsjuAahqIsC+grcQay1oWwkGqBIqAyXj1SRJNao5ZVwVzu+574hApruDGVg5jo0aN/imgzcHs
2EzpV+A7INEVXCF8xCPKQRQq+MF3A9AWMlq3j3GfS8/yZVc1ELyV8OfjvCB8O5mlfNIX2/LHNVxS
s5gJy+GwQ75DhRKbfe25WTHxxx0lDZa1EoL5nARCVKxbsEevF4P7qeBB6LzanoH0EJmehBK9pBcj
jrhLEQAXB/EGj70zeEFC4PC1Y4j3laM9Vk1QJw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7616)
`protect data_block
PJeAzFx7TG5BhaIQ7VTY6VNOdXm523z15bu36XoYNoWzesFpKWs4UNiaqeq0QccAlpsnLPYe6oPk
EO45sKFQAvSVmZL5bZ1ym6zUeyKLq3twbRzoAmilgef4th/t+d6WwrL28GxMPVgERVa+cZxOeS/E
Mo2HAQWPsMv0RPFVIE7x1gRUL1qSBaWe+eBD1zuZ13YVLB1FfsTrIXn772ywb1UUdpLubliKuwR2
+KtjZWEPd3Lwkcb5TLCtuO+CEbylhnq/+Jn3wS+gbWYQ3I+lBMt8HtVHCr/le1+89mMWe0hW+mUF
gTvAkmQDOo7eQgw7S/Ehl/oaTzuwQcvvw2RbnI24+3iyGZv4babtohvZK7xAe6OriYxBITpy2EGC
ZHngkjPFVPTjL6kN1G3Hl/oh8nz7BkdtFJdbYRfGCJEwv4Bk5Dtcrk0+yPlmVyQAhnbnTBdRj12n
RYvezhP3Ddrl/mcOInvCfRd+NJr5/aVrRRh44AcGzUIvXVKcm3UiZlUcrYc6Vk0+Vf+Srxwf+EWj
XzQb6YNTBbrEIWLnxDkLzaPd67mZInilnqlkl2CneLqma6x7l33F6DKI9CCjHFTzvFHg3mDluTTj
GwFd5JbpHU55MDmHowWpTJio26c92nfN+ezkCr9qsy4ctDnp2025cmfRKKcavHpcp7eM/WBtqhrm
R5+L01WN/8mrL2W/+LkqM1W4683v4o1gHZvT6rDzGgYSLGJrMfH/U5MbbchmewZtm93qkX/8yYvl
dA8mZwpYTUo9EAzKxugvl0habBJ6lGHl7qUIR2cz/1Psx0Bb9PL8/PyKxytR4DsgqA5m/WoTExHY
SuHGnBAkhcTHpq26YeX7QrC8EJ2bTjCRsyZr6XgshtYnKbHJfJlXnIsuH9Dm2qYHUlVlVVw9HPYU
kiPrmzV+6ez8MHRF79oxNACQIg/APgr0TgT/dCIFDyOdfINoJ8PvECa7tzS35ZELBvgRxtcd4kb2
X2zk74dVO8mPh3n+Zv4dhAZjZSqz3tSxyXR69QUGRry8YFkf7khTYpQvDXL+icnKpwTG+n5kEjCU
leWQcerHFtpXEus7tlfkWqjl+cZHFP1TUrM5I4Coyq+xKHKsye+F78m7Hu1Xk7LLATNTSerEcEqc
uUpiDVrBT8XMEpD+t+67t/p7jIvNNTFhSbfgCCwCj2T+gaWi4DODd+oTlh4M8E/d0jfkPNLd8YJu
JLO6iFa2eiXXnGn63KB64y5ZoAGpn5+rFbIB7+s697XG5RHBKQP/6I7cXYu94hGrRabjW/Vsze19
FgpHdJU32aqvJ3hRZ2NRPmumnl+XT2elb2M6XkVzk7mNqkweD93pVda22s52LuzkVBG/SzhwmviG
4blMPW5txSJ8uu22OYNTbD8zuf/dYEtPaGfvhBe57Uuvr1yOR8VpqW8WBB40UKoD9jEwzU3HfEI+
qQmxWoBs7q5/7PXVwbERJcQJxp1408fK2BMRxK9d1LjzvcPMt6z50OrkFGwXrUtluM+9SFy9WPTG
tTA6eU+h921uQGnGJp71nvtPEo6eTnK6GqSTAQJWE1cMBspztNs+FZXmDdBaln93YIi+U5qG+4PX
w1EIy6pKRBxlOHwnEL7EjI6ntsgblrJvUOVZjGxj8Kft+dgp3ZoetNmT1ba9CTr6LJG9JF9wpBTC
nJ48BHZ97dFlw3PmEcqbSgYPOC5i1ch3RfXOhB+QcKWshi6LY6dpocN/HAA8QxZDuDzzQqSbC+v9
XJMNqE7ZFuN3ZomK/ytwR1Dh/BW93+NZadCJsNU0rxltJcDfpOmrIE5LDi8ftmlpr/Fg0fp12wVQ
rHTtrZZu2UiTaAQhxTFSavQ68tuBmmlxW5+lOvkCMGtb+2K+2s88vpWoFETfjj8ms0KsGndWoBAL
7CW6JpJu7FD6y3LZ6Dy5N4O7kedp21/+WQ7nGscZClrAtPC4RiuOtTrE9jLHRiyWD/5isoTjZt9r
awUQNokWzgcdzrIEPEQkIrUmpWWXprQOhfsnjUZifIMKNVhOQGShZ4BSEf74ZsdkAZXAe6OynXMo
AIaiwNO75H+J3plgxisLTF0UzlzxO4e3qGVMnpxYnGycT6aspx4IPqCOTNK/4I7T2RXLIPK8Vlet
uAOresSmpcjJXN+IdheAUttRXNrgW+Vj70oMQ8Yf8Ne1I2Iy09AQ1TRUVAVdw0AHAZvwybX1oCzf
oZfM4dvXKrvZgBRBJKgnNAkzyHxVJliUi7XehrPJliTqtx3nhjJoWyeNyy37BnvNztv1FTuAgbg1
zH+ptNH0svy6xfCLy22XxjMLCmItv17rMBHp0V2RUgzjsIugffOSdmektr/2bO3zd0Wc6mna1Dq1
xl/mr1tXHpSOn2+Uz9Ka2Sr/qr3t428B45qpAoLeCXEsp0TyjejcVw/v/UfahWjUn28S2JQWmyf/
TGOMKih69fWzDofb5+sIXR+RWRypczeTW1w0shCcAg6HDX0pkBi7H8od6NshfSMvu2BcDJ2J6WMU
g/AGi43ewBQeUJ2rfVd5ZLuzZN6FaVFmfcDZwKn5xeBerkq63jGHwgyGJFLkq0f/EMONtXKFfNZr
/TVd6lkdYGqOZiBY7aMWlvJJiNbyZO/Z58+Rr0CjqDd82bKFXz/YYJcAC28vQJsY41RzzYCC47pB
7AWdbiyYyTqdFm0LzeWWFhb8Fus5mnG1OnBRG0RcYMG+MCIiMP31RD7uQjeMH4UIJGQvlPRySZUG
1CkDYaSCIPqK0FTm7bU2BCPTI4JsMpw102CpI2Y6Ln16GKrD6B8Sm+QceZFYQtXhRJoxJsvBdpWJ
mquMCRHm3SpgSFolgAxuLByf6vJfKlDceBACD3a7SskNCfk0+G6J6ipozxKbWj4ORSm4f7SOYgXJ
ya8lysKfFr7hAjqfHcID4skJTL0jnCV3Ks8ZAgMF/fQPkpKKWflsHH2PeO/3cAir32u1hccNWGrW
RBPb33vfmN0QrzRU692ENaZ3U7PgMFaUwkwBnYIyyIPomlXhVJsRRBPsGw9dbWNTSTI8uejHamKH
BuZQunnM+Vee8vPcG4lt0SGMetCB8xxmt/1j2FGW3nma/cLyxsJWESncCH68T5qqpj7dlO5xXuW0
GyBOa15px9Sh+yNPQbkVyLli5EgKmgXZ+PkpQUvMGt6w5vAb9XCm0zfFKXAHGEmp5ymdX1PkPLIj
6JB4McGZBRrGgKagZBl8oJoB2Xgd941bzMmS9NHoPvP+UEdaoOI1Kf/9glIZd6P1KbN7tjFwVK7t
5EMSJhT6bnE/JrOZEABuEzXKGPJnro1b1eGHNGGHBEyvuaICmQgb1ttyb2H0f0oqIIK1Ok3Vyf0w
l05shH1/azjZf+8u8i5hhGnT45ONFRd+td1SPl6M9iE02xwh1sDH22KpL4UoS0W9wEL5nWiN7lYG
oC25r387In7S+VBqG+Y8UEn+2Zkqnqf/trL8Jcy3sjZSG0EHhlbDXsAa2EwHqJd84/Q6S6kKe1Dp
m4wb+/+YNtqpzMWmsEA6m1CjitaPWZJEUn19fIgK90ZM65X08fu0IyfNTehTfW+pNmyV7pwGt3/C
TT4eyV93w4zoMSbYwDKNhi7UE8MpXCmiXXfp8/lZzkmNLqeEAIY70juAofdY1Eofj4WSY8vKuboL
LrWQ+ofn0/CpCCmSRScBhk50/m+m5119a6mDnxdGvBxUh4LMmKDmGoXNQbhGJgsZa/lTR5f35mQF
mL8vFKu1d19JR+qTxZF/PPinbQdffENmu2QnrvfpEuoneMKBFR2lecmb2nn7avvhfmkcKOLyoEGu
gTbrvIDxl60bbtlDDA7t2pX1KzKLJ5Pe/4m+s95lpZMG5xdRBqY4A5qZPBW3feqeMB5252ZljlyD
XRauNqwMFoT1igRqBEmDHfvxM/E2+8GCRVEcI9mchG9cXqUtqVh83Y06dTcXMcj1osMcQlaGlUH/
xY2ehstL1+Xy6IkOzlOM0cIVw36Ha9RXp15G2O/UaO8Q14RBmnk8j/dD8G9SZskjr+ChU5z990hU
TnUzmjsWmtA0MVjelWMnzRc1XX0JqcRsq7yZZIjUyd2mmFdRuUYDOexKNRWjMKX4kEcJvdz0HQSv
sTsaawAfKXB906gUcriep63IMPIb5rxvpsKRraGcvQ5Nc62J6YeV+xujnXxniVL2LoMI7N112R2S
fkImnjLV2klcef28QgyLrNWvrS7yQbQgJIja3ghe1h9T844MaioEiRSTOqqAB+4j2Jsv4tQkFGa1
siW6da380yRfwDteCzP98waqq0W0YgLfXuAYs+wapSfnrKCMrTnEDduu1+EeynQe5/aNhkMXOriw
P4caVIhNM4anAc8EbJihb/kLTKYZJ8dBTqmIBYolWnbp+UUiRHQzSRS05/H6j5y97YFPronSq8i0
ihRmna6USxUGNWAZZ2QlQw6ujti4m/ER9OuhJ2iykqXLx6dHRhDgRR693WDdoSekdY+fF7A7j3IZ
TyvhvH63zitUvAE+UAe/sqYTBmR58bPBmkDpHFB/uJ2mIsWK7+TxuNQgq3xHq0omMMXLwTAbSM8X
Bet95LmzHHDyOknKO8TPiGiA3PnTMNYLWK8p+vgC+UVp9911x7d7ajFfhgq/fz3HwB8qKHocg8aF
GxTTt8wq7kQtFG45LTwMKR2pjOTq84VgrKKD8R+eC74Tnerl15eS7MCkYe6H2g5rLxgEcXHcO6fA
vDVyreO1Sc9h/XT+LAr0UGuDDFT7M4n2JA6ZRMue1UlgUy7jSAgkQSOlXsRZ+9va4pQLvkT8n4oD
q/LeD5JYgy5meGkebtPDW7unAzD8ldoBdi3vjV/y2j2Mzc9h3M7sON6A60ktHXEXDot1D22KL3BN
ah/6GQKEH/tfcAxridxgvxhrY0MYZFbDSNLuh1BR9/HFn8+uqmc3S9vpFEv0Iq50tXCf6ShcVPnz
1RzKZOQw0V5jkVzdbjYw2WAIxox39VOC4kQ8GFi/lYnefZfiPPPeGGn60PZrtxndgcqn8TItM6Y4
2yqWDO+7C6+cMZVB5zBYwK2Yn9yJO8a49Gfn9MiNmLnB8dC/PeDMw33ixb8vEGubl+TTm4AHBPx/
3U33Nv2hxmzB3uX2jk7QHOZ9GSZswiaCZi09TA2eyycYlWTlWaBmONIhxeGeUGchILOfRaIlS+4C
NBARaIedSs9nYClRkB83nfMXg1YLmm+MQAY0BSsxp1wEdrQcEz7WcBXfYpBYcL+JyCQ7AJmCc2a9
ZE5TruQIIMYqxtvmU89PC61fz4WhneVGksWHvuoV53s7RnSMYQqqG/SDyuTvwi9cpeAGd3QoIPhB
pjj6wFhQcb//Y+BFONFIRe0sHMjDqS5p5hYPIWTF1AdShKKNeRdv/8pgrL9jLXhyysODA1bZ7tet
sRPCkgbOJPqEGMhSvJq8GQih3UQXmdgc33QPn20e1uWS7quniepU1jMdtd9PQiYmzT/aA4sb/HLu
3BK/g03A3Tw+lM3m99avGkMDAVRMBtcrA0aXY4vrLmOjmszN4pkqX14dNjdXY7F2x5i8ZaUBH61A
5SfR8wzstXdRZf+kv64i6/tWsmaBRDiqt9zt3MYZy2jBogK5+5iIjwUVqFVT34pTeFuffxMKN3NV
9VFSCHHIsEoVnQnuT8TQ82RcEkcxRNBcBq6sBWDNokH/4BVofezRLvQXzvVgCY6yDA1Nbl985+vn
JmnNRewhQRIBe5OKcelI5Gh1RqYIhb9YqqZqIK6lhZV22WmlFraRaZC/Dc1ldC4Szwc8zvQlCcV+
jszE44eeXnbaNEyiCtsdwV4iTNWCx0jwuk+TYcRjMEI7zCtcJQnHwl4j2OImEBuH3p//OYAOmnmN
M20P3FHuZ81h9LcewFhKNc9Am2NgepeZ50XHf6z9/Hytxtl1wIIO4TafhwGek/yr6bDrzxwwTKap
P411y5s6XbN4eTPAUafSbX3lVU9riVngc9gzYeURnHG/JTBAjXj3riG5hJED5qO1bmwEC39r38pS
IP2OrB7EGWZtwIckdOVIT41KkZ40XQrTwrLwCQ7V7F+UhWcQ2ZpYok763yx82X3fMqTIsohW25Y8
cJPOfo6QRKv/TcJ/jgzFEUyfoyYmM10iwBGo99F+Nw01SrwKO9WUfH8LqjUkuykGRKCV33dmwj2a
f8A9louWPtLe/EYcu9UWGQ85cm1hlfCv9EBNUGiLKGSpH7yEgSMvGYyouIAf/8tu74egTvvIfOD+
Y8yHZAv9rbz77jrg/N2Kz9neKbxw0FC4XORKojMnEMyyLJujuT8f+RPzNWSckEa/+Ss8DhGPt32e
e0w4whnyKj9acqjBXfUdm8U/W0lEPFtjgs6qt+Li801Tf7dwMgf4itzH+zfy1ubzex2+6H08joo1
DyiTs1+nIv++artxV1Jq7n+aBqzOyun042C857vOxzE84fJGSPdEau2tr5GkFJWWshyC/ichdy/6
AyVRjZXrWomgCzOYUkF4VqNxp0lTWDTbeCeDt6SVhTp56FoeNdkXAdwIAYU3U6ScYFgQc0+BfqyF
ak9psxy+Poe7hBbOy81Cq/DN00GHshIY509K468/ZAX8eeYgZD90YaFo6rVmfuVO2vovRgGVpnrh
Ph3sHDJxMNUZvJeVQpVLv0c9XYKoeHZShP0Leg04M6nv28+yknQxBnDevHzVSXijUQXXBuT5Y1a4
lJLSeFuHOemANPrkw+oj3i/o4sdjVbKxR0SFLWfBQCDwDk3mMm3xJxNeJaYOMFwkeKTVo0A8ZFfA
ClVTCpHrH9X2VKRs9H+jGecx31DobHvWuA0GzjUPv2b0b3Q7u3UKFL3aJrNQ5akJu9qZZXmkX7PU
mdcSFdnGwm94O6MA8UJcttBJKiea81x6uLO/k+oETvleBfy47SWSGPykgQ9MGtLLJ08RE2mp7fyG
iaUpFZR2EAi5AHDQZv8G03zYfBr1twbYmJ1kZPhzPQisjqk020J0TCtE/g0Km4exvkjBwQNBxhfh
RHGE6fXZ9VEwSJoiG36FwZ3+SsUENko6vIbJbBBXiYm1I/b/qwKh02QdLxgMKcTh2/WhXbSVc6ek
A/u2trvF3Yr+lPuCe3ai1AYUoxCh8Oi0la+vdQNNhDOVbw2SKrVpS98vz4tAfbVrS/tnuCz9g5R/
nFsaJdpKsTazonpUMkZo2Lqy+LCUU1FDa3YMm89i4hlVf9Louo0PcR6WwzH7WvPRUM53ToSvAzYz
Fiu15yN5zFe6Pi9spMgV2uEqaX8jHJxAN5PD3MKK1HdB5pRFDp3u+8EVAYqIGHIwLWkAsrgv8Jjo
KgJKhqfA+IQ3AwfQ/V6HaZRz06sBBdIqKfW9N9FFRBIXoriSb7bjugAuKzy6et+v13Y2mBixopfY
i1SEuezAy6uamL7r6jd+bIt1DoRoR/O8yQPue0ypA9Wq/v38RWS3jOvRECUdJWOJm5ptwkJRlVZK
uRq1A4Ktb3GCiYB2wz+MQ1CieSP3jVHJNq7xnben3fBxy1P3l+1UimLLF73lOmhiuOlav6xiSof4
2DM0FqMvyHm4S3VigBjLeFjSG+FA7pVCpFveYijOuEMD8z/wvA7+Kyst9g1XhGe6ajz4V5/VKiIP
O/LEZkzmvbQmFCsfZaJFnHA/PjDawzaxEA4DgxcY7qzkcgsRDhoMFtjOkgoIZyL3yJe1QFS2oFDS
VW3mEGYy6Z6qEjoByY8759vIEOmu08KGBayxnCaZ6J5wNxgjlrIGeXnZQKi3UR5wL4IFC9Cm4Dgz
DZq8H8B/NpBc94U449NRkHv0nxfceOjgK1KBa1PmTNeogAjCWgrKlH8Q0igJyoK4NY02hpB3Nvwo
7f7njkhl1/WyCpV9HsrQziYjza6yjq5KzFqrmaNxWgaRbW7nbTBBYG2us9f3PwhK4EC8VEEO6L3Z
Bhd+YL/EpZkcT3uuaH2sgVY2ChS+W4+kV0pjjvDBRQ50kw2rzWh708iq6gFl8HhoTB4z9fuGi5Ip
SVt5un/3J9NWR6hm7wE/At7P2t0Xzc8DPwsEE/DwDXReOQ6QSXaA/yUHAw5+gade6r/+mPzjWE3+
jNk56aWATRsJd4RcqsQg0/Lgy6Tm5KPz5BWlyHxdJm9W3yeQ+rlj9YiPlP75tnBKNLqu3dEfCMc7
7kMsocatjOM8lwoPm0ekPG0laAtN17Uqaqw4oS9qhYmiYIZEfFprGMAoCLV7ATjO+4gF2xf7bl5a
kDVCozeQKF2PqKaH+6mpz+mrlkePIkPcUR16AdnDdQzdtfyPBXse1nh1iKmOSyar+Y2V5bY/wofG
qr381/MgUmjq+xFekrroadddJQ/HDO+yq2CU5pM7K+OaX3dgLE03VJeq7+FIXvZ7czm3bacLOVap
qY79X79ZUOijdELwYvRd/L7sPlG17ZtIgS7rlVRJc9Eae4M08qQgLBmrOZ1saXBGng53CVG94V+R
B1pnxaMwvfmjvQrLHuGYVBhk0b2Kje4psOovlShk8rXy6c8kbOsZH84pzgKt+o6YMJhGJ0XSxl9v
d6zbIa30U3jLX7QNl7dZu9UsQMU2dsmVYPA6hh0e6nvtDCDSbsnSHl62VakNIAJQ5+rOaRXenlE1
6R3fCBklE5aS+hmZw3q43yb7lkoXaJH4oIITAvwJZULvvxawhctJ1caXPxe48cwF6VDEGVqZVVkE
eJ8z2KrLpnjZRSppowSbayaOQCAAu/Y9vAkzuFZl+6CrPj7V0NrSCGekc6AbuG20F/2S5ouxyuoj
A26fF79xZqO5XPsFtp/Ief81OqpKZA79vamsWvoG/xpqA0lmRyGVDEPgnvE++gjxFyaxMlZjNdKH
X3E7bGdLPrS/vMQF8HaqzIXewM6bSe+pjoPnarB1R6YtNXSCgvrsNeTnLoJQQLSsn0ZS1bdQiBEA
Yr1zw9gm45tDv3umDCjw7VW17op9l3wj1DaiziJEbEA6H+7P6CPYHiXMzAbXgJVKO6Q7uMQcp9zv
zI4TTNhnrMyuyB+cJfcfGDmGeAd8L94o/gwQHqGd6BWqMLaet2Ze1qypap85OREAIGCXmBAqjo5S
RWqk6r/9JwGCnNFC3k3E8p5Kag1kbXTvcU0eZ2sJHcYSK9D2uwK+NXwygIT/Z9wDClS5TGv+qC6w
4xYces544WZMlJaZc55+Gf8+xIMqLFeXTIiKEmZtP9JaG2FHXOAAxN9NuYJ0gytL7TWC04wSjwaO
02d/od0PGvUR3eD07Fu2B3CRYM38403fhg9OwWLN/318FKrpYkcCWo2UnjFAFfg6Px14WjMJvRVW
OpDhhygyo7q0ht7eihsIpN0V+20uNKQQeDz2xtKmbhwffW1hEnvDINNBe3dvGKtdhiJ/88i7PvX/
iSKOZr48LNv0seecppxXXYd8Kr3L+bxuEgzwJH3lnUTxfucaX5eSNI47iELjjDVN3BlQRn6IXUHh
ay3bV7LdJI7bYVacm4HDxmMY5F9edwjEc2S4qAdSKnrV5Mb1pzBn8QyG8B6Clq8LErX8d7g9vR0D
DQFTlQMAcWs7Fsq3af6hnaeT6IM0t/T/r1QT8W/pYrrpXX1+y91IFjcX1Wt67GYImzRfLTUKfI/G
p9+89cNfSZtA7C9ptsHH9YCacco6+9BaYpxS1f8vEkfpTJbBNuwCq0EqaFFTpfRU0sSGNzvH31/E
k/9DVr8SNfUokaBHNRYZbhMQw5OmfkW4AVKvnOOOR801btrJ6h5+0S4ezp2kIKRaq1um1w7TZVyL
NuNNUQm1y2cTr/9nyYoLTii7gcNxeZhGJUeEgHSKwKXXBWbDOoejxYWMefPc/ANpKSe3kg/hJ4oQ
QbYrUiKGpzxZJpFpZump6Kv1EwQcprMSL89B/t77ovxbd0AnQnX3bikhu+zl3M+f3DokG8zPPP22
gex3GhIMNH0As8B7jz+g9BPzAU4NhmKSRxlzEtkCsf3Xzou6vmkY7PwGml+ZtRqTRE1lAUsE4470
3mk1ypAacW+s7GbVQr4+U0NwgSgv7RmKPoeebmwo5rT8wA/sv7E2+rELfJD9o3Cc4yYffevlve46
ckSSkdXY/LtUbhg7ipff0DyvJSm1yQWCaYqyLgxOR+7+IiS+ieZmwoNp1yoBaFwlBGOoQucP9jpW
j+A6v5QizLVYqoL7E8vsxn153zgFIRox4/2htGANnrX0kPs=
`protect end_protected
