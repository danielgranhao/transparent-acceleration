-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
WVBh4Vny4waW/PS2X/hnvy/fnSO+ezDDkPOjYOCuL/OC2uzq4P8poSPPMwY7mTnJ
05c4FmTsXSGbPs6v6DqdMvj5Rzdv+JWZ9QeA10piAYbFYarUg5Tf4Gi5N+QhBQCa
gjRAhNIGNMnb3Dx/JHG4VEEHumzzUg3kskYIBK3J9ds=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 41973)

`protect DATA_BLOCK
O/18yNdkF3Mit866mYl2+Q5bgccCy004zp2V8e8Yoxx4OPvPgAEpjEqrn31V4Iq7
BiLYc7eUzLbd4hdBjTfdQhpf4nIWacYN1OdiuoF3m8Q4rUb4W0y+zyMKCnX9KO1D
+xfb+smrRgTZhMWCjKPDYgNkj1BnsIfkksyAvKmEu7ozIXvYV+hUkMzk0lXfCp6P
SIVH6C7U/w3S7SNKcxRhlyZodI/Yyi+7f3pRvuZBv7nnAF7CXg8vIFs+IzeDvYwd
gby1aDGtjhkZ0ZGRTZ+a7hJzRbW2Zsm8T+7WB9ueGnSbVI5Bnh5GvNheLfLCVI15
/8bm+FSHzpzqts/nk8jjhX2jLi+uIn0DR3PnKORRlbvejUojpckcHksYp5YvlRuW
t7K6HLU53RiIthja4WjCp/ZH56w3uJNd6a/9bhdin/NWVDzDlvP9u7B+wj8Xco5W
noOwi1ucxQmHcTTP2lWoRSjsfkAL7cpCm8RHqI9eKvpv4WSDqqXREgaH1kLF9jI8
7aowidOwEeY/jSLJ0JqZ5GEgyeRWrjPFts5ulAztJmosxp3S0zihVUk4K29yvHT7
1u54fgT4KPI0Pxs3mC1lv76bCcU87pT2eC7iasIRehT/5FDgOqqEe+Q3PYD+L0OP
cePeh6kcyKkgf/MDG8eMzX2js+On3/z+wvKMJjZtBoWmGxQ6FaaZTH+VO6nQiHpB
MRlV+jEz2mQKkV2YfL3nypO6MCluJapxhBK0Zw+K+LIYvDVIb+KknALVM7x/ExDV
7SYffhXKt2A3heDdXHzFu1ihsAEbaemKBK8Qd7t9Y3aV0mmHkuMki/1coB2l2Vct
qVBOp2bNc74GhLdt4rBWlJvtls+5onNjgChr5j0V8eUJGsSdTWs5sLz7JnZg5CdH
kd/lwJvYzdLbmrLPAeBKfcHJtJzrs0BnZJaruW8l8sib7ZhFtKte+rnDZjLi5VQH
Qu/ojYfpRpYzHMsqzyaC24wf3AfM/5YDondwBms4hJAdksBaPnwXclRpev7Uj5QT
8wf7T6P1Wm1C5DLPUUZjQGs6TVoGegP6XbuA2ow5sKTexjTAhAEqSm6VMRyPldVK
Pa9OAwXbP0lknPQTcIwvD9rP+MTHFb4Y7ubzHKp5Bmerxq0YjBUHY8LqYpvKA2sW
ktkjhjWrMV131l7bpcV0FkkqdNOPachgKN/YgidKdYggOWD6k9rL6A4jXceV0mrE
aYTu+aY8GAdjzRqnePfB/fQWgEECaccmHdATtdlOp6vl7GZoklJrv21RaZiR1She
UQfwdAhc32l9fl9/EB4+2V2ETG4gjNIsVYnTyWgbR2SKmnHF6pa5Pi0bCA0Wv35H
ACbZwqOAjXdS1PmNll/EBUQJ1mNPbp/2e+g6e+gNFWPXzApnw7gYFmxEvFTjrDsR
IB2bj/OZFG3qlZ22Ghx9jPJzG6p9JSEOM4W8R2lVn53YmQ9X2fNBcBt9XLubhJx8
RrOwMGhKvHlc/lefyXLVc6Pzw+9W1SPVhXnsvYL6XJ4FnXGM/ev5T4cknF9Bz45V
T9ZImHZ+c1bpsX5cXk8IYZdWeek3dIFX1h66KNtIdSjUH4PSPhUuQ4H2DuE1nlgn
Ik3vRhIColeLQjDVXO9ia+kVfMWHwqQQ7/r1xkxkZNkM2MoBIux6ue4ZMuMD/tEe
mag4UoHXAoxFPDRaW8h4AoTDcZ7K4BIpOYnZ+GAuGB/PBpbCd35i+NixU4NniZPI
YQVdZqfKigcIcBB0kmsDIGd11gMFNf/0Riw3QqFKE0Vz79E3YJQi1bgm0VMuTq7E
0lAUYvdJEJH7UmUbdWIkogRjar8/r90GbSmDTaEEXLE5aAIZvWrBOEbwS5zCG9aE
+wPbQTvYZ7fTfRTp7hb3viA7fWOCf1QQNI1Qjlyi/RVbRYstVW/ENkV7Fhe6dQs7
Fr5W/JBBmwiYdH893QtWahbibMvI3kyFFq2ngGH1xxd3IPlv91c/UlPOFDhRhjmp
axp1NaFCx8c2XUkd37ufXaZpYuAL4kC0MJh76k9ZNvSTbd/HEx+MAnvDWZxg3aec
SoXstfzJVGKwOfj5r2PAfO8OO/a5cCo0UmYf957U97YJxc6d7xoIrNSmDSKnhHfj
KHsLSlzXcU7yJ7BBs5mjYb0J10GMmuZTfw3DjUJOi+c6v7FmUy9mI80QuIYxLoyu
dxWI6cXFt8GsHYUbnqse39HtCSpG+K165Kpf05FX+msDMR2koGH5Ze99yRavFAEv
khS0d0bYOs+Sf4HnzZF8HoPvsIMtswJkMTi8yrsvcUErHub7IlT+8yCo6nlw39KR
22W7a99dYOOtLdR2jiZUS+rFZX4cgsYjHMubQAp4cmmtIX4ykz77SIrSkS57slmg
plkV3xzeo8RtmxZnwKPnju/vohYQoout9udtMEiyAcV5k9bCPjprwBDRvN1SO29f
/LSzZ01E9P/KPbz61UMPQSVPh9XmNj4KYGOYXKBgmbI36CakkI700VAm+9tiWFQC
rrscWp7/kLqfiTvooEv+aDLuz9Ibhwd7bSKvYWjh5DjzLt3F4UwRhRs52It68qew
OD13GlmEkVhYLQFb2glx4l/jCMXx0ISvvK4NRl6LR/UPaD5wY1OmUd6NyLzldMQf
hYLiSChGPVhaiLCuye5wHtTIS5fQnlSzmyJly5GjEq/BzqYPE2ymVa6qBgFOBg4z
JVgHrtA5F5aptUwkZTctxF96fJhO+2YklR7J3fQzZMP2gFu11WRP/4tCn9Sq309p
3S2h0FeRoBZ2MSHpDZtrfKGKtwfY7BCcR1v2815gLXtexDJ1+T4jm3xP+Jd7A/L2
cB417u/vm7zLW+ivK1VLdIQtyNC9oyri2kx+YbWXdmL0IzGcJMu9eA51GjQpTqa9
fyDfswshLgn1gPYzsyuRIMPcG12WnPDrlRPrPjFqRJFPgpHLWRT5J6w/KhEOlpK8
NDLt8LkZGFFvg8GExmdfMIev3STbpfsJUR8pXv1NcyOYLeYTQuNcFzWBHqcKXUxW
6tH1mW6NuiqqIyx4+tsuJymXaCn/xNGZ4SSjzqEm69WeQ60XOIcWPpJmkrHhJ4/H
HIl+KlrMPuW4ze7EyI2VQRxSG23zRu+4IGdWtwOQJVGe7lRKnFrgs0TCTfVVWHKq
1AkfxQlq6+pd0AmCq5YCiSWwVszba8Hb5uCLPLVI4TANNsLAAktTi5y8agAroJp+
95kIV2vXcykejrg+ZBnLtLyFL3tFEz6Zaa+drxpOf6e1Qz90nIjKWsI5HxceqTxR
GxeTvgAw1/wCXiF0JxQJpXzrLuJul1UfFR//dUYaZ3MiJGXPhQz4PVG0VGOKqU0n
UhlUzzzKDbGsHh1/ajc0vRYQXlbZwN06op6QSmVnIYuAf+JHUI1YIvY0eS9Lh4vc
jwMgBmx7Z9PaYjZSyx0rR7HVLAhHNo9syde7pVCdFxfcj4kdgTRfYMK9FFDgMlML
E8dItb30NoRWuqJuK+xo4tesjPI5FJZ+gd0lSK8qLt+CiHuNzeoyHz4NDtT5Z+sa
Qjwfyutbqtvfk7k07dgghhYDVjlu1hXOGVya3I9Bnp6wMLqScmLI6jDU0qJC8evK
CQsUMvBhPbHxVuXR4LdTC4Ulcl5iRO90ao8HwZhZJcTSjxXj6HQSAEcI2aujEkGv
Sal3ag3KdVd5kDpy5fLSBc0WM59BflEvNpkEbEjRldZmQHZTC8VqPZdQOWku9d4X
vX5GbwbyVWJ9LEzIIwOC2wLNtGQrSJS8ob0hY9SlQrnTxfFKViIGfQX4fGaayyP8
1GFoYp/PniAVyWFUFjbEnote3cv2ETrUNTTq5g14ksbknUMcByOLX2iufylg+j9J
/qaFfw9jeAFmuglIuo2vzLEP9hIio7c6PrnjPjOMfUTjepp2MRFapZ1T7/BMPvth
dUAqzXo1hfane/dk7mpcPcPgJOdl4ZyQRGERv8MTFBsP4bUTTjBNMa7Gmr1eJdbE
0crh+JVlZxVIr4nkm4LBKzeT6VwblxahjYzP0Oky/r1JGTOpEMSmmjqGOTI1PU5Y
JBeDzsBby4ofy7+1D4Fd/ZqrIXAzSCdPm4CMwGZsw8QodvxX8my5++d82bzQijiU
1P3yEr0Dc64pO6WhGlGPT8bgnmyFsPMwcEWl27n4R1TLehrpLroT2cEjxRR7ZxJd
jDb/lka71kaLqJecxZC78hzpW4QunHHmCMzZ0ttUmMQDvARvTF9g29jc86CS0FQ+
R6AVpjYXLnrPAZvTbKUkrhqJ7s+xCby0bSH7jt60lRSzG+ZPUbCVwfct1r5QVAuc
QF1iP6N9uVxckaIe8dnyLNKX+G5wxGiL+VUDIluybIMPaWJQBrNuweL/392xlFlw
aLMXs11NDsDyXRuA1rXjesSIp7FP0/amEd5RTGPS8THGyNwFhLST62YxaZH/iMWP
EsALjHUvHPNJbwQrZV1fzw2+/UK8hZksR9Jd/ro5kT2z6Pa9cWsPDGMcX03QJrb9
rApfoD7NIh1u+4kamFhO6uULRON6qZSISakWChxLAsBW5TwmPHBCcTGfTgdaP6o7
dw+Z9k6O70RCWhCIKWcBhXR4zPrGydfXvq2k9ABEzPSk722c0k37FsVOKIVMAmDq
zqvnslnyaJGhbZHDsW6g9DhZqx69V9dRx6JEuT4bIon1+JO4GNwnektX6pej1xBg
ML29vcxnuVcFpEcmPTIEMEvut0BbuawfzoVGJtli0iYUpv38OZw/oMXn8l0V3feC
cK6mOdBn24+UDcc7/GAU6i053RULMq+dSgOpPnEhrJC5ywvJI2AKf6XFoWEvS/dv
B2cNLhlbgR2lOWNyR28+E/A9zl3VTL1EWvQYSh1O2fQ3UohQ9jv9POYd7QGniWvd
q7IoDcdElp6+rNpjbal5T8Yk6F+1aZn9yPRxEczuq/n7Nbe9xT4j6ZuIhFPE7Q5f
zURDDmcycU8r+qmqXcmFuSDt4+iH/N9QBrSbK17rF3m3RHVwdXV1q4cZHeNMQqkc
6O1SoPAuV7xXi+Dmf+8rRfMN+bKgqCTOB6O+44I1AEZC1p4V4RHOo6/wPQy8TzGs
lVEZrhUzVq5IlxxTypmB0eZJUaHA8urjK2neIHQTEvzwtnK2EtVHnuUrxHQJ2a8q
zMRfQJ7H/0jpfGusB55tktxgty3gNkfdaarZEwXCGF8aUIwQ8arEbuFgenEw3piI
oEUFSJ5NOZvdjLqJcQa9yLvKGggCb2mlpgHO6XccegA9Vvm2jnD8svS5g5+XH9Ib
FenFMZz1YRBSv9unSsY2DYDbJlQSw19xCmNC+ALcRxPsDlSjJFxkY3KJhvJ+YzGe
X7L55wPe6Pr9jdLRUR1/kxNHtOQbtsqjCF+SshSQlcHl7VJS2P40rO7/q3tEG5uD
NdBKaEuYkMqYx2ju9GWVgX7gHN/8DpAs39xgG32vmuhCwP3aOLSNpdn2fDkPaH6j
DCzcBzL1bNWVG23Ya2PMzsc6jP6x7e/anmz1O631NSRvKFNnaRLci/GT7sopWwg6
VmswmXrSyF0yUwa1vKBufvnDj0Bx3yv9lz3RAfbdnigaZ+T2mHqNIU21LLgU6NXs
UeSXHisREOjSy1J4JrV+RUVS8wvVvT8Pk4BX4b+ywjgEJs9SkYXejEn6HrvXPqNi
m5egeOdRjtHbBVd8VSohceNUIIkJx/MX9zzRs0v5fVuT7FxHHUy/IdB+Jwgn0jXh
VFGujYbgNh3peReVQTlhyiemjlNjkuWn99kmMt3xPcI/JS2gLNXzXVB/9OJro0l6
08H775xJ9opHlfSYQ3cSbPUoKrpREOQzgRusfqNHLEaozLtbalW6vwm/K3Kl+xAw
TRIKUae1ZgGcY1Vj788GO0TnX4xhWuvR+TqnhWVQ36qNcTdoON7Y2gOJJPizeUz8
j0J1K7tYDOsOSbAoxmoeFA29jSEf5hrk2qJaO6pKUJxHUKLlCGLSQiWKyL3DIIhv
/2KZBtdnoj+sibENZfMXe12K6qAM4LZSiH+YX6bbcLzW29omnjHAbF2DmOG/8VBA
7BFiB23iHDmKwH8U03l/8s9+tfui6mHThf+2P6Gfb6GEbp9EtFINXW/YNZGA/AwC
sK2BQQJydDTjb8p0VVrrKoOCx/VJvkvp9skCseB6LaLX8lp46vH3xYSdgQf7poBm
9EB0cVz/ZSJI/8VC9zq5ELKCo2r49YyBbxE/snXi+bXq0Auf2AiShiIUffKW5gAi
lLkVibAFwveMm49HLmTqA2XGiQBI/zWuupEgtkaOEiDOWzyIpwnU2E5bGaOFrrkg
wgnePvKG8yWhUYzTDx1lhllg0nW97dJUvZcDoQULwRMIw+pWmtiaJng0nYVVU3KV
MAtKz9av+ZyER3u7pT1GeGpcHvap57jaDykkNhmQOu6hoCLlv2bbbG3Jo9ttXHos
+u/brJzBdszDYoO9qzKx/JKgCQaMFQ9V/VwndICbSRevkQEWszFBD2R5ysCVVey2
0LlS5PN32Azr3op2zX+4MSo/0Zos/thjcnLrKfI0VcBgdXCPksjxqLjORgLz7CJX
9YEJ+XlbTpk12b734cQKxwFz7rBHMi+d4HTS7YzmzL6GAywlIdItqYzb1N8uU/Y0
7+FEDeAxLF37Wo1lFYrxval4NkU94D2vOLj9crwiClgpWQpqdV1I23Rqd/oRvPxM
26lpjXuWJH0XWmWXmSYEi4D0a0eS3V3/NbHUV+5YxWa24KE92d6ttrda1Z2uRaSN
IiWxjrWg0d/AZ9WXR3zn2fWHamOHhsc/FeEcls7JzfvmtNiLClkMnxhQcMz1e2yd
T3LA5+3RpqXBzYmOEJyzSVY7p1h8geG+pz48CNC5swQsTxepZZhnTcIxZ/a2Jp0j
mx79CdHhVrUGtlh8FrXeHuCKxgVr5DxqEdyyabMUHd2KU299ZH2n66IK0U8To1wu
0ua9uKOYlpxBcd6wmbNDCpQpV6fwaj9WADhrUhoo3/0gIm6htg/Lm/AhqkNZ7WSx
AbQBIXCXX6pBvOLkFrPhjfwdqoAS66pgCi3coJE0kf8qvycYmBHP28MDPoR7zLqC
ESMdv0mAX7qevcyWHVhT3HDrPtbcpFmB52w9nvIy1daurBcsVZLWmlFzgRMPq9Sn
98znLyBDmwdVGyS8mqnCSvpVJ48GSUVHJUvJ1Tesecvp1rXyEVD5o3JPB+1Wn8tt
HJ+uvwB6zwUgKADyynbf6wxf2W1J6cucZxPXLx+DHsjieCkYE63TGn1TsupOKHJY
dEHFjnFzWROSGpvhgCIQHSGjj38N4EtqxC2wxkgX+blftcIefoldx2JeEfcpTcOH
FjHSvnw94+Qn7vmGJsxO3zcdcyji5twla+feZrD66YqDle9T3nFInwmNJMsxbF7W
0ZPZo3IU0Adf1f+/40aCSeqXl9ASnqRabzmu5SympYUsXArlhr749YLatfXJNgop
G+8B/IDvk6sr99NRqEpCUkRk1335d/oo6a2bZDpe79o1Olrdfczds4d7c/FBUteF
eMWBg6OF71JNxLjCtMyQlbiRymoVn1mgHK1JT5Uo1DpWXmNKbtGRdSmighvOYTI4
2N+QMyurWYKx9j2UT8dNv5d2tAFwAKEpA0jdA0rhxrtOYxmW5q1dYY6Ck1l1AxXk
YR9i9uESumRhTA3uE+OSh4++gO45wPQuvcw3DYeav3R2486FGKqTfEHtxEhtuDVw
2TaCuGL6syu1FnBEYA7WSHb7goJFVcVB2L7jpFRVJLDj9z8HUPY6u+TS7iJs+zLS
M+z0fWcN9AoVQTeLukr79iiBOYiLdmDmRc3J9BeQjMy2a9yi582h7MDpqvlcmaeL
irC+rDd1DV4OwKQN+qpW+w/9x13aDWIrzJ2HaajKncjAmjtM2uMEDBChPfrmAJLF
Hozx44Q674AuPkfQ+kfKmz4a0+OxJXF68D2nVvQtP9Y8ONotimTZvNeMHMyquT33
lopgQqdL6otrj9U8W0hiUS79Kopg0esRqAacZSJArT+dYDCaIHQUc/FPne+outgQ
s+jzlqSxu2XZqSS+KoNQhSR27mEOr0/K1t3oGjLQ0caxGMdEoT0lnM6A7WvjWb2h
ftBaB8kf3NGDYa20IRZDuOaREDb2Fufhzmp1kq56ief8fRUn2dDYGFHkzlpFw3m+
HcZE08F+vOL6e1WQQZ15ReoiRFlw9f2NH8VY4n4Rf+rwrtBwD5gLp35OeQy9wDNV
znl81t1En3Y/lOae+OZXd4Fyn1vUqmtlqsJbwokP6YDWk3zXaD1Xe5VQaKX3DC5t
/5M0zErCrJMzT1eFwAQdFJaZZuMnIyHxJOZwJDvEN711CIWj5bxIssYDf3qPeYgD
uxPcp3Ig0eZi61QXDBVfk5pLLspcf1WDNrurs+oaNfBM+hNK6F5235QWHw0XZdst
vfjubguZuJxa6DtacYGD3hm1hbO9CMa4FFH8wySpFHJh1UxbtZo5urZHO6ktstws
KqXNP/h1G0v69sionFlBjkjnuaqOdemYfrkb+4nqV33DKRJnVO8JhSQXKtxiAiOe
HY/0QHXFgOtAUyxQNgSTyeLWUMmX60j4xLtgc9YxuDM2dSvwDgiUmhCbpv7mDyt2
KYb13ANDw5cv2Ta3ieoLuo7L/r76LUbaSM5aMf9xvMjgHvCX1B66eOu7WjPvWcP8
JS4rTfqk/buOpt3iZL8APIEqEe/5SruJoe84+wiawBD/JItCw0lgDxdwqyX+zfUx
XLegClzrAGKW0VIZsVNaTPgAkiLKtNAsBQF/Jqc2dls1zkwjpMvsZ9etOUZmpcSV
wWirRAL8yIKBefEPT6dyXbv7K4nLBpMEaS/GKmIzJhZHZwc7Uh/gGOjy6cNWDQVb
PuwDAnC5V5VE7zY308GHOjgy0K8RuERpNRWaanZhQLVy3Y2cr42CpWOwiXHYnYTH
ewSW0d+3b6LdqM51/0TMbxdbRXyUIpnop8MOrCsLRjMiCdjGyp17623M5/FDSffX
GW1HhQ2JD3V3x4EjFOCb4aMc0gFAmsPW2UJQ0jIwjN2ZyHng2vwdHKv4VSUIMGCG
z+rVOfsRbC+lC5qt6AmI4cOqQCzeHNUfO6iAtTIeV9quPK0d3mNn96v7iqc7TWvJ
E4CNRfmEaBnTY1EY4g7R4bbbKyWqkC19e6rAl6yTclokmBLd3UMx3JFfzLKhu0PG
kSE1po7K4r8EBp5oBe68rPbc3ZL6inXi/Y84QgzgzCFtQqN8QfELsyu6QG4MP4Vz
DqwoSiTxzCkGawUNsc9oZN64pTs4Gl+5GAuUTAyAXJyt69FkSHIHoMaitGLfJAfe
59+sagRamLqYtaQddJePF/tWP2RdeJTNTfMI06zh7k4ap5DeYrRU5qLzdM08bg2c
mlqYfBXeHS5qE/MgINa2piKqLUw+cNkrsHmPzZML2v/uE+3D5YfDLg88taIkR2P7
qWMTIEI0A73TeLiMo+bI2BvhuZyY44p6YdGMsAaFv1tlrXkgIGIkcyli1a2T6e+j
jRwiSBynTItHvZjzKuR0gdKUtSWvqrkRtKVjcAv7StP5CV2eG+7Zeq8VbBppYMOz
ePPZ841hjceJ65ceof5Y5nj2ZwsBDMdxMHmvUEfsLu/YDAfjGJRWmJ4ZUmt3/EfI
tQisucpkNM3oer1FzBp0/dfwVUKLfTkmcYrOL6PcGLEbQlScZdrdyfVtZP+oRXg2
ZoXxwLGh9jJ+NktzT737+Z8HPsf0ssXQ4O6tZi53vx+YFzbszdhoXTcRXZ+02aAn
KumnVayUmodUUmAg4iky237mVW5LhP3P5YcIfw7fASIXD+VTamiKd24ad0qQ1xRu
0+dZ96crvpfIWzws4mIYd7QFimViAqqbZxrucb2O0S+oGYp5SBigEGtm6d/rKbci
PVStTG93s6pAuEodQHSUYlvTF4S0cH8i8/5b65cXxuOgQx7CMzqNCWilF69lVR7x
c31i5qxbMIqmYuZxV7U210nAdRpNdPZNdGxiUR+2A249iV9pg7D4US40/GmSl3Cx
HH2BWXRUkQary5gN6u199pwm09psvDOUMEgC/fG4OB+o7IldmtIg+lMmdRoMNvRa
+SysVI+SpH4/ZE3qgrKp06w+PTVqLiOGPE/9f5fw20/78NV1TO3r4CH2Y6R1YDty
gZ6wLRj7iK3y7N4iXTA+hFPqAmCo9IhpKN9/SclL3xP6ro0hgCDTfCAJEaU2k9Tb
3lEDezAh5WXbWCS1k+HOekcaKpB5Vx78Ay2pzpk5FwC1GhF+M28T/GnxcsyMIvhl
CqeYoj9Q438cPCis3vxm0oV4jE5eKzPRIe9cJsEnor0xgHFLsoFY6Flo/voRjMMF
fZN/tDbR2w6yAl7Gs8sE/q/ymZ7QdV1D2xZ6eyzGBVsHlmQDvjSZjedlf2roSmn6
tmWXUA5iCMU/wnVTQ/s3thNzq90QV9M3weih0Ktr39tUEDVGkgmoQ8n4P+oQSvJI
2YtijgGQ6fEqmxa+g2v11PCntI1OE06YcUOeOyHm2h6WSfTd0kThtG3TZtGSrifE
3N1oDtvIC+gu9RschCzjHPWC2kpaF3UFRIlLRFa7SnIiMR6WE81+aJr3wUVQdore
pN/dZe10lEYs9lJojUCtoaJvp+wg3qDRzxJPQFSZsPXJ+DLJxHt4DuqxY0Lj+pcy
WxEFUmX+k8nFG4vL8J8uB7urX6mWQU5KhwRpp8cjlYSM0o1aRCFr7OhlpQBATuhm
hIsTE8pFi6osZmZjmVmXhxt8c68BVq+H9KppIdQwyfUbULK387qzgwLSszfwEbjC
DMgs9n3qk6NSbAOUW6zycCagGZuRUulgsJvj0gfFYO8ibDusKYA0u5qScrykKtKV
aMTKJS64B60yveL11PBbXTwQwqR+ZN2VEukNDKM4Reywj/tq7uj6XKGN78PLB9GE
i1GAI6dpgVPoyNwyQtSsBCDfonP2iPb7CWyN0CaG5mhyMfdyYtOGPFJCbFe1t2dy
yUzi7fJkMKAnTf/N0LWBzjz5Tp+7eYMthzSlZ33QxYOdZG/612bvoVP/zf2+WrDK
Epx5EjcU2myVWXWHavCC0cVqjhqq3Mic+ruoua3tVdV0TXV+JEeSLC0ZJLJLrZbl
03/auWer68eThsU2czK0yOTTtHasO2tQ6U3jEaonSHrPzMhWMn8GwrFzUuRoa5nM
ViFelEd7ade26GJ5f81P1DDkq3h2ShNTDxxYiW5hLSTmCrvVWPYGa35UI2oHTsnT
B4ItAq/UFox0C62M2ZA5VI5iovlDWSjWCkZX4qQkJEDCRm37OzXxmdWBYowPgNxM
ibPMmBpkZlTa11vd1bJeTDpDWIH7MEfi1+7BDzd86Z7uvbFWDoSn2Xu6+NngBW6U
emAVqFJffubLvZPSRLHfWdU6178IAOUnD4fCzO7hq3roiahDzQCOYbZgTqKEwmvD
Kgt41SVutx/MqEnxSRljP55+Cip377RejJrgArd2xh22xN7PA5GN5sPfCzqcwZKc
xFPf98YjjHIu3pvFIv7+4EWelm2arUMV4DUF/yPqUe2FKL1FLQ26AGoYwm4NdZCm
NkxyH8m8Z5NGNPPBQyRvyl5lXgQ50ncZN/0LEhhmXhd91OcO9L0OqPrjFrU9qBaE
A3UJlKDWdHHfxeOzv2iFLSY557U1ArpxkEusMZeiw2oj9qdQk8mb457fsF2YPYNQ
GzeMnGBnsNkqpFGDdQ0YYuIIE+Zp/5N43/15sjg0rWQgGeZNdVArxTP0pdht5arq
ptrDxUOwiWArc3ncllCS+GB3etHrX9+uodV8iObDQVRvw2Th6h+kb308wjhp9mbQ
fkQpUAWXATtZicEO+lsmbT6Yr68T6ZXzEFyea5SzmpeIYUggKIE9R/J4QRJ4KWik
0w/2v4EOgGBaikV+6cmgfEEj0MbE5d06yWtvkMAGmW0hnfHA3uSnLLG9FvKKXY1r
+CTtiR2frFpw1oKpuYPgJIqlRH/Xk2ChDpoDI00I0+JLMhaPWTYWFOxGQ7AXx3EF
cmjJKiZpb67NQ2cNtmrOZ8Lb74wBaZ3b0JbdSoif3GAJykvwKsOu+8Nwps++NrsX
+f27TeCECZfooooilqbhc1qi/3u00gqYMCKWCg+tydorc9lcchhf5g9Zg7CbvkHH
Rn/0laoHEdDb+TnpnFteUmqsiJFx6GOMAC1L+Fv95OhqxZZxJs0+IB+8+1Xt4grM
tfxBWIK0sKHwYMv763I5ta5rPCsdqTwGcek/JkA5bM7pY2wbqT7J4NwvSIXoaO3Q
xjWUIHoHGoQufUzpizGqtztUjz9CuDrXJLfe/6mOJxaET8hemz4wJPEw/bon0upc
+3p3FyJnzUix2+kqzN9tyHyPlzXd9zk98L3O+OXxEr34OOmk9R80IGdsR07dCMto
guSIkfANX8VOeZOOCJD32wZnh+ORp/VR0F/6fL33yDHi8D1oLnymVOdKOQawSn24
GgbrysWpHWCQTiljZT/Z3OJRnZXctcPaJe92f3GgX4mpuNS3Xvb2WqF5vd5IncVJ
lMxteD/Q3rttaBVazJb3LZ7VecfrL1Nlx9Z82WORzqHMy6yCFI4Ph6mopiuflQMa
8kjYb1wpxA4+x2esUPoK/QRvKyVJrMkW9DJjPxD9kxUWTQIKUWo6S0UMEIL83IkY
qg7Sn54TFiciuSn+fmirpcFJWO9oAPb+9J90+C7oFHEfKmqjTCB++sgGXyyjOZWC
ZCJu728y2h6VIMrt4pf8HHRj34WiLzenpDUfLoDOuJudqiIvr5UDZip82/ePytNK
UFQHAPvFQ6sdQ+3IK+OzjyZv0dRitzs2FPBvvc9n6ss4adVEBDj/jRq4+rw8DG6/
UaKpmZTLUjx7+GcjLyv110KoR2NlykCMk04QxTZvGiZqSxM5cyoVh8z2mg9HvczU
XgbHp33jZSNqmDoUTg0EA36SKv4MBh1rhYqlGD2xTCEg/rxgWEvnq8G/CDbfnZzC
sCl+5o7RjSM9VvcLJOGMIMwIPxaY5EGnzVLYlCK1JBFUsim8+s+Nd9VVuVUnuYj+
u4w6YYnqJk6B0+vORGODqebG4NJiEaLiUI9V+I4hMog2cY/qbwbW2BqFeHLzK/It
gNBwJUDSowI1NaRlJiFZqtO73qaKrqe+mAt3jn6TX2Fr+9AuhSBRhU89T024uBvS
5oNRqhEEHGl9JtFIoq04dXa6uzB8S2BXJzEPTatxV8N4WwtgkbbwXdrv8uS0XSty
fk+p6XLlAWKqz6EUTSwZFGu7vW18ypTBHcp6JnlWUUeyOJYZbnKwIZBlqWZgiUS4
mM0QJucoS4B+qjxn0latfdLvY1EjnT0c6cl+ZHzD1gBM/MNkWGuniBhB4wweRgsr
jXZPW0xgzGdKFrHQL717JSAVL0allaivstU59OWxZcSzw2Par77IWlQldYWwcwMB
grUYyxFWhfNQprGlQNXxBDAC5laMPfJzpGTOK29ogTorEfq0XSNgQupkd4NfAzBy
P7vTEZ7jxwk0ylcmc8R7xbecDmu3FFMf1ZJXPq5uui7UoO9GakiJZ0pO0lH/4Wcc
iMoPyqf3Qtvh0FEIB+4CQ0tOyWA4riclyfis0qZFxAfmp1Ijal12zCKxoV1wLkuk
DX1N/Y+E4G6EVQDdFIWgnNvegM9qXsbT88rf1P5/rc8hHMrW1z+aJXHh4jGtHqW/
Cv6Pr2IkkKWB2ZG0CpFKqsNpNkNYScdy3URFOf/sYtJU07rrxklzlteDm3a40lP8
FHK22WNLVMKLkWm/2i0yKZShJYO9IT0aFDNwMefb7y+spX3AldpRp37avPHxu0Dz
2uLCVgl6qT1vgiY3zdpl9uypdTO0GdVTbeE0/xe2okhtGjOgWpyuoi9ceqWr1Ma6
wXNNslB7eRzwxXsrGSXdQUm1ofjsQOdW+Q8rBO+W2kl35p/++UxIkXnQvSGzaOhG
RZTUwj20IpyH5RjuV9s3Epf+GV6SN1gLH1CUxS9+Zll79h8P7uildwBS3HCdUTeg
/jn2kwFwkt/CQ2HihKEwPsDcOi8gOFx/28kxbcfGsVKHT+dYeYI9CngxOBbzfYE1
0YdLbaOQGsNW54JU7d4H6mQkNKgqOGDYZBn983ODXoRsqVzzKETJEU1q3HIX++Zg
4qkXS6QZfnuwcJI6pgAUk7TM18zRNVBVNTvd3qX4SeB/plsFLjVX7YcMn9322aFH
Bqt73AvP/bY5QRsKagXiFPddtaCOto8AEP+Nrk9bjkAguKLwad3stoHHHT/I2kdt
0j5G6mCNNK24WAdMeoTvKg8IZa5xsncvAWgFaYyXpoaCdmPD9ll6vQrStV9DdEQv
z4eIExTxf4edtsZ98yrwrLJU0m7DWR6hfvgh9BKMMXYptCHuxLio5+Iwt/D+RutZ
f1KG4MhiWR2gmH/rV1WoN5OYNr04VO0iXbpsPtyBObwgMC8ecRPNkU+1O5dCC5Yq
Zx3/M01vuyqO83BSwkfqIUcB0r3qFgqU3LcK2mDTUnFehEPWKIqnD1lkmHuHFIDc
7omV5DR9D07z2fd9DhNvlT/fYIPPRJLlylvSg99ZMPS85wza9eK9AE9ZiLal6Lcn
nQQnzRLxg+TItMXfmUryCKYs0i9Jm6SdFrawaaDvgpIvXNDlUpI2ISJQhX0P29eA
EaQEnuBtXXEn1WoZ8NNIi1bHUhz3RgH119GwbbQ6PtC4IFGNyZ8zKt1OX+UAL7F5
KSaAKnfrzM4Du9wPja34D3OMtSAnpUi7++jtM/fjjzvVLoNVRmSiJs77lka/WUzX
gAFtdUywgHUAjD5sxDrG7Y11fnaXbV2hU8Ka5YzO0t87M81iKPc9Wcp+pFYFOj3Q
NKtH5ozqQFYQe04Jmiz6IK+RLk9BOahwEvw2UNL4bDprVSXxgia47cNcYVdIaF+9
+DR4h0NhUiTL9TK9WhThkEA5GHyhAHwEJwgyti+irXvUsOQKQmP9Xjggq3RBGrJA
V7zshVfOKpAe9G5l3WXEXg8wFEqQc//93/QiI1VWy3bP0Bys4OA+yJI194cUcTEV
Kr+zT1Gwo+zrj9Xn1usNL6BGb78oGLNFO6W9KwR02ALild4cixHBfTK0+RIEIjaz
XzxxqABODUDT70mZyk3N0i6wX/ZUKVIQGwcpewKiakrArqb/YisnmgmUZ6MQcZu0
Pe+kLesIukiAFVuHIbPTnP2Asa194/Bx31Qk6sNrht6AvTLOQdpjfTearlNFSYHs
9p0HI4+C7iOGFE3k/kIRRyr4NbvGAV976qZ5mmmwBWJA0Mavwq3lvTpzVso/2BHJ
1Zb4WJdEuK/WfkhA62ptrGqN5fW7JdsONzeY5jZadF4n3knbqY6ljmCS6hROHKhh
9lIYfdq9/55zUQTaGzdIHo3SJFijs9YNpBfmTW2W8BBjua1frtjqhU4oW91DzPiM
UB35qCXLa0UxM7NxhrGlpasqs6qASC+rvIIoREdjpsLV0MTJ04Nq7ED8tALqo8ba
CybXhac2cZ9kRz2mrK79N4JrJaIRorUgJZd+sxhXtmHxEsneNlI9/Ld62srtavQV
jC0PxeTz6a6RkfJo8dERWV4Xk0yJ55oCdXuhRC8g7W2f4n8jiBGdRhOBhFg3Wm+Q
O3mTnwcS0TbFWXArWJESaQkTFo7x86X4HKkY/hn7oEX0bKLll710eyDk7nBwrg8K
NB5rsgIZBRsTgXxOYQCt6DD9qqImlgfVyXRmymiFXetHY+9P7PByhepV0PuGLXb0
acttPiHhOYQg0LAFaVpXv8nZIm3WGo5zhW3lOAmYWj/uPVPVdKynJ7+WvVyckNN9
6r6g/yGjtui4lUnpbLRXLexYiRimua7hEWq10yj/0u/ZxBpFOolXM1Ym2d0kGOJS
Dgoskg4jBIyKhbqD9sJgWyr8NIi9AUvsZa3UNKCZwNKlzjM5yWKHVIQpbNP6u0JD
qklrPgHf8eYqO4Ay1BdHsB/V+Wgy82RHCTs//SCL6bjbYTHha8C/+J2pOZhWyhxb
dCKOtFI6vu+BXe5Q6NX4AaMpJtI6ynyTiJH5T9x9e+jiDxDMC22lhnb1u9o6JR9z
roN5QmUBaugez6KQ+BtJd/GsITP/R4Z32aDmovRCfR+qA6lFRD6/2V3XOoUi/NXY
61u3y9Olx0YbEuQm1rK66pwmUnBSlrMFPKkMPx0aDqswwVNqugcBR3Jsd1fQuFNP
2gawNlorhgbaK3oH4/EsP0eVsGU9kTn5zzPBFANEQ72wS9yXDISY5bQLpkn27Hnz
5YKBw8Op3fi7Q9nBtKe9E3Gp2Y/sC1KYH+cTgAmgRS6TyJ9O/zNzWV9CDNdrfI4X
+Pl+olvqybCee2S3Bof+VKbCfz5apUrbV6nHiZxa3Py/3zqCl6oJsAA/xCu4xC27
ut13K9ZRkvoDttJIJtOw/HoCJsM7CE4r7UZ8XijOCNbPVvsuYKAMTpuoCyN5Hz3K
uoHsH1h4dhW3qrwyi2NLpZ25kUWqoBwILc/Rk+Wh8wfU5E2xyskoutuBrZFrkUiS
a3yQGkDyL1nQSasJw+k2JHU8QAdGGNk60XsU87l1mIDLGsZzBs01V2W2PtdBbLVV
1ovJW8b6JnR3chqaGrKbAFe2TrLLv9x9WgffzIDmv+SmqBtvefXuyfCAB66zP9hm
yx5Syx6pNbh3qi/VvjQaNa9oCkRVcgBGXP6oT+MgBhLrXKXFSn7W+X83ql0V2lPw
mmnYsV/8wGl0sg+6DThOGy6uL/2o6oYmTZkxYE7IKOP4NohPrbbobY4DUXw9uhGi
ZYY4oxz3uwbvIp5UBKTsNZIGJhGLR2CyuL7dsoce/N5lmpxHnqrD2OjRky0EIzMi
AqoP84NP3aDfM7MNmVyfng3ly/RycviOdcOAHCYrdi9F33EiiPPEVUNR9oaCZaFt
6JqdQ0I5jfZSkBqMKIp3jWZzPwIc+1DSU8EaGjqlFfHFc0tbLv/JAc9IOEroNBbr
X23RNdDhQRvvXULAoKS7fgGoLXOKUXAgmCK0Lio5OV0HnVZbx/EGM2vV1dKm2k+/
K9KansmUeWAmbHk7Yu8YxzcW0MxDCHVibOfX8uteyDz963lw7MOS0CiqM/fsYFVa
lDFfzJS1zqSfLx04c5WFHdTo/iF0r4b1+kkGUMLxB26x9rkTPk/E6XSx6SWnRBA1
lWJQorvS6/bDzsHt3eFxTdWaGpzbdg2uI5tSlcf82j5bo4O2LBDACv89iZ4jE8AO
U0dViKWsYxkwBb9NTFSwG4JH24N1K7UR0gAgbm1atcN1S9lWmPjtv81iRVtZ/gzG
8leDB5sLYwEwP+idywqXggLvYWom6bDdsFI0c0C45g7frtOvch6a/NGiGJCJZW/K
QYU670QgtYUWT65y1Vd1OuoxMlw7TThDFoyvX5BAbBKsDOZVLF9DSUR11KngG8VS
bdt/F/UyU7qQu+DIACOFGaTU5LzRJNkugnjYjYYQVdV3FgNZE8+I911LaWcJinKa
ofy7q3vYiyl8mL2CcSwuNAdQpj5lJxapG8EQPpTK/4w/yCdKrti9URsLy3BVvS+b
B7fDqFFRwGgbq9We97VALbyzRp6iUPKc4zy9JlT3+fp14eknWRA9WFiOZIvVU8ZK
4e66weIdvx4fLBtH5PvluKWc7wd3YkJojUuQ/QDDg8HTU7rC4SSZbTismsv/kVUB
O8ccSxKeH3WDt92mF7dgwF+HfWv8gTtuJ5NAn3DB3NMiLoYcLnCmnVvDLGq+6B6J
f7Urb8Bwwp1JQ8J6OV/hCacz2B0b6I2+qpzSBEn6Xg3oVS3rP16GquRAchCQSp8k
V4LFuqJicJYIAJh9c1ikRmAjzk20F+h7n+AHq1rHouEn4XPZBeQHgGYN28kYvNu9
cs2JQLlNNRRdKbvwwg+dAZWRzbTgYEl0k3jS4DsX7/+MKOjEVhEq4ayFF+HXDXPP
IBOIkknD1tx4EIby7M7z0RjXBdRWkwh9O4QeWdumQB0a5gfP+3/VXbiKzybg5Qfy
vV4STVMpWcNr6IdCPlno6lkdVj5nDcVsbtirN/e0a61weCvkZtWb0uApvGni2dy/
+nSAEZnAZ4BofeC2N6rQ5wYAqIzpYIfrdKHRCLwqnbNxqVlD7Gh2HyNyVvkzMu75
HVu+gcQpuFrCyLh6Z8dbnfOIcdeLv2+4aj7DpwpYqQr+V5LI2in+JyvPHboxQOjN
BxF2MP7zGFuXgDxjgNxmSxviEfI/dLENiylmUwuudfyoWxzvOCtcLk1KLnV51zWk
ggNEgePNm/KJNS7bnemZaXGg2szVef+oTaQDoUdBqCUS+imNIMxLOpjkAYMkbK47
BjBdQLhNZ+xRBq1kkyCXgcawLvEKQASF636AAWdH6UXGerMNATPCIndtXlmiXl+P
o7Gcp1frNY+tcT/BRFMOqVd4ClHLQ0ltg6SupYcz5QYqXqdFWBpY8SidSP6MlEDS
vuIdzg1R/CYnre/1VsILeeD+jzMP751Fv6AIdfZ4dyr8m01pq6eH1rvTbryBNwzW
fGiFbDzZ30EehSFzw9RRRNFH72jnP1ctA3FQHz0r75O5Th0IKYPXYfWymzf+YVib
BvsS89lHTqo0pvcWSNKuYAE2lvuv/L++ACeR4IbTbL72XrntPcqjuo1+Ogfg3E7X
e0Oq37CyHjWjG8z9Kqjd/ZGy5lvX7Rt86HaOcZwGG5LNVQt6LILQWhgHK+rdBDOA
4wzaULdDtTe6t8a83ajDpC88ps230GdYYFdoPiYPiVpv6E1OHOHaRsf3K1m5yQDI
FNCmDNtSD3DzgEkydpGABf+3nuLfAvi7ht1u3ZoQT7HwV6SrTgvAm0MjsMA/hkzi
E6EQfBx3PucSjjZkkVilvd7Fm1tN7am7kp8/PApUWRJcf+Ce7r4V6UPZk4kYpILx
93eDpM7X/e3V7ywIwUiSzsvRUgj6/13NXJvTTtNQ6H1FTVheG9f4DvZZGlds9vey
b8RYmNgXVMvXkowNUxLGF968buxdGNJzPiz2UULC66YrWoQYXxNb7c5nZ/bhFhMN
tmaNGaZD+2ci+uORKsY24yiU60YAtNqzCHhgDVdvqYLMUMngDI8Rm0C4X8dmjHV+
9J4XLGwJ6ZBSHKBLu9otayTv7dj1tGA8V+UReK7YfV9afFwwT6jQ2XZRzOR/bO5e
QKum/MWMi7otXWsu8D/nqo7/xJLVUyGBWJ6GF0WxbmTCVNah5L/Oq1uvr9ZrF8ap
CWCYiDGvpZMcL0ePxbwmv6EI4Orc7cTRxp5QpN5yLUeGt1R1C4t/M6JB8SXOQD6v
twxumbJEqMN9b6VCz2OKHbvGtnMW7bPl4TWCw0pp0ZTAGo3Oa0P20QLzo665C50N
Q16+rQXbinVwN766vjnlmzETZD1xXga3HLqc+2MyIjEUMfl6hl0PEsmZuK3XOT4G
S8bDHeEISLubkowp81lLyqy35aM36espWb0YtnGSpwQjgj6GIW7TrxcW1WaPpBL7
2L9wSdHeqkYgnOnQH0jnHwCxa5TNWGOLONb74AxsCfgm5L3fM5Z+64eXklKcZxI+
jfBzKfnV+z8K6DBxkOOEALxvm0aAsPsooD4e5ro9SQt3f1h49REJIZylU9JUeCGh
lU7mU7/ajdwcc6olVXYhaemYXD8BaaPybUEch+fRE+1OKr2lfiCdhqAb17ULiXxF
C9lrZo6+a+0x2G7zOzk8sE4bwMkHGvBDEgYkpKPMGIMAJUflcsHgyPXvhSm9DAe9
aGvNBrLMXI13HH6QwILYqBq+AMMmQK0cZHmYrsX/M17OYaBVe6swFpAGCweWM+L3
0IFUobkpVE2HCs3Ppi0ZkWmZE6a0kVY+DDvAPgd8w51YUlfNzcvsp8uf7247KNFw
PCfOTGnCrE6o1oHghNuAZHXhzLnAx2EfyuZRH4Gvlv5aAn3z8n3RVy25wyDhGBjL
Xbz8yYgLALpCetNK9N1HkzkYEaKYjXP1uhKlux6GnMZJa5Dfjo75KGvpeoLxd4hm
8fX6JsZp9PD2qp26JgjdfmS0sDWYGE4uAo5psINW/RmncKxMA4uUsIezzqQg24fk
G/a6IjRkDXxtsiFIZlI6BMJm0iG49LizOTRQAJmERokIh48/IilgEjj5abXJ6093
EaM2rAugv6zto1oG6FHDM6WX5LlbnAB6+o6aBv+/IDP/xZz6qWH+qizLwhTJnizO
le/Y51PAqjF+PQtxoGL8g8o6WwVJ1J1ajznOSQ0HNDIAAqKVQhNAGWqr88lrM7QR
w9QihVTsDlp8gSL2ubaoXNijGWeQQBth59tbDI1IbF2GODlbju9ls0PAvu0wi4ot
mLV58u7FkjISfGarRLFWNqd59RWlAADvJHWfFRkUtZBS3G/6VA3m+Shcxq/+iGAp
9unpFOkFWBw5Ioa6ozXDXZX3pF+W455b2RNNzQlvKLTH13M/VvJTDcRtA+Ca7tiL
EvqoYdSSM7iDOO4pYK8Bp5VJIv0DGANvm91yfqnkdDmuPDdfQadEmrjxhZQ2TrWQ
5dgQNJLODDbWJBk8oVzxcWfeDg2BzxVxTqRMThNvPmq8kzBNZritRkm3a4ko0F3J
8gdux/NnHUXrZSt18AOWy2MRMlA1oCjVGZArLz7DUVm3YZUK3zFU93IAff6VkMg5
m7yYvZho60rqPlzVt/V4tGT12UBiWPqyfFiR512n/IECOQLc+pXB4e3tjElhe0Sf
1aZdT0g+c6GGg2D+89EKh4UK2b0JwZRVBAGZG3+QkGD0LRlpUHU5RfyDUiCBqfJi
t3KUGVnrkXThUF8hlMzpKUV4+F5E/tuGC24a+9VoBK+a9bmwyeU+051AUU9MKqN9
Z6ZCFRCPA/EyvWS7QUABYcA9yUTO2E2qEkdhrFh779IxyAFUi3y1zvmBTDiAbv8k
eVJTc3CuEcYgTzC8VS7OcFd/70wMVPH1l5SENxU5nWv35ZA14uerDV2Q1sgqhctl
FfjhdoNfbBnMzcXy3zNrPCXaf8GMltjI0iPTxYPa7NU89z+vaSPHK1wyIL1U0/gh
lfytUP/jEhZ1G7yP/hy/0bKDOEzjjiRLQ+xuPLaYLRr5E2fFVnoEDrTOd166gYZ1
RgxQS661XlUaNnoOXvXr5jcZSsbovTd6FTcavHH19lk01FF3Y2bm5G9MUnpWSpCk
TtPFmQTGIjsgMsBQ4jjbYg+F+ygrnvGRkMlJkjIxcaPaa67cWld4GpKTP2PCGWpS
Si066o+XccwWn6vbzH28RZOUwFzTyDHXvG0XXUpmAGZ5PI5rcAU0Vt9jZ3Z1LeNL
6pQ7sQCAbU3gOYeJDfa+7IJGDnP9gHDLTW55of1x3e+a+HYJsU1MC4PIcfSr9p2f
6sStRgMQqqBDaLEN9l9go7O07aec14jGAy90lrJqz7xVx2CbwR1p4Ad5EiPpS1cC
pO8X3jdp65rj+ibvxpNnpwacVmDo5+jaVTTiM2KGVEjsVXY1pzPzUVs+Xtv+f4NU
WVoZEdqXUXwRVjJ/WTMaHODlFTZcEiqirQ7xL2J4gxh7bBCQbWShkqdkDXTNIsRY
FvmX+NqTVvJUxZ9cIO1onUUrcREXG29OeN0uR+KpQsAdwmhVAqLF58HOQsKvshHm
VyrM273x+H8mSxnJUaby4LyMoKcDBlyuzry6LTopd+nWn7/uLpv3US7J2KpQd6vH
6QsSYcQrJ62eCmLoUfh619RYHw6fLkdagD/uFesZD7luV2oKkG8wmCa75S99CycJ
WwMAsGnsS0wr9ZfC41boE88XvztG1My/QHRb+uc1gZOFolvmRZsub1zBQQeIJ1Sc
2TMGiJP+lkInWVnaUWrEXsxsICeSlDaXkdMW1c8CcYpMapom3PaHWycIv+2K3RDr
HvEINSaS2U4pNSoT47wHujNdlHMSjObQU+m/Je6k20Yv8xArEuFHYayjNq93ai8K
MISS6TNoCFTT7ebYB5gRRTHLNseP48w3YoV4FxspxLuoZJgge1Bl556wehI7kpFm
nOasI4SYw7Rv4P2l0fzn4F842B62fo0OKHVhVQY3mya1o4pj/ynwtpIVArycbD/G
cSy12C8Fgiu225073nBVR8fkmqRR1v0ec4n9zJKfwjegWs/TLrdpXx86THoBiuav
tBRIA+z6s31wj723GhQe02bt025+FJzmNJUwXtCbhbcq85qGiacEkQtovCFBrwSq
NzjOJ8IoZFzhAWLQkVDPFbRPmTPvtr5gaRRjObb0Tnw9rHKxJN5z5IDz3Lpkz489
jwF+zDl2eDE0qFJKM4oVR8DkYr7R01/2TQHXdrtiMrDQfK4EwR6nd9tNjKHiA72c
+mPCb2dY9+2X4QkauRDrXvBGDXqCiM+0e3/gg0N5GceTRMDbw4b88DFL2mFIHUnt
nlahwj89KEK2WAHcocyT7hKwErVupR5P0zxzyJwSOQoCG2ulvFH+s54iuuTEmeig
xwKo6l46krvCyoOAQFGO+7DrHUjy7jmKjf/MYlT2CwWG2K/YSOrPeJ9jZ+kc17Jf
w9rhII9XYx4LW+bpBUAvQxa9c4zBwlu8R/BtWFJq34ZLudIy76OYTsca10R+hTAw
8mH7YntoxtCSJJ0XtkAJ4guKufXgIijSabGKvITKn9G+IW7RIYvkGqLYMn0lvcnT
6J0gh9ed43odbxgzzR1a7QdNA00v4AE+0l5/J6FnNutGY6GCBKilSIHk17yu18S+
QvNYuyNxd5sTKJWm6tDgSltUHN5iFSfUw2exsnxz4Iw0rEDDcZ4srb1YAu2cLN0F
XF0k72leNkbz8j9JCM6cpcbaC6/hYlD5MntZF7Z+RvlNYYmQuJ6VHDBCuTfeDz21
bFlbk7pZrYyGfOviHTEMtaIR4jEnEeg4BYH/CDZ+ZUpeUThIKBQeGCpZ4qSDN8/n
TCYx8I5GjLEtqaPHczz48+vgyPD3H3/tMN0R2Csn2323dEnY7X59Qi8VjgoRK48c
2e7QOBxtPNJuiuKKEyZG9bR85qIf9rUEwJiDIkrEVJr+9d14qPISspgNYo+miocP
JOHkeZBZbiSKE4ZYUfX445dSFpSLwI2oCzfUjW1I+vXkoDCvFKm13vpgXQL3KCy1
JB4KJsb4dfh8TjDMnDSyX5MeFuqknPrfgemd7K1Gs62HqKIwYorPKwHjZNgiNR9n
haTZ7tYjRh170vpssPc3M6Frap9T57pUqffSVULW387eQNidMTrtR5VewqK5+4an
8/9ki5VjzdrYldy1nrje1n/peIliM0HNw/5LdfgNXMssqYNS7TkcguA+IvYmYwxu
D+puTXIf+/6rwfv/npUMnNDAuyCSRtDin/HfpT3kaQvk4AGC2tIBbXaGbANLA3qF
sHADS6jxlve53nUlva7sNGPDzQO4wfHiE4u7xvWK+LcMJMyv0rlZ9fn7btk20EH8
w8SFR8xgFunPyaqO1fJktWljJjjP9iA8qkRP7fzQJ6i6riRGuW0vfEftvuYCbHwY
5Yqqry873UdZOPZ9zZ4rbi7cQ2bxz5/o0wdQDJBcnJSE5uNa12IZ/yxWJPOHHpLE
JRaWcs+9UFDgcgzOAb8SzpWK0N5PwvBmncp4RhbMIFKSHAYx3iTei9tMccruq0yg
OSm/kTBy61ihL/bTG025S1iMMjBUvvGVjtGuvbnFoiZ/4nZPocEFwcCGz5AE5J6L
4o0vRQ4saqWCJVx3FUNlqBC/4nJs7XuBb+zAKvQhXUgMRrnacx/4TDAt8p4PtzEq
RsGsYAVeHX6uVKeSTU1yFIVhnnCjA78Qt4U0hO/cU+Zru7tnbeNy7tHPSdPIOKCU
bl+7pe39Qf3L3TlcMTBLadDJXdrEVYOKyN8XQ7KlA+rsIPsqEuC5yAWwjC5q3YAn
zR1NCaWWX8NocaKyRpz2LoaSfj5B9ahLh9F1f+v+IntnMzQAkWle1+Xe7uzx9+3g
2oSXsIKZL6EMmSKPkcAwHuK5fHRTixevfZdtZtLszpHNPd3Zr+AVTPxO90dEX9HB
fes8BUWfvfDidYhHgDDnM6/EYT4BECNJ++OBtTqPDg+07DZnJPLvUz0BekiItsy0
+AhKdbcunyfQ2FZNHWajDhBYWWH7zja3ABZQOLXmA7+i0t17bRkTkQT5aNuYKDnU
X5hAmn9NQyecvDzXNUaX4fcnMoKIbqZtuy/LezpUPw0jEP0PnOLK38LCN5588BU/
pYo0ccsrcmVME4ppPpTxULYCVbnUiqN8YnU8jNC9l1NGY+41xcOCNNNfwBfsA48U
IzM+5TF1eFbI3C0R8GJIBHZEbKzuJCjpBZ4N1WI/8y9fbBmaBpn826m40Wfc6Pw2
lBeU/yhwUkPvry4CjNUPCtxlgC/fZt5u5P5loWtTs9PH/4+eepfNqUyf0I8+E3Ej
6IKdypOFfI6mF+WeMpy7050wAD3eOpRhss39RMf7jehjMJtm3b2yJ4uYRiIenMYb
Csi5zbU6DTKob8GqabwKGTvLIRxyhaa0VX5XWWzZm8VlFQnBRUi4n38TPjr7icDZ
Xbkk3JFYpdnGr9B83Jp7ChapG9VfA/3GTOr7C/05O0bN1MT0obwCujh6GkoXlzxb
ng6FEMBlZWfBf8T2DYW/4IHFMc+vFFrzA8qDuea1bo0m17gcIYqdkrrVa1B8wUtV
YPzZVEQO6HFcTqdsZs9TEMW+RC8giyTR8c/jxuAgAKHJ9Jz3B/Am30rSAWe1q3tv
doZzDbR0Hb1rph8p8BQS3hfBmgamlDHV1gAE4kVnDB1jBeM3/IRRcCUquGE0ChKZ
ggNdYElyey7TEgzE/6mcjuCs4+hlDxgWMwzTXIk+LrQ4sDAVGtcjPwM/bL01bLlP
lVLTUNJ2xCCFtJpQ87f3iD0MQbiuzV4VcbBmrdEX+bdNwchkfRO8BgiDeZjqM5PR
osdaoPg39uXLYMZctGVbtxkCYRrrgzfreQKr/Ute/m3wZqSJO2RF9a0/M+FLWUg+
7jIBbc54CIciesE77f33ahFX9yTMzRBhY4eAPQjzLy/NznbMdaTnwVcuRgNDGbMu
8+BewGC/y6YIYqqth8rHRY9bkD5KPRjydf7Ev8GNdurVN3MkvICEogAi7JSeEfMQ
ONmMvEq7YKRMUuJYqlV+IS5+h8A9ipREPuBgedoCQNlvkxNbzv10P5+5emKoVhw/
+YqILAUbaaMyOEEc8hmNgewfweV0jmF2VybhjjhALztYpEWHgVMMKrn5ut9uHk5S
Jq+Cw+0ZlIDRQZeXgQYxQIpkn4K0HVde17b9qKBDR3XihYbcp1GYrncW8f23HUKc
CrKINm1lU3tXOU3Qky7g0km5Wd/UV/Jp1PNWazRtphHhGVErG+1UOWwmgyjDZOMi
Qhpqyhfm2s9N/5MJQhCLz9cAlCumXpce6q5fX6PWOqTzpGsz4GiYjRKE/BW2Obda
YqRCpHO8Ao7OOKrF6G63nvC95PmAMfXyFZgwnAUUqEzh6zQIkO+O58qoIFZc0L35
u21eE93Rji/wmpQMGKNJIp0fURZiRvP78ZKheaIocx1QktszdefLiEZodqoIPAr2
he9BbsODcrMEmpVtXTfo07S+zQzutdBbVZPM0Y8GCyJeyWGe/nYGNjQL6zP1wRtL
RRdROcO+p/5BDS8bIZpz6MlUH+TkseoyJLZ3fktbTSGu8fMTxhmFqOMYnKIpPIhd
9WtPeLvdBmcDDHAlsp8f/a6Gb5TPbJB+Xv2wF4EO0KC7AQCgOgtK1YD8gbVOiReY
aJgOeRiRuISEYpYwIZm+drVzuyMv8ZXpDmF2QhZoEVRw1xw8vHX43oP9jLaZQ8kh
t+CePae0QdBvMwxicUOy1LCOiI46FKWBKwD86fMeRnn7szSKf5zI3C/dsiASUoCA
qi+0MQ/S6B38sW1OSZdTYpak8aOpTE14HBmlz4fAzIqX+sFRDF3uDk1Kqsk5H8AG
+LdxW187HFIex1flBdXJqijHfaC6fjohcqyHSIoLijObfWUm7SoOeHsqabjxinah
28JOn9PVY7y3dEqChAVYg6/F3EEQXax3V5VGmw4DkqQZN+CvSO2apGvosTTF37br
XBM7Bcfe4Et87oCOCBJKgv6QEp7nvgQse6RsdWRHDg0/kBnq+CYkp3Mrz41/Ak4r
KU3YzW6ytwNP80dqpb01Dq8oMXs/hn71nmOES0jiljcLuDJmiOCVlvLHLwTk3kDY
JM+L88Fd4mNpD5gx9i+a8GW6+NhxFKQR2aYdC8o86LZYvY8uspxNXwI5deGIyiB4
q29ZBMD4bHbEK5409lvi8KYJ1s7nTt4JHajAvVKS9H8R5SgrENkOdXDrHbryUSw8
86ITz7A23Prj4FPXcAtZ8wZiuRxqMj3suCvjkBfuDTCMs4A3TpsUp5P+KGK+r39P
7ECr0xi2/ILpbbN5UtkuaLYZUhh3ZqFE0L7QyHtTA3f0rddg87w+msfRHXvYiPri
pPtN/No0eqOZ+NQKfa0KoPG7fOZ3Dli/gb4cEhUORUBR/Ax1LXTRg2AHtiw2Zq3p
EmL5A46JdHtTWXmUDRokticHSvCVeE/3Wm+gM36M6ZIeaPgMB6PqJPBlE3jIuiDv
3NrErCDprFVOqEzt9X/PZ40B2Qj23DTnV1INEXPK/LqWnm5NFThBYsEbglr6uSC/
W6Gfsu+MBf0LdishmuuJy8pR3Z/5GbvK37bAkkY0ZyXh5BcfmUhoEpM6cDjmom77
i4ezSwvpBNv+lO8Fjl6b7Zo6g99XcCaIf+39VLnx6QIIJcES2I55SoITKsciW3O+
Ux0lb/akjC21caN7agK9K9A4nLjlY1/MEiKYyXUJEj711QaccozDvB5jxalwUj+2
E9TgM2I7Z02Ah+sVSsJwquT2jRiMtv9xYpxA8ebw4gt1+1ZRaBXG548UcOJ/UErf
mLxzo9T4hnPj19byp5KDixSkhBT8ZO4unfdYvV5wCjQMBuQn2JihyDWze15t2VLu
M9SddST10azMGW+m8v6q2Dl1Uo+aeWc6HU7fcPrNaznxFFgwoD8S/i9IozmOPqtb
9yISpZpWfWtFw5lAgspFK950TjhhwUROkgkJjim/eYhsq8CpSbPIt12iGc1xcmYv
5kvZqDQ0fPdPQT/janzvGXminmKR2kpf3pQ0Q8BQdoAXg9HsWkhZFF8B5+WvKHzR
i7o5qVB4z6OyT007yf4AJgtkbYGvCpvhUwtQm9SVZRG55sfxBjbl8eHL66rAiloL
b7/0fhXlcYJCH1MbOII0Vfghn01aOpvvLro1DGEf+TZNz7EjV3UVm1dCxrM9e7ev
OIOi4toFzNS+6O0sZkW9HIl0MKXb/O/I6elKxjl/ONtNi6d84PApLnAofSQI2AyL
BfpffF6CNko/a+4FJ3V48YZlpgXb1BvXe+tcCJS1nijJqYmLO1sKx+Wf1SDSIW2W
xD+DryEGG+0zYKlX3o7e01s72BXn3dKlmNQHmErQN2Ah3A4ePF6OEaHEN3+cTLDx
X4ulAfdPWhKZPeGF5tdT6ZGbtJlXEoqgm66vmOxTZND2wL4LY6bgNt/vSKwhxC+p
Y/yWcBEOmHmcObYmyG9vUpQJT72TB5Pkdy6yOEVf0yk/R/5dAfMaiZHJ1UjEKGTw
yPn9RfjgjL3qhkW5Mbfpd5FUHg66M0FuVYvEV8h6FAeGUPBKQMD6lGYLxsJ8jMUO
DH57j3h1HpSIji8YnS3UOdgqX5iI2ITj55FDCnRYAuDAGUJjwYqsjvOfcpXnOTQK
oQubfiNmH4yDz4ZWUqeldHHNvA6tCqot1u2ijFQ6zcV8LRnsb5aAQjEF12Ost8K9
zk3dL8uOim6mQL//1aDqWtT1ht8GlnnSvH5JDY0ZlLDAgwpLMAunXcC9aszDI/V9
o1T5Rg42qWzngNKJ5DAgoJyH66eKt3tngo1VNKAm9QAGRRI+JJglp1GDhGpm6lGy
zQCenNEgs6+gU9IyJbABVnhejBRvzxiDSoaRaA6rb9p/ikcN/uLUEMnJS087Irsc
hJwgV3nqym9zCijaeqkcLJutlDTWLwSvLEnpD5FN/o1x/MB3cazLiPFNmWlhFDsO
vaIDH21bqbvjQCZ9F7wKN4K1cUC1LpUaR4enm8NfjqOP/rOcBOgy9mkwZwpqOOm5
w3q/l+7p85KiJeW7TTv4vIR5n5azuzaVzWDWzugn5Zk2rM0GW539tajCol6RCWvh
cRgGVaIuAXmB6OecW2MT4CHRv6boCTrGqwIPbzNc2gGvjyf3Khaccg3HOHLBt1i0
9AVnFFGVZI6EgWt4RXOTFzHkeix+zPmHRCVbnfz7o18zfgq6yu+tQNQhb2LyvkxN
cUcUFBmpKpjSsFSKgTEg8mqgUZ63sqXdeRrO3EvBM2mnGj7bmV8udm/kRDMT3AJK
sIeR0Cn5Is0qOwERNKlT69eqcEjpbKitwr9m8mETuaCdkscTdzd2fJXsweUI42DE
wx59gOe0YeA2PGfrEcGnCyMpViPtgVkCQJCPlDsULE5ugJFIZ/Fbx+91Ll2fPGyN
KsWRd2DsZd+2SW+zuCRWT6bZAbxanMtHJh/29RVopz2nDCuiImBvrRBfysaJ29dZ
MZxMSiQO3Lt/VYNU2gp4occzM8nigQh5fHDbRd2atRIV8oRR4q2Wxzas4kzzXP62
2/3Q3y1L3CJjZ+ZbC/mJ3IVw3qtfw6phyy2NacxKKACjQhlbGMjOv4J0Vn7Qv4nv
UD4siBj4OLZKx/b46z4oDZU52DgPv9OjtM4pmrHV49P1bDjkRD1ogfEhLeqi1dVN
YwjHROPubx1qiilKUVlO5K3d8i90R4gqqtzFVFrOzjapjAGxXp1l/YYvsL619xdE
yLER7hI1nDFDLeKQM9xGCBlca0HUusG6H8MIRnqNrGob4dKLB9JSfYXoXTGJirDE
eoUxNO9z75WePFF2afi6h/6bWnbz2h4VBx/xqy/LNymCYhK5ycU6i5hRpDY/8vl+
L1c+ofJDayDg8GLPY7vA+jiWokuH89qF2qaEHWGQbcqG0DNg7rzos6UjWIgZX9p5
i5+Fcf01TPFTlAG8thoqEvF22RWRdiiJ1aqvTNWApye4Y7N9YirQo8c7/rrRefE1
Khi81mCe7NO8p99KpAMsSsXrt3DMXMvwuJLeqvQB2HCvaoTxSS485TaHVVDGgBPO
ae5x9YxnBFweDcr3wzuVh/zM2hRijFBUuHG1kuFUQCDYvIcIAQ3fc3/eF/dZkR2W
rKza1G5sDVNyAiXmhXMVIhljRhUMd1U7j7eyGLGUqE4e42oaiXmqbfciq2oynyt+
03gFgY7veIrlwsi+AKI/U/nmzGxNhcM5w23DS/SEKsVq49bMPBSxdmaWwAOvmcCk
thK2JxKw0Z5whsagtGMWIAFv0jGOEd/UlhGDWCZGgKfES+B4QDv4fXl7SQMOopsk
hY+yHB0Boidt2AqdxKfJy8iXdwSWlaYQBuRIqjS0c/NCKbzQZWJ5nu3GndEwsO29
09F0FkPGVqspR75Yrxgju2u6GsOW3UG1nN+AXO+51Ww35IGDLPVRJsR8eDL080U6
LvaNgMYXjRcChLW1K1NiupWFwMZ8vBmftKVh8DZzBi4zXlXBJ3qFoWCXm17oHQOV
UH6hJa3gH4W63DHusSKqyVU08ZwhMXTtvLTRJ3GT/Pjfy3mcWcqSYJ3FlfOplVN8
nK+WFIqqvwjOzElhpLrU0l53dujVN43PyRf5CHf7ZwLp5wx5Pf8nywd75l33vGbY
p33oondy/hVXyZDTZl4CYYAcgFRywOMOGux8oFJBBnhqVxqtdnlqiaNIeXtL3Lab
m4+S3xxhIEl5DZkNIg/1tekpCTli7wevl+pi/50iwuuzHoAvzgf/+GFoPyND2+GC
VUpf7S4RDfSssTzPCB6PEKZliSKSnEL+re4x1Gzy1Mj30hzVWxwnm04gUFR61tmI
d5paMcdl5kt7+envFWGsB3mbDBwOqbU65EY/PEYnkx5aqZBma/67yQrboHaWEot4
ffbEkrzZXKY1f4cZ67F2Nyx6d/SEqPBKKSizp9CeKatwskcl0v/+MZH7rOSCV7kV
1qZDv65jybs3yZ1+Zdgywr9hHZaQBYnhypIMvWzPSteArgXGOO+b4Z5+hGcqykok
B+VgME5uzLUEt5gYRc3ozC9yGPKYKkw8kVN5KKTsE8BcCP6lkPtjunuChYYv4Gf5
Cm2Pm7vGc/d4m/gW8ywRkjHKjt5NxV4KSxrGzEzWvRLCN2sOaO661Pk2PZYuiQ+z
/dgqHd57YELnRI8RZZ3VE7XoGCkIIgOcFN7uySwAxXjAhuvJg4Ig+TCY0T6OimDl
0DlwGObHXRUdrFQepWptE6RhjyG1fuZJw48IaGu1eVTtlCDardAyYPB3cj7UBFlm
XH4BHz9YzrwelCHHVs24PWU18TGXLYHBsFoUQ/oxKM0XXMGL2EhJ/DbptKgTObzt
i2HjQsuvI2Ad4iFUsef3t2w6p6tpK1CDS/wSHx7OK1gjhTCf2Jdb81IgVqj8CgBl
LOwIDOQTf24PYUK2ctFISJQj7bPnBVRTXcrYbG05Aa8iZooOGuacg90g4skU+ySM
xOa4evkOZmsS/6gPWzpyP3fV60QGOxy4f0I7fmXjTXPXJ/Mm6pjSRltu7naypisq
ARIgDL3kcM0SnMg/yL+JPtMAuhOC+eir/WGRwGFU8J5qYpLNFGAepUpWgI/9/PcA
XvVmFSKui2+hhJ7atnNDy2bSv1nSFp36Qi5n7XZ3JivWPJNQEdPYGVbL/Lc55AVX
Zuz2EFPBP1amULzL7SKeQaTQAYNPJ3cGuUzJjxxZhFQenYYPWOmUWcWdWfLdn94Z
XyefOHYY2qzIBAKCzw99lToqBkyX+EAtj5cMr8Rdw2gOv2vE2g0Z4fdm1dlaRzV3
0bp8ons/IdMoH63/U1u2saxjPKpj2VmX+RKoAxuFqe4VXXS+Vqy3WyMO9jE4g426
SUa5qq+/jdUId2v7rD6qdvI7+/hJYziL9iVDft7Vu11GQXkXENzWW6pCizpfoyx5
fqmA5GuHCsMgRAAwJLwnBNo0GTBuf69B7y0Sdm1PKY6DgmGb1x0LEOrBDKCnhk94
+r6dBLxtzOVyFD9fF0LdbX2miHRnH7pmwNwhOrHNIL1zjO4s6MdRqEHYxXLi2tsK
RMXxiUC4CQfmyOOHPM1w/3LVw0jwflC4OABZi/5vRXfWZBsQV5NA1HsanqWpWrvy
UaG+PKQskkO0K8PgdWXeO35Dn6l8uG+5wrHl2a3uEH0wX/XqpPMz2cOeWxKlY3BJ
bqJLpwoQW3rfbjRo4/iH96Y+Iqa4mKOMs4BL9anZIm7nptSUelSZv5luLi9/E405
cOD4q3NVi+ljMxf7FreWViHoeHBi0qEcrjMXj46v1nm0LjQ9svLrJcDZv5+7ZC4j
wKZvHxWiyK49tFmQch4R8yryUww/zzY3gX87IoheUxC4uczVj2kINFjVJFyjoufr
bdeaW3AS2yREA9TyY5PTQsd7blrctinouGLhtfNXpSqPGZrRv3pQppHp6iSMAvxM
H3W+7ltwZ+bdUYmTIsTqdjWEXErR3RUeSV92bjHqXmsywNETHpzdpogpzihc+IPU
bQlu3W52ZF00fnaH+Ww37eFM7Xb/nVCdHH91BkQkcw1SDgXQrQt7yP0ftHfbHGH/
9garhQzL97J1SVCfwDteew0ex4G0IuDaL6UIXN0fJbg4PKZrL5CVkn9gVZxYvDCl
vRyWOgwUsVdAC0VrrlSBV0QZrJRPBaTETfIrnxwRkoaEIIMwyJNPfcr6vTbSY8HU
21R34ZRXTk4WYXETPnPbOZgnGr1KlOXI3jOV+lyjoI72rmSZw100Vl9HWUjeuaP+
Px/WJOSRjuN+uaY6bsXS+oBbXFl18zJsXt3M7s9iWgU/0dFqa/zVb2UdUQuzjlDA
dRkfxzDm2pf2trheKmmLmCL+JbFl0mm7fboAAtqxZC/PM3wPN2MvKYBFcGF18dvN
XACVIm8xuZ3Co2hubITvuiifqBQIj9aAlXbeFXlm1GDejlC9H7jm+lJst/z/3VND
NWiftVbS+USIgq+SSph3BhAP+MRqu+iWWKHgAjlbZvMCac5awM5nNDOfFz+dwXZ5
f+a6VVlkMS5gxVdB6Qm//lhjlJIKmiswo5w9ST7A1kUyIVw1NKZg75lHW6RNhPXv
XoK023LSonMcafYKxEA3iejeUQ53n6YpTZ47lz8HKrKFdbq7AUM8fYbK1/PNthi3
nQviGTgQe0iYU88qaQGLOhQoLkf4uTuQHErtqlnpR/cqQyoACslsXZl2pflLAmrh
mo/hlfwxMGcvJdHc5so8fpH7qKbD2YIxcWMjpF9mIOlFd70LvPvbabkVaCAXmIob
eTHu8vzvTFKyjopxLfOwzYkWCoRdzh36o0FyTuY3eMNXu9y3IKy57Pj681PcbnEw
hdrq/QOhkT5RZoY82ocuwXiOI8zXnEAtpDkwCFMtd1ioZ56UXjwB9D68i2MPX4Ag
iOQSnBkb7Ihe2T24P9UFFkCfUE08ikreUEudxUl2LI1oSNTW20VEkbOB1sM2VXsK
iJMuaQBbM77ooVR4+n44HUpwK71I34U3yeJwam2ZwXGA/dLGMYAYuKiktcmgZb9C
M2JXN4ApeFH33AZI31pajco+Ad1M9bqRnh0UDwE1C4cQ2J03ci4egIrIrobD+rOb
TyBHbtOXp3n/Sy1draTrfh5wzjWmMGu4MaSDBhAyTwBKSgxNS4incymFh5sfxSfK
xZu3ODvumrikkQw9B3DIh2HXQ8yQil/QDVkFtNhnmYBOKJS+fXuOXvAP0XUPoREx
JrzVurzHiWexlc0kAudX5toegpzRvQHHk0ybEJfhcNbVLejvgqeQkKF2BXS/zFF5
Vpk5fVgDyBdp7MqQ8K5uFqp4T1ziG+Sg8pO8vsHwSRpyv8Q9e7srfYtWnFqwIgsh
WyNYp2V/WG9lg5Y/zkR9ZN4FZW8bgbMF3LTPUalaQ/5d/HK19/afGyAOmHPmDG7p
8qZS8lpiNryyRBp1fLEVS7TiTFW2hjw+x+H8mUWXSlvQfURUI/TFrHaDVzJ/2jVO
/pAD3wYubTGGxfTpVuq4sEvVrB23HBM42IJtrMVKJGYsCPo98imr9xk2WhFsNOwT
Rusg82UqdNybTCsIxyw7UnuwlCD6jiG7onA0VuK4NC7ljzbXKYlPScmRfG/2URag
zi5vApYxxfVK/1sbSi2B+81vUHsluFurWpf830gxy2W5FDTcuwJjkCWk5olGKWfM
mlUFFXtLkKJ6h4X5LJUjxyr0FCorWOBSYrxgDWOZjMBrWXXZsxen4eOb6vmPZUfW
PC+4KEcTYbH5JlZk64ZeJuEgAhzztTLIlAovXzPVGz1QDoB3FHi+OmMEH7ZCVzdZ
Zh7Tf7dtXW9Yf6U7VfSx2erU8MVn2IaqelDmhIx85LsUa5wVpm2OHoYGoYs6DXbD
/oFERP0phKLK53HfrIUDrCGREDFIbdNJ373YAlNiZjXM2a37ImnNsGj5ocsPq6eC
7QXP3ARkfjK+ZoATQCDbvEELZV22uMc0VBoCtfH0cFIhMPoGZ9WFLU+thZ98rSP6
zwukzCTeN2xVgNvndttZfwwR4Yxgbtyme02uK9zUrzTMZVbFsBuCw2gdD9c8hQ/0
XJvnvRBYZ/paXGuoMzIc8DRRkb5kL8ofZOFyVvVUjN+3FSQnxP0kdeKIY1XVYDXc
1Bey/gPR+voQPRahP0GhDxVRWbJ0UssGMt/Eq687NFpCehYYY6jwq0LARU7hakBd
C6IF9pzXGgRNuLSRwWfjj7g0Ia+PP+ySo5lpDnb2+51h8+hVssfyOnsCEqwJZIHG
trKq+k3lDm4FImo2Vbs3OjhpacfDByo3WNQH8EVATwT3S39MpH+go8iWobjiVG5s
ar4aHrteGrgRH3SwWAuN8fyDZ/Uh5Zj+U+rGLkwpUpnRBGvhAZ9xrHTjeBR7hEb4
3ps3iGmBAuxeYGHmC5FhIg80QdJilAQEjL17UHK5FD0W/KIHe78bC96ZJV9esY77
bR1r0K1amsdGA+ThDBXyrni+FoQiWqwr7qqtniwGGl/fCupbS4JuYtFc4pFsy7ab
xhusIXi7FKNJYl2vGoZCnJQhd+WCo6ZwVCXREo9rt0FK6cAi3M4+sK7be0Jt7zvU
QeObmnUh6yx6KQOxANfi70fftED+cXkLg1YI8oE4gH9V1LOO9ea71dYShZlh05HX
0wfMCssJsK89gUERW8mWpvNNDlBgWcx3fSM+E7mQ6ZfsRaseujxE2knVLiUg4Phm
J5QLj8QRpHLwqfQe8csz2WIkb0RWBi5y9PPK1fMR+EazW8HBd8teJ9NhFveLPUrZ
//UgkYh7ZaWAktXhHDZryla8xIyuOzLnE/vXZxaDNU55rLPh3zOaC/zv+CvKnKJZ
nZttAfiXZ+OgJTu2bWcNA7zI6bSWXVvyg+SxpnMxrfNFAIQKkexV7lA1ZpDbt/Wn
GoVVUxRKM9rswiTdymR+I8zC3NvunLkcBSgmvZZSkYQf9cW4jlmP/WKqkEq/YC6z
BvRlGacgIRyjbJ/hE2NM/nO8wMz7UARDhE+rIhwuPGn5cf9J+JI1xa8J1fxUyz9j
9mYStZIS6JyVUSIt9ffBwHApa/XrZw0LH9hdf2q9XnYTuPvgGPBDj7lNR3akWc5u
67oyDr0McGOMcl6Scel0FythGfZX+CAUfpfOegpVaVAgbGNEQk84p4T4ZfyJa6Ci
VzJgzwyl4E7DW79FmajCaHmy37zhE6LViYH+9Pr7O8Vfz+sJ+1sqOT5Of1fnNqHY
pTCDSoiKD2Yf5H632CTpdxevWERNdF/j4e99CFmgXmgRWXVtLWNiWq5vKw/knk9k
x2kDoM9XFcRMPxBVGG2dPnuwA6HCkJ+cPWlksJB9j9/VVQOOhEwyC2edlkaQuRJI
evy72rdaMkiX7V9eVl4KfRTmsIAWdTlwwmpnIRDMRxB63+TdpFkKB580zDxMPA10
kEfH7JlCn/PRCh+cYwOTsMv4MBXtoXa9K8grIIZS2azk0/QNDy8gFB/PO8UoC1Vz
R/77hGxM3Itq2ZrEVphexyAWvqymH2tGywyO1LX6Ewk+s2pT+PhgWsewi0rWb2Zj
s+INcqCZcbM1qSwOFcLJAFbU8LPBZxSMt+USVqMM6PK3GSwJjMrH6xqYngkdHxOD
4n+6JDWe+aJCPf6OSVUBEZSyikN8OPQkVKv7pyyq59cMYS0o1Hf8XKai84nmoRxY
96/8FVd+GzvNviuEFHAbyV5GiLOF8W0ilOcd6GFhYWYQCsLMjIZ24HUazsqfyv+D
gMJZF7TcDKMg10ZAH8fDHfIo+8GjM02YlbTmFdGaSjCmzKZRJGIajafG+acjvEH3
SuxxA93bZbC1FDr58hi42pG5txlp6Lf0Nt66MyShVoXypVv6J5RJp3woeZurbYyT
czHxUPOZVFNDicNFtAu9JEeANmSGL4qqiBew4l3xBtwtMb8qpeZEFtXczS5ZmQCA
ZTE+5EZT3yGugPNZbr3RPuxyYPl9+bR0Dbn0Qmja5OdtYJxPJ54UWw7FZ8sYZqAC
la/rCU8HQEucPNZ6wCil3F5QNpsw2rJPo9FXjYmhQQqqcYdw+sM86TwG4jAF+wQN
EY8bIbdiAJUZvuzom/SI4+Bb1HrdM9F6A7ekHiQnpLsuWFgNH3QQXwB5cCQI6dXl
A2CvPmpgV47xMbrWed1Ys4PrjZjSGRcz0qgPVdc6wkhTOv9lQvzaO1zD+VttnYWE
8lYphZ+0aGHxkrl0RjQLKb8qrjmU+spDcAl398SJGFs2xCbcGue2oiJCUuLHjamq
wacA0RDDdUZ4ZTIIiMQnRa0KxTRhPa6GcGm4LCTYK4qtjQ3u8zLv5A482r/L/o4l
p/KVbbHctHbczDUYmlUXyhQ5f0YmM22kDU3K+GpjQFmRwxEZex8uO4SGmCNXYQOh
9aX8914v5UThE+J6RJrx8peG37Is13XJvoU0PCeHwO60rr104xO6cbXNwEKLvLkX
ykQliyQvLnyGnx36QRPgXQka/IJ9DRU0O/zGggUsEglsLQ91vSns077MI7A4V7/x
mefIvGkDDQpAXIKxdYquCjd5BDNjuRvDAkRdfK0jYnbLUF/1KIbCewBWYEyDzf4g
K3oldBP3HHSGbs9C69u+PdOsxKlBJyu20IoW+rG7BrbzmsqWCeaP0CzHjAmMwXLc
V2lIkqSUmkG66S1Io0f/DRiGrnh5NQvaIHwvBvHTXZQ4W1RpqxaSp9ejfKhVLzvT
e1V4D/9syxIqwI0+g9OcGrdTusYp11xdiXSHKl5jibqhBIQDSIah3OWNKs2EFcg/
Ilb0gBWyuU4nQZPPRg961LzkA5OCueoez7+gy0AcqZJtlWZCfWWcK+vSTipqNofM
8PvesMfoHkFHRVDPUwuihCTpToCK4scvzs+ZeoInmP5nRd+7SdgMfwIRUuMmB2jo
xielb44y32cGf36uJWM0L6SrQAYRJp8/g2U2sX6ZWip5IxfEA46zKtdvdg1XIkhm
bRyDL60nqIMOm7Y9rs8Wdb+dAqRTfJJ/BqZwtfQP8QljiQwEnREKRpl0XRIyM+SX
ulVB/S0icby2YwUiu/dvqZ0R+KH0+8sNVigQ5dq21lOQNzZXt9N6VRpg+U/DExsJ
zv4+NuIKjwVl0V5PgGAA9nTyIQld8gTEtVeTXpmtLKtme2cbjhE+EWUlI3wkBvhL
kwVPXtXVSYS2Vx7kr2EMRWcXUpntZSzyuEdmpjeF2FURdFwL/wrhCdX7BW+hh8x/
w162dUBeodAzGJjnpJBZISaUYNlWmT39v4tsE04+8Y/W4YQJEGkDoOIlc/6ku8EB
6ONhiYwNEWfkWOgNTkV+lH9e2FspK3wgcm2SJ9cCqjg+nd6v67MqNL5WkPa/WHXV
bUBgqb5B/RMokNVSKfmkTSWB478ZQw3NKEPxHKmx8E1WzNE+15/ad2PpfyWyQoIj
sfMif6XYI8oNSqmQxF0TtqAhRsvURWDDwgc8lae+QSHrsSUjdbQyGGMB3L4psMYL
NCPVbyHOzlpSdIRI8I7qQeQlCgZrI0EilsOmm/hKNeUoIwNrBd4ZpzQsuz22aN36
hse84k+pXD1JnJhnK7jRbIdGB2AKKw+kDP1Cp6VN7HZivZtJIAVhXN+a3pYRxKOw
A2dqHiU4WTln5F3XYcbCe14wB8bkOqQBBk6YkvlAvjfza5xDsA8ETOqftGq3L+t0
uvSaQ5z5FOg8nCvy8VQxoY92wkaYizHqmnl0cDzet6ngOixc3VpZhFjseJ++XDTU
k8pmKbLj5gAnei/BcCidLnFwEEUbMEDZW4WePJ1apOpwaEeB6Si+K4y5ylxjpBfo
kAYanxfcQj9nmWlNB3MxmBGnYnUunpeUuSzEF+4ekLsurijlsnxeBio2kKfLt6Ix
tFfckSW52xa4cwC2phw/IXBVPNCet2vAsIvUMzeFFBx4zvdPnXoPuEq2I22SZtz2
epyyZGphZ5asKJuH6KGS2EvvKmBgVbmIAneSYhxrsaNbWwrWi1JS9m8Msubq0P/2
ntjt2ffs8XIDKspz/MRIboudRQHV2fP5kqd4nJYaZuTofWEpdot7psGVXn0fl8RT
4ZIlhheCbZpecTZoS/eS8JIeT6ofgJumsptm0+93OCtXVFH4Nkilzega0wpa8Bzb
uvpKf3Vo/9WHgrhynfWy7GXD9nVSp8WddjDl8MCJVO17YYb6D+24I5A3S2fJjVh/
6lGYrgnEWWv4m3On1W+UzIbrIFN+TEsZ5GJ4NNS2NDCE9EyN0jX5egWS7+5os3o6
aAWl/76z/NcYh15SP5ZAZ5zy590jCNDA9QeWWdVAF3XXFFJjQmaUmMVoPrXFFHh0
vyof2AHIvs6sJAwNE3hUOjyuCD1XOmQ+lWYG0vVsavMdTItSnYoxeBc4ersnARwY
9D+lgWsMgVLH5EJLEe8mZB9Y0TD1H9v/GuGCgSwoqMNKhe4OWxhbZtFkIS2g623L
8XzBkY2K2Tjey1rYNWJI7lLquxey+jlnZusTY1JtVKJTIFNg7kXO+73wUF5uxh5u
bMWddEHty6qMbD3FAAQsO6O6437sSz+kxIzKCxGqs34xtgErdW+fmDlRFjMCU7n4
H+oZpIZvdolWTq666i6FtG0TU5sNEvRWcdnqV3xszG/ZAg0MvLqar3/MSWK7TIUO
ScDun9AL4iVGfHtqa0pZbEEwZVSixrSZiCskyR/P5FH8K8GnoNs4KV+PVc93Zzc9
Rl5nvNMgw10FdtDt8jLkwtRhFsDacUfDUrG7Pr5AyPSRUEW5hBLG+fmPpDH9LTRe
FN6JuNFMMZ72/ZC7uRQuYB+xyaM7jwztSbf5tB/PAG1DzfHPkkXWk86L++TmGr2S
1M2qs6qXairVr4wIac5S+gFUzohoNKeNrEP+tD0p0F8OrNZO+bQmYHZOZK7GZFk8
3sLFxOl1j7CCuZoul8P2Em89FxdD2mvgOKBjYsprXYvyKEibpUZYpZXpfdT+MMJM
33CqmjmhcoGdjotlWhSSPXeiXGTPDX0eFTYxaJGwvgof1ojWip9rXtVnMfrAyWWf
HuF23Yyez05PljeJHGhA2PUm7cNrDoZvgqekyxx73hUU+YH4M6zNo/yYDkmBq2wY
smHySIf5aV7tY2uKb9sllRuUCcLB51fY/ejCJP7/Fa63oiP2HBWWIBs28pABAHAN
JInDevvayyNi2dKzoXDvuZp+CzmKSrsAG9IMrJzea9e6gHEZ2xfsXbITmSMmvxFz
q1DpPP4nPMobV6DNBc82VFf65jwh3L71JQiUrHcwYZH5XJXb1NAXtwnFczKtMUE2
28N+PBgxnjKjeH8qTC/2rfCHJv4ILLro1h2dM3ihAUHDnY4WBJGyqNDzfXE8qcSu
IjRLUn3NJh0fXqupaNCXMKKulJy6pEvxfsvjWe2f4w2WIhlBaHtbTtcR+GUMbTbW
msc4LXhBfyt7SbBB12FpgUjc0HdyRd1DJREJuoEgPdXIF/a6K3fBtVInslt6+4Xk
5dzbQhWaBOBkEDx4YFb3+De2HzCfXN3O86TANCzA9TSs2mQ4VLNjzZm8Z+fJpEc4
2h4s0x07FfULmISFR3eBolgCyEki8a0p6iyZR3SXf7uYALOZWnuP4txwPAiq8ii/
YFDFklTZQKnNuP5xzOM8emDfBQ0YfI4M17mh/0L834q2o11RhKr38Ck0WNwUMNee
B+UnpfGUNK+ntwOOKtINY0X3UrOjhpwY1I7UcRHe6t8Xuh60b4zAMiKvYxehYfpD
QTUxe3M2ad8THhrVakRMkQQ892uMbQW2fgivockU1D+TFqwbX3c+5piIx1VU3UC+
Azd3yiXCntziiSAMuhBlv43RxcS3ylawXDb105nJHP/IvM/2wTEif9p3uYqn2X5F
1LRh8JhPaRnH6gsT9UIDZqMczNZWQR8g7zzXN2BvqtSCCnHC8vSuaxltuvEwVLBb
BnpSvqs4EfdObfWKh62O8v5rsMjHawlcD9unVjt9jqilXgyHQlgHYHpgZ8UNa/NA
dwv/Hn1U1ubDe26A0EqNJknh8kwp2S7HY3wz9z2VQ4WGVyYM0Ht4zdRMNEtzuY5A
B+QKLCIr56xOKR0LsJIFNrYWj+r+/v7oyuywqto4TagC6HYT0qvUSF52BiryqD/A
xJNphck+Hu9uR/NXP50VePAF9OfEP9asyMDZ/ops4Jv6gFQKB7cmPw/EFMP1lU6F
u6xNeEKGrhDL9n1QH+N3XmPvi8XEdgLlMITdZsvPMy1b5ai680R8C6af1SEvOgY/
M52o+uLVfwGLhccgiGdH/2bxYex3VbbwzMPA550XkQ444J7is4RxdtToKBR22wPV
5r1HIy3sop/8XSAjbkmpOx6owz2yH0PtFwxhNPbLBBfnjTqeokQouQZIIoEov8/J
SDzC1mjhpNSpSb/DFrZqPNnxhUAtWkwz2NFL1tD5EJGqOEI0vzpxQ/7VIRwkJlC0
LBrEJ6Hcguw73ZuTCQ7wJGlB5g1hfiev9+xn4M+qXdUkqvFyz5Ks5z1O6T/SkRw7
51EO9dl2tFBV8TIyy/I66YcvitsUafEeJtVAGiRhC3eboup8khyLeVH5BIW9WC5y
l/BdX1un+3HXlGqR8r4WInmG24HOU3agrXp4E/zznLLpXoluSLgH+ULXFi6PrzZY
nBiMLkdjGY5QCYVXpmYRUlLQushkzTa+K5xx2zr9GLKgBDsBkgPxfDcBP6UK3JWX
E1iNbXSgf/O13o83pv1lKNE6vAyZbbqlvI654jOW1yGLJzTejh9/w+d3Vq2OL7Rb
LlahQ2LwHheZqMW1WPXbY7JElKfc2xaJ1UuAV7+GCQEn38FED9iOtOONlvUzdqAn
e3+VsRcvzT2RY6+ihGA6rNZAYNWZnLXLAhb5nr9ax+2wb0FdGUlQPiZWE8uEaQHx
GgH6asTx7oxH6W368y0IUEJv9gG9DmiF0L0NcTD9HUaHuV9BTmAJ3VcaVrxr/6I+
FPGwp35jKOvEDAb3d/Vy+v72MJz+nXZoQ4dlYI8heIC2tr+mMSpgX4TdT3X3FvQF
K/ZeBNV9bFh8hvURw4ftZSldeB1mQJmnAHcsr2pD6qR8GVy0aa//6h1zHXEojA3C
/PokLjle+HLPGysl4Lym+SMGdqnF4ia0EK0Nibx2nAH9u+0mCx9JhzNbC1Y8sxVn
DVX1Piczii5GiwtulIJz7ei8t0pCtu+QyhY6cbzN6CnXckzEWTdyPghs4v6u9aFg
n9T3DsmcOlJ3MZyuNh+UTzDt/U6lqL9OnSd7A3hKM3wflS+GXRo+2/oGEu68COeB
fvC4WdihZGudrDpzuBPyDAsV8Wbqspkxp2W3A92FZRuauIfrvZxXl1HA/dBTuVss
fpiAIf8f7+Ad98pxbjPUkM/7qPLBML4LDutF8mW2mCgWiH73KFh5M1XLpTZbZ/Ey
Ff1LDBUfId8Hvbb5t3xDR6AJsiOFLOpKtvX7OoXenL/ABYS43iGstMu7rrHiPtPG
pVKOBKXFR5gGwj1dDMQ3mjWlUO9kYYLWgTeml+8t4TTPsVqv6nSlORZi0sdNELZc
tS4I4yJh2/mhvLq1SIgV0AEXsD35xwNAb1J7Ts8GWgAKl8lHcA1EnsZZlWVzO87o
Qv3nJ3zwbeRf32h815uoSTfMgnz/6EEALPl1v2KYXUHJtWYFWJpB+Fs5+JwPxLdJ
0Pl4pTv9rmPDJeU6Wp/Jwxl905hPk21cbW09dfFWdbzwXdiAtDGcUzPLhhvB6uBF
nfYuocvAW74uJaA9+l0G5MXp5wNIB9ZWstvfOq3Y5IOOM4lkFp+mfDQ/o5yJm0+P
DRXym/CDlkSINP6SABljJZeXnJ4qgKhazG2kF1/2K8RgNbCYAr8ZZqgboMd9ezRr
I7SkWcokXP0i0egJEoqMJXts+WXE2Y315UY5tksN+8rhkzqYE+K27nLAQKI0tyzw
bZsk3+Yvs4w/N3JunYjvQoGlV/qL63bjHNR4CqbmCXLBcMPMqtXiEvi+/9wN0HAn
5i88Z04utG1P/lkeHpm7bdLrFui5BJ2uhzOnrMa4RA0AgOTNj368wttdMsDeWlM2
X6blBOwrQLpgmZHQsDOeiXoncndLJvLpXCwQrjcWUss/KvJ/AOryLiwGbN2BtyRc
tFchZW2mPfE1Imfwy7hIJtzF9dS0ibvgv5AjHHj34lXAb/ztGDUc42SIbRa7mRrO
ORmXceUG7RPNEZAOSefHe+qqldjPZMnoGB+kXaYdYzL8DR8vC4KJTxDu2RPX8Lch
bX4und6B+siX8VBqNDp1dudURimQKys11Oc9W4JROcpj4r8NNrnIZZ4IvCx1z01+
Ju1AMIkbuEcTLtl/Vg2dmomyO9cAP8BZxfOb6fQh7/xoC7Y6WTiOUSwHGyO7jZGF
eEh3gejCPPa6TN7Wl1UDBlhDLPmnqNc0nu3MZe0LpL78WcPURaI9rsuR4AnVj+BA
NEBsU+smGYzDoO1dIZkmP4gJCSpcgMrm+RkGtibnQaaa1nhsE70mAFOeTyp/MJjF
DkY3vBWerh9cKSMa+tNUsyMwscx9L1ztEiHTaFlEcK743HTqvtFVWiGDnZ4g/qQJ
oimBk1vlmm2ED0mIS/QxaJ1pTS8v+v8Fa1FGp+3CFciwh1i9IciVrlNBMOJizCiz
QynswU6S9TovcmA5Cao4LSq88NGtGhZcdk+nnsoM4Ka+s8LtLVN106EqhDiBEbxC
7FsIg0sCj1CRKtZhoJkKy1UbfqsNM/ZRFeaI9+dg0nHD5fxlSpJ2tjN9y5TsvcXq
p4v2mYUPJ1kDtRttyUTCUqSCxM2WNTJ3AFvxK9ec5SwSzVfLhIQfsxBDYbler900
zRukYyPHTq70NFPQMYjmFIsY3jmJ0HxfGyTbT/TCMjF5BWwuPo0Jb0Fd81erXpCI
dauH2BZ7jvBdBunJ/N5xCvM8AME50czh5R2CazHfyv1e58nBiTLWjxiPmovLkfqE
pc4q94G6AGwSyvVb08nw/Gor5QVTlzCBYok2lAzbKheAU+HKmQXK2fjO9sGrHAw1
hTAnleawgTBa81V4wQdjD2DSR9lfWnf+v6/p4B9wWzwAitnOnjfCoWpkvBPCv8S8
Zw2tYZM5oYZHmbezonO9uXTOUf4OVCp5GoDKh+1H1EoNgaSLhmcGLJh4g1jvp/ds
WLFn+saDqgmEdy9aObIjM4GnTuVlZJ8u1/IGLru4xQ0yu83LaC7qfUNm0Jd1Ugqx
HOoNtTqI1zzU9y7emZP3qauCSfWdHuakz5GRMvi+bLZfN7vzexbeXkLDQ4v4EBhd
8co9d/t5lV9tH6g+dfa68Qav9aGuhNB+vyL+XfLeNtobhAVk06g2UEk5Nf13rUIU
YvM6j3mGAlWmCdGcTgPjRn9tvWXHjapDBnoUw72e83FRa4OdNcdbaAkJK98YOEC0
gCSzAszwSJiVg+MnFdgLwcG/o80l/+zBeFP+6hCTa4qlfhizZjbmQTzW3I78m2tt
Gk3HGXimxKJLEeraFiQP0zTx+5RsJUio8VB8L640GUMvXwsRFsTvM5OeFqSRzBCI
PgzPtQVUard57i12HEd2I3DyysrthFucBInfnmP38eadN8DdjoYs2m0vmkcyTPXI
eBHvAzJWmkUsqKLexFMC5vio+6imjVzZXVgp4HPZc4J8DQllsvde764URv4IBc24
cdD5xcVp3eT+VNS4fRU306ICx2sNulG03bq6B9pm6SY2TVuhIsGjFJwbq2WmKIDh
aqfEZMrtA5vLQ+VCbnqzwQemPBRTTsbk7059vD46S7Jyua1z2+vSjVK8hAXyj0Dv
3i1Jg5+1+ml3nGU7uSFX/ikKD8KnqhIpTnj0XcObBWW+yhjhhZSvDOr2hFDEzQrt
ecBM5ITTOFPtBBGM3spGPKucyAxeKqNwN1rbU2pJxv16sw3L/dvn2IEKeqj8qN4t
1xvDdyI1yH6R7cqJ4V9dV7td1gDt/zOamSQGQ/fGBuHvf6fkKs9CrCgxJM/HzHlv
/TPJv23N+qkrr7YPfn2wg8Sk6RmkxKiSFJa77z3VJFNJwEEJ4ugLrNGZJornBrww
AeiNSboj8Rae5CjQIG6f5n+JanGXEIK8QzL63DNpUgbYcdbRmgFnPI2s7EQ7DfAI
xqaTQyppb2TWrOrBztKMOHaiEMbPYsQYKx5L2IMjZcP29JiE9cP8PoPeFkDsZkPg
88MJkZ2Ystp6+kDH+S9pAiQwFhkkWtIL62TosXwbPbNHB/qk7m++wALvZ28Ruiye
zzMT1Q11ukEyr0VEOqSSahzAnI7XT7NJpkPyE9zYsXXkjDWCIpGPh6y7bzqEHG/5
wfzm+Ycsi+HTXFAcYy9/Xgu2ZDWrGtLUjGFgdr9VQ1Sm+24ye0WbEt6Bf1WbzF32
Cn59tEP9TNGu+KeClwbA3WxOBD8cvCTTAA7wBMBJ0r+zurLqAc4PnGfR33xOuOsY
WOQ4pecCg/Xm4cLysS4g5Uf3V78gVs5SjtSsESM/J1x/UqblrzRNhuYSS/sbjvXF
Mdkj88Zc2tDsbbi5Yqzub5teFkWQpFO1/Ye2LtQGlq9Oj6EPmnyTginHPEpkLjTG
3oU09j+LfEwoP8W6yyyGNiQw68VLm0EzquW2aRQn7fV5T2nCYeFtxaRb4d2Dod7y
ZoeJt9mLCaMUeSjtQ/1LdFTaVdJzTI/9StkvFyQKTJUCulnULQU8aSET/iR0bBtZ
/oaoaE6/AV8kNp0AhJ6v7hCDvEsagKzzm19WW/yQVroE6zdcSyf9ECOXDXEXtD1q
TXT6Olxk3jasATSF9MjkLnn6R/Vkn02kURtf5nXbdoMfnrWAZPn3HcAsfRUmf0ZR
rIrRk1S8qBy4L3yjwtrA0iWaNFXcLeMVdOF2zbO24rUGBk0tyD9438woBOPw3ztb
Vy1U1aYloaEzf5rFa44nQtC3o0D6tmtUMHeDQ5PUFa9BUP8AvmN/rk+76AX8oa0z
qLzELmKS1o1gCdx+XbpIgVX3ItZb0+yUmIieZgzx9EhFzpZH/pnqhoDGLH6G71yW
THxmpwLNgg2xMsHsMFRpxZ1xfxRyMzKsg4PG6NLYcZ7ia86T6BGzxMF5ljQCDlct
Evvhz9yTg23yMg9YO+8WeP456kocIDIouYxVvBCO+7XwyI/QIXgECEVhlauHX4rg
qJ7nHXc68Nh5rtAiAR3By3vwaqroV9w74nRboXWINRmtPBmzEg5iTkFc+v54Tk1i
Tux/P16PZVY+6l7vYK/tnmQVpfrrkDiL8RCOTgAHCIGc4NFp45FBTjHQjDH9GEOc
ic8Oqz3iw2u2P0LYpSuNzmZoTKWq7Sd+pfKULAJrL3du0/oxbQCTg7KwNmeFPpWE
ka72k4QNQLRCGAio7FvxutA4aASQxWlgh9pRpPMzVMsJPgWIUuyA2vMQ3lj0PJza
7gbp3D7dTxUC86QeoThxfeMlfOHEU3/ubLs5TwpI295yPBQu8GB7gEm9M6kzrjME
2Dh0K1djDONNJmldRTGFxNvCO2OOj2Ii0Yz1GOT0ZWD8s72RixsWAbUtH4ZXntL2
lMon0Epv3Zg6U0Lq2BudH2NRM56784R0C3eBy7WEavwMX3h1AXKy+5pEuRd/XWGc
hiEG7/WGLoObISVBKDvzxn2ykQYyShi2Xy2MCFlzU6NtI1O1p/saazB7b2VQmKcW
UyHolWUea/IsjBX3M1Fh4pSkxzLROLwQv7jJtRC8uaMciKyKZynJn5rttDqVhRca
FozEQpMnPPnIOgW7PsncAt8k92xgM+bYhoI+O7QFQtdte7kQ3Bg1lBAL8uyc9QQt
z08gqcYQmxqc1l79Y6Z+kk4ds5iE1ejOj4v6RcQH/YSmWVZzPflWfZnw6zGqiR1A
tqPoIDyh6QIim+aBsVscMM7VrtyBncwBN3ku7mGyh9RpngKWir4kunkXeB/Rb7GW
Xg9gAUWfksY7B80Z8VZR1sbR+UvVmL/7ESLrIlNVIpsx/6a7KMHgdMgG/G2j/+No
FGqvr/Eej347DM8D6F+BNZo7DOGcrboZbSz1S5ESeV1Ga4yStn7W+jCOPWseezpw
pums8rhbsDF/AKcVWjNxXXLcmfGQGTUqsgxE4U2teevrEAknTPruyIbUsWb/NZd1
Mmv+QSj2HVmAcx9swQE6fBKSbPzSqw+BYQxaR9ukDyGtnHEK9k+51R6fcCDxH5T5
rU2ZTHVsp7aynU755OzFrD0HCyNJvFCSBQGgCRwkw9yyMfrc5BTMPZ29WvA2xDbC
iX51rbpJHIQ1FKhH/blBb59FgJUrbp33lHGfbAJQ/mL/js3LaTu5fPI7PYf/ekXB
UbffDlWLhM5pDI9kRjJ2Urb00RqVZ8wN66506tLArO8P7c5q7J/zze5t8yfj3NY/
zvB5INd9EX12HRUYBC2r9mTlz4TyawzOzzW+pfrwEpjGi655+gAGbdfRkj5lzXLr
z76o9sxB9gBZ2SzB8TEVQIuq6a9zo//+KaIO8hheKqSuchOpl3ePK55/PM+ivKT8
qclcoWEgGM1bYZzfRJp8mH+SwXhKPmrHAtGsEIrGkhZO0NhqauYzb9ieOfWLLaUF
nD7qyvvjVKk5E3UOhPCmXsj9o8tQnQQ2mlRchRcCgY/sfhmQ9B6KE0vrYhKOLcHq
cRLzg3uZOch2k7Hfe5IOtzhJLTGqqp643WkxKiASBctu28MxLZRUuhzEZV5sGQA5
R8+NDTweuTdLeH6lSa3LE0wDV/TELoSsWQhFQxO5KJJ3Igllyr+jFZWLO/fCTaZN
8e7R3WJ9CoqZtzfkoz5T/Sq24GK8qAThsglQTGDKNeqDRJPwW7N9cuCE7bz66gH7
M0l0hWDkna0xgeYnqXdmCGhxYdQfJwVv02OGlVBX5XQ/l/jKmTRqWg4lM9oCXiOQ
D6Guusb5Wb5qmImqRzEJfhk9X5FgkZ8HUhUWT7R+g95XACm+ryWy7QG3l+AtWsIH
xqMuEti8b2wl4nV7M0Y4aXTTvSTfL1k273aSUFcaMSmD5KwDY8G5/WLSqqkhmUvi
jOarlxfsxu0AL8hdMBZEnbKYVqMaBfLSjqiLpr3SNOBm1tyxmMhNA38HKyh4a6w+
AEiagUluMf1Z+SMWmX6GQh3d/az1SFITVvHKNruNpHuWrVcDoruPJBx7pWYn5e64
br5f6UiV5nldtnaZe25A1iGq41rfTVPhHJgL5wc7norum+lxfuFj7HqnekgsrxwF
zAT57MQ0A8s9XSplNzqQk2CNd08atKAsaMqzwv/aSfDpSwqUwwgw69tZGJxlVsZx
Efq1GVvvag0DitcZILuQUUSWjdQQeP6Eboaw6i+R8wdSihvfEbpqvZwXOwgJQUx0
Zav20me41PJhJg+D//ko7o48q5gwYGUNPYZm76e/ee39ZXYuYFHs2Refoo1u20xQ
yxGyigJZoaY8AE/WaQrzWB2uFvWSZReif5QsFzFYVDkRvTZhM36KMMp2qCWQHOas
W1ASetuuaF1WWY184+QnUXVt0kTgro3nVclz4pjMRgMdxSHafsTInkTIL4/zaB8A
ETP2/GT160Ppyz2cw+WbXwQD+GZR11t1crKHr9C3ZBiPxTWWApvXOGQxKqoEzumd
DmgQ3M5MGTYLhD3vUu/0Z5h6M3xzg6RkaxLwhobSkpkY9ZGfuGjUr9ek8jXW98S3
zZVX4VKxiz6XP9hbwBJqVIjcomvwTorDi0iC+9aBNUP70ScV9DtohldO4RlUpcV3
Ese4HMkY/GjvbKjc11dEpAes6xD1D4iqn5YYHe0lQH2GZZCwHetCbLLxHHRVJRC3
HYBzUwVqwaDiNJTkUOOdM2hr49vINgex1EBnEp/mPpsklrfD1QS1t0Oox/s+sOt0
T0cScQeHm8qjfsLZYnaeX8zA/Uqa51WkHYnPl4Fk5i3RkmJzRmBj9LrqVGRCeXCG
9aenwBPpctk9pOloEyUL5gBfFFxcvAAxY5WMcKQ8GwFWymKDcuOay+NnXWMHG3YV
T6m7ONVCXTiFsBpzd8Xh1aAzvZZmm0hUsi15Xq76wB/jkG1+6qWBu/5dMihXmgBE
9u+5lcsasey8xxIcMQ1aRyasNcx2+hnF4erggSazI1MHiTIdi6tn9zmFSUj41pPf
nRqmMrh1mEJwNHZElXFhV8TFzrzv/Y8pN4K2UMgrhJ0BRsdFe0uz2Q7YQWwY1gkT
9MDfEsBdEiuGGkzZmH4ENSVDfyB1bZ7lxFPu8136fGWflic09LTjjMnwagCQUYzE
xni/zmVKQyRx1QHBy3DE3mN+aw8Tws6On75cKXAY8DgFI4CTme2mGjCmjSBqS1e3
aMJFVIs1UjYxVvnsNiff5pPklbqRRkxYFhxT+C4fZsVakIftg6FqGGO0tngo1KjR
KL8CG6dRuZwWHSldnlAXFlaKxWWVnEUW+uLE0bDMrS3vbQH27Gi0Q3nNEyfog5YT
GkcHjygNUXgh9ENoKUXS/3ERdeizVfYYvT3imDNspCAs3I1KN4catztW/jc/QeaR
ti7ICr+tOiVPP2Gx01Pn14tXg6px5KcqRWhPkV5UwwU5hrZYzoUwinBcIF6ml942
kmYqEsPBn3i6kBSpldV/Pgg0LQa9/DwfuPpE7TeEKZ2jO79sy48jjwix16YM0Omm
QCnqaTvC4dvbRw5+GkL5zJEebBMy/Egbx0w7/Hg2qCw7lz5RHuLb+rfrP5GAo99w
R3xVg3Cm3y126/QIulgW3A8GUsA+ET6c3TOKITDZkrp13hK9f68eOR3N5nhaSUzP
gMKuc4ow7A4c8Ho/zKMQCuQZK4rX8CODn3bYd9EZCsh8tDdvUf6jvdML0R/MrfRX
4PDxscNMtyHgZZ0A7x8QuTFF+0ThlJb0JMvsMySh2nt76wQrMaFx7ET9zr239EA/
KRQq9+ZYEQEu6kWwLbHGhVyO5cMZYWbXQLY2JlhXOac/PVA5dgN3Ja8MriBq6lxN
TSRpUk8yMqaXsKrfGRouLyuD/8Jvenl4QbtAzXfWpEyfgXMnu6LS4KSrvZQ5gHAT
9HMuAbOPrWiS3adtNMzAOqk9dp+c8Jra60SQXNnKSKxHw/SXNgqePdUSW3yL8mn7
kOBCOmUTyr0Zr4lCPY/u8BSQKsIZLFK+uBE2Rl2/Q5jBfBJi4H3Ecb6xbF5ZxJA3
pMf3iGOfm5CvbkCSi0rXlpWRKjV9hUhrsonjjsrZiL0jQLq/oprr6miCbuiu2aYz
wCXvxtmFToKMUlbzuFYHDB2epGXPsoDDPrMDd7eAbESVDxKX0Ex6UDLrzBYYToVf
LTfwws0HTAf1vitzJa61Y56wtDWdZadcPQhTxSGHGVsdy+cdaRSDxUQCIdmdXg2w
fOv8NfTDeEpESEyWdblNs7WAML3izDICqD17ep8Dnw7Y/55wqpqtTkc2OeTwnHxp
/M1HdCptzcoHojv9v/6Z5VNmVuPJx7qRGAqvDpFP8+N8+iS7i4/xFt5VqHx09BLy
fqw/byCy/4W0dMdFVLuhA57aM+eXaY96844pTFBd5NrqsC0vQvj+Ldsp4I7k0ckg
NXS1QhLJwhpLDql/2AjHOHRn+ia5zWZxmJWT0pMp2LNVtIC6iaPeGhivP/gDJn3H
jmVRFcw49mFUjnBnaeu7c+38Cp1Zgc8a/da9OB9Hw9bv7TW/v5RDo5oB365DnLCs
tcOKWCs28tll2Icw6Ja8G9OhKNekuTZp+V8KgLqVqRsJNtLlC5xf1L2giwnkkhmo
iR/h70GC7dqVPlMTEldA5RYstQgKsA22mn21Jc4j+q08FibxvJz00VBr3epuQbS1
9n6gGqbiYmqyporNL0kJv3W9JGPezSR9+74RcmYm7aQZ1DTvGbF9cB5zcHAweBxP
cuHea33zlYtda23Kruy/PMrjJfk0gKWTIbanABBRKHx6bbauWldsx4+kc8keI7XV
mf93omLHO/W9k80rFj7zbMJhBG+fwpqeQ1punGbZobb5b64Au/j/mntHyZ/Ek8Em
Md9HdfH9AETKorufPjCbLTJS1HyPEcA+SgLoCy1dSfX+Go+Xf9gKxfErbCIwXH8t
U+KvXFT4C8pffzKiZRgv+7xqovHcmwe2UpItr/veLLKUb+HgsM+Xkv1PUR9TKHWn
xEtG3WsReQSIHsZ7cLxrbMZvjVz9RySCNLpYGLXvW0GxX2NeLzJtq5tJ1v4KD7Jn
8+JxlGOv+dqz7mcNwQi0GmsM/IrOZmh3ahn7NVu5yctFKzKbAafVXZ8Dn99BDBdq
oEz9HHxEtxIhH+ljv4BXGXvhCdN/TtzyoWxOcct/SvND68XUjDnw+FzM+6Mrq6MO
3X4rA7mTn3a0sSJj0gWfAh+i2CppEWeIZ0eiRXHw0Fl8KiA498+Dm9ChID9vr6QX
ELqxfocyJgQMKnivlMojB+UaT0KsiD+81MQHkVxtJujzha6B+315QOWIMDQTvLaE
S2DFEY+VcSYKjZ0wzeAWh++987Cp+FMwTOLDIbE0W+zWiB8XN2lOpVy2fwojb2XD
/3TVreTVL/KGW2dtsxYu3ZVm1vHtR/6LQaxPEdmoGOcOPWAlMaoM7rpAfAojXCYZ
FbCPDvvz5rigXar84TRE3jAFd3inYvIXGqqne0la4YBVJ3mVj9byntfmlmIt/af+
edKa/o+6oaJrIWZTwqyALXiPJVFr+VKzGgZvLKbUlc9cEO4g4njbF2jtRnNKj5EK
I2IBOrjTnh2UqvIUpL0kMjCBBs9dvlHardX2+YSG7ewlYeW2a+WzBsuTxzBrgNlt
TM1IYg4fsGfy/VNEn3iGzZqsmXm5d9vm7cL6O/TleSzbSkL47D0QkavuibqJ3MqC
/eCF95xXWRaJI7k4HXX9C0dSwkA7kt0P3va5gIwM1ZbMzGfnNfGbWgIJKK6Q+4C6
WvaVUVNn/a2vCCRZvTE9axOfqyT9v44MnBpixcQANzlfV31EorMhr+078cc88SEC
kZbLkY5Jk7YlxaE7lz+D26cQD8bl5LVePIITXE303EHw9Z1VTd+1viWGpwnBljNG
4oTZKD4LJlRKzy+U4MSyZ6MiG/tb3UZisgxrN2ZypFIZSID5jhMiUrISciRgKzH6
Ky8a+4QKIp3cp6HwOKr3fu2DroN4CjK2B6YeFzSSM+g5JzcUfSbaGxsZUevi4o/y
RhEAlo4vYZNW8oEmGkLslHFOFDZfA6i+AszIWVxTjJYgQBHWgS7pSTS+noo0Mmci
L3m2eVdjb4t5Hv0dfAA8wEBXKCj9N4JYH14dCP5mswy1Vp2H6fhNnWLhHLZbEmWV
c6xqTV6F5rFPwzG8oec3Mdp4cmtdyIleKOc27E+eobreu6NeGiCQqdRZoGq6HxM2
TM8d3VCOT2uhOL6t0iSFnWOpusIpjkp68C1oWTMEXx5a5d50Ii1dg/wgHGf2excR
cVlgn4Pcht4QYJ0XPdnUV3K3+9vx6WQKFZnOOlpa87hEYLMd76tam9tgF/L8ZX9M
fq2akxYMLSIq77RqGKB7WB1zNPCIXqBT8xRDVLGmzayxbgD+/pUbpAEQiNAYgnW1
R1uSppVNIhS2gLP18QXl8HJwdMcwQnzfkJX1libv2UAvWmltxVoVr0aZJ65DLsHC
rSyaHfYzbP2+EUjzSrkaos4M2duimozS/OJWcOvCVGeO7+ygNWOfy3O5rDEY8nPH
tfAgKOWPNUul1822fjqBMASHh+3Bd1LXJrG+N3fLffBHwbiVtBVuHM1gaMvGB4D+
2EC82LQpw7SWocRsFrpYYQFgkNFaB7NGAelC3tKkOXV0vnqfO4jMDG8pg/KNd07h
L9GY436YyIrC/ZG3QuQ7dlf7b3UTjqr9g/sUwEtV80sDWYmWwL7ylnr/4qn560o1
LXJVtKeXqVYMsCnB+HQeXrD5kBBBFwtffI/f/PV1PDmSCBhlAPpcEHrsAMu6iqHV
9i6HZZUqlTO9l6SK+31ONJW38d7Wwh0NUwF2re2whyH/i1JLdBhmGOXa4N11Ubyt
e4pZSl3tdGK9KCg01XV9hry7XFQlbS5e9x+kfgoPpg+c2+8uPmouwIUldqW2F/ch
hiIOejEbEFSf8jsKAtlX0zbemZOyEouPLR9EUcB7SmAo0nj4rNs4H/FdKypJXr6b
BbIpLLD4V6ezg7QmHHKVEZg6egermYUtU1BcxkpXvhs1Da9RcV1r3GfhNkINLH00
MxXxEoe/IoMF7SK5y4wik7cVkJEbXtguNb7o8HrfGwQ4cxyKcR7qoGGgty31+LCT
IOyeWlaC0W0AQB95jgR/hCFSnrXFE4m2hTqTpOJbbKmuoruqqt9tHeit3qgt7/HB
YRhiMD4wpzbgIzFW+e28KXu+5LCjOsU0l1XazQFMqBOQgkTyA+TQ3DwCKmY1238S
srMEnGCgiYx+oPsVtBppOpiL1lgH1OzIRa9+ZBHtYaTYOjSo1Z4WUlOmQAuxHRrk
ZqbmU/IDVK2W5LYeIgEcZXybapAVuxIDzEuhVVySeDPIsdGEQyiY1jIp4V9fKQPT
4H0d2cVN3HoeNVZFBE0U8qUXaod6g2oMWw4sUmAiBJotWN0022YbkGthDuJQgoTM
HH21jc/lz7KzYk7j4BXIMMVJwdY3w0IgdW7lOcoHvq6TX/GPdTNjQlWUbAhyZhUE
vtQ2ZW8alpS8Oxy13e795wUnBV4SqoQc5eT8UJI325dAlnPm8ceUepAoCJ4IvvhU
IZ8f7vytlqbAdf6G5feyshLS8e8ExHcl1eNJQ0JALUHObblod742tqWqrA3HUgL+
w7Gi83HW/s8D+ur1nX3eIsOxt3pMs2Re25EZE3yzNr1hyEicGzKqVzH7CuCTyJeq
s0Q7ddGNG2Js9UOZwDh50UD19WWRrTDgtczuivtcAoPvHF8ryTkR7SgB5xszKddw
5bhHBG2MB5I37Ka9+eyprFirMurnAJzdE4pSzCRVQaj/EHXK73cFWizeAhpmM/j4
vrOQBQtH0jYMdqyh6pMFarfycikwhSqxRcL7HVpa2pOS21JpkLgS7em/WwGDCaJC
QttOYAvqxsip8BFsqeRoSgMogjVsxrWDM6rA3+0PnfzPTSlFZ4qU26dVhWaHtVZ7
GKvwY1rQgtVICSCo9J2V9odh73RWdUuouSb3dUt76Q+rXYd/WXQOReOs/9PeEMap
uhEF/5qMXKfEKNMdU8PULtmReAp0ObrBP/O23fl667ZgyRUAcMXE6G0U9mmAuC0S
mrS5LszXzjIqRix67IhfLnt7e7sgI9xBF915d/W+ufogVXJKljVN8G7a5qX33Leg
05lfnxItqs1fpUIoCXA5XL9N/5dy7oZ8JKF8L7XW8cElKwRK1/6dy2N/g0QEUGR0
/dSoUqXV6yPI7tQO4FtEVwsJ90b8lbG7lTzgo6bQyM/w8L0h/FBnz6vs4ZkcJoxj
KhGMRexGDugsqbUWZCy97QTZvk1N7LNH7lNkasGqd4Y8/XVzh06OBO5N5EKmDfCY
PgOVS0VI+l+t/AFEoGepsSl6pYYFqLgqFNEsAuNYIjK1IJl49FrYxDR9G27tkVnf
+pXePyU8u8hFYOAxzKfsgCt3LChAdEtxVA8zruf4ZT1d/GYIX44Srt2SiWoJgzQF
wVy4pHPfQAVbdxU0B7RSCYb8GshDpZStVt84c1i6ZDLEgcXaET4PqGjpE2yaU1r2
7wVywa3S88ol+dw9+i2G0xFdk4es2s0m33gT1YkAlGAavGR7NBFJqfoSot4Qgk+T
uYPvczLJprZMchaLl4aKMqXP/Iw+LnP25x/XNdPjw1mWisiXFKvujXYlj019xurV
2qx1DFZ+IfdFiamrfWZCNS1DX0OZYGrxlIWnoRkLUhYHO+j9vHO2Xjl/eZ2h5R6g
3dMHy9pZCfYFQkCU70COFUaWbJgX3NcEbRcrBt0IRqdQ+mwn6ZPEC7Zvwe82rLmu
6I4INPthAlwBSmm2D3m+pn6nWVoF1c+Ub0ezcwaITf6/SB2uLEOm89M6AISlouyc
Mu8NxIGMmtQacduccofz0JiqOrQw/6b8cSx8w074YpAxIhvlt2iWUXm4X/d/wlSY
yQqHeonRdf1w+IflnMVrBFj08KnLs8R9g/QGTBb2a7DeMe2zWhP7F1CJqaWixsZk
QfgOAOuy+l6o/5lz2/HhOJ41hvlerJXUxOPZI9La2CrOLtncaFvplEl2Hm0TREJp
yv/+TXvwcqyHnFerznYVC6zSyToEzvmwyhVa2qlRQgINZqNG5eNywTpJ48wsPe4Y
Ar5VSoybCk4iqgYxqXqawg333U+kIuganq3ntxJydZBMwlbF4NwwWcmR+6GqXNIu
5smvKWjKav8AitznBzfM+ttV1ATvVusOLTRgVO9UWwrW7oTLw4BvmBeDXPv3ESGT
wC+L7cw4C4hhTFm0WJd4+4xJJjiv8nSPOSmFR2udR07VvHVemF67Zv1BJX0BQyfD
FHLDg9z2+Jx8GXL2bOhqtA+iP1sAxvvIVqO+59a8E3yZz+1PpudcWnTuTnSxlrWx
BnRyxK32ZzbJsNMwO/mf6nJttjTUBl+n7fhtDYz64nFbmUyR6MNsS1yoceXjLGEP
Jdm+mkmLs/UAXa0Xwr/On/aus2u5BJnC3LzEYvu95xitPxG7Sz5XbdglZsh6KuBT
o7Sp54jZTb65xlFBviD4JnuhGNGwYuGxF5M8Gtnh0mEP+qGdf1tbhjAjW833y5PJ
lsq7+KmCpBu/0lWs26BpHtXC4HYE2umTqSDlMlCXNnSohwQAjevzgf4OwfdkZm4M
BAyG1Hk+3r6w/ed122DCGcbNHTwwRDatqlLd43PYXjpf85/EAKPPFxejTeJ1Xoga
hm8gQ3oGw/aFZtXbzLW/wjLCWjiE5gdoio9txM2ev4kkxTYbX12eLV6+Vd8vJkX6
j8fk2RbLC5lMhekKclwyZ+Eg8DzoqPqnaf5B/Zbv2YQmXAqgBgTfNNMRV1DuJ/wc
Yrz59hE0sIpE0+EO9w892gnDO5cRB7WkEQokupptDidHnyhvG3M+ZSG+aSULcH03
H3SzhPwaSEoxVF8gmciMsFQ4REDeeFAYzPG3Pa6Qfkz7BsZSPelzgPzuUy2v6KwB
iuyBUcEU+BVo/M4DxPY2u94CUkbOe5v6DjvPXJF8/iPUhEt9osF5FGez1Dw/NGRl
9FlPgBcmd6Fxc/NGyBf44ajcundBPznr7pq2k1rsFJ+YwuqdzREn2Uzmg+FJB1oW
cYDA4NIkgCBNaKAy4uc/NMRELF0LFvEJyfhjPda+6c9evKnpWCVovxi/mputQdAH
PokvrRv56muu4QMH24PzfzTtYqRC+i5n30JfVy76yj9bAzPgwOnppCcscwAq9r7d
k/xSgzGAOcJyxmEdXMntTmhK2AkZ0hJlBOvVRTIawTUY4/4bAtPCw+rcFv0Cs5dv
EgccugPNMyAtN2OocW461azmpQfeR5V84S2ODMwVFlPpl1aNQyhRv85mrvCH3ilq
CIGJjdbqMPwk6yhgb0YIYEiDhvGvt/zGkgheC89xnWCoEYmIG23v5uYvSeRD3fb0
vo8Ob/AIUjIL6L+SOX2Dp9ei7DLadG1F5uoazB8QcOLzxlQvSH2CNNXsItdGm5NB
AzLw6D9bKMV50m6Cl7TdNuWOdYb/kSntRgTPr6kIYbUrB8tGSExeMpZTZlWI4MrB
KEHPA+8WJKUIvdLdxgpnsThSQLUBSyql3hbs1uIgsZpE5leiMgfEpWkqvXj/ydsZ
Y6wFocrsVI/vd3UFU8nyrfTbAU+MG9mTzJ+Vr46VcqohF+gPN7FN5s4C8J/NQPqo
Z1IUrhGaEMKmtasLm7tkPUs2ZIcf/CuAKvgkiQSjZrqKoShM1ZjImRnmfP6Xj44/
uVB0jmODh8gNlqxygGSatBEnOdNFAI1HNnC1oLUR0+FPgEISn8SXu1dDfgUUtq/h
4OcXBGem9vk/Ui5Pw8TmXgptuWvWC76kpxVjh9weZcuK/VXtr7VAdlzGI9FSUIzc
eh3olXw8+yYAXZKfB5JO3+i90PRvuPN13EBS396oQ4XMErydEOOn92OIJ5lkruFu
n/UTNEisUUjz9xjFM63N7plRCH7vKdx664piISyHeW/LJ3bh2esdcbr+sH8r0z7S
QtbsaKP1uD+GPay1Oq9ODcjSCwycPMT3mXyqY4fpHXG7rLSxAlsWWPrlqkUhBC1Q
UhSKv/l5yYqw7IiDOg4H7yUNQ1hMNDl3CEw5v1g1slQeKxlTV9aVfb9MJGTb5gac
UMhEBLSZ321pLZ3zVLqQX9HbUwtomh1O7c5V3ktlYYDmCrsGnXD4+YApeiUhI59a
txYmrtG5M7qQky/XSbIR4nUYS4al1VTHSXBQ/WuEx2iRhjNYOjFeslHNA9FvrUP2
MHQkK7vXA/HHuju53EzR8llyo1KLhqv1yYaUSMCorScKhL93W94Ga5XCJEnawD21
h5fmylTnVPPjRwCcJSWHAY+Sta8Fw25uyMPRDLPvdxw9q9DpDcaZ0W4BlZNIyiTm
kohYJ8SmEf8CiO0elm0yAVfUYoLQ4S3VK06+kW+af9MIXzI0lue901494p+Joeyt
4WwywuYeSyCKKk4xgmw5lbgsbLQADv66R0/gfKO9uiTf6cb0FNbQCV/kvU6DdelO
PB1NkHxaC3ebyof6Lz8obm5C69m28A7BQYR1YK7GxeJx2n21JR3qU4AxEbVe+NXY
sfeJ/VdgUwixNk4p7QUkRHk5m/ouHyVSEK5Dppczb2EVbfU5OI6ZSZXxmwKpf4yj
`protect END_PROTECTED