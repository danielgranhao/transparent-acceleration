-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
KQsq2yU5wZgHz5O0j/dbC6jjEzXG8HidaBKU24Guw2+SjdjjrlaCT7/sfK3krS2x
RFX9/4u+PbyqRj+UkZOexugas9DFjiNhXhVkV0RKROYOaY2+VNZR/PJlh7xaSeRK
z4u10XUkkrLzsD9nBZxKr8ZFcLXjp/fepRYKmCazaiIdsDcSwL6Q6w==
--pragma protect end_key_block
--pragma protect digest_block
R/Blb/jazeiHJcHQNyxaykP6L/c=
--pragma protect end_digest_block
--pragma protect data_block
prgD2VrbVoq2fYI1H4W1BDK2wQdY2wd8Upd+lxBuRAgmLfHs+/2CVKa7QQrF8HpW
Nj5ryLmwCZQt5NnxPDok9d3JGPhIjCWxL6gArux4geeJ34E9yXwIN26JGgtqZO47
b4zg5xknCY9YHCEhJ6NriTPP1TkAo6TDHIwZmjTs4iDUBNkbhqtiHqhLg5tl9wpk
ZPMM0Q23TePiVs6334JtFdiliLEzXJsquJ/6DDu9UJIgpp0UobcWTS1FnUV4Bum+
qAtGx/K9oEfr4izvSQrn5QTVLy4K/E9eQai9Vq9hEVxhxvQykz8VkOrMFeeWmuvW
XaOburv4U3pIS1fO978FagsU/c7e60mUnExhkozwn3vVwur7ACjrqYdSJZHfeD69
lHMvEfzrZm5Vv3od9T+fqUp2jsf3fR3RZfdm7Z4LK5MUXLUqx/HKOj5OZMs8aWqg
Jh8tMRBCO/gucY5H6sse7K+29qGWBIt3izDmeuJm4hO1JwZBnGLNpqBZe9Xj9Wt/
I9hAvUrM2l2PTlQyoI2JgXbwvku8EXuVucuCpYI5GRFqgeMRw17hvhxgd9k8sR+k
SND0t6jE8gwrQHKFLFzeJ/cL742e5h4XfYqptivX+9OB7CX+smJgfbaZX4rBjnXn
EFKSMwLtuxrWVH5NbP1TYEGil8MjHEGYZTJcuYDfSB45cWkCYdHEjEREvAx47iuu
yQxlPMcZl2NiZs8DOM5Xe+GXXeBSQX+TYKDCrsanlJ5Jz6xi6WVIJMi8h5ZWn//z
z+y+aBYNILKC9hpE9NTDriBLp3vdK8ngk0oZw1gFSf0fhTYnewK4U9dbJSSuVEfv
Y34m045bE8e0nRemZ/oXSrx60vofFph5GcvjOgUvULsAV/JujfJb8sT3zJtkyYvF
HuH9TP4kJq85G7KaHn4q77NGxnSztDAiiot8+XRN0Rk7uz8s0hgAeh0BTUiZdU93
Aq/vbS7j9uPKlbmWdZxZhF7cPPyNJC3tSuz6ug42/JdFXwADb3PhjADd8ti2o2Hq
s6Ti51fQqBsQqsuBfccx//xeUX+5WNg7kSkBzhA/jvPVXv+Ovjt6uFvWOEdmR22u
6zXLxpKojDqaKEqrSUJqquZyuX4NXwYwcKl2pVCELdpctRCWg6WQ57EWXUoHVzo9
P6T37OEtaiWwthcMb3wZTStSe/TJnbIw7CsvV35JUKmTMbYc9a6ocD1CRGtoafbr
I1K7Qr9jPYvL2CiKWbCMRg3oFekPrEC/Uk1OPGf+55nYocYqj6vER6IVtZoBJGje
syUjkVCWp/Ol9D9szEOXLY0bKkl/lWoeZz9c2OtXRzgGrkRFbiBWq9lpDbuGDSHS
Bx0RvK0vqHh991RI0rxnkfM1pgYQzOnfWhuG0LtN1TwLOZGWkYa0L5bBoOPl3Bfj
GLE78y4KNvo3f3Mss6TsG4xQgOKESVoIibxDHSgptu/jAT51S3qcQIfKwAt0XufS
4zrpidLdZh1LUqEaTldtjNX/xMnXWH5sphUtEjuaFavN/g9JBt/HMqiRG0kVpi5H
WEZH6vpqYQMrjaWqZfzG7y5dnYBc44hYyk67fqXx5AVEkzOSI44AIq2JTyd7ZTTE
pzWJGs9wXJMz/mavLMQ/Ox+zk7rOW5OeUwOpY9D8FWxX0UFo6oyuOtTbC3DIjs2M
+oUUOVQ4SL6JHKz7DaRTU0ihJvSjpDIu+USqu0E55He3LPEaYUVq0F5QB2VS1K0t
MKdu7pqPhzk6pCD/Ud6af+pg66vwEDScamFfVNz/mVCzTBkhfc6Ek8k5OB2Z543a
qJiAZB78Nf7y1ILcLaIxvC8phhAcedcbB5vCn0gFecjZ/f+6eRjqbo6c24KYZ1NQ
UCxi4n33nbd2mUJsUvJKaXuR5WYFmcSmxrT7hxKIbJv/HlmzF2P4/nPLQ7S1REMr
AV6i50fzncVLpYMgm+6VceJ7/AHLYe22+F8FxjZniRpLHjHniCxHzUpwJEW570KO
D59tijr3nfKJE53+L8pVRUDA1Imlh5c1QdJLLI3Uz50PCEAEH9iIMc1kMaiEGinx
7YzfkzoTclgj4xxHXSnx5XSFcHOAnczl3xZUp8Cs7h8ME4w9xqgrKZSAk8hgidjo
xj82e2syyoTp/zTiQgi4fpvJd6IxJR0FqQD6WXVW9wO7fTvcWvUB+oCs4LeEXxd4
+5fSxTquiaYiISNyNL2z6+rIb4mb9HNmUV/9G+KfucXPdTb+MpbrqW3VCjHQujqv
b+7P581bVA+daMUotjzbdq4Msuf8yj4uQtC/iCd54FMWFqn5KvWjWENrjnha69A6
amBSukNjzvcB3zW+4+XiADzLfbd8m7t15aAQKRWJUKPsh3MYKb5wxxNlicedpXpJ
XHrmSe/hkUauU4Cv5qEshXrPoy6rDemES4jWAO2Fqq2M8pimXR/Lq/vrJGomkAPg
2MrRnRl+6FRAoK6VG5gYb2Co2WsVrzyETxDuQtOEws+7EO7rEuWA1l8kl1Vpozx8
LvQWhv2upuY0jZXBdLdbNHvPFeFpvPMDcMdF8uI4xTsQEhdQohG5BG3Nk+Yhpz56
gxL57iTVu9AJcKLeuiZaqnnXkxyCIu6GWd2jpLwDPWCjdGRfNnH3tQTyDRXmNOaz
DEaRjbtf4H2vUS8VQRrXXSRLPTgsJK543KlJcBZTzm4HxS++b+xFWjp4UVSLJwIP
t0pFf2LZJM7tLsdYd5izRZshH3KAOcxP8eoKsA5q4ImZy/fFQkQmzTYd3bsquG/s
JTxK4gjp0eeqKB8aD4QClCXiEYWvEkzpRB46TuqxmjJIzgyTLJEtuFWqfObnw7HP
5+AZEp7DEI1rj/DM6qkoQpuMlYPSGVnI92D9bymI50AJaefyeY/9l5cgi2d+uPUC
f7aiqlpBsqXxl6eirtm5II82iebhmciRN+71RFHL3yl6yp7ZWU5FKJB/Fd/0BATI
1mGi2Uw/esmhjOzizhSEOmV+mpmonxm5lsOAPHjGxKQW03uBjvsJQhNbq3sp52lp
siOHfIMI/lgCded1S3hNAgEW3FbtIHabVs4GVTu1KRsjbeidZnuwMCnvfOy9IMt9
uRGBTZGF0lcR6IpX0wyhbZnQ5Y+YRjHABf9V5DJdFe5Jyo30sR0sXT5WfLQxJLPx
n3GoAMEncvlIiO53XepmZcqcFEe3AtHVUFigJeu+3w4Z/vU/NJ4NllK5o+5I82w6
ZPdwe2zVBvRN4y9U3hFCTl+a6zqLiKVvFO1/nxapNt/+CAJg/PPI0jYLrzJuzkzm
j1sIUqMeG8QuKKzcilmcNOnK7R7CR8QFFnmBFTrbJpH7D9acvIB/97GPaqsV3cHJ
Ry6VHsrA7voH1HdR65Kg3cVAHG6RAahkjbywIMFeblPsGjy+OaZNN1S0NYfqsnk0
onPfUblF/FEpwHS1mJF4MlZY1723p/YesM0RwVUsPXTlCtxHgIngfLgbdx0lc3F1
sskeEdxsnKG0vYmM8caGTt31GwITOmrhg2Gjfxk9JxB6AK1qvTBaacqXQ5N78Hzd
Oh2bUThoBZlkFCEVYktiimJMIRkXetH5pPmC5+rsd/x5x8iG4vTvyk7ssSbIxxkl
IsRelfT90hnlB09V77sb5nISccRfzsE8hgfuid7QD2ZpJqCY0utROlMbZ5wNiXKS
W/zL8Ltzqp5Of3dkaGqWgngUgLSzzuPX1AP+iq9gQ1G0QjjzmdzF3cRUK0DvNddv
b8ojCcgdQtcdsOutMQa5UIucR2ymFP1omSNBYjpiSx9Sm5EK1EodKG/U9BQHE3Gb
q7Qv0RRsSEbH3H0zR57n/AmW0TbSdHgPtbO/N1reLTzn6DS2TfudnxuhTHWWxmOb
uYxWp6OqgzT3EWsN2kS0K4y+T61sGSvvUexPxjabFtByNTwscB6FVuUfpUlkXyr1
c0oPLXhBIWHuTRqJsu14FayP2ZM362ytztenYW6CWU9RMOjuW8NWZ9ILEwFU9fJt
wsYoS6didXYmuVCJgPIKRoLIpeJI30S07AT1ypGQD3Xrytk7ndE7Kh7bXaXTiQMa
IeRP1ldZDK5wXK1ANOXhxS0V/FdlSE1gGO46s5smP6p2fmMb3eyHBz7kNndSAM0a
U5tgc5ZvrXP05ZWFoR95h5On2PlMfwbRUCGAu+0iKObTiLLG4px0g9hrNiIWwYBf
szjvPLav7DHijyheNzqZJn2ZOjUR8gB+OufBxPJmjPQABwucwxFDz6NWm6KDozG9
kijPGNmwzJP/0OEH/jeyt0Apmz6RX0ICDAACWz5xnN/oz2SdRWVAPew2jl10cJLx
1ciMF6BFXPUjnFcSklnM4oEDDC54w8CVLop7bsWngapiH8/fMSiwUVH87qWgrxIO
y34N2XYl5FP3o9cRYIox8ypdjsIs94znLSWiv5QGkBqeke/ajYx9gSQHGYY7q1Mu
ELs/eDgtRoDPNRAP6CJ8X0M+TwnyvkIZooqBer1OC2GunUwSQwBgxon7TCHSw/al
GR8WDjhhVrTegirP91jb8qx2bs0TgX26c0nW5XnnfAS3hbzysDcJIwxnxwa5350k
kvBaP/w5M/sJmAtRvqdh+AZppcZsTvbw9IIYF39KBo//UhqOf8eSnsqGCZ2D+9EF
rOVr5QZOFjSdC41O8tNF8ERn/SJCde5dTYylMJ8PRyHuEDbMDbUDIhVQf08oyAy/
AQ1NdDfb7g3W00+CR1uYmD+dUnSpdqS/HNc6TzoaLof80O0vU7ywL0z7ZbKOmJ3z
wpx8aw7BOk5qVrSnVB/7UrtADk1/C1l4EUJavG/ddQPT5J0gZG+xmdKImjBrgVw/
1wIfkn5VxQrQLRJ8CZpLzbA10nUEkQWL822yC1KfF5EoGTQa+tUvJeBAb/AtJqZx
WpbTRmQwrfXz5qyLulsGpKcOth2M5dCc2iwSFADE1N7eXPhSMg9TKaQPqaveBJbx
f+SpzXch9/nknjFfkEIj/lkcHQqi1d3pFUz13VO2f0xuxbZKGhBLfp+fZXkY5NSA
APdVlOdgF8SRa8B1G0O1U1gNY0jjSHhM3Aac4iMlGCPuPf9xwWPz13HEWfgKTkcY
D4pAmvClyxPm2+k5oAgkc9/dn1MFER9L5K0RA2Vg/4n76uyzzux7aKhbMW39wyCt
WPPzFNOPQgyNFwSum0qvIYcYntm2V/oPkU3h0r+YyP0iL2p3qhLEargG+Vh1+xsU
4FFRDzmCyUUHwXBNU8juBoOm6Bzu3Sumwhly7BM2RttXOfaYOzUwEOiC1x9j4kCY
Vr1dmrSk2G7YqHBQVz3H4PtaEqgr9cWSKFWLeu8W/keVO6c65TjCo6wO4Hw+ve+R
MiNnk8xBayKHpiv+GkVjcb3nU03VJiWKThnJUGmrBb2zi6MfBFr9gokXg1nRYX9i
cHVzlUQ10MZIEM0OqKWng97OLyuvy85oEDxM7904vzZN5BHDyAMv8hpcUcLuyPWD
diqNjMa/bELz8vX7PABJIrkzHIY+9SsAtRKismY83UjEZgYToP/E+TW8SnJMIvZj
+8QeczyzYhJ5HOaK5Xcle4ll4J6LfgsqvlCBOlnUlfQ+O5Fm0IrJwCciZfgwDeUp
kUfiUrBxm0DTWk7mxoGBB0OtWBOd2moFCBp0nZPjXb9YlBeDmsDPwxNmMffcj8s8
dm2AV9WhbOHCatfJqzK6CByDRUbpsWu++pA4rXBBoiS2KAC3zwGKm6M3xaSSnENw
vOvFzro5e2+lWUh47T85oBvVFH7I1M1GabfovY9WvVfk4szsj4sEU9t4xJzZvaG/
vzd6wl7WbnVkctooOPHdVQRb9DdNm1i/Ps9T7+bplnVK93rCH2V8jdG7+ltdMky4
Yv0z77z+8+uoKnJQc/MzNT/jmwzxkoNsJcdQtH7KLY7AZqCUMJ7j2d5YJ87dvJO5
r4cG3jPas/O2DsVEX0jIWPTFJbVaSkgnGUErCZKEOZ09zM4ZIBft9Y717NGEmamt
/3YCPig+KeV+4k7TxYzsgB92Te8M559As+0IiKYLLGBFiBXMvxcvnbjziL5ybaf2
HKe7mQLiWLhpaiBUVl5Fk97JGcJ6tgrtyQFXLk/9LdYt484e+L4XdCLs+dDKP7gb
D87evnJRehgNDTKBwM46wItfH7KFnEFWPnN1mtzrSSQ7nyFwsaS4mbHNtDxai6qi
Zmg1FnBrvSlmzqiFxocFBft/brrhWtyDcIj6CE+fm391VyY5RG67mNDwnfBj7T9Y
9DCphNcOyY5eF0q7grKPr8ljjIYUoKHXFIMXGbedaGUvbWjvn/VEAYFlyl6W9lH/
w6JkZ9p5gJot0BpXTTM/RxRahy80xMdvSKsoL1d9QQrhDtVNVr3aWGjktb5KuN9F
6jQQ7CSFY4/xj0+86feHsNSstSXaGsQPwbd1YA+/oHw5YKARLmWcKutqUB/haz/J
kLD//wZkMHD6qZnn3LAK9rWD3hXqxM5DQ0PYFcP7qpWzLHFdjM8UtNEUc38Omff+
Al5SZKqfBV0Sw4Yzv8EfjPRmFfjGFU9TnIAKIseaz34TDvudzIvz9hK8L0UlPNWa
qjDJhWJJxXqZ1RXysKYpodwqgL9qJ0gYMdur8AcVU8/FQAwPLghV+NuNYJh1Tzat
ejhBPDYIiLrzLxjMzgpMw0fLB+a2Ob3t9iz3QLpWY/9AOxc+1PMJ+DE4GE/jrp+J
01DJrThgeBQrRibW1CUOCtVH8SP+heoBBnv12ZRGSmZyw7KjG3c167/kz2zm3hNX
I7Ug6YLWpAss8r+tdJfMbGQT0jSMF38ersG3P3VxWUgJkaio5oF3BOWbAgNzoWZJ
DLdjQHYB99srhWtETLEU2yiPxNe1aO5nN24/pksdVXFLGJOj2fcCGb6A+Pxr6yFj
t0tIPY3xzZhogWNEw0MUfyi/h9MuQkJk8G5kyunmAI1WiTn0Wv+HOuIS1MvDZq23
5gNb/IL5NEJDFKrof92cZ1/w3HC8XCxbTQLbF8HNrtjrsUX3fcYejGFJaS8wK6KF
x9aTlsjp9D5oZkAC4gN2ifxF9kgGLCC8nO5nqJy6wXX+ADaG3J2kIFFGSiBjJrI9
94KV0nLs35Bmt+dbVwdjw5NpJnK6Odu9OVau5Ufj0LnHHNz7rVAhEoi7D1SMHPXA
zhFnlH1yDimshOImbZu1qE72mHzx3SKM/kjtFQV3gPK/1zPDCiqz9cl8nDvVhkEW
dvfV+DONWkfS1EIdcR8yiTg/sM77Np53ARQKpGJQLEkwEkfQ2T54j/4EaGt315LZ
4ZfvO6Ra79NeKjM5Qf/XN/jTU3XFj5nyXga7qDDUGBU7GzmBP4Gg4vk/jNxIUuJO
UH6uJ+Vj9Elx/Xs493PrE+O2TRkmRsVjoPRROYVlEgcPxPnBCGilUl/6Y6PfsLOI
+XTvmDB2ECXNoEQz1VPGMhQU2IvTY41uZ68yT7iXAbj0T9G+Qwq7XIYYbcrCN5FE
tG6nUmSstoCIciBXxf9LVfmBnAw7SmYfz8IKDgFc7x5VWq0EJB2zz2i6qQuNKwx4
INFSCW19KlTHIKwvTt98bVmLEr/S5kk4gzLpwxYrMyXdGngn0aHOJ+wSpRz7y9Jt
779SxJ3Wpe880hhwAB7A8U4D5FzwgCXK3YGmKBnEUvZfWmog3pmTuFG027+35ec3
n69y2OoxcaQzLubgWsPes1yQk3UKtjgIr455NtCBAlVDNGptUdFAjxBuTsmjOXTB
Nnv7dcKaAmwkytj5PWz9ErZ74okwbQStHKTuag2YUmxOhZxQQxkYsCK3Sv6yksJj
rEfixlmDeHqpdiRpE1pHGendqaiUH60+O4wpq8P6Fxekb6qTH04vQjVLI29JdN4+
0CqKGOhfH6pBLpxQ541QofyEy6YIxway/H9GgnPjYWM+MVcxa0FNdFqMfUKX07rJ
4Cf1Ihc6vJAwrQldEVpm9hvM22kDbbeAAnzm+hsg4vkE8Q0C6ZgrWQAclRMGaMpH
Sq34h4KzT8SxsRY4IWPAZgMLUqZtoqTPFcc/ybgzmC5gEOBCjE0N5cMgLWJ6B3yZ
spuU0t4khTseo+SqvP36qZecWozhWQNfqmvRysKPjfUy6OLurD+lZlzfaL6Zlld4
/sZX0c4ouxz6yG1MfxAmYy/sUV3B63WIYXWWUNoU62BvgFTocQI68I2l3aU7K63F
Jhg3oYHIcu8CvQ7Oo4FEpk0qhPEanVAdcl5HcyTCVpCnqYFzjZodb/Eac6lQIi8C
u2z9FuJ5MPc2z5iQQ95zCtmGlAyxDvUpuIkX+xtkC5+DZABUNH/0JRxDDpMivMoD
yHtNYv+XARIEJElyL7R+rcYb5DVRyK9WY1w+JJ7hoRrSStfE0Zdu+QLVP6tSFlDV
L2Z8FanN0yLLATNu/3vafRhXzJQC77vTdC+Exg3NUHC4FVirnGUwzH3vcyuBYhwg
YPtvaDSV2+gVkD3CrBRwDPVpFkMXSHm0ys44kf3TdZaCFqwygIgtlPbwF/xp9Teq
c1Sr32pFX3tPphUHDyc5kDPQqq0eTleOxfHlwRgBGE07ivUZSEJ4TLf5OAQyIBpC
Z35XEy31obbydkQM18LkxAAhRKu+lOjfHeDPNsFGbNK6son2ER2TcAyLLPDihzs/
fvGHnf2QH7uuOmCOu3GPd1mJ3VrFlmBR4PHqvfHYy3U1q6WE0qOklm0mjB6k+Vlg
dEdXoQp4OLIxEGypRMTntxAvPQE3eyrhzpNSU1QAxE1sqdXAKcyImHcbZMb+liVw
7vCROHakx+BsWP1MSqHeGGMojQMOdQUNB3iK76iVF3RMnM7LkcFuwqKlXPhO/2cY
3eIYdfpbHUh0ZL2fVfvMIg6rlYFySkJDfkctUmT+VGwPqQia+NHkRlCd82+pG3qU
PN1pzuqTpeb+Kc93ejLVaayE29ZngK6WlBKGE7yHrk2PlfnqbhVaoz2/7ARnlAnK
1e6+P+E3qq+78n52DEJ/2AGwUv2TDVqIKC3EiMlgekro8aqU0XpRWB7vSVF95wxo
GNlvepmHcMNBefba/HOcIt4fnhvWrcSG/PXMzSHtSMeTS6uv4p0f3ScAkSJ2KB6m
6W+Yh99orjjwxelCT5HfRuUtzeELHHNIRY19pcbS6ZbEkk58cq59kya9JMBpUcxx
8akjuGPqHK5EDSKOjW97MgDa4Coyat+USBGWhiBM6AGscJTv+RWw1CRuFNYhxF31
xqG4QmEVOyQDuT6127kPWeCQH7Qo6biKWXen/7Gce7YyV+7S2noR+tg25HgQp2ps
BT6soJN+M0KU9SjYrrar15EAwxoWTAGJce9vkqJdtCS/Zmz+/gwa/k6yld1E4jLj
abKW96rjgYDewJo9YN6cIrE0rR9WsQqpEwEbUvWXVgwc1MUEzZayGhAK78bU/2zT
lIHxZln83CH7YK01EYepTpQJ3j7UWVcLvmyKp69b0E1tpadEuAj/p/ERHML8wGhe
DA/S6Yhz57rBOnydrNKWCf3Rjr07tfdD7h+41r9qXEzrYLjaU3wavAToz/2CP0T3
xA73PUgzmpKeqZDVNNakrxgEPzd6aUjYzh6oRjJ8bdmUPl0qrXwA/H3aQFOYIv+h
CmOwGx5s5cauja05VdVFXAz4odgzWQ5hvFHNjGrG0w6E8WDggXeON/hZ/Ac/D+BD
+GzKxEK4mBow9/wK6lcz+hYEe15tQqImkSCu/f+8I82OFkV9O7+APWJzaVybaSeq
bb4iNGK3weQyANOMPOZ7uSExWsMj1/KgWjLFBFRYuphaLgZ0hd9pJ6MQXHbx8Djg
zihcOgHUVLKmmhX6/KeOQRii90WThgvpHQ9ffXOJONhkUfPxWvi999Gc42pviad+
Duo895m5TbXYj1HMuylUxH3ZXunQZC02E6CAp9640dI9XHy2XorURrIvlzcZjtdT
AXOKKP/yjaFzkzlsw1NKa/4dG/ydouRthsr902yjAFgwjeyL5uDrIWE8So60MgUH
t2MzW4Zxc7X40MKaXkbXy5/2OE1LyjZUaMWRxmcU610sTFOXuLH7ckufS+GG1Oj/
XmSBjzoqtImenVJA0lDgpYwhio2nVNKPeRUWP0H0F6igBRgMxH3m4EFKadPLOMXs
gvncUyuv261i89xNeEbDH87o0TAetNOMkAQqy1lZVUtqiDXwyvp2O5EAM7IMbJ8e
VstTQr1tbQtzKEFv72nlpe6tuZWhKKf3zF9Se4Lr9Xgwocnuqn+13kU1HZpn35l1
mDMcn8XTS4pcYqD9yDGthASm+9DGtUsPsvkPV3lfEz52RV4NxJcDZzgdcPL8GZST
RMmc0JMrbUct0csZs+odqi7QX35NpcnWQ5QiQpwR4HV8lS8Y4o2/RxwEoqfp4ar8
RGsHQZYDbdXYE7J0YOCEPpG803pWwNhTv3mlULJOoXo7IvWT4z0/x89sKvf2641k
WicSl3GQUkvUXdU36li102bYdeIC2BsQG70gYNfnGrzSSFfRMNmNkGk92uclLA/5
XNM+58q6SxKi39UiwAVfpOnWfcU6DoSfyaHS10H0rZRAPZtMJky667+YDg8GlRoB
JaiI1KWOaUh4t9axQ3oHzkW+cu8hg6hljJ3BN5o1BCDiTQplLHxdudIcaFPt7KoN
C6bWp/lDS7dPnqFlLptHtpphDcWrJBTQBuvbzzxMKTG8f1KXhMx32NmplGZZuhVN
hZgqr71l1mesXHNJEfopSpeqrdatyw0dQxYXCLIq2hwUrB8nO8grZob639zxFMMp
hCZxu6miqYP7lPwSOVONIN0oS2jYP4GeDerUdtKVJmpEinxSHU3TX6pm4P6RmClj
QRiB/eDGKRBv2V42yS3B0wpj4/6jEEeDBTAJH2iDkgwq0ImtiRjiw3RE6TGyojRL
Vy88BvRiRcmgWBKQU2YgVGsMzHsMmsTKwbaCkY3TEboaCyndVk4Ws4Pla/KK9Fpy
wGeANIwpS1qHm6ar+uDtqfcC5n2Ez+QQxPZdy98xI/Q4JgmOJyZlu3fK0o3EikTh
w+Xtzt5tqcWK/sxNVRlZCwseGL92Bv1i6jS00Nf60AuP8iYYSdoNuvBKUUGcRx1d
dB8XDRE80cGop8zD891+zsd1ZIY0HBLJ5ylALSwvlrRw0MkgJKMqm3aKItAPllOY
eWJb3jIVBwDdbrXS47znKpwXrFLmq6C18us/AobZkUd/IzVQH8IZ/EP0Qb9Y495N
IR/HNYcSfAB62vQFHrQqyj9hd2oHC3Sv2Ui8KQmO8VIP2yy/FKhZgEzOGWNQFC6w
W86ZgdssJSkb4YhpB0xxanyBNTXKazs+cfvGsUfuzRBfjjFTA5wc/FEuBZJCaOnW
Ty20dQlGsL9K0eo7oT1xkeWEvCgslXjA3fWGyS898otGhco9UjCeQ4/ktKfqbOin
BlgcIfu05wQqeIpSrWI2Dd1AWvAuaw85sNpzGqIBz6Gnpyhwp2jnEG0eptZiDnSk
gPy+i1oj3txf0HXdJ3WG0C9g6rO19tJSSfkQBdcwhkJLzOwWYqWFTAzisRSaT5MP
MmwS0qCahXXzEzVEv0WDuSToU9zMkZfGcLGKzh3flygjVk/dT14N2KArnirDVyS0
rpjJYkQeTEJMgxOVG71sc3e+1IEycq4J9BsJ0hkKvY2EBn39MO7sZMv2KvYGqhNQ
YMB7OIEHIoYZc8vzWg7eO0V1m0LukSRXNPAX/gFOrXfObq7qLoOJSXpLj26pLPun
XFIthLGJCw8tRxl1k3ghcL5rh6dsmBdgVj19mjgHU/nB+f3QZDKu6Rn2QJgRGvcR
wPL1Hc4ysxKLhd1MAkkXKmqe2X/CNfB5fj9kmTWhzQnOub7tKZrnJUzmy8xraiVQ
ExHzQzUrL0wCcGnm9IZifYzTFyAdFyPIGbN+d12fbL5+h5z5ywzcSkT441n3sgGZ
5EnMXtyzVkCZRPXfWh5x4e1xDZ9icksWNNXCLmqSCZjbXiioU8yllH/GA1eALVK6
tht2crwAciKra3iOV2hwHzLVPh90LlLXv9ppyPP3IexvLvR8vvb3+HP+TR5vt/H6
if5M70/H64p/jp0fNsRZ0IIYHHpOVZiQVq1pS6XiLv5OCkLzqVlmDEL6jfNyebEO
ZnMu2Az5UV46C7r29TOWMqn67SyapPT85vw3PIu2Ant3gYXjxxw85lug7Z3aI5xJ
bq9g4gpGIR12T099yhuW/syWFhVG55SnUoLoUWPjqPKbk8TZEjcb8DtXHtYxKRae
nSLYhbX2BCKf2ub6NGdpRW+i9T8ECLqE7QuQPt8UMBf4hER3lOuNTgMvqBk4xRs8
9r7WNH3ZKOSTLWUPj2K5W29Hy/RxjP2R5EnLDP39AU3cjF7GlbkcSR7UFmSzFlLG
tHGgtzG1KiqSjt5Qry79tM2wJnY8FzHAtkzY3lbuDB8Eju5iG7nuEbyTzbetjpom
teBf/X8ulFjgxlbjLCf7EmvsM4TgDjtrXxLvgKZblvkp4OhzCA7QJ3aPeegPgMgo
YTuOpKrMT9HilaNyUxr738IgI7nNcR9LVphjPQosg64Q3NbdU2KQCnCrJeQieMyr
apBv1tGvm8IMqKH/OD7hV/Pa+XwlrYWMmkHtgUl5t8gua3XKyVfoXuyy7qO+JAuR
YXl8Zyca3YGU3lY9Elwxk7N68HG1HO8q2HODnccA2tKj9eIW+hNQ7LRnFdGCtKiT
yX7znx1zhba7s3xxH7l/UGXetQ3cXY81g4lZtqxo/s2jvq09UJydB9WK/y7oIdxQ
Ze3GzXbCROPzlMk8ITrqDiz2PDrCtDG8Z+GaozyQGPDkXsZYWP5ySQZgRP2TFcJw
HFM6yFIH7SrEJvbG6cWU7fKpoCRwljD3jZ/bwhDcG9GEDp05wPvUQO+RWPVCP9s7
LR3wakibVv86iatbG1lamH6nXXfZr4wIrJhMolHhSV9MHtcU2+oXi/awCwzlECJB
E2+C31EeyiOQAdSJ19zDRYNFLtZ4w+XQfoXsHITQ/N3hrwW0Zy528qu/i9Azy4Xm
r3Ivgj26tIxFMztCkNqQoCtGmkI3AEIscmiHbZTc+ZO6fNb3naqQvQ5GSImfkHFh
BOi71QCHKMFxRPuygnjJ5k9H85nzhnKcUNVYh1GKn6Kv9ZcgZHMcsgAIxQ81Peqp
N/UxopxQPumn7U87qMJsjYartcphlkF2KnHCc525yuM6kpXmM8DGczvsIf/scZyc
8QzEcQg8uI8zcpvuwzU8K0RKZLObAJhdOtRlB22cP2v4tP8HnoC7N0+uxocr/HxC
OoWAOSbZFxFQLUGOqZLK6vWeb3M+d9aDgjlIDEGNb2IlD7R/K02YQT4tw9RrtvrG
/jPp0riOVTf5RkIK9Nepi+l5hzs+d2TMOV42tmToaq2BARB2A/eUmilN+qZWQhYO
SAPIBHsZRL2M+O5i5XPBYnRn21RBf7Tweq6HeyVhwWriM9gCJmCqniHJwLRM9ecY
kWOSTwGe0By2jnB3e/Sj+NITB21v8tshIkPdBFgxmuGqG7nz7ePw9venaaL3QU/Q
x1k1lBatS21FZejCF3uVXRgWddPTwhhHCgnXnxpztOt2WoMV21Fh180blJBqKfrN
Dv16wKX7Lto9kkilMPBQyi9URLzWyJIq7ZzGnAeAbfj1Dcv6Um2SqAPxcpa90wGN
ZGPiKVASDHYGQfP/aOh35QGepEqSx+XB1BDTiTEG2tkw1IWmXEhh8oHl1ekOp5wD
JU4GAjnuabT/fFMbccYsKt0Z/MVgKTJ9J/96/f9uE08cn9haOFpS3Sq8urpHaxuu
ayqgJipw41ZYImQOIInnliaXZMzsiowpNF9p27j7Ptpw26Ihw8/ycHB2O0/rz9/F
KlYkNEYXeNnkV7y9f3OWCSbjQOJTAsP2X23/0qEvbtzY/7swWrA+qZzSls4C9USS
lK76OhTM8BP4MmHpdkkVU46OcfzEnKIQ4yy/M25jOetczTBKlFR+LgjpNRERhDbs
6HGN4xx5lRBgxv3f+C4PK0mqvt4nb4WD4YQF0FeUCauzghNY8EgdI4ITJnhS3owu
7uVkuJa63iC9jeoVKPQfU5SHw9X6OH2PuIarW09G/P1crFUzHLQTNKX75F3UMk66
u2pEVEkv0/fkYBq2RGZxuhCGd2RBvRSgfAQygMD4mQZrv6EHKls5DFVUSJvldLF5
hLEVWrT9nnYWbZ4oKc/UsfT2HA0VsL3WYtNpfhQ8+0ND3Uj8RQ0QxeVwN54oAyhx
4o/tzTAgvQstw7H24HU18wv7XPvEPKFK9uNYghErp21zj/HNR5wuAGdVwVfJ7OiO
mZ77z0klS2vGyLIpKA7n93fKjDWIs9pfs13uGanY3xVuu1uMHGIwafF1M495LfCU
ES57US8Ucrigf93GjR+TyMidA9LyIEHcFQ6qMVNdJpUBQTN9zcSAoWYmURXyypcS
WgP8Hsoas1/5XEOerAG1bmnTa9ui5Ik+iypy0Us2al9KJqw92EZZpF+oAp+WRotJ
GSHEDFKihrVUy+SVrV/6zoWkzldFnppubFCRscCoCeTNFztQiDSXmpuO6m5W4cCR
s2UOBGadDhB7L4ZlKYJhxNPe7N2kyFlyZCAIm42fqNGyGBxSZtcVVAIuiK4H/YKo
UnHzKxWk+R/QmtdXkX3UeV1BZPQIMtHHotRTPu/m55hBI4j+2lOAA0QbIqMYasQr
fKnCG+Nwc2/QnOyP8IHqZohKEJI/5k1HycPlqUS2aufeCpTkdwPwKbA+RaLn+Pao
3riGZ0AjHSM/VKvZ5zhJpoxzikfMBUzkQHT/akIWvIHlmc0/jzB2KBtLpWOI7NSN
/m3xLcir+10uGjgEoeVz7Js+Tr0a4YR0r+SxQfbLkZfZUTRkenXdEs0ITDrG3d5A
THhhHzqU3Rl2j09aIUTq6DAIXBbW0BDMci5QhjyjPARfQWwAS7c5MYCRnZIG0VFb
8RH/XaPiDL/mUAGyeWkrdbydMrjlotX77Gbd2M5Ox9vlxd/mC/21qD/BRUgSlsVZ
4GdN9vu/w2ur9u2ucU3MJkAxB8WEoMLtw3EkhnSkafF44rYwsiN+jFyrH/QBg2Yh
cX2aNtMh+0bseZq4L4QsFpLpt9o8Aqbj9KR5LrNhLcxmONXwy0zXd80fvKnOCdVq
apXs9b+Z9KJbdQNOcnTuyxtBkEW+SP3CBlCXaFy0VElHpb/ooVsIpcVLNCgUl19B
L4jBBhelRMX33AFYLrdDp+/pj1BCJz7hJ3ycXLj7RYdZpvyL2X07M4RNzBaiqcpj
VrIP7d6PAKcsj26ae23YXUOEqB9MXUwtpi/C2RsT+PQh8vGoQekZSTh4dfd4ognM
ma7XL90dyp9q3bql913YA7M47txGxGklNlYgxZlYXxKuPo9EeyFKMgh6F9qOApGd
x+pRD1Tr9OwdKNunwYgre465/jrOJQ5BZVZgbPSHPW1ty455Sf8fFXsl/5GwTi7p
4ujRy/02Hpq+rfe09IaQ3ORo1a/d+pXo1e2tl/wZsHSArBA6lzhAxhjQpqyfMEDz
4PwfMZidzRlybrEQ94MmkacnUvKVkbvCslI6nyp0DP5pZzAAghcnpemMgtHpGAME
/FyttoBUqtSl+QNR3oCqLnr92xPRr0rqB2PAQigncx5ToYaCZUjpPIxGIV1U/29M
nylkK4hKJLg9BRPNPXOeWo9eNYB7Dmwwonz3+IXljxzP6hj4sqhJHDsD9oq53Pvg
yvkr706ZxPTQtxypG925vMcmA2uhGVuZdU5tLsDz6BAGzY8RvAClvYonec4qCuVm
WFEZhc8XRvBiZoxTSyt9j7YfNC+7fTdfAjH2N6ZLkPcBnwCn/lJN5/mNtsJBTSVm
3Fy2nvcvbsNht7rOZV4KP3U3cRdIikqTI0PKIEJsjwShGxTETMPVIVhrBfJ8MGGd
Zs8WiW09IUS5yHeYg5a3ny2T/dgmiraLAjYVBErNY418b9cMRYHJowXaWR1PhMID
z9lSkAlKg2MsqU6v8ODyRxf4lTv5OpHaStmbHRi7fe9wI/pEKez7WwOSFrwVu0tx
Z9noaRDmKO+Onuwue6cBlVYLjYDKORe6r1DVdQ6TPijJ3MGAyXgRvMXlfkec9Y8m
M1os4s5MZJcbK6RnD65WzgkO+56iF600JeXfmSeI/ww7qVHdhkCYbpUOKcUBJbUj
z82nuI7snqRxkXJ/pPdEqrzP2/DPWf1ou9nqjAPsOIuaEZSquCyaHDCG+2D6mfgf
1sDXc753PxNfeerG9+GBqlasSEzuz1DEcgwjpNX559H600gIEHf21Bfc8FDSgPGC
p24qdvtPXBBoka0yGb7ibRFxpgUMra3BmHhjfq179yGSG1Tkn03o2yhiCG+A/Jgd
D3b/N4rgcD7Q9COrpd5NZoLB4YFAO9nRyC+edBC4dYaUQApL5akOXCD3A5zfrwEI
fxX9h8J9wId5H6YDy1kllJiIv596m4Ek/4IE3ouZ+EdibZO20Wd3t3JSlyUXq9Tw
IktIcDaB3NUQ8xZ5kyK1/dcK9hO6FYGO0ECMJfHHY4YYPhwUvCzFdo4FY5+TXZ9K
LWEraEhNZnOSJj+HErZIqxeLLPgbEJrg1V9iBcuh0EQQ0ysJZCzgbC3BRtl2BXh7
lmPrMWqdmqnAvILKpJQVCsITeuA/NV40afyK7NUbFiXB3fpD/uOMt9xdiNyCEMYd
x0xUSLrKqr6xRJltj458smb3Yye/oXsk9fcFd0e93yfIKw1YoHF/J0UiWMJSmRpO
TlMLMtq3XQJx5eeYrrNW95roqsIJXfkPWPUkRrF1Mg3Jyj+yqQSDj3e0QozInqRB
g48tyOFD3OrxMmVm3dLhZsEjcDbk4BFCvG1Nv0tpV7vLrm/ty/OMKl3V7M7Uj8yQ
dY+f1qOO/rAJdgS3rY2GA6769V6mNRcVmKJMrA+nFxtQcUscJoDlSM/gsnz/g6l5
oMq7q/2rnXGipd+x9R6PQe0v14Fu4iycNqkojF2I5Sk5HbdOgjeOPhcubX9O4h6Q
pZ43aNXoIkF6jgZNCdN7HzTMagNcNqwRS1b640YzOTYQMUMrNofdXt1kY+ZVx73A
PIRydokxK4V8ovIQDxSAHbEv9o12rSpRbe/BTYFHHClp/6zgkU7walouurQkZTIa
EGgNZQfzggSaYp2myLIlm1Bcp/GtkN6FwGgNO4EZxtAyAjOnG0EIuA9cBWXGp9XY
iczYpW/MpgJ8D7xM8K5teEaq4RmrKxP/ml6syEXxiuNGaOcW2cB8BjYw0aCKrA6y
TBbAraz038dJ82nb2WmhkmAi844KEVh3OVYFn68fQXHc5lRyjaflFQF3BBSwIYiP
GE07RLP7pSXK0VFcoKkSMTGPD9omhyGf4GmA1oGvXNnM1Xeds5YlW0xUDHgNv4I4
BSIvjAgswiEY6TsvvtRABSFPLEK5QmjjiwEmQMMav715t0qz4XuFbA7fvyNEOBPK
CJ6NoMpPhdMjlWQ3pfFKSdBKYNVnFWYipEAebDnfETdrhfmtBtqAYsrnARjl5FrG
ij5HacTtP19BZpuBO7zZg55nSo16UaooC+HmYVXtP1JFhYKoSp2eghcN/DYhd+BU
Oky8JMoYExj5xjrGSFMLjQJ5GpW1GrUCgJEC5SSTxactv8hqnGrYimPtb8i4gzdg
iM2CSyQBRm6EQGZcVTJKXUuFi+HJgHFLYaolrPwsN+EgaT1wH+xTSEX19vYy5EAE
2wGHWHUVuEVwdKvUpjHF5qxcRGXtqNMynTXkhfhMVIPv8ZkGf0Omlz+ugROFd+7q
xU7I1ICIBBu75BbYKTOmFQ+8BnCxVCQiN/FMgNt/aKNQWUAb+vEV4dlf1ooBlvoK
SmfBZTRGb7+SJRuFw9/IMnWslgF8bgvGtQ9jITpvs9rPqGAqMeGcIIVLGObjRg+H
clJwFYS4XSZYDSD/vOTerBsTOLdL1MC+czZIqiXfchszT6xKyHordSGwais4Caxv
etXxlYIeXSZzsxiH8psEE2vDMgyMVnFnztgE/Edu28glrxXSMFxxIj5uBiqjyYrK
Mn51xA2c9+2Xbc56i1zrlQV3I4uYGE1ZH/Iq0TkPokjH01ZKUubdzv6E3yU+dOPy
xJREpUOrxXQyjzWvRDc/nWo96qI+emOAAQSCrXOy5FA5uZLfujTYfqzjEdc31JAi
PyaHUtLq1FRwtqFLlLeN5LEL/epq4LMA2mzYvwQayPzBb4Kgp7RAVXPXaG8+PS/S
sEZfIOKxl3Vm2ljURu7dhXNkumZ6SSAmxdM3sOAN4xeM4bsLxF/VqseXhWynP/K9
Q3pZPE88a8D+39YfaTmN1BsTdpaHkY0KBQ57jbRjmXDjOp6bk7cl+bLu+0l/he/f
lgsCJduKkoZNq5riko96cQIhjM0985XECgDaicJMbUwXxwdUhq5U25u3os3i4zF4
DPj4I9ERVM7L+RLqCvE4C5GH/U46xh7Pn7/ZBq6e3VEjq2PGGml/lv7ysRr1lk4O
FiKRyT+hW8kwsUN1bhCF/K1HsMRa0IOHuZ4FDWGmiV4XsrVEl+4qnYbUo2SRM15m
U815IsYLZCclJhmsT2uZM0iLxTiLMhMklxD4XwVhC7kB/FDRd51n+AmpOW9k+efs
FrM4vgL8AoObeUB1uLBYTXB67OlWH5W5ZVvxvlnAhVgllq4Efs0YoKGqoRywxccb
USStOtl4sa61b4+3NWAqIdx1c0NAG/DlApW/7EdqE8WP2RzLzkVrMGL0tXKMnX79
/oHjDih5i0/Kd/Qmw5cSpYVU60JevEmngmP0de/Kzn+i/BeTI0P04XXnwrelI8by
hoqEdrKnW1hmB1b7WT8wXOf4xVtcOlvVxYaOYLsi+UeNEQRH7vwQNNA/Q44Fxe6x
CKX2v9t630SuuvEMVO1G/3ohhslTnNvMJeJdFZ1LhxAAHGSvGYErp0w7rBBemOzk
ej4RnYmUWmD85/V9oxkv+GbPyRw8CPmeeXY4tpcCZbTMBguQyOd3zIKfcVcnFRrH
GIg+mGWkTT6ntD+gRFox1lWThNkVozzTeWedA4lRCkDkJety0m4tA+G42X2cTUK5
L07OeSrHra9dPQsuOjctAC0LHcClapl5JORl/kH2Gn8NuBdcVeAmKWgRQ7hSuqfH
t+4QQTsWfJBAJpzkhhG2WXnT7c3GsmpbaBBMMZgQpE+JMU9R4smxcnjCaU6O4489
38WoecWXEp4C6OBhWc3Hpw1ri57ZFse6PFY6m1bNB5BsrQpSsYPBV8vMXbZXhSlt
a0jl+m9+J24MLY4xNlay5WC2MvbwjJ1eBUxlSiFt1zZRWt6EuenVXpoJ36qtYI8r
iWud2/M4aEA47uZH3bJl4ZQVq83tRCnRsUT106wPTimU+QK77ATVcxQGMKSAi3X6
oMHj2jTFOvFQHCp4LouBDTOW5Fh6doxwpFLRibh9egXbVkx4cu7zYdbu3nRS3mpO
4Xu6UxVUDvxVaaLBLVlqEpg+P+L68NWZJGC7g91CGIjDpjlqxCIk24uAv/r3FuZn
k6eKqYzheuZ62VbBV9VQleyRm0JTSKATDjZ4d5E1K+mQ5JZKc7pWEKVeGPrU2ZW5
Fs49tAGpntp35NwqUmzBu6WTtzPJpUvhbe4F7OZxB4zQ3zsZc4vyJOMu5voI6H2p
nUZDEL4wJRWJU8PYxzfrGYYQ5j6XHZ4Q09Uw4V8kQmDipCkC6cFhFM2AjXyoPYRc
CiumzjiHRa4TXFi7I3MB1lJearsdF2pzhHl0DxLQhtUfRU/11t0lm9qiMcNgvj+p
mr0y2/bVOMJJKXMlBvNqm1TkdHupV6WvCP48utRfVhavKt6kcoiGlcRqU3IhgnOI
w4HhFhDfhfMnKy+fYbH1NFmGiwnUuVuNVppoulRQootnN/dS4jCdfSznJl/rbUBo
dZlZB2TuIRQd0Rtqm2ThdM5V8lFMrpyLPIvTRmsaJ9uyhIl8/gztFgwGa8TK2gmB
5MPVdkaJqw2sjQHNUamsJF7aqVGFqJO+Tf4uro1IrE1iuZoGejPKThVVOjFdTvou
INqArbT4zf0+EFJAZjFjKyV8nxNvIocBpDHKBznblMdSJD1soPJQ+sxc1vEyLUlq
UfALeiSNghjxTbuYBTlEWFOU83b1iptTvtCnOlt3hi/EkW8LSncNO+j+NsH5XuRO
7ESMtfKnFiG2KnqOcznCNp2cjQAv9EeeHurkhrha5EYFJ+F782PofFSVXDhOuvrc
gdETpySUVCKCYsd/Z/ZJlJwd+8S1UjtCc6D3U+tNWriQ+opqMmqD2j/dWR2dzp+S
d22gYD3Aojz/1165bEp0otGgciTcseAPqZgWSc1cfjrYjWW3rIH7GXNQLtdoKsjP
GNOEwjZ/4GX5wZaubcIPBJ8lGlpIJRnhcjEt40tTz8jnjKEVKvqkcWTxdN9g86jD
10OTWYoyg6fDi+Z1X+4QQ0D57iBtBB77umCdWKPqIWRuEEquY84+6cGr4B6K7XV8
vQcqU9QoV/ydxYHeoBfsiXrLtLhqlLStdAT/48k33QK1ZrDX7Nnpj5jy0e/vx5p6
TvfKxaFfCmkaTVnI84hplJ/M5aoLlFAF/vYkqcWTE3cW0EN9yEpX4WqVB19NAsJM
R3WNdRAZ2YnzCiN1vMqKJxgtF+zkuOZbeP3VOLwcU/a4lkqvnXYna3bjReSR0gfY
ULq/USngQee1BP6nPZ/Zq3tg0IhfbIuEellyYE4AIEVN+b/WEa/GVcUvnGsn2IWL
i1fZuDVEvrAVy2BAqGqEudmYmXzz3kHu45NdHwHnpSeModvZ27BFxkdZbA9T6YGz
d1q+rWcrAXK/9WtBxDpYh50teMX2WRJjytad7lA4YtdG5Kp5xxHOrKIHGbOa+Tdf
OJFzTSAqzyvR15pbhXoC2h20pZh1AwjSA7rLSJRk+ac1vWDSJkOLwT3UZm0XvNEr
WAiu9jImCPBdzfE0n1azQjXBG4f0QBhs6CGPO7STiXFNxQ+P7wZXAJgi5rZ9CGXM
LSS5CB6BS+/7onsk+7JQU9tdKetKW6dFCWE2Stx7TXk6wkF5W+FE0Dj5ov5YheB5
vR0wE/iGOB9dmyTUeHzgLgch+FreHiz9/zhJS/VuD01RXQindkYu5Rd06DYtM10K
CukoUQ0d76tEO2ISd0u+RoYg1OkeIPLI3cNHHMqpYOK5Wglz54pX8vCzF4gMHyvr
+JQmMELjBegSHL1K8rRVnXsylkV1riMHUgTNp6m2G09SPQbXLHm5sN7rATqqZDRt
I7bsEERnUbakn9bs/KhhU+bGRqN9v8l2SZFO6G3z0uqoWQsL5CSVWK/hYxPegF/O
H+wWN0KOLb9oVEP6wityo6Ydw3NHJbuiE9RgSh5gJx0osbSquOUmEWTlyvUzL0Jd
u4wTcQde9uqv7wAlSNA94la8EZM7B7EgCCoI/1hH2DZevHv9eG9mRQ4mKjvAJytm
iZ4IP9pjnmpnJzTNQuzw6E6n68LtvgK7HjfIGmfJWnSSK8hkmrDIdCz6m31J7rdw
sDJJiBYJPvtqx1C3FOZGLCMzaf/4r1+EDkvPTeoyIrh3v4jL8R0Ma/ErpkGrt+yK
bzb+ThUwwh3BFovRuzMMhxvolD+W1C+SaYBI03oEFa4xiLD55eC8TenYytzJ3Zxu
+7ULCssSkbj3ur1tqzLg7KRJun5PO2ICUtIiiq/347bkJE2V0WhkMatlTvdeX8NI
2yXF0dqtUYQtF3a66V8GFa7LYe2y7fo+2ESrIGSpqWQGhpTVwvOdwlLmQTGam/BS
tvQ3oqeE94EZUK1bwztSrgLEfzv3Po8CQ6MNMZjPFnSnr8zl0H/edbUzWCzLEc5p
XfPfFKhGViKg2wxo6hJYi/pvn2lPJNOvBTphPBwQ/LflepD6W6Q8WgF/DW/VYipb
3Eys7CU5Ca0YumynwloJzrrJbyO/DaHoVILO7EDapm7koPX5do4FGJZtjmr6ADw4
eWzhN7aEe0L2GZVxUKPGUEzOVdcMZ+ex9uQAIZHE7Yb3Hq4XejSzZc5KNYwTtcSc
axPaivnXqPT7kFcQXgRNq9REA6STz6AOJNrfbvNOqifsU3GlJyRHdBnDxRLrrWHA
Vc4H/FHEJzl42fAoTUQvY7pgcm/nPvk4xvZsCIX61mZpCluFt8xnZp2IVmRhaSzz
SbiKmPCRunU1Lk8Dq5+Sjpg76DlX/BJzWQbJ/jfGpDUWJYeS1IgODbg5yWdTpzZT
lxg2ipfaBSddzhRnhTgBZh6b+rFwB7Ol4U5GH5p8H7zAhbwEc13VXdGhIDcm4i9/
Zi887cOYwJygqbgJ7PZ0nbofosirC9Ly0pA/xgbbmETHgBb8/tkUb0EirUQSfR1g
mm9ro9nbNw4Gg/U6QvG309KXjaE69wfr1P8I7ExEV03Cnmqo1rw79SB7cCHI2IHz
z61aovroTeG6GV8GUUARxH0w91zJSOLG6jc4RKJ5KMK1/02+mWe3NZ5t6Kl3uXFO
H+zAhBGT79fZUpMjc42NCBwvfpMjUaS22BWyo9qjDUIhkOJYjqD+lkRbavC3tgc/
CGy5J02l0kqaGuWlKQCzZW0sAiqcFahzoxEdsX0lSOrznQuYqrOcLJu5kSdphUVP
VO1mzr6J2mUXZ3T3FOkwEZmK2gnszeCsoR5mnjkppWAJ1RgvjoCxF2CE4F4DCz3F
p6QCN/ZjPsRxOYYcEGidV+rk5NeNpsfB3Fviq0KWiuuuRrLzBPJRz+CHQIE68SP1
xv64EAiPe/EPPzZQNMFowWZnZW31Mq+5fmX4/eNYWZpveeWwhNBR+eyKnuPHjb4J
T+LhFYeSEFRVhNy0ekC3p7CkUlosuT3jkfmOEN+99l2g3819Wtn9lHIlioGhEBrA
iqAA9d3NamCegWnt0ehYGvGL9WJEXQW9pYT4q35QVX1vqxCuOfC++133448VAYtH
MMlmAbffIKqRZHcoonaNIArhy3EhynfqW9hXvvdar1N/ZzOWgdSrrL7M4F+oMpWc
InF/fTgAQz0FpTlVb66CaD/AmhEt0ZEqklZQ6RBN4h2T90JN4tg7dqCim7jA4ceB
mqoWLMrkstk/3JD8zWOUbKikIhNVdaNix456DJrfW60r2xm+flkIVQdGx8zjvgyy
EXPXme8H1biM3gv8RljaxfAcSZw50mngoNdEWcqLBD3a+qNUr54a2Qfkl049YpaV
SVi+GlZ5zDAJ8eyVDM8AaImGaNxrpsp/Hnk7W6jAN6KSBBICMg0cPj1+2O4zCyN+
UfPjJUNEwIALIC8LqmlSbrhWZcHsOgo0vFvHLJB1HHRZGyxP4G6wOg8F+BEGYMZF
WL/pdS3iDWERJ9K18l4Ok4L8Q2HqJwPDSOg09hYFoUqKVz/ofGa/eqUE/KwbvGtq
4Jupiif/ER2ywtmsFMMlO7OQxHGqwVMlmlIDDASnA1tyPGdVYDqbHGsHMP6afdWa
jiBD92JZT96KcqOVV3itC4jcgfYIHb+VM32pvX8TmszM8Ud4gzvEOqqY4KEB1zrP
sSrFxI9t8QMaXjL1J66vMc3j+z9q7mC39MunIa0W3eHmEiqKQxBkuyUhtRDScdje
b7Sdqs+m37PsEeJ17lpCteUoXODLuDsCkktiddb4J7TsoU2Ct5I/2S8/9+KgoZdj
g7xzp2bCH5DXFVOAD8h06312rXaNrf+bxyDObTM+uF5TVGXKlTafyqxPKUA0i7+B
EoD0Hfe7NH9xORoad1+7TdqOWVSsJtKFd46vu5yrRe8cz+b6utYrmALLm4i5VvPO
p7Ofse5mmG5Lo6F18YzY15cz+Et91W4vaL7YJikMoK/Bc4v0dZ+VMRXIuIS6huH5
2oIFJvrxYwJ8usrtW4RYuWkTvPrQeuT+i6CG0lAAzEo96W1nQGyOWpybTWYsXp0U
2LFOZDl+WHUaEqiK9AnLEC34GmdfQdETu4YF8HoMG8m6aX6buxHVLZ3Mnv3iIGtz
niBeY/EJGbI2OKTeNf0V41/tjLVT3zVkQQWE6+Q4UCPFg18Q/Hmc2g1acs3tZJXD
WuZQ2+Ez2elWlKZ/gvVdkfR7Vpbuyhd1b3nf2QlhcT0FHh9En4MIdjoHNshQQC0H
MKIzMySrpkE5D1FS8BbJNnHsg7iaQBU2uBD7cJQsEk0OF1v6rZemXQWI/Mf+8kWU
ykbz9w/qd5csAn3sSfAFAu3RDpcC1sXwYv/G2B40d+IK5C4I20p/4xzDJfkSCpS+
DqfKKmTlAbSJt+0+8hVGzvBxE4cmThPSBuHpEbxJXg0wA2xg73Ng2F/0p7QyiX4N
BiXTcuzuW4fQ7G2t1wT8pKVf1ShGon9rGtmkWxOB0dNlU1NfhmS3k38Bidillvn1
j++MFEZkANwopnZj0h5qfXIdI18HVVn1p/D9d1VYGQqYWQ85i0Dr5mP+6/OJ9NRR
IvyfjtymqvEX+ZcsrHGWpniiOcwcBxh3ympHZ6HK89vXGcvR5MYS/T39t4k0uSNz
ktwVf/Fyh9B7G3r8J9CebrjZuCzJfp15aKKcJ2D9DQUH7/4Pf/FoiuQFNu4xFaLY
uMng4syqyW/G0QeDziWaXrwSefU10XjYqc3h+MurbR8bwm+n8aDvL8Am2v+rkbRo
tTXtySGgWd/wWVi4L0XpJwsNqY8QcwG6fPNUD1GPfWiDg3oWOG/rlrMmJVyS81Kz
9JVJHGL/JOPBZJiSne/6e07eelotFWz75gfToDJ5WiCb6I2xLf1e4GKajuy7+ukZ
vFhEhHF+MwUtYrk36W1gHtUlAIVJmfEirNiv7yGqTzbNPyX83kmdLn264S11JctC
HGjAq0y8Tzns9EaQIHssr7Jm+Y3q9TT7hryrMy0990t0d8nNItg3kRVkfx/Fm6ug
mcHqIIL9QUOv9iyw7aO73SUfEKx+Ec4efZGsbBOQpvVsx23wn04MTcObnPsS4sGF
9xk9Mh/NWNH/3hr/lipUVAaEdQfTa43exwj/Vm5DBHamRYsDqlTq8YttdhV1cb6k
tglEwoVkW5idMnC9IuawnFmX3dVCXvlYAFzVDFDT/A5Ou6e9I47Q6wSNEH28EsJA
2WLqFCcUfvlea77RtAjyHKRytOFwXXKqBjsoNVGlFKd2q6I9o8wzyDdLyr1p5T0c
u6hMTwrgcP1p76/1q6oB6s2Gjd9ONwaasbe+0JggX9RqRTcuMCY+OJn6U8RhqL9k
FQHFB/zDagnsn8/eCTCcZbilk+EJaX5VJ+/o//9VioB9SW4y4faKYEyS489poabz
ye3tzBiwN4gUYHzkObO/eXRjiaTT2g+plhL51JSUEQZsMxZyt4mr2EX++ikUKG/n
H/7ZrlwCANXBz+WHEeu9lejj2tzjEf2Likgyrx20cSBgIU/hq6QNzhFSaU65I9yv
lOvXzqZSyAPofFS0xJzTad1RKr2PkP49MKXV1desC+zBN/Rw+yhiSrnA6/ugGpl+
sIaZLEs4ZXK25j/40mIk44hni1fMUa3RsrFuLZfHe4lky6MF3yOLAFYhY+1z11Mz
YmoJ40nH4R1wL94E/Zr39alJ596nQmsykvB0CcXMLIY5koJobX1mNBEPJfxU6fK1
Uxxbrk1sfxD1L/+WWo+n4z6sRu04pECDexgU9jVTwPHR6OQlDl49iIWlmuN9Ajhx
60dgS4C3i7evaPZ0MQCrdPPWicC7NDZRTJTSAkK2MD58ypDbbnxlGpDIdspmjTpS
sqHtVDMl7NUvL7cZMmsAPFzq3umqiZyN+KulYl6pVho1hemFdD8GGrb3NGBhvZxr
3V2/F2QqtqmiGctYXw/dglUpcVHLbQoQWs1jhskfMy694F+Avl+tjs6zFrOi1DnB
qGkcFeDu/R3UmpMHHy5Sc62J0JkmYfF+TMGZV3jaBMCC7rk9H8rQmCXPFoFuc6Km
H7OyWYNWk53oyyZrJS+dwTUcnbrvw3/+2BDMDvcsDqJvc5ZDpOO2Mh0zLMwfPeTC
N3Jzj0JOMdzTjdRWqZkD1A21Okd5iIzRPsIVCA+F4P7SKknmCFX3xrmT3JH/bHjr
KHJmqCz4AkJJwhKu2UVa+9ZLvLQ3XKL58c3HTqqjVotYspm1GNZZF1ccNf7TFTaY
AZ9RAIse6+02Cpm18YTl3hiarziROUykoV17VwTIuDFCy4owA7M97cTbXojmwXYl
rF+VBpd5NSCSRmIvDym+U6fk46QR55JWdgu/42uTvC2q/NUEztwn4ur0XcHazy/x
ynaM/vMTHuOVw8akDxQK1aUAFrp2y8EXxHdBRA5d1+8fsbqwiDBaiGfdu9nMrC4j
9k/oQ117vZYRi1pxdig7PGkZkWrF6kRw+dKnJVKXAE1d/9J80H/J6c0wRanid0Y4
OW8UBpnu2IwmMgAA1u+KDqcYFYNgfixumBXX2mPzLZ0mPn7tHZcVp0LMVWUMnCIw
kmVUsEHqbb5+VtpkZ5cTJTXnS2nxfvpXIAehNFRP9ZMxt4NDfJfGyBUglSEllRtq
aUGw1E6QajB/fvt0fDabiwx08iqeLN0e3cF5pfaGsmuR+UCueyITpCg35A2km8hZ
qHLduPPAq+a7rVpI310AUTZyePgApD1rMzMd6FtmBFEFWp4WQYp1krVIUMzoyc74
07AX2IBI84PVW+QrzyGq2EkiM3MCkNSqgxDOhQNcDB/RAoofty/ZkPihlvvmqgpy
O/pNXKKWVMsV5nh+JBUMeVXLLfSR/6hP8zKkpUBBSZ7P6n+hVFvn2GPIZMsWvQcO
jfXGyQ40nlpttz8KSDrAXjNrWHGSMwZqfAy3mrbtqSeaJRqF6BJojlUPLu2N5Euh
ITbuFSqbzXKfK7rthH/lm46RrKIp3hBjdcxxe4QaUqKlk6uH1IdVxWx/9H4jYjKZ
23TW6mOoECwLezUA16JXKmsvUPdbXQLd99K5n6SL09wPtTPmu3NWP8WC8T47i4rJ
/f/Yv4IZOjXaxByU73kVHzblg/UqEyo4CWPnXgAtiGAuwrSZAnSUR3p+U6PdaKST
TP4a2uJWHgWWEO9+HF3m5u7uCtwtolyHOOqkZj2oJ8O86i3sh811Y0GUQTtJwFaG
/ysOW0YALUEEhEkhu7XIi4t79ziFfVp+rmlBWePebGK6Wkm9gsDRRh3cSA/W6hZc
nypnFx8SH90Ls7y6ADGPHIEmetcWRHf99LIFhRVodBKRi6WQTtxSWdCFe3uW+le+
e4KgLlnUiU10oW4nAXGa/ZPJykhzPPvMfELIxKUGNpNzMhDZ9nbO5z9Bk12ZHhwc
DYvfXWnFphCVIMYq9G7g2IUEGwroJLy46+d9CIUYci0hgMT35efpMnwLpXaQ4T5Y
NTz4qQVIU+xEdPTGREi6t0mLBcKO+xm1CdYlLHAUC7v4750tBEBDA/hxOmy3WAsA
G/UB2b7dIZCndZMEq7Ynrl3d5IF9YRftc5WYpOKO/VNTvNKVI8iDkBnxUa91L9UT
0reSdEzvxFnCgwA9LBkc0JyB6zYVw9cGAioSEid4pGGRKlcUhldKdM6vJPioFuME
uQUgqKPZed550UJ9mujjmf7rMrEVHcsHFI1hC8eMudcWdMcnhTJK5S74QyJe7JOi
9KTKyaCPHYYVLR//PrnjlPZQxtrAKgApxpkEjfGyQkrrseVYYJWIELne9NOLkqjU
iqtk9x1bJxW0dU14oHCLmNYH8jc5Wx8juKbM7tSB8EeAvZ23mHQuQNzrkk7ZNkdX
EeSL/MNM5eyr6uIOrO3AoGq0ixnpy6aVRbwAe1IKF5mOFkknK0HChAJrI1e+tQkR
qC2jMjzN0BX204YfQkO2nxWlA/TV2sJXp5v/rEGBmLwQwzqF+4jU3nLTzoL0ujSr
IH3SOWnHsR75R/Aqgzm9VU3N4KbNPMiYYo/RLE68JwVlGnOZJuCFTrRLjwCjoGEz
NEBjUVIb7uXvDXwUGXbrOuOKBCtGtc81EC0mnmkxy4jngJBWhGb+v2XEk+qsLhxk
UW3Rap3pjJ2ncliJYCeN1BS6qeonlYzaILV/xQDcpfnM0hDE3j0M6OAxeZg3aoXP
vXNP+XYGYU4IQIuP+9ct/nEzKertDD5K+cOSxe9hEvLd/gLFglGTC3TCvOZPDewZ
5JENi91pxIrZQu8nKKugtsQPZhMCATzPx4mTSAtIG8BUVkTzuk8xpYm7qxH6kITL
R8FK/hRs5fNOsShP8jBLTA5FwxZ/IothShHUQ7qiBe7Jhf60YNV3FvN8cab8UkWc
EncqQi4a39EqFsEHKsjG+KX7ER+Cnj3HxFLCB85nr1SagZsUzCGxYzNlQoR3P/lf
6pk4ib6kXynP1SXYbR0EtfZuB1ydvI2V4jHVBKlT9tfTOgxfYrmwqFlltqXHVLpK
Ak+JYwl963MhIzL5gVyybpQ2fAZq3X08Ho98Jcn0dMCDwwF36p1x3J/KebsIC0rh
bRx6Q7S0cZQnS8PYzHW+pNkQGAd/LWrMBl71VWar6BRiky3RNp2fwHPDyxacjYjQ
MyODb8ry/QJ1sppP20dNS06N5Kzggpw1mhOLqX8NU+NYhx36Im3oTxMnwTu8LzUB
VxrCiWTiJEpH/+0FejLJgHVgjPvpwMUN3VNRY+ecbX7NDGGt8nrrZfPUVRwG/8rj
K/u2AhlBttYR+RsVdviL7TjxzJ29sqPVPyKrsmsUuYzTwk4pMfFuhyGAKPc+czCI
nHJG+PIJSGJkAhaX/xIQ4A6DpEk47wXL+3iYb3qa3TkLcsUjRfiszQWNitlkc8l6
q1hgbzEE1WIq2mjLNb+1GwIWue5OO2Z5CiP3QblE19NMuFbPRh50wNOisAYwzoFS
A59UCfdBPg/Az/PgE51RL9dp4dQBBes+1qxnvDMXsn0S9ZlhULJleoPQtCKZnbAe
gxQXjFtaBJ4mIbdeo7zd4AD3Ynd4FOFn74VCqJPOFgxisVy+SW0vMmMn6KjXYDph
az0PxwqBFxLRPKXIfo7/Ix0YMfwyyOyQeWnusCTvm2WVl1pptdVbz8cf+wGWg2db
s1f16i9so95RuxrreJnvq6QAUTYzx6UXIlTI7ybmAGVsAhE9XkhR6QODtA3W5TZf
YQDw5/Mso9C7XPpIhazT9DkocHAc4ovNAK6hoLAcA1dPjDyv3HZSMV73nSCDusfG
ko4ZIKVChE9HstYxRT3FjLZrTlcD5DGs+Q9SxF+DHwNzRnHVknLIHPlQITL0xsC2
2p7ZOkqv9JxsKUFPaYIotLHVa0euMUL07iYkQO7TsIrZouv4qwW4qolYaEuTay2f
/CDsDkmqo+MqWDgIx3ND8RCgSBiRNtPbQ/yVwA3mMW1nOvqYzLCvmlUdXcZhbQH4
Nyuz+QUOzUtaOtBh5wFbb8Akzn+lGcWrcL9NGSqjlJU2nyl8BI9EjV2wZ/wfpcWZ
bdfVKp5Ghw0yBbpGiX4WCJtiGCIviUX1bgHZSgbAd+rm2G4dyhJDK8pu0tqcQ5Il
jcP8LGgNA27eSy35F1v1DaLmZFSfw6DgalGvq+ZzyKU0jv6uAu+AysY22xllbNUz
1yzErbtxeAmfOyKJgyH3DyLWFKvyzXesLf+av820krhIBrbQ/9IIFlcyNx5xlt/t
z8ySftJ9V9AHlnrPleVTUKuWZMWAffsp9MmiBkT0W+aX/x30x2H1tCZGlPIJQRbN
cu5OgwPTdCWr72Mq18t5wn2OgVsKNu7wOsIy/gS8/yRbLOGX1aN0Zv0DtUW2Eg1K
Q42odNOelJEMpZxRo/jlfj9Xpkb+8tb8uaIAypKF8vxNNRbx/y2CdDwp3wJw90LS
uxAQIMEZ1qvhp/6Euj8VPwycVNCpbWVVrdhbyXxrZlscC3RUrMBIA8HK/62uxHW1
9FZvqhsDIFfGObHxVZ95gZ3/DN2H0K2loQElBT9zM3ZxjtNow/FYes9Ieb2hYlT2
WgwbdzGDKyxfa9vFBebVnbP8YtstHgtE56E2BUmH2nZho7r+dAF+HtXEm+2SjURv
O48ORsutY263DesnRiIsuSE2VSiqwpDpdWltA0NdoUn80jELqs7x7/4PWRyJn3m8
V0nhZ6ZqKPZzH9GAFbwG4s8NFJhQJ4QbcZs3JpEcS5xaHNsOgKLNSAjb08rJ2Tmm
ZncM3CrotaKLhrtNSrrcc+u4B4Ad2VYR6tA+tddFhexImr6Kd1hQv/+3faBF6k6R
KYzsfu0ZNb0kPc7iUnaBzZjt+b/vT7qfsFk1+2VntjkXn89jB0zxDmBHEnDoBa8R
A/wBkFrII/jJXKA/7gRWRwf6xuRFTZlPF24fg8O/pVAql9L/swqFgvzAW0VkvDuu
E1DrTEKQZs5WLvyUockxiT5F0cMUmDmSBVvy25hkZIlqTaxuiCnMmo12OvQJVl4n
QupeH6sq+nA8S1WPcdmF/EBRiNfgvo2Pc2kc0l2rri0b5GpFICcVyeXk5rRi7kCV
GcmNP2o4uplB2R+BkIpiwEULt9z8oCGPN6cFjJ2B/g9H1XmDL3/PnSqpRT698SsI
99yEfQONYA4bN7S8t7R9QXeP6T0oyixDSGOVvyn3ZjDNsvl2LqgUshzJ4cNsLG3O
9RVIHg8fmAnHBz837Zbf/mUZnvRcx+/QN7s2e0Y0f8goZG3Ha0+/fl8tV7YZJ+LC
apELwTk+gRSwqHQO123rizXyt969PuCfw/+JC3rT0F3FzJmYa/wNwwxlCxhl1g9M
eM7TOrPSPsE+S/nzN9MypMEOPaguuhzkTqno70QyOGnWJKx0i6dflsUOY7Ab+7m5
Yh0Ih6jdTZNkaMgb42m1LVZUwVO4Uwh2tfv7w+fWc9pZXeqoZvkSS1RdikL0L9gS
h6nUHV/yzAOJ5vKv2X4EhaU4QsJTFtSLf4F4xbTC54KF29EP85yqrVHw1B7TuZVL
L2d39Wd9FNaiP6KLXl8vo4KhFxKvcDgfpuzy+MeF6tbYdOGkcKDX43eyVXWAX0yT
3cJgP68HyFc6aabYst0IBb9ZWkG6uiiA6sYBqozywEsxniBvUNdv106BPGCTKm89
fubUwx+KmL/PizeAHJR2BiEwCCQx42lb41GRjHAkwZCM5/q/BhWMEXOqouS77YOt
oA5r/Hh5mDaqFutb/cLOckL9BYEolKxo7y/AZuoMvtt/TXBeA8G/EzKh7RABle3A
dOZ6BMpSaaAQW7x5v1AKbwJGEVJBCr2bo26NGxr2cVgySVu+1FLdHCWXC3H++AGU
smBgx/BTZzQUCwmxKDLTBLu5LmOYAgl9AcZfEDgeUKbE+Ec84/diM/qmSebwkQZU
iic1BY6TNmux+dgGOp5Cs/Y/ZZTzrZ4Z2hk/Yrb1ab1WJ5Oz0xkiUhbXIDGsCJ7S
pu1nXCeOsJG0UTA5kIcRK8pSPoUIz6ukKrY5NfW8PFUY42SLRoYpOdBCg/QtNhHK
Qm0v+YbH3UVwfYaU0DGpIyaZyDOL8TALrAcOOVwc0NAdl3qmKxNTuf1MgyPN30Sz
dWA955GOtlCmqqWubAGGuusGK2gyorL8s9NVEps9/bCgndMXd/IksEwQEXgb02iv
ovEmJRBKajO1pXygdt2/wZ7QCdK3cbNZo0sbv9k+pG9Vr2egICzSko6xZ00vxNc7
F5mU4zwC+kfhY9GQCHwxIajUK2Lhv3P6yH5Sv2iIdM8OgvfpzrHamQyJHIjnpIxw
9bwHxLetLQr5hYgYSIPVcRU6YZi3AhcQKLkESHWZQBcbgWUMCSX2cMVNgOSmgJ08
C7sh+IZN9Bu4k6wPyUHh02XgkKFisOkRHLaiGXukV9teXgie/Dah0h1NxtQql3S+
K6IbjmQVkIEbPb9QcvY8sRg9QkXzY9bUeKoZX0WuZkKTo0xn3EbQIDD1rTvYewOQ
tb5E5GJtK1Fz1cL7nJWOzCwAZWXTOSxMsOpVdXAQ0Wp/9h2fDZvAppi5+dLHk41T
0x+8iUv1wD9Bvpw+c63eXtVu5Jpw/YBWxPzDa8VlA3CEm/fmSxNik/3YUPVMSIKi
BiED4El3mXw/iPttp2TJyOi9Aoi5Yrm2NBSV2eKCMK48TWUiocuVtCT+xQu+e4EG
pGqKatVb23htI4Zf66G9ui8MTX7KVigAkPwEt2mgAK06BEtTQA9HXaq0XxMnVkCf
regRFjBi7paOrRJgfhoFx18BCht7Wzcc7ZzD9rpSvsFwTJpYJwnRUC0Vtknup/IV
RI3gaf0IUL6ID6Ut4UTbFLG8KxbUbdZ/H8dF0ZO2LhhiAJXNkri02GKikfENJTuI
zEVNyLyHyYOMUj9tk7SNkXtZpx4i+ehBHbzhFKqJUn6+Kj1pwY6klO0X9lutmuSX
CXzl4Zmc7UrczVXYDB2o7B9XsF0bgCzsKaaVMYc+tLcQA7l2kEc0HussUoo0gsqi
nvclfDRoy0a7CFTKzIbXoj6QMkGgzJhqh75cmASkxvjvvHmcfxOFXIof4tt2XNi1
+qWQy55eqRNOTn6jJdg6RlCOxkWe8JThdI+1vJvxCKYlVjl+tA3+AA0DqBenXUSN
RnsDh64AZjyKH86qRfGlzvlBWwE8TWQ/8YJHElX7IcuwH0fA7o9NB13QnDoEoXMh
tEBCjdVI0YIJ613bJkN3PIoMGPi6SXEn4xIqiF3B8OqMkRJ7cUNWzzaP6G3o75WP
S8Zaq3vFh26q9iY8IsxJ0unorAhtHsbkBIG0G4m3ACc23aX0gTpHwgJocDAXltuq
9HzH0/uVWbWpRtbiFaNY1cZYlEqzJFp7e4SnjzlXmdP5bZ+wadlMhJx3+MuFttlk
Ifq7zCFWpByKYEVr1WUdGh/dFXeXHjK0sdm8R8vCq5kuEqY9ihLxYpFzo6E78s74
98XPhVW/mBRG/b+GTCsMVk+V6Bv0wa+xIwnJiGpP/6y+ThDaFC8gdPIvhYKJm3fm
amBaeA6E4CzEsIR69VMty+JkV+q/LccCSakfp+pPtXJkwSCKrfHMS4mBw2nF62pu
zSd35Y0V9pJiJ3q9vBsxCEbL0MHh0SXl0ttJlZVonWkU/EJJl4Ovwq/5/Ww05Ne6
cbajM01L63P5GyENmzAjYZSlVrBxwMjfYbv2E1QCQehIvdfDirWW5Soxoaia5C2q
hdbeumFIeYhrUpnUY885J72OJL9Fmc8rIOWsWXWJyU59BxULY5tJc5TpuCllszfW
CALwW7XARPitCX3osPYc5agclz89iWO8laYgNZzEwPAXZP+Zd+hJEJ5bA0ZTRSf8
kZWkG5fy9RnFbAU/JnYszaviXjuey3AxewKtpbh/KPAS+Uw2WR5Sf/vg38HPhVX4
Xx1Uf6glrANKr33/yzniHu2/3Nrt468eOFgBY1beV414RgD0bWYngH8IPRqWX2MC
YgSQgVMAQX7hPkbzaNKPDUvzzkdJfBc+Dy+YEUhAup5/W5e2dCkaszNO7OD/H62H
oXBdvwwA4vD5ccet9rHqILSD5kiMn/I2jvYsqgrL3I54ty7KFlUUZ/5cvwZQqMiZ
A4F43LgCQ5vCK5N7NPpaM92pW7+mLi3WvygK8Z9GEErUPuOMBMLI2/odcClAhETV
Oqw5ux7xV6pm8wwNQPvrnxjLD/fQKG3e5LqukPoS9Dg+kb75tK++sOYZN5LStN1p
e38jgXgPYhS/iqitQPqZoF/XDI78cyytQj0vFMNObkbeudV3VVPSXBqU3WAakaod
PoYVM6BoJpvMe72iu0Oo+3oaK03AdUNduL/nTyjAjmg4w1Xpr42K1OySAAHxv/ID
UxjjpP+ZXLvTKVg5B77lJ5cXQ3aTZUnhDh6vjdRcwpMgXOBCnXJEIv1ddG2RpKh8
eIj3PoBthpzGY5Pz6iJDXvVZG1IKykt3TCu6Qi7I7CKT3mfpCCg7Lv8XyOZVDqbQ
ccGrQxu4FKwzCOxIv24+Q6Nc40k3/SNqzI5epsQGYyikazFdO/VuFUaGV8NnQwpe
hvRFV0ABVv9KQ5dkjpDGP6tswlKzuOWqzik3C6+/dIbhuQbsuQPtMTk0CaU7gZkP
0bkiOJEXN7hEhJa5cShGFTTZfjfYlj3ynHK1REbZXqRgkyC94YJlhQqGsKwpfu5K
of0INiuVF9KEIe5s4FglyjBoCm2/EDiix005BhtKiDr50E+zF94tHGgdcf1Ym4A8
NFAa/qb2IZ4B8UhRkiiKiQVEwI4oGuuHDSS7u/ADU3cSLLTZ9pt7Vj6nD3XGLdoF
+pGfcsa/uk3qdf5PP8wlHdyRckPh6JQT1bE6RctFASZ3TH+N7G8I2Em1nS/Hl5sJ
ej0XC2WKUGjtNs11CT/hClEx5j9az8aaKbyQMANUbApVScaxS1R4/nmjl/ZZIJLT
ZDCY8fP4gB0pJEkvJmGVmFoHRpjW6lW5qq9ckK0q0t217QQeZDpAn3Chmzy0QC9W
b2+CiXjrL61EebzpcjO89PgHX+xOfrnJ9kEtStWasfit/uhQCza9s78nZinqUAzo
du7/zO6nAHV0Ln0NrKyJ2+ToSh+IUCV4oU0yYEzSKXXWcvH9185diPgLcqTRW9pQ
np8vGMTjc7NKEboCJMsHPfWIXSwGnWKctPnH3B9mJKQU2Ukz+FmGDj2pyDpSrjT2
HH2ujpmqHLY5KqHhbAvaXuKECSQhHqqQ6KxbvwHe/f2f/iSFRxhZjZ8sOnR+r8ur
y98N7NTmT6VKROAHX70MtMjGtdkp0b3IwpSy3+fgrX+sKl2MQI92uEm/a6dPzjof
yuVvrb20Gezxgmq26cx6Bp2l4B6IvhYDgYAKNC3LXvVx1LbG5MgdkPBarPBp/Zza
3BfT+KCf8mxgzKdEAoXnsq6xuI6F5Xar9Zr6sg7zsfNBaMuqfBjJrMvFhYxbD/Zc
+JgFbssPOSrCIi3N2gpl3ukK2KiQukdEPN9sNXBFQrLLX5U+Q0kwMxZpz/CPdvs9
/Lwe9R+lu4rpugyXGiXJEUuzVveehGdO17yPvr+pWp+1IhoyHfpRtGYP/yuLGBds
+QCHLBSlqW5r33M9fiOA+n2RY7TOb3S8xViMTvapUUllqnreaTZaovgsNvJf+SDY
nZX02S9rvd+Y9vN5Ur6BZq6S9B8EbPfQ6lvBO97F20xccHFS1yzTrr/IwY7rAazS
grSJNfXnxISi20WvUGFsdox19kObEFWi2YTX2RslXPgUQgLJJUb5I0qgJKuOIvRx
oC9klckQmIvqmnG/it7Ub9flJYb76qYJi6icCsw3WLNKVmh7hKP3U/JZm6CpPgh6
Ku/8oBrotveGHjz5aayYBE+bl4dYAd7nJgP4xXVFB4X0SAXL/Q9X9opl05ZC5GY/
gIC19tZWo9Lgh2WbcReXK6FRGJyAv0dyfygAAtoejW9RNdBrKpNKpKe6OEcEZpxy
xBTP4AZA4dLCWwb3Hrfxstpc5SacufqUnJAXu9esJqyyGdYvRC0+WgRy3ckuEVrl
8NCOHXfu87uWRL1L0UlQORnD1btvZtba4cimOziig0Sub45zlTvMgVDIv8MiBW44
5HxsKvwg3hx4lVQ96m6Pk9bFBU/PPZ2KaN3qvmZRK33XXz82m7noW+rNJo3hNW8P
Ji0JXE5Tj3tQ/yT/FEVngGCiLnH22M5z75Ey7nlsQolODc3oeJmeD8n4o5AGDITF
zN1uJdt8AE6llt4BMS0DDxvOsrjkpgsR8VGoK1oMhLVWt9NZhAWGPzp0t4qGSVic
Dk3DTtQJodKRbwtvEMssobtLRkqFUvOOPkwPkouQEmYEdgFzS5d+FefPFHlZqISw
kudP5wiZYMDFlkwk6QpBc0Zu3nnaMNG17iPi7fs7QPVtes0nPIwd9JHiw5utnBL6
22LPn0SUEzCGE0faq+lFlmXksGIpxREJsMXFvOcemie3sY5xGTY+MO7SBFRoRPLr
yV3ugxUHhtgAhM3h7Fe73fyhOjkKJ7fMhwHIb6BQ6N3OWw9fi/3V8N56Xx7uYPV1
z2Zz1/pIT5T+vMTFQBBPs4fmKj/QrPvvQEnv8H+2dZ4P1cEwn/UmtnxTlQq8IyxB
I5OfLrWRiwLjTgTecwXt1ePmIWbcQrPFoOqm14ALjDcWbc7N3SUTb57fwoRIGxuv
7UPtwkAukx339WgCxPJDoyV2cfeQcW0Xp20eyYB0VSWLOwg+Tdk2h9N7Br4RIiZT
S4AgZ8VwM3dGBvdwMRhkak5g9FnvmV7DOs3zZetnoTLD6aEgsnQ9lxw5Dhha2Sb0
Vxtw4QVeBuX3W6zmbKkf6H1y+6BUDXUfvEKQrWc+0jcuGuSMi0zjkeiQNPdODkdF
PNwRCFdtL8hn9FvOaxu4B7kEgd88kErJB7bn6qcStNveqd96rwt50v+uYeXTKrY6
fKfBbptL4d2Icsvdt/0+GHlDfslV9zdwgFceCcWAgLZjUzF5MlhRLd7Zv+OZQ1ai
PUR3d4FebqgU4Rp7K59uY2hdWgF9vyDZfqCr6opWx1ln2Kqg0HUkx18dyb91wlV2
RzL/lzi7rbgOJt78EFJgg7XInUwmqPsGjE20Y7OU/squJz+Bo/w8DAOix5WTQc4q
/ZxAKXMHnr3y3WHKeFFRxfz+bqzrrcUf0qN0oEFEGCbdC/E3kGo3PVtXvixFFab/
OIBpSVhNOtELH8I8i6rXFIvOZz8EKrOiuHc6ORhb4HnY1q5BVHLdVi3jEy8vV4U5
YhPpx6ggfhR0kIsNdmwoteME50+cv3TK5P8lfzvtRoAYYvjokp7Zjq0ZZ4c3yNph
NaasuuF0DH8Tozv5E3GTwEUD9EKpWP6zr6Voj95cRw7JUuwmrVYDsiHWBfB+71li
Rq+orViPSuoxvfJMSicgvSTVSpn69mQK3a7kD76PdMNj2lnNT1/Qi8qgHj3Ph4mc
IHY4BfVDBHeAWRANbErPJJSoeA1YlShOWpi9ZGCXHHTQDICJNcDrsaflW9U7NAWn
PG+ipglLRwaqM/X4lLkO3JB+YCaIaTpvX+dayLBOarkNWPtxTniJRQARAVf8gU5C
44OiLW1yVSM6tcYVmwE1hTleAmF08tW0zwZaTtbR3pWomZ0lCamowL5dU0/HJZCo
8xy473Z0Bv39smrABy5DhFYag3jbjLc2sL684fcFY6iIQMnUpVXznLVkYPRCzqGm
JcgMA+7/F+LjWnlfqVNoj7qoh4AACfxFdUgk9cZEYIiVhut1nfDvJMtk21BcdwRH
1IA794DZSyrImiyRRhYtdSX6QMDCZDIjHTVMSCU8jrwaurL+Tph+BUle+KjWtLa9
oqmB3AsuwjHuGsLrjKx6nS82g5nBALWyEd5wUfqUMRKzLYBhwJv5yuz1x9LUGfgE
XiQTpMeBOd/JbSBZDQbzHNucAZR7qpLrptMhZlsTjf3afEA8oq2x/lJDa+2TwRQ1
bBI8MFKXQSLgJh85h4q2CnK6qTI6Z4GH7craH32fMgjJPoSRU5hk2O+E3/dCRf72
5FH5xWEjq7NTsO8QwvUhvNT76h/khGt7DDxXfr/KnBSRJby9Ii+gy3FjAPHN4sf7
olH0az/bvdds0wQSAmGBH5wIIKBBzrwTCZeAvrLlHvCZf2CSbT+ppO2/ETiBTDC2
YftCXXj+Dz1xtky3T8wi3beJD8ulypP9tE2MGbhtSeOABeNy+lzTycAcQSALTON1
nrb1/cXYU0Ht3n3bKPHz7FbAe2LWGkZvqJ3X17B/e65k9kM3bRaYw+TGB4UMjtkf
5njAAUgfPo6t1gqkPgfHTXfMaaoOjNxXg/3kCS29Wx4i0fqFMS+VyY9/M3z8SHso
ma/YmCYMQOfQkXSn67EstLn8Uz8eFRHQXo4sx0dML+UvLREMtX6N8YXnXAoxIeDQ
ax/CevRCxa9eEZc649uvNbUtZU0+1SOF9AcWNOKBHhbunZsgSaCMoMMRSUD26QN+
z7t/o4UCHrW3mtM4CG4v1WbbVbrGI59HWogscMu1Y4znzYOUjTuVSsZI0+Loi6J0
3sX+rTjSwd3V1qBrgPF2HYPteiOGZzVYbQ7l/1cBgKAiiAMDPurU++GDnxVIJ18U
CCj5VWrWGRtdf4h7PzXDDGenpa0eWMhqPfwZsJPEQJTeMPLYHETNhYH6DJLCYd79
LVXMAJWz6TtKrsqeZYRgvMzJoYESZYTR4Gi6/0yQJGeiS2aHaojdKa/tHs6LRSAX
sH8S3cOkTpHwaM/zw+5Bslmiq4iJzoA7Y3PzkwCMqkSEM5bu0CV2c0OxXS6h7YjD
01noB9u9lgmm5lUciOwAehNVhpvtriyVEWBtCm6kVx3R1n7vlDoGSZPkdSmpB65+
KeJFcGcxos1r6KTkh+N+gesltkTyB5Qw1LQsKyIQoUYhC5yHRcYtDmGLLHf1UrZG
ozntX2G9gsGeNzaY4wKPetO0s2UYqoV7qyTWC79Inx7e+a4tvu5rRbAHFytzTkSL
1SlwmaqpPH2mUdid70t+789lmdOnKd2skqDtK/r0JgW9Uwb/G1gywzyNVlTsX0dk
YJb1xgGFXCX/46eXkeelJ2j8cN8vzv+dpFujj3EyBmsfxbarb/7R8lxdWwHAt2OE
3iO+U0IBYt1a7c3jMoV+/vrKvA/9OUQYiO1bQ+vX7ADzh889UT989NwHWGJ+ljqa
9ZOhQNho1r4arw1tnsZfvApUzIV7gScD9cTMDjpI/E4g14Nq4kKVKGay+i3Fg7U7
8aIFSqjeVvQASFvY2CAL4c/kTP2KOXhnqLsEoUZKK5JO81KvIzyHYjLXPyir+nB+
Nxb7Y7xV5LgnAcWiAaosvIfSaMSzDjZFmX2IrJ2ugPUniYKdQSq+h/JK+eF+SV1C
SM1ASZcUCBrccDuIL2WqEQ1EYnjDpnz+tWCSIxbJaVTN/6nHTpQRwWZ++ZUNo44R
TTykTwEM5vm0MEetOao16bCjODiwQ4R1NoycLXTLtQK5pTjcoOxL3PHMe7SH8EUy
p34i1VI0ZTyWTDdzpo+atNo4+VEUWBcP+945CLk+S/6Amzgd7H7/zsy7BQ1wJFdy
CwvXoTOX/6XNb5jwZj64I+7OX9fMmhix/K2fNhWJf+oskfO93yUJBjG+6/Nve93V
sctWLKpInTyYvf07q1zbxhtrT4V6jmsqmbrsLKyI9OWCr+07a7PYS46iKEndfwIN
iB7o1OEQFnzvmoyEpRZ5XlkdavoCy4udE90C3UF0PzIHownWGZKoOC3dAYv5MKWl
VtIJIyFU1yxDewrcwqr2YZjI8XhOsJH2HPsmhL05ld4Ab7tcNUzZKdplbgsCItnQ
yv5GYChcKUdDtht2dIiJtUyH2mp3lMRAu0uC4qIkspH1jqDVxkdgewV8cl2AVLDt
KBq71I7nL6gJw13xgSuPURffJ44QtH++BJQb7F5IsLuDk2HEZrjz1QmM+D9Z+spA
9ZCWh/V/2XNs3DIMwTZsr08OFac5rAfStJqX6Ca4aRSXHKgfUsPotc73ZypmYiZ1
iurUVhN/c4LWJq9NGInGQmXGoRcB1lv98GlWdykZkm1mcv3bdel+NjobOsQg4PcT
eI/qz9bZBhcuECWuDZWrxmegbgeOZe7QNJbMaQBk9BWq3ITEGGshnF1iplxmfAVK
pHnJd45dwmrXriOBZ82iizlg54dOtOuTLawPtmJ6Z/890n8eQ+jJqesgjziTxHLz
ZwhBpTreviRuhPzqSha0V5Aze1VfXHrMvjXLJ40mMaGIl89VLsWbxC0kAVFL2WGk
1hSnbRMiTdK6qZdOxoRQKEsTfSuR7XO43TcS2rQyn+wohT0jZpxQweMzChMipGvK
89XYBAzsGv4SPtflOtrtBcvd24ZCCm8TD1B2wU4osfaXU9Z9gUHCyyheNuZoiSoU
Q39pQpdQRf2qasfn+8yuTnziNvmEia1TbkdJAoV78VIeWQnoPKUEpd2N+otQ3w5l
Btqx3mXu8cfIOKnymBAW3gW/lAekRdRn4HUwQqzFmAx+BJKsbY1jGYgv7wHzBDnG
G8d8eMmbTT83fy/OnI4iY0bWvMntsbpWlQCE8acyBVv5eXd+0CJfSeI3a4+aAECG
oGkYZ9lxkDeAZ93vzt0kBlUzoygi1n1FcVIFRhNNKkok+2VRNZExAN1bYQ9b8BxH
uqyKLbW/FFDKoUFjTV5BjSm+u6CTnxfMo2i83EmHl6hFLYtaWw/SPdpXwEcg722L
NfEEx7v+CJKKWOa7wRQYR65k8QzGA6Z9PKYjlDeKKfdapysguy2x2Zin7otE5Clp
HrK5crF6H6buKAp/VcQlZD5RA4gbLDwDIqEEQRgO6sqwEAmTfddMgsAmoibxTifi
Zpmcm7WRU3xDprmfaiQcXEz5JJ/Hq6RYl8IJTq11I+y43E8DAp1laUGrGZrNzehy
zsbETSfDUweDrTBU2Blo6XidLIOcEqtfUKjLkUBOA+mccXMyj5P32daZ1NhAQteU
WgBbgpXKARTSndCmLLobVcvDY6YMWCNC5SSuwnH/rblNSWOH+J3fRXB7lV+Bb0lK
uQVhg0TVEWyCgElGT9irweKMrmxxb0xsxfRXZb7swBU07M6vUcsIhA59mPfWxs+F
wmXgAwgPrueyaekgNDoYITInjZgp4lXxmbR2XKBvCv2GsdTduoTcyJbKRtx5nRhP
1lGcFsyDiBD3ziOt3GQ5NaIcdRuklaxh4ErjwN/x7essIV04bRdIQSbmzwTMuXAe
+OO58C61qUfD4DYf6WQWyTHklyz3Px/s7pgUO77ofSr5Y3m8idlJZ9AgdSs6yTjk
rjIVY08U18gm6f7LxiY8J+RqYHLlqdnM2Q7HSuO2RX0ohIHeWU3rdnkm2v6pAqdZ
kfbHWj/LtexT54SlqEo7IzLqOLC+4W+FUQNslikMk0oLCnrUJCY5Z93jMHQ6z2LP
nuwLl8MqKh0FRYO6LUlP29iKpZQ9T0aKQeYrpiQKjdv59jdIqRVJbvl2SEFvRiu2
R9mymIfZYibq44EttNWsaKQxVAIlT6wvEIhzPao8krQLrcq8JDWZfUkxYHY/U6fd
zt8DFrG68qV6BRAnzwIf+4hsXmdIkYO8cD2BI8grGwnBFO9oVx1lZWH8b6MClmdj
hWgPij8+n11FlgOImmVFV5Gg0+c6dpIsRlYR4fTzBqFBhEZ4i2NtN1e5xtFOiW4p
MhdSYNVlwTWxLKynM47Mp0x3FsEBQf9aDyuKGpMKtuKZ1SMABanfOnOiXpJrFZ3U
3flKoi2+Nty/CjzepLh0eg1uMTsWUP3q0gW3xxZLRniRmy3CGrFTabCa9uQpDM3Z
8nw6RJZ1oOaFPXcNfO4xC2KjpYRl2LMYgkPrqrmwWTJaxvXA2/7FQF866aelpDoh
hON62GIV87cadY+KI1jYiW0R6TJRpqtZa9ZkZ5uexAV51OLaDJGgRCYg2lJ4ITWP
pAWIWKLNSlmE/2PJObgRucp9IBYihKEN1Efq4fO6mKB0S2H2DnUD6ToQebNO5zIa
IOxsJPwVf5DcXZS+/pw/5gvZHKt4kngGRaFxxmC2Qr5ZSi7SRQoLo8X88nIaWzhQ
Hqt6aZv0yEw2rk3lmdr4ZL8ObsKTnhICOZSVspsZqKbRZdWxkzFUWvG4cogtQ9G0
dUlhNqZwSC+LfK2JvTI/RTLTiIRupC2SV5+QuuVPajaa4/7tYQMU64nEQRfhdWuK
BcrKavX+2YSx8HInN+DnCBGKVSmsh3W0x0ykvyknCX08aIBiu0/liH9A82NuolCl
lFs1tjkTVjlysJMVI3YHBi1ge4W7Y/69v8GVuMg38x4CEwefEteGUNicYi2cmwgF
WDB9UWHYAnnkGNoxVkhdcP9oVejRJpioqduA1E+7PU8dmx3PND6IoPVtU9U0bLjB
P4phghsUQuj4I0Tv9dXMb7Lc2YcuB0sPCLf9JDn3PMxBLi7kWtusHZ0vcfR9LFpS
9e742vkHlKl3nuoxWqHNro/S5wYk7VTd0UpdLDRSEvMax72+h+/Sq8S3ltYnWLJ8
jpKVvM050wRcathanzEWHey+nt+uoBylQMKpdpNBGnGzIOMAY3yJi4vBQE3TkbMg
sdSd79ONC7pHg87/D2TgSNw8lK9Aiim0srhV91n7rlTOZP3Brwy/Q+tOrLIK5HbK
bz9CKREsf8JOOUGPu+B8LSPNYGs9FE9xc9v9sEvcy4/2wY1u8ytIouRmPhVZ90Xb
tX44dtsYW33c+4+Q3J+P9M6Q9lJ14hEBiTQHQsnoQ1+gYl/G844g0eMWew4858bC
QIIJCPSHES3w9NpUQ0kZqekqW7zYPybPCNO57AfhAh253NsJ8Yr4ucrKJKI8BYSf
2dWMU3n1n0l+aH1K1nCcjTeHrJ8RFj31Q0M+XNYHeU12zSgsAiVXNIUgr1/JkhDH
zRUnz2c9fLHJAaw5twRAt4MxajnGDjsTXlkkiBMEJ5nQ6JHrLwdzhUTRdl3CL8UI
OFi53ZMZhCNhB494OLNkN3erP77gVsw0Ctib9++4NtQg1Qir5rbtXKL9BLwbr+1x
m2G6UfuwX23h68AEsIEVfCdHxzcQjOmnGVWcYBAg7gPP4dt6BctXuGb55IfD8p0X
tfxQLsx0I3rH+JUFE03xy4BX4dbjE9aZVKCvTk/Fwlm/MstRExQCH8MmOtYoAEDj
OYgfe3UBsJlQ7H3H348k1FraBEpi+rP6z6oWQCI2Hvor2otWUUg9kO5bS7ilu16H
FREoHA/nDc12hDOp4zLSOsusZOB1HVti8q9FkCJJO78r9y4N/8AAoDeYDUiDXKNK
Ftj/+XfJIpCZyPqtaueqpRNY9l+fUe4IMlyrUizsLj3XSbePEuoEoOk1J65zLRU4
Klj7MFjdBTKKyFHtriPOwHBrV6/TF70u45HkwnQUms/d9m6veeYUlhQDG7yE+B2+
NkUexM0T2QsAMbsJ2dWPwVvGW+DsiuzaZ0Dnl3YySCzzgPf6FRbolL1O5WiIPXn0
GvvA1Clgaq5kglaSW8+rnoNygNNO62sND3iMjWQC7PFKOjkjCUyrISX4WtnOuNpO
wscFA/og7niGhDdTqEhu+UVsO8LFB3bW0t2REA0r7xKQoNgfkL8SWaspCNz144L9
gMWA0CcUW/ltzWk7xMjWv5E8V9wV95HrvVlaxM+lOe7vc0MBsIm3M4d37duroXnN
+qUY1viSJhcw7pZGh6DD8exXfrl4dFBIXY0VKDkGyIxHG+kdz80f6C1AY74QCB0k
oTuO4QdjLIfmYVxzMW3raKeJu3yNdeOdXZXbXmFE0H3uVzh5T/bPWBzyX7hs4Ods
7CB1dclmDjJIiP0dVxEPPBlHjbOQVSbZR/j8t1A4oEOGvesLRmck+45I1Y2bifji
n3EQ6FID+NwP7u3oYCWcj32kLX1AqNm56EGcK7MPxI3fg+07dsaAIWiBcrLySON+
8xWq1WLALR4nqEfmoozxtrxV1ELyDAc6UZJvp5SlMJdklo7XWA7Fv/Jcye8uxwvR
Dg+bgNALq8P7vjAGnWRqlE+kL2ccWo7AFQlnEQUJIFmK0ZTZ27PHHH/kTVWn0MBT
W3tyDGRmK7pQNGoWgf5BD1uWcnsq9HiSdWjUatDn8TS3EtziINmE/eaFyVJjTdLm
HmjYoOZGQ9FHgGssZyCQDNLZK59CLUsx+GhU50YVWDqNIQnvpUYcHPH+bp00SatI
cG1y1Uqym6yBWSBcXRcgD2y/Bqt1+K0MOwEURC1MXwgPlSUNtQw8eueYt2kb4pN+
ZclRm0EC6Z1xWOu5T54fbP4rwogtgtyEusu8ytFW4hCZq7r1bppISlOeJISN19a9
vbiL/OY2eny0+bwNb9ArKCxUe1/q1ziOvMJAbxZBAY10xZ6egGc4QyzbYXQEXtsO
MxOSDVNtvme+xU0RcgkqEPqMPQ2R2fCpDchoOgE11y6NJbajyX981KSltSQ04Dd5
DJM2Pxl1YkpgoLLCKkjtfK2i2ASae2erWwje1+/QS4fIwhIsbnsNuq4gCGk7u8oZ
ucF+UZH/qcjuZD6+UCBZ/NqgO+ccl5N2t1XLnsTDDnRLFDnxROAe3rE1bnk3gVds
+5yGxMVKMMJao6uZQtiLPa8tcAfgEBGcHdCf/HFr9bdWJWSevBfCrCtZ8WWC629h
L2u5jqQkeXCiE8M63so/jccdD7d/+Hx8QTZWd9ULX8MqU17zyEPZ2ei5IZLyEYiS
WDvDeqTH97UN5/CCvqaXcnXBY25FWvAxbjf9YvZKfJfi9JXsjZf09uzajfvgfpN8
keXbCDkZb1FMH4HdatTZquc2I79VOtJUdpensTJgnxixiDWetM3s7qwjL9oNMZ6c
w/6B23l6FcWdB+Bp0SbXF0MaAs6mdP+3DrueZGUhmMA4B2obcnK2U8LoniTMR56t
pwdjwZaWGfx+H46yWLBdnYydH/pzEre2TN29dNzW3rLRzRVJlDWGQhk9k1uKMndy
bz5bVCgYgMRJML+FsKM4bzWk72hWmugVg67nEJc5Aa9CHHJxc3y8Sb7cQmz3xW3j
YAh+iIPdBAmlxr/rVevkXrgTHnTE6H/qPiMOgxn2ZzUS2WToMZwx5YvLCbm6AP+F
stHD8BTOvaP5hX8HqFR8IcH3zlKdQrAUOU8GSONFp53nH3Idha4kfgLih9I9Je/q
VlXDM5WIfzUX5V35nGzU1dA63icDC3JlCG+N36HUC+/nZi4AV2IuPQzhs9kCmCfQ
j6FVc43RGr98ZGqOgFCLfiacAkxTVsmB6SZdmvV+aRTdwMvjd068/0LsihabGhQZ
lkdJozoHgbRYp0+QHiRJHtHB9qp3a7Rt+JoKXcTaWb8NWboLVyQbEHV0y5StAbQO
2vx+ON6o4dwIWyKVJ+KcYJWj0bJu3Izc0TO2vhwxyH49EGSBYl18Vly1JiswZzs/
Vtnit1LKcdbhUuylrpmUm53E4Jp62QqQ8jy+lfbE6ro7g5N0Qb72fDJ5W7zR/Xti
CURWs6CQykDlk6VhYfUA1UcC8v2sEGX4MtaQ/QLVR+0K5QoFwjaxPK4Eq4ulu+0x
a/cV8WwoNfubrhruGlcXN6WAZzn779fwidCwwfMfPv3PmN/+N2fM9+T+5a2EBDQM
YzfhsIy5qLazSVHIiZ3Pdb6IlZDo+UtmQiHDgMHduCwbilScqKXECLLJ1ablfKS9
Q3j3yA6P7gYL9fyZdZfWnjF/xFfp+3OycNjo6Un1mbhZaAOF3EGTRTKUONEMu8zz
D29z4G+yQR5mHeRqtHuKXCa/qm+9y7IQcTkCXIFguC3SY4j//yTDPnrCEFnAB4k7
qBgWNHfsDNAxBLxMyufI4NnTsBxhGtYEvJXZt7w3Q2AaHn9lmE+7CHkMAOD5hakv
eMnfImfjC6nmiSUzAaJzVKf75pEjj+MWKvsATG1rxEZSgZRsKdybWIAbwkxiszxF
pxL3E2W0mMFf0VrU59glh3N251dMIpNSDnUrwVfUgfhNbFY65MI2PQTYIxoEcbU5
3rRqz+ncKKw8iPQXPg/71S5TTPAubJeUevXqs00lfrDD55asg1rm7B68n8yzNVR1
sYWz05opgB2xVh7U0f8dyTNccjMFyJg+/d4CJwNHa15CqinUMLfG7V/OOlJzGLe2
EonHGV35+bJEBybgLwF7mZGeqsHBuEIahpqcRuORQf7Vqj/3m0PlvOD0+jUOI2Nm
f+Pm1Ml+I2OcXoqUmCjqqnFG5WAYcOHpxA/mkOGsehhAXwMSEQsLW13JqOqAAi5A
j8rE3W4HGo2mLZeMUnKA3bvTHDlY6b2BcPU9QitKvhVE852QDl4sEDAFx64ZWyHS
zmNZVYj4vmYiMjjEU9mrs8D1dE3m0GYOqV7X12BeRV9UauxPpcn7QbXL9JpGcyrz
2urH3qsRELgpFi8SPZC3DDaVwdpv8yFOgKS8ESymDFq+MWDuOjADeU3jcnDaiBjm
ZmSFShbWEi/oAQzgVu+Le04IdL22cOG313mxbCs3u2wj8cFk+8kzKnUom5iJKMpK
siTJuil17V0OZQPTnPtu422nIrvEEi8dol3DfnBEaFBe8tb57cOVNCOuriGnj1Ho
FtX/IRDzY315KP6q5xoY5q9MOpdMuB0YJjB3SPBLKVY7Tx3f3JodfXeH8Vb3PbCL
N1e3bM01Q15GnVKCcUsGPmiiyUNUIizEYWFalTUt7pOkJI2zYa5+oZUxXtbenT9Y
ZD+nc2J3pi0wjjJ3wTvG7dAY8gI5IdtP/IeYHvGB6MzBOmCqHEwsnE1O4X4F7GiQ
Glv6fQHGrfXrQ8Q7UEZSAE/jIp8wtgY1DC23zRYJ9DMrdA+XlMfzpGRI54+6k2Ot
bCfCjIPxaNT7IfhS8aJZ40OsLv3inWSavZx1g9Ikd4f2Os1odB5pWuKjmJP5q6X/
mxPYk4I4cAaqvrAScu4Lku4y2f9aGYrBQ5NvjH5n8OzIG1NUoi7+JweRbHM3Y2AW
9zn8GZdg4HjJUQXZ+PD2q6WswcQaXQplMqRovnWMTeTd2tlaPcXOo0D9l7hKknHz
wKKhPu46Za9VfHQSA5uTa8wtj8KsKvRcoj8M9U1T+mGc2NGestVWSg6hjaToDwgQ
5mHH2ze8097GgXJQbtRTlkV+IGkea2fY65WmkXhyaIhnPeqKvJrYl2dQrAdlqjdv
B93H6aKGRlYkViWctIgBHZDeBOyyNjHPNHzSlITf513Xt8AxnJm/44AgGzdXkHgu
rmufm0kc5e2/lYB00kgjUloiNFXVGzf+5cCVCzZ8hkH7d2iPejcRK4V/tF3LPQfE
Y/Mc4fnexJEj2KhxkTW05u6v8kJAMp4Bx6w9WSDU48UYytSvCKVPcS93g2c783J6
vT/m2Sx5XhiIKeLXEEBXNGL72ggH2OOlrrGjRmIqfRiZ0lTslWa+ycmiFXjIH6ix
zP66H0i5aXI3fREkknzcX3zb0Wqkqv7Ujtp84h+HnuWneFEdt+3wRbbPjlZu+vkL
T0L6V8t36zCYd1S7oQWdN6P+TC5zPjUREvvqP4w7fZKLB0mYvaFop8nMfypGOLdu
AY5NDL+zB03U28/dAEaCppbFifKacNaoGXdVXvBpF2N/QA6l3AE2Paai165HlbBR
dlxHv9IUHfGn6MEOBXsOCxlmZLQY9x3fCgLGQZypYM9f5to/gBy1AYUv12sS0det
FiIi+sh2FX4fvrlV7a2OWzeJ9WFzwqm8U6Ya8dGn2MWr5hf7TCk+L6+1xsCI5HP0
ieM0VqKZv55fNV8iCj2wcAhvtH4CeJPmvgH7pVQ95+RchOEVjgQ9hYeSYcgoxEVu
eVkCRSOLtHM8UsJ67nwWSa4l25fEWnTVYMj4WHq9cowa+HS04s3VXpdAZn4qC9QR
8EsVWdolZ7Cd/4MOlouiGfE22rOWilRJVVL+sHkIhZQyxD8PKAqMYoYzhm2zR8aK
mo1HVu9yDleiNTH/w4SP3f4tCKdjirHYIZQi5BiBZF2qVv0nx/QXH6rWWy7i36kW
zn6lciBomHEhjKtY5aQ0snlkFqScJL59+yfBCWgCnBajgGJ3Fwe28pAkmvVnL0cg
7s0w0FKK7DmY80SPwUpWlKE9q4WPb8J9rnu2oxgLOloFM01a37tzzsVnZrAUmmac
WkCtycBuZsy0kYFqdzeZxuw5Lev60JA3XuQ+6Mm11v/XLmdnHx+a8SiS01cyUnQM
UMQsKB9z3jeiOyWU6R83dotZffmW1t/8xhdU3H+UtALp3bGXGZwr6W9dYgODkoWX
is38MZms5BC7e/M23pL7wpKBP08ig+auWsMe97zz7XR7VBjcTIltc0/UtaYqPs42
4+8VuUz4QdP7BrXuEmKMRqX5L7vb/AYKi2LNqTjlimpBMWjohQROyAvsry7+Vvza
eNkQL6F5izIv+lypnlD+LXERMCqrSs/ysyFaStlVp4QxiBFmJ4cjzFAYPst4N+ji
qfSZLSdynoJR/l161zYy+w/WJo9fC92tDB7aF+bPEapwBSWeuEKhv5lSLYevFXB2
PwuJYbsIcbIz3wCjxaI8ptqb4zr+zxWPdPnCUPG3ZBf37w72+SlDWsCDhfcBQnAp
1KbGFPoRI2lXr4+XjJLm4CAtCu+btVCylLGk9rqXS7lmRffMO/Vx9yWFTQZwN79A
dFee2rC6tIx7qigydbgDDU529atYwf7SEq7fU5SrqOlXxNM5U0Pf5DELCBsxBYgK
pwRE6Sr9ZwIo9lqf1Lgb/rAp+kukokUDYq41X76GFE19kz8CDTPOYpi36o3jmH7U
YLzML/x/TCsxjWLPZayM1yfcF44aXfq7YMszR8JlvOzyCYWN1IAZqJ66bghMWox2
4mkbiRwJdA+fd+YoI4qSUfhKVQmsaylurfk9/jVI1RjqXYjtB41KEFZ4Y5lx+kTw
rG6YlK4HJzc38hbTgWyQssgBdl4GqPRJ2GJyjDE8NqcrqqTelZDOCBkDWJwzrWcr
tyALbKV2vioK0kNcF5Fdy6t1CM3bkTjR4zv5nla9+xTgUPek1powy3J1ZuT8PrSr
G6ARMHhkrWbg82RSMmXTP4HLOGQVQvDbo4Yt250Q4RuwWdOQpHdKbj9z0DsRIJpa
UEz416zStAaFZfGORO0x4BovTYudPbLTzHEvUEEEygI3tk/juQAMB1L7XCpzkiJx
X705D8x7WdnA+/EvH9/Lep6RdpL+Y5eFUpYmBfxX8LreoHOdgLegk9ecOoa3zL2i
mmArZ5MFZpiWbRh4auBFJN0xsWesna2cNA4ZtAM/ULMgkEcwCcpPNcO9dAv6Act4
pMUjUFxX0f6WuAqaILodlbrQ+E3YDrv9Auoq8vxkRq1rrN+t4kbmDQ6utaCc6SE5
S2bECkcSXIhkWUtf0XkOwT58K+J/vP7QuuziztYLk495U93vIT+s/WonnZelm8dw
Ib/wZ0OvAsZpO4gtUW+xAFdi8Q4Xw/sY5SBeti4AKpm35zhQsb9cS9W5Uo61Pl/y
i/smIxiQ8qxWyU9L9BSWC73qhGywPQJlf9Eiv0xWFmuI6+7Y/VYqK6HIZbbFzGAu
qBpchtWiKi9BGZprSr39rK07en0hG2/dxL8wPk+lPAVfVPJ3QE9f/32pjoYCdi9L
Ziw/nA1tcF3v6D2mHtBMNvNiyjzdilnplqZ1IQNQVr3tqTqzhI42Nxk7wg6gCovP
uf6OarZWC13Pk7m+PJ7z9Ff4ZRxzrQaHIJNcqgje/n1RnlvlUOopURb4NbHPKpqa
4Bw3X4TKHS4Dd4zKl4RKb6+6+vwigU1BwCFsRTC8Ihr16/qRYpMPOnyKVwsRu2na
nrJszwvnF0dvQRBx7gsZae+EN7vt2ULufbhTGFleCK+6Yd0U5SD0pesAXpdkA6hw
YNqiLO4UxZv1/6BEInDdyigJDZCX8pCA56GZDgRoxEAf3cS/e9M1KLZmvSMUSGZ/
X/uUk7TG0V6Y3TATxgyqs/oULP+bV5oroIzCD4AtTM3lxZccJ3S+YXSw1pg6bi5h
ZUVW6viuzxL+jAqCSr82yeR3S4/rWzCHFBZO/tRRtGUgB/yXY0sCZtGJfWXbHgK+
vh779YAT+XzLmhBZWZNUmteL4SnxrrK3oX8cx88HDHWFh6Z4b3AaIC9+LDnMn0Ii
Mtnf/CWsEGSboNnWLiMHPag7+PjmhowmwWh3d7gKDNOH/rNc1IWbwo3rxfIsIp0I
6/qSNx0t6ZMg8I3zLpLkXrx/JkW59PE9wTqqs/eBkF0tbDwKgh2eVKhk7Ve3hpjM
dvWI10F0X+0FM8E+c3l9qlYh7Fv/8Nnb+RM5gH2krhmEvHvQAOnTkOctK7g2GkJx
e8LPfacWd3mJZeMWbpVybnjDc5ueIEH0kZZDEOyW+DxRfKhqpsx57M28A1SLFWNR
TVOr1lIN9amZ3JTROmNEcKjtFTnIJgupvQGL24YhdkUb/7otbjK/oBaijzY2jqJ6
JmnjpN8p6vNcZTmlDcjTeZ+9qz16vEeXDebXsvqzqeShMke36MsyupSSw9Iynuaq
FvbjPHGjceJoia4cXtkiYOlHlU7Z8WlMvsXv4ugwKfNBVNfnPVtANjF82IPjX6mD
pzZY3yjiX8EOIamZZVKJkhGv5yXrTgSvoMxd0QxWgP097mGi8WSF8gHM3GFvSOdx
wxkDqoL9gs6x1LkTBlBGyFN1QjNSq0pNlfIzUztwZXPRKnt+nVN/DztzKq9lu3n8
bWvp/MOLoPCJFaNy5h/udB0EqEcoT1PZj5iZAqyPSMsC2XZdai5pdtfan9Z9BtxZ
SS/Yw0oRFJ/EfMiDLBK/0TLrdQdnNE171jozLAZj00H+IYUsj8u4jMZ2tz9Ngo+x
BUVatKz+1f2JZvZfzK4CKSe2Ug79EkdVCZrhZHznPSwAVwWRBmK4LOuYcz9yGHAx
pamK/I0M7wUCYQOM0EKlypN1KC3nK8+Fzid7tHt87dpi0CBFjuR/T+IQ4lSxQqrD
pU854mGqxbsYIbJut/nwnWvtwjq4EQe7LP5/Ffz1MkakX2AzCinv7qX2H50OKmac
3DbeyWP2A8itCp6caPwJwyv/X/PvhgnTweaUXxeumvB1z1syylm+4lftCCwZi/PL
t87BiwpwDak2lWpSgxySun8I9RTHR1mCGYtt5h3uolQEPPjpqsEOoDXLd+DsqWXo
GChtvhLXXqVKSOy8fHgaEMOQY8ycvzZ7LlkKMYLSxJyDdSJAIZDSugkMWlBDHuD9
uYAHd7/cxdrwbUuJTgJMo7IYnEBEU2vhp+4wj9+FSo4YOjRMroB82cZK/Ud1bGE5
zTA9ALlKHfMGSnRV4+giu5IYLr+/bpTRUULw6MywsObSlNXjKMPq0RlaTIdgXxIF
BcvtgyQi7cb51dZ+tdfasXxXyZF8utPgmIRTS91C4NCglV0TzrTRDmUfVMtSYzgT
vAK1hlQwblECpui2NZd7HRkX73456sdCXXNslqj5b4fYII7QK+cZznqYjZHI7egb
9vXHRTpRX9s0I1D4+7T8YKQ/M3lLss7BQObMYTEglTC/sSgYJWdyixdv1In+0HXU
CC6EQhpN82FLVKdZ2O5gt07DxI9VeNE/9obCVo9GAv1UkqUMY+QXf9f3PPyM0K2Z
+2AdS76sf78fN2S6armaAyJcKidD7H3ZzIJ0XP13lRe0yYjOE+tyQxg+gDZCyUEz
E5R7cOUp2qGoPGXlwURaHrDZMshtiGsas4H5CmhbhlWb++GqD4H5yIm0Wez1cXx2
27v9gODp8cLGiWAZ376Skmd+FDdk6JzzyCgv6vgk5TgroxvfPeQhUYs9FPqKcCOP
DZZ2suOlJ7LhRPnY1gULkiepdOXsivTH8Bztqe+qeHhxWVnwWltsHvCfTX6UAOi2
uXH9nwRaNTvUj0x1HvnLlbLR34YTUN033r9oFItQJ0qXqDRaOyYYqZQy+OEIthSE
dR+PClOw+t4YsruK8HVurljSnjLzd50Wqf9fTw/30c8bkRDpYnMLe5sbK3/3qmkf
OC2ZmvaoPBrx8/lRj0Imnd6Z1gqXQlL3Zy1uAVF6vnCNxXPO38aCwUZCnbbBDqwj
v1gaxZgJ09PK2g2jcaO8UWOEWYVMrqPBTY8P46KKdtDKsRoDnRUYXbNoDJrO+v5v
pxQXT2wfQoeh0+FbbRt7IZvBydsSYMYkhQl4XgUoPst5ZvUMvmdVefc1eUfyqgA9
lYbZ0Q4ZAgQRfteiXlHlvqeolsvigWJPA8K0mYA85ga6y1B9GoHsr2HmyfaZFkZU
1zCoEw7ECQDQ3jo4pYJR2GNt1cW702yL0mT2iaKR4VJ9TKATIhwFnMeC4QVmHhAC
QE00l6xsCdrFTj+vxbe48VowAMJIbhg5O4/gjYUGLYEOFFY2SWjDFF3vuivsOn0W
+PIniuaqM8m4T9/+Z12KndGWfmZJ6mPeoPt9SA3xhFHuTCZ6XzoEcRdr9OPKEl++
G7e01SKXM2hb43bWMJ4E4+42bNa40x9O21MunxxqM+/Uig9O1Yo+C8PeeuQoOpbT
i0861t3SXyKdYXJGRvOfg53+jx4HQKNZLBbv0vyP8oaezZ8ixzuPAykRJrzKADli
KI1hdzBamgUR7gmrcNVjUSa7Y65Cv/RAqevpEsvhtONvV5LSZ+skXg2tCcwAJYuK
NN2rtS510p7tx29fnoVgG42Z70b3YKOlML63Nok9NA0Ap1tSOvEsGdkwogk+Mca5
LetFFQPDS7xlj0NOC00UMn4O0/nsnWvwufdckZIYZjFoY4u0LKin81cYQYSa1Eeo
e1CAqbujsXpLeWURVXaSMGJgJotiJlyu/51C+CSK98Wd4nb6UHoOXCRqJemCssaI
d22cUDJPq9HcbazXL6EkJ7SyUUPArIOOzmUuubi6T4kgWe6h7nedE+i5d2IpgJVR
UZMqGh0Grw3w6WnRF4rpdNMWoywCssCFUcEHUQZK1z6Ig8jp2/BHDroOjcpczXms
Z6/OHQC7AsJGtFA6kSq6PiOudVjNNLuburYqLRU4bwNvJ4puNBUKv+ucD7moHt+G
bulajUy5LIlP82lrDDwVmK3Pa7fzfCOB84fmMM0G1MyQZjk8Rbs3zd/QcQ1AlPnJ
jrjelZaDkkmVT5Ameel4dE79/NAMpk/yFVRAj6pROQ1WS4w7bFsTuJEVfzS/AD9C
pfxFzWo67+PA3K19e8FbLGnJT4AxrtGqk7EDEty20fdIZaO33/oC0Zi1uDu34cU0
mrKk04TobzKW43eJ1K5PK5uCsmJa6PhRic3RdrP6LEHASPyvVqNiwi1EvzHt+CtY
XEE+RSmoHM39r/Ld3XgaVgiFIX5Jd6K0m3B84bTUwDAQGtQ7nlqgk1Eqk6fYOSNP
LdRe+rzDXccoIIVIQwDjbqDZ/0c1TBsiacfTKC8lhFeAb0RaWKdwJhudaXiVsvy9
MgY03yCLMiznY9YmobjnxtpNA7K+vOs6UehXdedmWKGw3nD48/bOXlUAubh7mXEL
S3Gey13F54bEzm0ct7lKWiC2yrbS96zuEl2zGMEDLvtCWbzNCciS7ESxrSxZvUuX
eHcsSli2z8a7NWamu0mvB4Kp+mBBz8Z/RSSXiE4VK0qN5GoGk5LcMKafSka6KQQL
PpNKslK4AuI1tvaMMfGxiAcljBAamwiK/dJLgT3OBXk5MnRutbReByoyA07HISxK
HDohE8y5oaswjDUwL25ouTciVcZcpOFA9FlwX7UZaWvSbux0TwwFKyM+pIhXJivW
3JJBkG3zbRAkOIDYs1CODO3nBnOI7B10U+lSiU3KP68efTNKFvO1xQ7ZuIM+ptc8
VjcUmxms8a8PKTr3anxDWtZ8E2o3NSdNlsswrQFA0dGn3SUYpcldWV9vJqeTvthB
ibCuMAmv1Nqn6NvLZQdlQ+A5bsS+ZmqzsgZr0TczLBHBeTbgZAE7+ZCdVBLPvrsT
DALJydkj5f+lT5EBaSASN6wsSZTMI8RmiXDn6MIaRuwJ/dgj8JM3vq6A2rS2t5F9
7YoID1itxEFu4HbhXARYCLSRODw0F+yRc6036O5ZJVbz4lr3uUGp7LLeJ+nh+TA4
oX8HocMd+sNxgKDNlinOuYG+xmPwpkIQQLoYKTV6qqnZbpYe5b4hjvKUPSyj9Mgn
hCNUoK2eunMnwef2BzixQTINIilBkTbvRpOlhdyiDNVCwhoCS8Evh1YzO5TkS6kw
sUFGnVqywjf84TG1vDHMKZ3OyEjq8jDlO/k+TvEBR94IHdd6jxCXg8uvr00jUSKq
M0fKfYy6O/2Pi6VBs9X0nJ09SCUk6R1nviu0tmBOBjeyQizTaco0MNe0V159h4G7
ONfmwir96nKbkuJFSOxVC9q1C9jPECu1le91FtHx1PB53jX/R5sZSXtv3NGuHTDT
W6W6E5Wq0uEMmEZcMaUAu7KidkCVj0KFbDp+kdvB1ipLDHs72htBBCyUlclnMXIe
aQ1JD/bw71Fp/gPjD+G/E+VJH0qaSeJkJ/W9/0GdkoR9nO+GzdsHk4xt4i50drHB
UOhepLY+TkxxZzzM8PXFbopYVYOwuYTky95+uZlw7jOBwpHFLG/S82Ax0dFAcmiD
mADZBmZpFdVZVMuVesHnQ3H9swAhTfmHJv8h8I1oX0RCB208rqBRBeSjo1INz4uM
KI35YK1XC0sqQ3zEWtxww9MSQOMRb9E5r9Qw0T2sU1Prsm4xCxiBQkw8uniST3R+
Kk+kZgq72rOysrvPGqcEMDqxzGHDJ0LIazxcL0RLBDm+3MDVsjokca3rWkwRm3il
39lDMV0iylpoGmyLu7EvWxz/La7O5OtDaelNTIr7oRYX3L+Dj0P5thBJ+UiZEi6t
lQ6APWYRZ5vbeXqd+MU0C5aKW6hYZV4hFht0ZXlgGgkkXGIJDk+Af44WV07pxBQE
B20JTLFAt86D4f1d65hjKuAy2oBDBiFq8fVVHyYU3zlOttRCk00ASUWX/MT0U3rX
k9ZbEkX07FTU4MFpa0o0V1s+2N7kBtIujKAWw9/KJaqzaBluZb5lxlo4f71LORNZ
ypFCzRd3On+23nsFnzxE8WN8lzHLeJ/jPil/wzAyNPbdycMdqvV37aMynRtn3TCc
KBxCHAIFxAdk8Z5NX9ON1HBtfOhOuKJGdEYkz5BpPrUE/EntzPtgS6sb8lZQMmzy
afPZMX1pPym7SOi8D/f9rmZqbciu92hbxJGRrkJN6eE0bexgjEoBuMikVA8PrgrC
U9gDp3lTqcny4geFDoe+Q9qGM8WsYEOLwqPPzKJ1vmhVQZ3e4OR73DFMVldtI6Ji
N0Hh44+evMS0Ag6kPN3yoML9mAw8Ex9R+7RyQAIARmH+0PIxm3oymMYeuqpJRK14
Khhwg0UsSpUBLmiFdzfgLfqOWg+S91jnrSG+OOf0yLy4eTD/98ORFM6AB+5gPEMq
d4x9az2b4qmLxbHyoRcemUW0Ce/8yLNecs2O+VnZiUV6rF6bfB6QyTgQ1dW5Y1w+
6F7A1IrF6y900CLY+5nAUZ2gRIY+AFh3l6WnO2aiH9Wg9y4r0emQn4t8S/EsjlYu
lkivFDQRAF4gXgIiaBsd4K750x4gTBoCkhSiSUQt77njz12L9ykJV9bBmvUXVkTM
T7gvmZvFpc65mxzHAkxZoSIyWtA6MyWwwSACO7d8q8LAeN80lR+6F5AoHeEoCS5H
H6ob7kiqWATsjGZmwRDr3fUwsue3iab5yYysPCNEcMj1qWbgxEOcV+yku5X594su
Lwyu4avBTZokj6LTdlvQI9C8D68R6LLaz1wFZDOkBwk96Md4cFo2FTaY/Yt1eUWF
CQrLnDekeYS8ScthnM8zt/79UnRvbjWP8dlWbncqenZpHfKku9VHyX7OfxGsdPfT
CGTPQT1DlBve6e1J/vmznxDoCdZnGx8/NJZ2uc0+C3GsWXhgtFZSVmcoF+V3TbUE
BuKt6LHTVTzaGGmVyD86dKC6xsxhmkNX0IWUTTZ/OfdBeEhRYxcDczIaEox3IpMK
CE5B2Qeaf0rAh1X26WVSSs8qug1Dz1exRlqJaIwQnb8qdJH2ctwq07uyZv75KjuV
x44wblMnP9heWS7a19JIGLu9JsTHE9r4l4vOPvRBZjqXQ/F5vFee0vM8/emXkMB/
yMT9EItIZ6RM3RgeWu6M+CfMOHw0o9GfLz+dxWVQgKsZJCwZcLGCzE5SbWMWoTep
wjnUqD2PDiQRKv3mHx2RE7UUvKeeu964TVv0ZFjgW6ljCtZhhRM+S0ax0m8qHKG/
m82a2gFGAXG/NEOKn0hHX3RWX3rCvifOoJzwJersrCdz2dAZ4/W41HIVwSa2YYa7
DDefBpVHa5gMPZicLMAIu9n9Nnp9flzITdY690YAs7sP22Zxt++RglCpdAWn8lt/
fHkxXPnJaJctSAe71TkBN3qgNGmWLQRsAA9ak8NTT3Qr+cHD0s9sBPc1z9USLhzv
OuixTRAg9Ow5KPheWfPjko0exxdSsYrCz2VSVasm8M86XxmXC2pW/6MHC9QnRWvV
sbhyVBRSoWj1I8NDrN7nDE/ZsNPIiskEBe2Z+urQF9YIDV3tITwIGL9L3xfRnGOn
v7FXF/lh9TJ+9qSWGriuO78D2fAu5eybY7GnpNIqtsoqwZyvwL/5HnptUdV7+iy5
8itRk0OKafpLGL07oOzZzo1WNn++Y3mG5DVUCNZBMDGhzhrMdptPdeFm7iHhkQr7
/OjG7AJgZubKZCTrPhOimBWIGHetfMgiiG5zHyvAjfqFA5EaoZHR0IKGE07c+Rvy
uiuPzad5gE66PaeRjiBVS5n5Xb6k6V/uDTPCd1VrK45BgkefT417ry2hdAHYpEhW
efPYz13oX7qG8ud46XZbug6oQYDG66P4nWwxyPtFIE35ZkWer92sKGBVkapgLkYq
NS0oi/zxytujxJWXtyPzOGADo7+xCIrhVIATwvCZVqqnxHgaYFrH3645FkpwbJcj
S3GlVnQ04hlVvgSt+KYKH3BYboSj4mO0klP4XSJPeWbIdH+J0NqudiSJ5si2u3s7
GsMSvvdzaUVC+hFDwJ+herlenRqsvEKb8o2s0BWIMrgRggbR2BAAIlUaGozVlbU3
XzwuluXUNEYPI6f5MJW0Fvwd0/Ob/9BRmg3ukggClaWXgYiY6Y8cGUmzPAWlZGw3
Iq3cnp5jLobf+iZcWW/x/rWjxL2ANDUchQyVKZyWeeQX1INSybbfyOWBuEHUIIco
KQzTRZnk9L2V4P8vJOCBP/qHg2vyxVGv+EzpZQLZSYcOgZewfSiY4LFgs4XapWAa
/8Rf1fJFdHCOj6ulsceh9TaI0Jp1Ps5VfKuCRKdF6E9+yUJ7T2TDJbupExsf4jzH
QbH2J4X69JFv3R+tSTibRFvucgE0jfrG4pNqNirVGsyfsVfvuqLtuGuOSqfAh5hd
o34PDnJvNhCR5qUMUEhOx891hDJ0PcfG510clkcc71X01NnBSUk+RreaCB2GByDC
PzOt0+SSNW6rnXxwEw87foyZ5mCwSakpv6wb9/Gr9FSkzmiklV+Bubcg2RHG4+Fj
F0S7F/jJ30MBsnuV97pYn+6rROo/LIiVCUd6X9aHSCEill7HXCmC+hEwRBgui/eS
nuNfLvUDpohTflEVUJColBzjhOUO/1zO5zy1+CVihZLhh8JQ65vAObneHxM3MF31
pGDquwJgr3X3fDf/x2fGlypWFlPUHyv7Ibbh83W3eVUKnogMZYNXX4wGChokf9iY
GXpb1q5YqxH9wyUSe+9Il6Nw6vO4GxB9Il1KxsJ+TYQ4rGeaMwo/crT05kqMtagX
YjW+jjbaNjXkBkoAR1VI9Hx1nDUro9/ZH72IxFe5BlEFyzKkKsZ8w/8Hdfo7q7YS
wXlshL602Cbs36MblzVv4kS/FqTZKepCTLdZY9vPnjGUS8jb4QT21qGJsq+n05hi
zXILVFXv+cAjus1QX+uh0N8y7zDnpqxKjXxG1kw+W9uHDtQh1lKq8Y18tVS2+G4+
Z3aksJuN/lAGHlyUlPs7tB2KwETdgT4q8fsmWOm5VYZwhbKTsIuelvAuulhxk46i
oL9/Gz+H+hoMRyLFR++svNOLYNPl88b1cPwYAIaU+0ibg2rM+tJxYp3UL8CdvcsF
O6cz6nfbPYtjeBFiAYA5owtw/oTOYyPeRPzkqOyjLSk6SkiBNu15Ig0OYiGv4Eyx
gQbcYkaTyVbCPSJva6iZajCpdgqeN79IidFe8mfJWlzG6ufbwC2XPPyXN0dVgUu1
frEh9PlpC6XgnaKK5lSGyYn47KFrn367pBcaGfvTfRp6sNFdtJaChFbHiXxNBNkP
5q/Y/dIZNxQJJwteQAWqOF1GX4r+4z/cffg5xFhgGPphx/FbHqyJgrlZ45eI4DQ8
LxWf3+JBcAsLKxANmyNMgUnUMl2EerhdNaHgDJFSgiK67i7jrEb7I+nipVZ0RJTX
XTY4XzFp4UqMG3SCSTvh8nkQNuOVAZrInRHC3qUPqq1G5zB/tLREsE9aklOVpHO6
OmMTp4UIH69hPM6KdHr3JyqKnRNz6Ev2tjQfeF2j9e2jlCG0jVlIGaREo/s07bMF
lo7rJd2pJprjq303b620GhnqZCetd7bHrp5B6XogGcTeaKvyTCw1ZwhnrOicMl59
23VV2o/xUdUcXUANn/0J6BdewLK5/Q74pBMDvxsh1sP52coZTm8TXdSbp+lPd6is
+HfgG3TZl8lV8RDqzyWtaT56/+cxgA1ezccUxu/n27rTXNHSAACATia/A3sZd9Ao
vaJnYD0vOQTmupwgumcXI8A4WrMrkcMEARc1DF6f+H2q0ts0wkNP30xJiXSGxYi+
GDwIIBPpA3tnJoJH3LCN69SGZoA0MpEzDPkaWOalFT5w0juP+y2sTzar5KT15EAn
ZlF91/CrEMVhRz2YRUjD3OUJETHMt8RdN4akV4cGX9BVP0aISF/8Mt7HofrPTxxv
nOw8Qz8exXDJ8TXakbE1WBHXYs14S90rpp53aOr8NzE7c9KHPOQJ9gFhDMbGa9uM
nU+2FIDM78q3ct4oyhe9OwziXgtaPeMhasM4VLTuZQfuCKhyLVV/SKbGVUUwBPMP
EPkO8ZZEYqlHL8inZJ0N5WQqw7HBNTyswJgK1ALQfhN8dKegS+YHpoAj+kHn0Ynu
+314VqBnJf5M23ypwKNlyXzgud/FircQi8f3QPdMD0P12Bv1orKIYRBmo2GbolqX
valJjNA5TqAIC4JeVGAKEqANCMz719VsZLqF9GoX8nsxvknhEwaTWuzDuHedh+IK
oXoSHEsuhBIs62ZG4iQj68FnaTm2eROotQ5o+Mz6kwEL4wwL/Vs/KNpEXDjibQFJ
r/Wht6PinaHMdLlqKEZO18powgJetuW1y+CyctyQkNthDYGorsaXvQgy+gqdl89s
Qd98EWXzD20OIXsY0HC8dDr7QkYX1ds93L+Kvy4u4XlvywjPYRxB71qWSyBaJNvd
sc+UZMuxNK2Y43BNe6ZZfG5FKedp/UCW8HGa4pBWpm75ryPKaZ5RpvJ/7MbtL7Ix
8s78coe3HpANxIdfn4PGwIoCjYLERNovMxWEwMPWT5mlwXiwnUwRCgb+dilYcTLa
l3Rd1BqyLxaiWPZovLWxy871WwaejXXH/l4wZ3FfQfwH+S/tqoOehFoP9zSsAQC2
hPlB6dv/36ojCjTEPAMjWBce9qEr/fJ9vG5C82PrR76I39ytAEqAMO95YPd0aSrk
bvyY3162yPvKWcvHf+lXEJTujQ71B+grBYE6zsxHn+C+LnZpv3Z/qWLRtqnbO90a
p5/y7SJhEEQuqD9Kr8pfzC6NXTQGhCSTRtKGzHJ2JAFHTllPU/BHwxSr5gZj4Oig
uxQZoynuMFprWdeYKrWjMpHcY9CxYZyM11q/E7UERnwQr5w9Bb8FdTzuY65YJeqg
Dc0eHKZUe3wla9Uv+l7Z6njZ2lxniDn8rN0wX66EpDW6IxBaR/6oGyPvUvgP9Kja
AxZmuh/QVCE7p4sOjSpA8zMuiUQqhqeS1fZQPD98CtpNIpIiH2Y37UqPaw6d6Roq
Tf3nPF6qvkwvQe3bPuAUzXn03LBPRFMYUI4Tpy6RnSQOwpviqMMOrUcy/kUVNRFk
cp7QxAUSHJ6zhpcQw2VJXejZbO3aPWLtW3BlkEwIX08tJ0nZTZV8cnh8tgLdrAaA
sa59rI2K6ZWEujcEzRPS0iC9rv7sIhAAyzqo+/G5+1dityHoLcRely8vKSpjy9Tc
niEsJpIlHgYo3Ltl9cmu7lhH50RYqbmHjldFVGXSrsWRWKLkRk4Ym96kIiU20FlU
tdC0phVcTCjO979UjgLa20thQ1maM8VLhfTaKhhKtLWyq8+Tqh2lHpru3w72pWPd
I1aVLRv6vocMFfd7cC7+pr8bTim8Lfcd91gGHLs6fGhCZnaXL+ccD6kcF7Dq9inm
gpaJoZEr5WYMPF4yhayhKjtj3aiwJSz1gAKVgL6FQsrfozHo1roJI63EtnTVEd5P
jncAdecjDVGVx4aukw0MyDQiv6RFGUhn2qDH6Ehk9OeABWC2nkSZZFgSr21jleov
1GCrTyMmEm+4r6JX4BZlgSg3vOq/5TBtEcun5HMf/V3e459962IKMI17+g20axC3
NRH9xV/lt3cKtkEa9zr2ktxd9/QYgprZUNJ9Z71VkijFvjFn28n0b3Zq/AqzTMl8
cOd+mT/oUvvc4qCZNCPR1vQlIlNGL5AvhRG0gmP/OEQFzEtC04ZfAz8sf5xNrKNv
rONe0gBLR2ljlXJOs60AWLixZoV/+7/g7yaFJqEqxB2a/Yte12KMqNQtLHGE2Bey
jPsGNhrOyMMZJ3ML7twIbJJHYi5AjqQG3FJhAi4nPkIClf0cfUlIqlJtS/nrSiIQ
w4F4tt+rPgKPhrNw5HjTYyj8pbqXDuy9dczlBIMOLRRiqJkTN1jvKOL6aVwbekvK
uVNZ7kmwt7WJQfvb6qE3brBWV3A8Z84ayckcC9hX7bCwOjKN9qisnXMJQ7+uOezV
U8gAd/t2QCY3LUCzCiim8QT79Xmzh2T9HXb0H9pSurwk16p/ZlFr3thwp4XpHn1X
Uy5L8brJNZU2tH3a6E96M0N/g5KjW933tV24+kTjD/eGw+m8fUW8WzLI7I3kDVLV
m/2yRdO8m2hA4Kko7DHr43JOyGl3IF9OG5Ynql5PiUeLGhFDBhfu7W8WCn3Gr7Ro
YYp5TbmAiA6pw0HItGsuyXemibHoVdopnrLS3PsqKhoXUTUfnyM0GNUoh9OAGiHY
MRtpMjS+ziO3qquptcAqQpaA1BV22ZpVU7gGYExU2XnGp97FRoumGYR3aOEY0hXm
TTUJt+XGaB0gc041wJ6CdgIHN08v5HUaIzNiY/X0B3RuHY6wGN3zCxeVy6mGnsuH
nBAs/+NsWGpL6S8aTrcqlgWghqLHB40zmdWEjo/EoRrOJVU1ffFQuwkF8WkRTHLg
FA5qUZ6OtQEQwZy/1p6dFNAVFftIjqiz6x6xxjuJPw8yydWFdRF5YNJaOMf4Pe0Y
FT0uogHx7K3YYUul08IZ5Iz8puMvyENpQcAjNF1CZQEggyuWM9RzGzRarFr2ZUhk
rM5zriTQ3e+2UIGZ2T1RLhIJAM6s5eGwAttVI3za95WCTJvEETwNLohH9MEmQVo7
teObU7tEtSgTaCcilG5MxlcGqn6U4BeIexSq+OzKofysLZ8tMf6nyBMkcFAbNthF
zhJG0Monotsf4yGy0i0QgMUEhfcCXPd2TXF43DJrYve4cU/HkdfYSj57xZrmKDZ0
nz/8guOswoH7YaHufF5lxn78AyY97dKdD4PluQrj9j++fdq6N8mh/fjDkv54cBEa
P8/bGiPnydF8wnIJ8o0LnB/7ktkzowWJlFFNSyqYLu5DdOaUiSvQvNPYaJVnuEj/
0uPKHImqdcQXJ40zFICK4USv+XOI2HUr695QzzjjDTQX6D1Pucpk23jaCebzhyLo
FZfl+iqwDr6odDk8UmBLLsOYBxmSFxJchydpCumz2CoCkCTsQAToCjy+uN01QWq9
Q10QNqnJqqmK+Md+ekm812mJNor5jBedJ9AK9KLcJA0ft/gXdV+MipxN4kMw3XrS
dNPFFFn83DNL1M/9bLAR8qSR3udQ+/BydjWhqGzH5dBCKO4RnE4hu54aCTXQ24jN
xYTOQnhYOttTKJpMktmhEMoCYne5m1Bm7iR0ZHsEpPpWiQ4cLHUyjELCZgq8S4QN
DEAn4M8FveGaonFiTSgRFtOwXzMD8UKsez+Oa2sdg2P/9kNRQfd6JAJ+MpB/yMMj
7JGaQIV+BhEKMlbIM16ws83/QVnSzkHjdBWQl4aFzTsNy3XS9bIanAW4F7W6GCC3
K1z8bhnhvHObkdEBkEYecp3JYXVrIq2AVQq2hfVCRN2470gNqBB8rsMjbpa83oIt
vncPHmbSROxhDB9X9xRUfIVu79lHZWvPR51Atd5H4mGlC+ukttegieVdWJ/HXw5K
zsCEPq6Bq3bRekRir193aSLpb/7Bl0jPhdglqvctNzNDwzVVbLXOixTanHYR1qOl
vNyI57vrQjLLI5hv3dTdzrnVGT5Fp0Hvv6aByluYX2tbZKa2oTzEDHatseMhQQF4
y2XyL2HtiS8Dv+WxKPo6kgtcTWwWBIs0TV5aGHGdUI/Do+K6U7R2R5gE34TeGF1J
oCqVENgDIzsH3BQGDBal4ZOJOH1jDqM8boRghrT9uPVzxLqI279P2fWZGOwuq3N5
1UlQbDaSEmAYCWxw2Kdq1XZiZbZ3FhbdO7iQgDBbC8yUAGeBOsluGVTc3LJlJnWF
aTy+J/nh6H7ykCAUOazg/w8DEUZ8lROL40+Lnq3CNh9k1IcsBdge3JwYD+1KT6hM
fPPoyXrZCQm1kF3hw6cDIPdnlt8h2UN68WAEE0yGhV0UCVj/0nI0juQFJEk3BBlK
KM0cnXe5pBFHhI3RNuuKf1RSYRTQTooKrd2j0P2Oe4/xs7zvGPqnBUJx709n8D/N
o1iMuTWez4j0R//6eUit4jy6ZR1UP90lghpHJCpWE0Add5chZsxk29bFuOleSObQ
hFVbmqfvR66i8CDzTSLFugt81nYMSdBhGReBQ8uJ0aOAmwdV8AymEm3iQfFT6lET
elxTdHq/bavxvGsL7j5lc0fXgemZkHOn/jhVfeR4DykPwE2ti/BUEl96K/JKamIr
pP83+ev2sQWCna3TdoX78erRRZHkWeK/5NtGD9YnQ9Nl5MkWpP+MpOT5ianh/WYT
YMicDR+nC0NcAMOXMQTrnGrJAOdcB81JlqhGWj2lKCRZCrdpu/5nr9RxXr6sXOns
76hlNdBpadSbRvKLNqKOiy0KemDb4sGxztqZR7/uD8Ea4pGFvvKcdSJXDY1s4h8c
iJTskXk54+77iNCAYDI+AyIN/5wi4CvUxXESNoSkdxZJSYTxsSGka91aPGyxUOVR
Or8a7yOx3M5cslahY4BW7EfZoMiRr4qedbZRiO2sgNzv1bih+Ez8xs0VS/H8AAwc
33rjUArjsFUcBNDk+YRwU7Ojzd4Xc8O+BBpsFdx+1+0Go64za0advn8E1szBj4Sf
q8uu0ENNVWDyIIgVqWqwdEAzTmOeaBcDBZA0H+gzSWXO250KzxWad9v8wnhiOaoZ
iF0n8nOyrE4UCIVsdExqiW/r6v04ASB9AqHQnTN3oKXaKO78X2nqFzUUmgPHgSTC
rZoqvKPeVl0D0XuNxvF+fEgmkISPmdnPVpt0sQN9KNUIW/ZuXzayPAg3dF4LSVbQ
RzTaMrLi2xMZ0W0neEJ0Yrury155LQ33r8SWu7Rb1cjTE0HvixsS51r9ZxDQk7+p
qV+W22ZeT9z7sjUE8BDSVWL+HpqQ89nepi758Cepf92TIPZEjxEOMH5owFvOh9Ts
1AHuLUCOANmN5G6asjGLcL7XtGogs5KU06jeZ3ARMjuK00N1pdL7/Gr2W0kX9bZo
C3pWquRpPMk9zC+7sCusLiILGGvbSbpgrvOo4icgWFhpqWAY+UUPk7BxH9fFYPi8
wR0B3dX8mjgAWLsrkBCfhoC+T8adLQMg4CSir82xburdiiyHvPYFGabPhT9J1XhN
MsBTRiFhIsKElupiJ0xyZrKZH93l0nIXHtD5XwdAz1yNtTjsLuvwDAN0sT1eTqcd
BGH51xCN0eJ3HJc5wMxFSnJ8qVI+94Q2RX+J+6saR63Sy4t+y3VP8DVOgN6K6N0p
Pk0oAFIDp/xiO9q/YGC31BQx8Iai4moBdcX0sh//f/jQ3z2kcG/3MmzBRfXHKGL7
FLblUdN3XFU2DgtmEgxjGj2cyNLAkjZdZHCoyhMBbtFF9Y61Brq+L9q/z5PPdLNj
OCsPSy/NgSAz46MwbV0KPae7G0LKzins6pr4d6h0DlSx9Vm6PWin0PbBfYzkUoC5
NzkbWJ20sn6FzY/8r9AEJBsZccDE/tWIT/7rQcC9q3eqOvm3DmkDh9QmcfIez3yA
bNfzEP3Tn2P4TUQ4bIol0FEaiIhbRELkkn5rVgZdSl9QiifUL9RSoWYmUhPxl537
sU4bWhOa9gtS9or8C1gRDl7/OqZoORxqrN8+jLdGFd4zFfuFqs68/Pr4BKLYbynx
eXGJhsbpvMbtSKgj3WKWLyRP4cadjT/IPKzrLJYZtxKjzMjKrRg35MQ+iCQGd3HU
Rd7BbXcEvmDSOoC8smwhSVddHvzGGiOWHbVEdKhIUnpPLH/hRbP1O/jHs8UlJwZ7
SSwdDwQDHEU4zbXrOEva+JvpXY2EOAijhICUTnSocse3uaPh+a0msMoASYpsrT8f
7gU5i7jNiUGCPO8yEKF/S7KjZkse7ytDd2qayY8QN8wtcN9B1fyvErDVQtpgDYGZ
ybEHmhqAJZyVl8lnTRASYqe7h6dGCnHldtj/s5y+IY+D5WWB0EA8FZ49cwg0LHup
HNCIUuSXgqIO7ZDZTIYfFSNAVkpKMkiB6Z3EdOiHGb36ydfsnOT869Nf23I/BNdr
HecLGsxOzBRbMzpl3Hr9BhgTW8JeLwpiQjxuSRdCZGviuJ5N84L/GPDeJnkLpcWK
V5vIlfqeqeZHr6XvP1a2VGVzFdGeVJ651g9cMhjdbaNIMScGHmKhZDgyH1KZE2iJ
HjOEF/mjMetGu42LPSWaXZi87yHts/eeNSP2m+jWy8PddqJ5r2MUNcj0YAQ9vG3h
rWmRIWOASHPSWqVred0/gJGbnNcwmaTnlWgvGLkOQfZLBG46ujqsNc8gsTGERp5b
nONvS73b6pD64p6xkwTrQJa47SsXdPXSj5inOWdgzpjQFrIIPO5cxP3x/yzfMVe0
/DkG1LzdmdBG2ge1iYj+ZjLvYP4Gaa/n15erFdW7g73vg6O9DNH320vsMf+45wpH
ER/uS6bR8P/sBGtKZ7YeLm2QU+YH+LnlwqXhQ1REvNujYvBpecxQ2tGECKT8PXX0
YLzvw3Dqo8FPX2p4bOq+//atM+7HOgRLaCxfWn5fEuIiTsujyIi9XYHHJXehtgzu
+IeLbaiX754ma4TuwMm4j3JWA7d6/0VUtrFKi2ZEX/aOTMMTSJdONbnz27j5CLax
tKUHhqiGRyYwzcsINAMUwjAeiK66v8JjgHI0Rn4InHbrMO6x9I8eGHhWgsaVaPsM
yl3JET0rxjGH2Tp8VBQ9f1I2qJEJf/2HXSxQlAB8L76samW2gC/zPpkyOSZnIUgE
WdLf2C0rHXxP9Tp2RtpYwpwUuQWmX8dqvdcc6qWYBb3frQa3PJM+2voYkUjfNtZl
xkVkLIFUbCWDOTZfZrmUHzJJtXCfEJ60Qq3/C7gmgXXZ7uWIVrQEQxRPcYu7q+Ll
QrPh1snSy1FPjvGI8obTzw4z5a2GpM99bGYpEkTraonh48XHk5/YTbitxYb4iS5A
Tbpr1HqVXxRycFWunYN3Z2H5pxUpgPpyqtSjZIf5TyemmwRamOG7KTh3MUDaD0/o
N2pm5PRcOl3ZWKEs8gvXv8WTZSPCvyrJJFDyMuWkbiU9+AoF7xKM3cYRMzs0BsJj
mUwHrrcnDIcprdVdwqPbudrjIPJuXCYSBIM8jiyhsiHhC2JxD3GsYaTfSEWoY4ZK
MZYlVtPgGrXAtkQT8zwBE32D5H3E34dSQed2L7qPFApe2hc3q7Y0VHefvfGPPD4Q
8WjDqsTpwgnc9YHyXkWn57wlBQtU+VB7Z01gJIsnR9KyP8IdH4lt9hCBpujs0+O9
l+saAN0py/+ThP+Od7Phj/y7u2kGqnUgDyyUF1iIS7Vly3SS42MOWY4sy8ieh3qi
wm2THWDH4OGeee+YCeWF1+hrkgFt3lCVUPOYuKFDnNCI/y3zNcOTN/P0krBAvaFe
CVGa1b0MtVSHNEWNid7S2XvMcgOyx70ppthjmrOoSgfPRr04w6oDRz/eS0cSuAGD
FApqAvgs2xa+sWlbY18WbS4FReFqSxkIyamZUyEY4oe4VRvptWfPEC2odY7F5GYL
kBj0q2Q1eY4Q6tGgu2jtz4Nss1k02P0qWsI7xpr/k1NC+MX49UfaKMoGs5vzGbW9
ZZzgjTucos5P6oOSiHYNI95Dp1cJaZICTs6jqksX7OmDlc3wwtxkQLEFh7r46M9L
PoBZoipkL43YO2D0CqhIMBwBtdQ3PfNay4WtHRAjYF9aHH4ybVpwHkAE++/BbMDE
aZhs2eSG82K8jDDXaxYB7NkAORGPt8M+4V2cudLJwsgoEeVb4LilljXtEBIajrzQ
dbp+QxF3v3nyTAZuxoxNiB3iqanP0eT79lDhk9jw2zcSgVfgzun6yU0nz8/8WGgw
oicqwEcQi+OnOGA+VX9OeQdlgM4nDDl7GYFKf0wcMAGOQ33e+eCKrFVTvfgKeJd9
AIwRGjMSPTqt3iwhs5FakJnGkQPeuiBh1hDpRIZ9xflb4qT93gGeDpRBF0S35L/l
vK74hKujI9JzfIKOACOLOWL/frxJEWt61/avK9EFoGu9jhxYP6+ERHyPbgPBZPgb
S4KYd40QTqcn1I1c8Jl1QUZrM/fRxCoI78RWR/3ANp3G+4i6lqJv7E4A3/RqrBbx
JDleSEDpg6xDzSK++hP1NLZd0gcStbyHQwb140XVOOgIiELd9x77wwVQaI6SLHLX
x07t5ohpmj9SNseAZvfN6NAIwx3B+7IoRHmNGN7/Ptg1/wl88/Sm3o0ULndis9fs
PpTMjir+m4xM264/HukVq5Pjd3txj/VQ39a+5E7Y1+dojXUM/P5lhxgqM6yfEPK7
xNW2uCgtRxObziy7f4M83ZYhmz4D+szxWvNgEa98tmTM7xo7yCZkTht91Ao+Xh9/
LmuP8tSrKc+1/+2KXxBMPxQ7Vq1PBemfvMUYeg/fOS/NmvLt+ClYM6a+B0yz0kT5
m1DrX8oPiiaPy5sUTNVkCVl4E4tOqvMSSNJBdAfaYpMJ2mzVRAD82D1bVVrw2yiz
14aGm+Q2kIQ7zxZJ0crgdsZH9oVNQNStQ//gVfcPC+8Z+JCWsDHKJRiPWWd/Lw+T
FngIwQ+TZS+mJ9ihN2h5lXOaPa1dwpanUpIY3zQaniiz4mQIZ6h/eHzTCuhr8/F6
OtioTZbjYDUlQH/O4evA1sBxwZ9E3ezeTRghEa9AVPWHEe5ZnKjMfNDWxmQ92e00
lRLT/ZsQOYV1pd7DVj0PX+gm2Ay70Aigjqs88um8erR0WtNFoU+9b0tvm44S3uwx
BH9PfbIOj0vHdr0Vx9jYFQKTwnXFCL+odtzx4RBkdGGECoTTpi1aHssiNq3YN0NG
bFfc0HCdo59LZEdrgAa+9w==
--pragma protect end_data_block
--pragma protect digest_block
j3WzPv87u9dITkW7SCAfEJX87JE=
--pragma protect end_digest_block
--pragma protect end_protected
