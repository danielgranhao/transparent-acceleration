-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
VuXN+5160RhMoY8MWppKAJS/20U6ac/cj25RT1hiEkgeX0pNVAFkETdgnDKCWNlU
x8PoBILe/uvgrB/Mh1EGEZv4tShVy/wGWh+VV6vjJLr8RmpVV+7FXxs3ZLS7Qs8+
2DTH3a984wtDVHUU4oliykEr2dCoJdEMcVz1GXUrOsU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13584)
`protect data_block
HW6alffehG94QMfJmDXi0oXS5Z181DMoHlKMJbhoo9EtnEVfjdw3kcGxMa5qDQ+d
mvYaj7w3v0uJljpRhD0mMHtjQlyeYwTPSEeDmuVO+Yf685HFOPf/LBHzPYrK96ia
LxiZs4WkhJH4VGzWnaWHnvN68y1LDcP1ae2TYmsWKt8atq0351NXhQK1kykY8e/s
Wd77+2YW0+swZ2zQFKA3s+3RwEwNe1JMQSjKdZPhEY08APG8qwtqMf7fsOK3jgXO
+uzQByMhzN6JSR60ESuPcZBpheVvHJ4yQua/CpDut7iNX/lBIpc+ghVonJXo47Yd
+zph3ocdRp2y0LUFyg82DsTIgjLPkzBy4hGXt7a6UJw7x5hDJttyShduQliZ3HYP
p62bMyiHAZeYiiaDljHnG1AvT0SqdOE9Ejj9B3PNpyHfo4x+nLMh/G2weEQqZppK
IRcEV/JSMOEuuziuacy3U38zebs6rzvX9XbyAWIq7bAfr1qMTCTZX2BCtVQ2faDi
x/5+1uyufRkm1Zqpv0gZcNxrvJ7glOEe4U+BDILcDOf/6pnvSHDrCaUKyS4zDm3H
Q8Io/CMzsfDHLg3eX3nQ6m6Yf+QvuP7nnAPyBWVnExRerek1SxWqqgB2p30StDZv
mR6nQrhJtXQ581dZMcKdf9GoQu+hrEwSrItDRG4LVIbxOqk19/Jpau2PIHhx/8Am
sa7xACF19WLDqJ/KI0pdSGKzQFP9k4zUrMuEy8kju4pcI5sU5ZrHc177e2EdMTUw
v54Tfp0cv4tTRJXn0flqD5XH5sBPZNtp7UvS3LxRuizdQBECD7u5eF8g13HTbQF7
oDKLvz0NVozJIer0JpaYVHPjfKLkThyDj6XmRIAtNBQ2ibmz6SxxvLELApGjz8GA
nP+gJcwXgFy75DKnl6VkhpwwqRd1SeWpACz6BAHB87wwG+fhsJA0/RGqPHOPEbE0
haG8NtwWfWCc+6V7NZJsxfarOOQmfVXBtneMOkD0ZqkXiacxFRtNn2wAK/qApny5
W1vfsnWjglhbNNJfikFPmaF3ZLWf/J1bJ7O/fpCb161wBBVMY+HPd/6ut3BTfIqK
QwrQDbyMBQdFZas+AdMo4nP7nQz5af+cftIA4EIkZqIJN3lne0ZeP6n5RpRS24ri
+40avZ9Ioj9L36jpiiwAFcWWy8hGZNFpo8kEVbsfEQg57ASWgNTgfqVbz1A4qyg2
y4cVZdH07+gXVxBL0leCz/Y9VHMROiE4hnQzkX4tueLrWMh67cJyM52FnSovgAtC
IBtgKIOKjmbdpmPPwiJIqWJguKeWr+ay8Uhq5sKF3MzP0p7yS9DQzyEZ447yOPsX
D7tCVz1frBnQSmVgUBlk8xC6fq17ZRHZFt+Z3pkfBvd4tvPvo4QOw4sXzVLRfBjZ
fWh1ilEmnxMack9DsUTJp6u+ECN5rqA6TZRieAebL/RreSh5qMwvC6a0QIYYJimj
ixMjnlEQiFsoPY2sFoIWDpRNnbvOK9EDoo1WC1w77UXWwvw6mXEvzoyMs9qQzdzv
zWfAI7S02Xv4TvuFxsjduuhC3D9xvLYM+CqQh9CS8722X+qRgGcspdTxgJVEherW
aNmcOSfQMmzM46RlJPHh/rN7+dVE8h1Rwyi0G5Dd1Lq+yqFoskzIjDC+Hw3hef6S
07oPuDh6th+dMDGojp0CnOxXFhjZUqjWSWzXpgEFd7JCPrSVShPIazCj9iFdv6WT
1OCpn00tNj53BwPqWxX65KSJdEQDV9dWrkLdKQB6EBoau8jkKPVPPAQnLgSBHCAH
KglqTTyCTcxtlNld+lp97jXhVpM90x9dIHqUo3uXC1X7OwGsrDop9aIdsijDZZkl
BbEM4Blj11d7azsHxRyCFdng7lPQK9vXNstoY36EnJlf1+XDshKdFyviV5QvnMrC
SOTzwbWYjW4IEX0r97z8XqWiOhtK8thpvQqB45kKq1Rx2nDHTRgb1UesaLSIvIyq
vszC2CE9Lpsnzk35whVEzFqQuIGsyKwMfgmGWfalmpxwDpcAT3pEbOsf6Fd1F3Ll
WEAVRAxIxwUPf7bvEE4yfUgsDyZpsu0haP1NRhWY4ORVHj5ezvJAXLdj0Q5jii8/
hxB91YEDPhHMy7QimH/kWQVs7aEbKHJ2i4m2zN2GjQLi0eV1ejBrir5dEyW8C7gB
0pD9V+gn1vtgLNaBTSxkJ3KFqGbNyC5ONTXSv/2BWHU5TOeRXlMoeD+M1AiNjs9U
Ow4ZRatVRoE9/51R/1NDxptYeZ0ekQSHMGl7qSyCnLXB7Efh+IZq/Hz9yPXHQmWv
K5XnBS70rs4sRXnjUd4mB0HZOO6Rx3F8MJHJX9BuI9rcqrUBC1B2ie4yxyORFpKT
yJW6ZJ/89iuDfU8bRmhMkKjBTA0VUWrcioMbjocfDhsyR/LNMS652RrAmkBDLXfZ
g5cZmAUPTe2wOKSrY9FzVvUOCZzqHqi7SfRfu+RH8ovdlZ0dSj7QPHgpsx+va5Fy
k3T2P9EcAzos0LvnZen4Fk6Fqiv5yns01Hm52QMLDFwrnmuCKU1dqvDhPzASldYA
1cRwaqPZkQwKjI4Vi4K6nHQztvDEuZwjNcfhbh8bVHbLo6RX4o1munL4aGHL7pOL
0Y5z/kHFOl7RUC8nDPcMI0C6Xo2ikiaNZtWkKInvg9joqmc5WCE7+zKC2w7SN1XA
3tgqDEfScEBeLKOcZXrdZdK9OxE38+1kjwf+HhNzIpR8L+6D1k3psxeFDy2PqV98
dnkn9txm45fZoAnTAYeAJouokJCmNUJncY7CFa4fixhvuZwXrvqGVEGmyu/8hTCs
9/ItBVzglv1tPljvoS7H72wDrj0UcOsC7vwm5ocgXSypofvJvTFJmQMsgWNfYdXF
gTZTRvpXLK72eaSYeZcZQ3nSRudvJfdpRIz7QckU5f+xsDSuj7CAjWubGzZ39wWw
CrZQAGS8YPQtVRYYcJUv+2nWbdy2SsW/tinFw+yL4gSuohl4MTz0VMAe77QjqW3f
wA3iuplt3vnTyEe+d883CUlUddManaOA3QpfKPfYNyqCGqV1E3U5evIy23JS+iTO
otbmzaU5TpTpw/q21JaCjW6mzwE/IL5OdhLtFUeh4NLJJBfig/uXl89YdWrq88Fz
Bjptip5PDltEagoAyxxpJJKJOOG8E6PyCXQC/qUX2ZZoXBA6eqIqNq1t+9BqziOL
pUvl41Hd1Kc3bnZoekVc5LVniY3jrt5cLJHlklNZlETLxYh1ltiBhM3xrTmh/8bZ
jW09OfJCpmQRuNpcbMNm0wIgvtW8MXR6Q6DitLNWGaEbsnkc+ZXO4s/GTfKxiIG7
yJC4e2vXg3nfrP6yHsc+hF0QNK+K+6g9ELFfPPym18y5Y1Ewfv9CSmwACFk8WQLg
4e3pFa2hx0HZujzlJOTRZJ1/qtlZCSus2Rz4bbp3ewbeNS84aI8zCIyJj4A4bOri
Bb6HtIub37qQJXTVRLlbT57PYX0eAyKtGNxE4SZN4ZqiF9cMazqW9PwBzar40ypV
yzFf7Nk68kQTLh9udNlxYMbSTnLN+zbeUyNUImOz2UlkG3PPZQDS+7R5S0GgZ56x
uRlJwLHdte5Hxq4ahQxQKC3VDByvvC0+ZZOjrJ3QnNyZbKTICLQIf6jqB6G/paq8
L4gWgOD+zo9ufG5+1pDkNl81jFaqId03VzKGo9mUZlp/wzheMM0D4kaBd4X1yS7Y
PzEJDccknHhdhrRJR95Tx79BYBkFPIF/iMNwwPiNJB3G9PBSMPmSOTgBUzzJHCrN
sDVsLH1ywfZoqkiMW76xIWEBp4i37pRJyNJeqsr0FsWmpXhBhyp80P3wda1g0dr1
H8cFypY8oGSICpB04+WVRRhW0ci/OJfTyDLE5sxJryyrKtDcCeBhOv1NNXo5goxg
HptMu6WxAVAAsbJ5PIszfTQKBclkWUMMViH9JxWa0BeZifF2oDG/4YncRLSnSqg1
Fx52l4KwO4rsxa1aJ1spB8E8XovBXJ31yV+w4ctxhMMuZzQrCBaJpytrh7/2sphP
SXKUM8NXYL6dRiX8k/un/JLIC5FbqHJssfJn0U5YZ2aINXw8G+Rgc5XWNtIm2zSm
1I+ABxzS986ghtmPGZv8S8u6Wq2sRBeRnlaZZ2SSIzzSE6Rd2uG4B7uDgBkWOdTN
9cFpUeJPle9EyIK6H9L/DuE80dMw+ecCnZY7ojj1FkdJegNQc7etGsTrdXaa/g0t
eTmN4qTT6x/8eeFBEY3EhM7IPGfT5HVO8ACafVkOAf+gitr39qrxXaGNAU9xxNxP
+P7XcT4mI1wQR0y3aV/YOyeINSiXFj/4SVMl6D9U0MOviwKm765oDxku3R0d68GM
fUjeis/mjz1h/Afv2kESivgt5s1qQBtfZ38LiJJxcM5Qn77E+4KgYTfwn4QswOMp
kQ/Kh6gTLK1wN5B46Rq5HeYjWDov0UtzX9bFSO1eu7nA/aqMZOESsnQ7SilWHreM
8+bjEJfB6agNizXB+IOBfqaCHW7ioso1NrkOj/lG0BHqtWjAgDRv0a9s7AcsOtkc
8BZZ4nEnx63/0S2jUUb5FDTaM017G6iTitjWAhaJacaO1n8NvtDRCdbQtdiocFG7
q3wg/+/BIfphVxlfNdr48DuI2FG3Dw1427AN7xnrUMnHNpMsz+l16pGwA08Y60Dg
DCzojEtWSV/InanbH42ZD1N5+Yh8AvCr6X9JawfXADbulaCvn13TAlwR+c1DlxyC
DqDBARuLsPaTS6cza6NBiGQGFF5Mzoix8ORzFUCX0LpY/lzygwnPSfmzmOSLpGiK
W8xfHpd872NKU42X1fEzXhDGiEdijb8HE4rn216QapxCCbzcUqsnMcNnr0fknkAd
cndaoPcJMlByOHYY7E+Evl5kOPPtyLmpuO7mDsZEJamFocqrhW+8d9qxKD89G3+J
EFVKQddm4LVUAcB4g98TBY0CnyIyiuvE5CRdzUGC45alcYV0B2r2el3ei7+7JPBC
rJdgKRb2eI1GIjSRFe2uXF+3IZBeonaj29ih+DzCsuYGmneLrw/9Wh8rMfD2FH3D
aWJuNkZuxl8vdtlZ9jtzEX1IY+kKZYBZJr9fbEckPpOSSEKpbNADWUPOyetsChgJ
1zgjSCrqHIFhIgRX3Y25YpSVAxTj1xWtzntE6d0lkC6fHZA4dmrlHURubBMB6Ke0
d3cnsXfT7HfM3CLNFcbRlyaDKB1c8RKGKCZAWyQf8hNLSfmP1ixj6KqrN3wdrCDY
ehBR2QGhsg5YsH9d9U7SrxZLsrSifLDbwrEOxUbuwSDURAgYf9LQYBuwbE+htFHB
jgx8CujqpDeqzyVYbdg2MliWbarUFieRx5a9OCzfQcJmeDV+yyUpPMucNXqsxCQ1
Cl+3CA6eu3gNc9GNdoaWtda9S4ct7JC2M3jzDs1Kz545N2Fasos/aRFbpOJmb57S
790H0LvUwV7NhuY/t2tXPN1bnkymb/n2gsAimTFftcOiozm/DyFVHfjV7cP8sXzl
IyExpJctMcwdteUuKDOog6EzJ32hjJ8TQd0o6UBN5DaHttzVoZue63Y3nl5yPoiR
U2l+f3zuCFB9tMViWSbqCx+Ydl622xSd38Q93SInAwEY0mU6CeJ5/vR52gxjOJo2
zFCQe1nibx+Ur/6dBq5txkBgyGe6sIKh4b0WDE/CGc7PL4MhDNxHos/Z5wC8FbPh
osyJCFrk/nHgEg1cPo9jj6tIMhg80oaULpMbHcSrRZJQxDkEuw61aE3nlnEeSwRe
rpOcQzBdQ6jT+WSku04qZKNEwIYnNoG56D6ZyCXtIqNXGrhnyeEqXd3fwHjRKWow
CpqdMpfAd68WeTclk6m2JfogDzq0glOPOOFu+2YUw9mCKnetp7T+7qYW1OBKqVgq
ieWC1FAAGUV3hGN9iF2Ckp0psdQDQ3oN3QaBAiuC/2sg7x2bTuPl6Df6zje47Hq4
0QUZYcpw6Q+g6qIs8Asv9BYA79mclUErATcGDVCy773KmIv1bqXBadfVQdvjfc5H
0fHNV5uTffheG6wehVxzTjU/dqitJQu9wqxtd4fGx7vt/gyrp7djuQXO5WQ4XMg0
ERJHDPUTii8iTPxtLf8xlZbQ0bfd670odD2KzSxwWjI97n4NsPy1bwZ0G2xPdZUj
HSExwR+eIzs8nrTNk7RDC2mAny0lUJ9n8bDeVXpBlVxVkmQVYZ96K1nwDryvXXZ/
ZfZ4L8GU/bz/bO818fU7G2K10Igp/bDN8yFy8bqul71T7FDHQ2UngWfjeLi9XlA6
IzXH5pIfrfUJtuIUo63ZjnKx8HfLcsbNh6w2LXKXdSQfels1LnrB5eCUKrrOS6IX
ne10eybrWePDEcgEK+wMLUlX0IzwIkbjOxMaDR7TrpgSmDCQsxOaNuSRj5buw9nO
C+f6AHcVT3mk/CA4fyQuK0qndKAbgcYpu1w7yq8peWeTY+QwNzqI0XToBnKS1TDf
Y7FOiwus/NM56E2m00H3blB7d0Z+/6kuSK6HlA4a2ClV3/IxVubXqcR97CxHHV9u
kRAzsvGPjxmmMQxPpPJeoi7vkjQiFq87rbUhzqLVBCEAwWCqM1fiHlAPUFQprwqV
3ChZRsO4KcCxAtMzJm32u6mJ0gzkPkFXIABD5essTvmDhgmW3rm2gMZ9HNheldbU
RXwHUV7D27Dc+XQTnNluAeInzjoWGhZnrGMk074C3JDPnJAoUnP03PLXLU99gehF
04on8gLKQ+XGEWuIet9pVB221NBIZhOCRMCcK4D0AR2fm1CWGTj6xNSZZjzTE2hr
Z6QX2t17b3x74GLPfs+ds7pOMhVDLBMoSXe7W/e9vl3RKtc3/shgSr5dIxPmv2Tk
6hIUIvLUk224dqrwQF9HIpBZsSo86y/emxL/edEF3k6V7ZrLP0K6jCaULSWpdlTu
pSwdc5JrAYXK5s0h2Sjd9d3fJ701Fmalp8AQ6SuT6jOii5IcWnt1Ny+eGIZbMS7k
tbAyTjsY8KHmvznlKpmY0LLrnURjcV8HXKt0D2ovkohIn6yznK9hOiOPzHURMrZJ
ScfbtWdcb3mIVX0sDBomQoaVapkZNGR6wM94+Ebq0AozacOilAmHKD+CIY20+r3h
dNx+E8i1U4XtaJ/JwKPvwArXNqYHTjBb826gmZkjRvtuSwU3Gp60wZw7zZ/UlDTL
KQC57DfPC34poj07pAuZCu8dlEzKBrdxmawZUnym7jWwtQ48tOS7llunnn2zDjwn
Lml1CtoYYi83xz7A+Aln2NYBkvAl2oXpceDVQmUwMC078ThOLGnycXGkhHsOEEKd
b9ytWKopdGpUszhUbhvEF7ZvV2vc906rAsUaA9Pet/BnRVQPnSpjgkhP+nvzz2U0
3xDpLLn2/IgZButNRAtTk0PRNNeuVzSNsw6zBGxExzYe81+cn7w0N68IxdEGIKAK
CtGC3XK7/G87KoBFUKjMfL9UTtK3ZOH37QCSqpd57UvKA5Pt0qqVGRM6PlHSoHAt
zKbWQoalFhS9bgL4BwfzjlZu9ay62DsIeY6kZ4nJtG/Fjft3zwmCLsHJdscfq5gq
VL9WC1c0xNR+7A2+aM8k2wrjvvxGyB1GEVIYxYXZIm4QSSyESQGREKggtmFqlgxj
+anet0fWoF1Pqgdu+3Przh3w5eRxGp4KLQoPUBVPnYQiQQrt/pBkC+VZbU2ke8ag
7gkPsK3LZv1LsPjqlHFoNdQpw6dr0vJVseiFbMhxglTj0l01u915gcELV+dUknPT
sDBzLM9OgT0dUsatYfrKUNuK4xdsl8PRVULtb2rTX+vmq1IV206r5B/OAYHCtKl2
s3OmZDbXjbhdz/2n7trzMT6ZHhGD0Sm/jWaNdzoNnZkMP+HnkPMMY6qcNfHqHkZY
MD+WfF5rsV5SPaVQ1KYfUNc2g/n/8d0NlElTupapDxc5ni0A8QdCag1bSPZXOvTl
uK/GUGAAY5fN+9watW33r8VtK1b0QilqOo1opgx5a8nzVToLWaOsihQ7bAbe0r/e
vp0FydLlZca8gMl9Av43E+c94PNSd4ei/n5N2gwrIXYnJ9Ss0p7arD95E9AvG3hq
Yq28RMJlzpi+tS1JTigQUU7SA4fY4sNun6GCvhnowdMkF6z51oP7TFw/T/ricTtq
4Cu53JYRSdgpHSFXwmr3P2RvCDHhbBarmwrxVXnqJOd9gSUlovAoJb7A7XEI9UQM
35noLyoFrPYpxgwsbwvfq3Hq2hqzrSZCMzDPAWcJjUtIJnxNzCp1JmdxzOzq/AWn
9yBxjgGVgxwbocQsFdGlkaKERGujL/oGI3XZ5U8Z5NrmRk7bUhByjShZeQEuWKrh
mVjXju3lqaYABm3nGpYKpK62/n6EiLf1oKWZgRccyCSEkdKFAjfu/8Y78vH4BiFM
Wp4VW+C/yt0yTR1qJmRXddiFMAD/yzjFOGIcVLB3jcWCTdhNBlbKsZc0crskZUAK
wkfN+p4h57eQ3Hx9poerEq219DgPU+wNtpBjr3WVTcYuDGnT3vcsTnjfdLC9hiT4
yUfaStk8mec5cGEylNjLphqgkAy2MU3z2B9tMeX61fXiZFvjgd5QaIjv/K+5NyiC
pCG17JqwSos5APyoJNUWWIWB4hl2gNfSLmVRxv64DhrDG7b+LuMFV7U4wIaNCdjC
LJ87gUHfW4NQWUPTD3vNhRnGWKrgXHA3BasGN/D4gd/3JcIVOb82aRdLMbEAbkkV
ftk9dlhXLEOLyZnKUF6DYCDdiTZliiButmAjUuUSj8KjJgROBOvbtrJ4s5n/6R5P
oKzb0JfSNYHsMyvycFOOQHJxy0J6TZRc0Be8LAXKNqWNQeM7bH0O7MCPkBSOsU0s
HGlpMTg1rhO7KCT5/jHtN+0Wp8ppZf+U/WgeIPq3m68rxHx/MtBfwfsFfNB6BYgn
0o6eTwVTR2hJUOhyXRZ32pWvPKX6+5w8XhsImi52fsKLNkY1PfOZQHRc5IwBjhDG
T3uCeqQ1Eko/6nLeu6mlzbl2GU5cnMVXRiddcsWPr8hxLv7TNovIo7SDwX9ZIdIA
hyoj3UtjvN18+YJGxLzzgSouXj6q6Uub5qkaZZFtYUe9cNrbPzBuyh0GXDH0bM4p
SJfzeYZh/Laq2gMwQ7o6L0Wa2YGNnA6DZl6Ob260jR0c+XxLyTnPIcPYjm+JfFhS
NEHtsWoUI5M/7YrFfhOW5B3eXN1WRtWyx4UMEmMmP4bBBswAUia7My/Sr7WV6/nT
aZcAemwOu3F4NvAmlXiqKDdcYMmwculehYsvzGpE+WU/T2L/p8+eXAH+/5zN1ydP
Bu8KJ/mQQnCXHM+y8MWb1ZXAmMHW0BKMMR5LEOICWIs1GnSqJGxgt7q94ecfO9/K
+X8CmEFhtAYo5e+RLGqecAUbYrp88GxX3IO2e+YGQZvFgG2kzGhL31RAzKOOKDk0
fSZiuhTIV24GyHjruCvNik/sZilkczY2KVZX0cT8oLzM+U1eWn9wX2UImggT3WFb
gSOH52EhlqoxkePj5HMLvLAts+hhoLmfRg/P5wyDa6ttDp1H/xeR/PfdJizlpe9V
4HXqS0sYut4q7eogMy3d4YlxGSFtk0ANYTVzuwxtM91mucXvdvL/jpvxABIe+vpC
DE2pnsGQeQafpsty9A+ij2/WK0S07gK+YNaNMUZh6+REK5gTyRgARvGPKfoEbBcK
5fEtTnUljTkMdGDuv2UTJ9wa4BggHoz58T2HDtGOQcik0qDuDZ3qw/dNl0T2QyCf
tqU3Rv7V44tuoegP/+zDW0ug3mMrMYFnIV1yyn5FbyL6CCXoe2sp9lQusIoE+d2f
wXh8GaEpOa5PO4eIl9MnbbcEJ4KMJu/OI01QhNPhJRH4oqFNMKZGYVGKWxycXR94
tTzArECjcYNE0lTchxE2pnePmiQnV+om4XL7unnih2a0Joxw0uuGUy0eFcLUVuRm
Vn9dhxJSzli/llxmEljDnnPVJWlUGYJXvgO/hlBlUQ23NWLTGjHfozTUukE6kpwA
ackVKqSgevtI1F9S6mgqU1LWhpj0I4xEiIdWfr70EL6LTMeiZA1GB4Ctwd7XZzKU
zfqJre7bGxy7BDtE/AH+/47/Ytxbd27tfBTBBINyJGJq7zCaP8oZbqvEGkgK0+Ci
VUpOlTV5YZ6omLNDeIT+hHQXK3GN8d6+gnUfBOgtbfjQmocVIFiT3O0Mdh9oy/WX
zIpd5Pz++pKL83fuxyC4Dh4Pvnmd2NM9fY4r+/juNyfr6vRGyJvrb0QUFyUfoqVD
9XwxiZi77GC+cZXLL1Wd2gf/YspZOWdmIP1zf5ix+ZshKyuMlgMHiQn4SVIWKZb2
XtEqFREQHtAd2SZv5210XIhOmPCuir9ti1gurGveN/rXn3oMSfPjNAH0/eWIhVrb
kWLIo4MZPJPRxt5CrzvJYHEt38mConFhf3qvYpDtjDendFkIf46SFmEaqLpUmyQU
5HpIijlfARQGEcqjIVUZUkoOjokWt39XoUZfCKv64lchHM7AQKkxRnGsdk2kjI7M
vsewEBYPchOebRz8fot2LJ4xNWA2Fs5HBafH8r/4sve4fA//N6RQB3/nLKjA9OUy
Kfy5A1g7X1eJ1TRtnmbcJLiai7GrYVSeiWK0Xw52cGUlK8OX4Hc4OSkqPUV1pGPO
9dCbpEzm75GHFqNIVuOjihCFj70ARyLA9hm8OmQJWRB2UxdW4phBPn9VlwMGX1L0
wT2fM5eAXUTXHckem8iUFbtIMeIsFVrDNRY4taCX72g1AoJtIKMeGWaMf6YkrO6x
0c5DVaAalIxFi0lqzGFOFSpkFirfZmrwZ8FMM6vZiEYZV01xk5btEO57IWaXk6YT
furO7LY/dYbYLa/kroLd12ZMHIzgugSDXrWP1S/i+dPSb9s4KEvbwHlr5ccpl/Ah
axuw73WMTKH/B+9o1iXcoiNVhBs25GZnlp+tbj0hEpjMjMInBQ90W/Jd6MrxJlu/
W/7QQg+WhAaEhNbEi4mjiIDl7jYSCAnl4kGJpaRFsVtp6uTZ3L/IR2X7yLaTfJyD
D19GlaG7pX1ncrOyv+ZJXDQkJtBgA4aRf1OrQ1ALuymBYooC5xHe5Ezhu5+wx0ar
wsTV3P3xuonviTH+nNwP4KqDs+h+A0VZ1slTbmK1n2+cYEyiu150P+tbWHoelKH9
PDeh8qpycGUmk/l7AWJl2DiEXMKFWifwYZqwcOsum1dbVt+r0b1YynszRYFoxVUQ
klvDqU2jug6xZYwZATmOeYOrUVUaxqtjX05t5gTVXQ6fxWwfIMk8z7xFO/EEJ3Ie
7R2/TBJw0DsgQShqDIwGQciBCAsoI3VY5YNnvcOQISqZqaeYtkiSNB8PxiPAMexW
w2JXgVKr+BVqETCNEP4A/6ubNnmj8ak0naHzNulQE02zGSZJvM97XNocP5hTQT/F
KsBWPR1t99UDVMrZtaUXCz4AMMHOHp+NV7OnhQF3wy8lPUZE+gwFgLxu7wTq0DlT
5OYKeE9CaRJRmfyMV/lmj47Z0PyN7PP1PMnky7vQX1AWjZmUFnOBSz0k+w9HlYy7
XkSYYu/UrscmPZRvOgr9A2CENc8W9SZ+oYgUUayCEbRNyzyZJhfHCkmOFkbDifYB
7mJcUA3UNPjfs32vOB69FICJt4PQGI5cCBV0m7cbc460B5H5zDSmpbDNld9kz94p
qPbrhJZO2DoecpoR3TAhd/Rccb0PQSwJ4MdCeK6pZliQg1K6sBbM5csvyUfiOzy+
GBmLml2nFuQEYibsza3OdsnzH1e7inRlSCeuuSu6+jgHXRgV3w5c/LI/mMyVD2B1
vqIM4SIwVl3uOhvNaxANo7KEKeSGV4kZ/3ioISRvOj1+beC7oLWujD7jBukkYldg
Sg8ivOWDfdBxKGZ7xqfzit/QyNF54MCzQvauSSIC2eXWSXH7Kmm/CYSbXQMk1rwv
Dm0THFNCWfs39YFPkLNwUAg9cKdbif2J9tC2mZ9ROTUOzp5YqetsuNQFW1H0cBx3
Z7MpZrS80T1xfWsc++zCVR31QmMHwZHWajSzHiOEvcf9A8eB1SX+LAtgaOUIalcy
rDwtaJ38n92E9437bubrj2xJarODbZnAWjW17hj0WmQpaxWJ06SWEJjoQalzRVQP
er2SfHXYR4Lygok/cHIuNgmT1XGlOo3orIZ51RxExfu5NBC8MhHILkbHX33sqCsG
TbneXbqKcJY9Bxly4yzEB5PDqxSRgdTaKTzzoy6Ian1xuhhYTFBvMIa2VF0geXh5
g9vqOAm39zc0+8trVGHEoDYUKLpJy1xNoaTQElaW5s6Sc79oXVCO7AjA0RXGEjqE
gPn8fPBhkRrzI2tvw87VQW1QCvrXy5621RupkRRYaoQbCYapWmUkEh2ikUeQat7d
3PaOA915Za9WqJiGZRFpSZEcDi6KHnDHk5zH7e1WqybEdipqoGysQctp8nrSaATC
strzRlSWJWF/LwrmPi+2kuTPCZpRS4YMjZ1/ry0tvG/oDeb0qoDeMfFhG34pxkmk
JdX3szgjW9WTLKOSBZr7Y4qBZyTcO9LkO8OmHIbQDMAQnm0qm5E+faQR/jj1iPgs
27dGP6npdjUVAi5yFln482AE3iXYxmS9uM+OsZAZuQPsMwdLQIMu4FngZelYh1D5
vheCkdCQ9k7c7HhkZHL7OJIoSk80l36+T2REKOBs9j+kV/IBTjS1NX+xaMwpwqN4
f7NiqJ8zhIn+5O0IQq9misGbms4QlX8O+TYLjqRLyQJbyUp61OGRBE2A+odSW8om
LLGvyfnwEVFHoZ4dZFc32g/sDZnRMUiiYJi1tcHgiJyTsrgQAIGrIcgSxhIfueMQ
654D8/FxwUaP4f6GiGT+2MV8fociNPeYiJQAFvVzGZO8xIQLIwKr2ZmbD/sSFwBG
neLJFuYMvbloqr543I8rqYIHGVDMUrQlyrtl4LT52hq7BbPbit809dgwDHz8Pag3
07d0IkKybDQzIio+oGJFjwpnGCjPI2ludK1uwIlQZMHjT9pisK4XpY9TPpKL6YkO
lrn89jkrS2nVuORpZ57m42yY5qr1Qoq9kXRC+WnYtrNBe0FGy35dDQAVzbLmKQFv
kFyvPGHiFPab5dmWQesM47kUHUtv+YBg9kANI0m2FJoYIk6IH9gtPv3Gv1MLBvJ9
Rcjr3L8ShRefJjDFgPoY7TEFpLGpnnxiq7uIydZEST/MyOtgbOTyL+9tTXiktuq3
+fI4657mUs8iD19y3AkyfosPleMhOEraYaWLMQQMACsv/eKFKNzRwN4BcqD0zOaJ
lKSAabRLeW8D2GOOcUWRWU4bdWRcQAraJq2JOb5PUtWSRlxozcNvpLTC2nWHAcmx
ROPZ7wjq4CMpttjlmECSC6LMqRuhNxNRhjQub/ZwrmI//BGtMIE6hP2zj51qmkuO
Crw6zX2lladfBdBf9o7bFiQvR/kk7XfedA/SYcuurH+Fx4h6s6PV0rb4aVCCREl+
ZAzD0NT4F+DT5L8iWCw69QCa5h/gWDttlhOKjGLS9vyq17fWJ6v0MJHctY1G6p3R
088+rBx54WgpsuCl+XBmYzasCqFmzi/bSCbtwComdWdE4L/LOzBPOKKYIpjhAzRK
ynZeicaJdbLE+tCteA+NOXjXnPsUp4ZdxbdIjVTzRWJa2UvxgWLwrcJE82ckqhyn
x+xHpHR9eKV5m8FbZ/h538r48SU/bJEYIsxnp1921URs9Qr6rM+j2D0pYdOdq2bP
LiNU4XJPggDvNY0YFgT4agDHkZPMkIvhLQvR35t8Ytiq/zhK+tkmhILfcFSQBy6y
dcO7bqL+VJMqqN1aFo2KtYDkGXzoKSdRe1XPLsmOUeqWyWXkRGb7K9soMnPzjgmA
uTOrBhg/xCXjAYp1949azrbZPJsnYPSUv1q/laE3OMs+FtAJKw6QKMGpqruhRnPf
4ctEx/2l0K3SYZT0TAaWNp28CzzHUrQOuNaGnxHSNDOJUvw0ZZCQIqQFQ6YXsPjY
cAEJsXJBlgsjpu+V8JUJ4oPW3b0IUkKrhdLoM8AaIRWnI1pE/vW4Zrk1jgXNm9OS
+4KU1MMtlW7Izffdr3jZlT9NsXZsteObKDYoyKEJnJvBPsno3/OAKflQlHzKqLlO
4SDGY+Y/WimEz6CjHe2MxzR359xcBu9e2/6+m9tDLmbslDMk2fcv+18mLQbRuVFs
SBTiNTf642jK70sGMGaQ+KX9ZBfl8C78MLwNUEc7PisONqBG8/1upxrBn3QAkD84
/8JRbrJ59P7CT/oGi8y+Xc27ZE2luC3FxB/iTQ34xwA2n/tBFa8DwHq1ZCSni9YN
6hezfdOYNo37OBBV9yTGu/5FapJce6HVNbNJnDsnZkgd29ptZWVxVE1cu14aRHZU
QHdWTYhINVXv7ONdIMQ/80oIZbXybYJyKuStmhHuVTM30qe3m4JjcGzeFJ1VdnS6
+7wq2GOsfx1JrQ4zFASxAulyJFp2gB2N2ngXkecFxymnJd70WKcmoYYJEF4ZM/a3
Tu0Mg4EnRl1u8MvsKToh+Wz/72gxhRV8vWCLaT9Ky1Db6o9T30fZ+WoW/WVUW3ds
dYtMW4YIjTy34ZTdLM2MpbPNkkBvcJxtzlBfAKE8VdU6kCFm4eRsh+YGj99LmNvI
GmSB9mGGs0dR+pq659a8w/zvRE/f476Rofhvv2HNJZTMy+U/OoyFb4NqeWnSdqU6
FsbeysLxwrJoXRJjBm8vLC8y0LWYusx7DV9hM4V9nWzA2/LkLl8sGgtnAvoFLs1R
C+FV9pV25SqTOaYHJtf0JbSfu2aSwRtIlKNXiGtBZyY2SJhD3jinJcaGQNkyRIh9
LLN5Rcbu1Qm7TL39klDN00omhE5g5MbFrcr3JJft9jIafEbV3p630wXZkVgnVZbN
8yP0dO70x71RaTDlbqFQMGoy2bHHv//JyCtFsOYUst+eqT3TpwVW4BnRbEpXBLpY
1l2ol0K8AlQHSH1rbIuI0rsA34TDKk7HAIE0lfY+1FrB/g5mujxQuAGl7Hq5nCE0
zgutYbl3vaRY3qYBz2dGZh0RbAFyDrUvm4BKW4a8fWG8ktnzVnE6LLopBidjeOF3
xOeKuZGYX3tK3yZjZNPFXFuwGHBBxnPAudF5jaTDbygEdJJsUFzs7HfYoLgJqSf8
qNWbx1QMmA9FJ9njG7qA24mcH2lXnJhQpJrYJxkK9aGKRbEGRmE+Qlu78hXB6Kof
uPhnO2lR1xI1fTquhXOES47qnmn6WAthL/uIR7Iz/fzJAoTkYVXrP33cVCDzjU4Z
jooqoWCfNWAL7VOxQ1VfF/6bk+RiucDQOtCUGXqCgwNc/Z4u2qid0hmcGrOftrKS
H//5gmFME4Bkx1Ix1zwCFl8yKOmrUm/f12mk4UO/4pEOBsR7p6pnH5GfroWlI6SN
/tLtNBKnDKFdwIxzXrFDIH6iA7UNC1cDrqe2C35yk1Nqo0H9byj1N1zAszzYXe/K
T2pnJX5Uf4VTyqzhr9IJ9GoRGZ3Qv8k8ivpX7xfSV4a4wYCnRdw9mPP9T85hoEn4
KTLkJKv7KTCowI/rnlB4FnvmO40A26cM+V/uyLpF3rpikxeRDV/lf2RM4FuDRjc/
kAa+/S2t5bLPue11Hn9RQw9IWT6sfk/CZPMPb/R+18QOgaAHYICjQzFKZC0BpJc9
F2gQlQXU3zivnSoWtgBjG3L65YsefNfFox5g9AVyx1mcAqbOiAgdcdozX1GkDESR
NbtYQx9XSF6Adpy5F5SFwKFFmULgjjVRS4kabIsz6XqJyYV82Orbmj19NSB9CnG4
RSfzYRnrWqitJSCEGpdnbru3BGhK5JezX+GnckKcX9F4uW6JYQQbEvUs4QjwyRX4
6C7vJJWS/5IRrJkw58EgbwTh/ZsVdnu8WAcbXuHDTx/aTDgcVNsrP7sRC8TSVLWD
6B0YgVErSRvP2vdi1v+0r1Q0flDRpcnemLa9BVgGn8wk6gT1CvSPgRSs85XfRarS
CjriwsCkSsxg2hJ3TY88aACfv/XG3YU5knqO9JXnvxuX2USBhbJDymR3T27GhBEB
OB4t63tai4dREpdyZN0QAGcQFu8nbAYp4GFDKD4/1A+cvkAAVWzIXNAkrMfGqSxR
w4u2jiFoOEwLAD5S0M+P2RSeqVLN620IFH69XZpEWSjdUJS74OpFoyw5ToTkqDbK
zZ2DqdlFi7ccCAZ+2bX9i8YPu0hCjeg/jUZ/fU/eQfYNe4hdgfoOlOde+HouzLd9
wV3dxZ1TFZndPDj6/BzMvAJFFuEWCT6Q+WaRM+Kb2xn5EMFKmV4vzoeoAD2A7rwM
ka2UqER5qwVNkv462evpnE+5P0C9PoBFzYOThjBsyB2d+klDZ1MWRvS9FWNHDsZ1
PG/6MhNYIrsXVS5owvVq54zics0+QpGm5USrppA8LKYdUWvNqqbSaNUCiVV7NVmY
xVUt20rtPVjxOSkBlaH8yMnPwfFzqRcR1GrVyFbN32y/69Vt8aL8zAkrorPX4Yi7
srnKndSybtHpzola0/NhxG9U83P/2FZpmpdxRw5YFZCoeLksHl9XMq6YbUi0Psw3
uY55QfmEE6F9DrTT8QjbJ63Q1V+A14i11ZqG5NIj+dQCTQDByGQzatGtTSInBJ1Q
Pn8urfPcat268+yZLvTIiBrLuYQt1P666tsCgNIWzB7IaopW769yUN6X2b/r8f+1
o3ZUGp6TNVXYgJr25TmZ2onJcfZthKzbkm+POgn5dH2GO1J8Pa9L9eiFcL7kP6Ci
FwxMgtWPQDacZ18O8Q9PxjcVtqzXqYh5UeISU6ybvKL4QkdVGB8lQhIN54129xNU
Z4ApYzscov37qHh9ciZNRWZd3+XwbdOfBotajYNHlgdJpVGdUJrJkSyvrTC7aUun
pOdHNQA1siLGsjScINqpAc5gGSMnOhRXli0jeMPNoJKJbtzp0lccdlz3Z0kiSBKy
wJ4/dZaVspApZ6+G3XDpyFLFoPBzgHkGrpw+vHxjicKg7xEjA9Wtg9Rbph8dtAZK
SJxwK0vcO7/HH0WCqO8MKYqFR6Ja5oKT8RfcDo8mvKo00u1Su9YCOjWQwmux/yZH
LqbMvA0YzxZWUp0gFznmpI1Sz2Bhr1c+h2KM1Vg4RD1g8o8xc6/9W1/uPJj182Wv
gi5/WQFsjbNScGl3mafWVZ99TzJS2mtmFZ26q0IdVN8QeHJr+ZWfQEd5UHF3kzsa
Bx/za4/fRln/zTwUCaRVe672cPv2DqCHvDF7YbVnjVdkdn4hoVVx0BfQXw/X3Rzs
5rRTu5yK/cogLNLZey3Np6JEvd3cJXzwa3vcpO6ryAxwPJej+fNzyXwFvaKCkkru
+T9oiwhANUjWmdrQtZ3WQeaa4CAPHdpfjANqpy7mvQYQjvndSjNcIUa6n0wlzBKC
j+0nHbmGYyQK1AwURVBmaGZiaeVWx/yaG/jzfMuDDMg/UV8r+zghisuzchgV+9D4
/CJFKBGpo9vRYoLc+sassA9NKdrFMN3vMwLZCz20WMrklw3NhAGtc2OB4qTFN63n
EkTSmm/4+YIIaECV9rfpWuOwI35h0YV1oqx3mFWdqPv5OpX6m65j10v57b6gsnCg
tUZ8fBy0zMNXBXt7dDKOEMPt3Qr7gCLMO4Bgoc6cB3awHav4tqeaoox4VFO4zQDP
e73cWMQAr/Trz/OMFgPRBLWzJacNI/4acGBDf+f4Pfut2fa0Drc5+64k9isWad3b
rKsy0Nz8ByLs3kV9UcvORMkCt0S+d7cR4Ctewexk+1N9FliaIDx1YGRhh0Wk/nYO
vVEuoMh26DhK4NcDkc4HeQj8ycxRQ2ADOC/Q8LktuGf9Q4Scb705MYgzKATeXJgE
T2QwBGwiGFrgKIwA1c1AtTvwfO7zlL+DPd6+nkuTaONFa3yvaRbEvBSYRGfVJxi7
WO6gsbJ6Y+wixqcNyfHKk2h6+ndghfiv/hzY8ZthDOdZlbvDaw9Vs3F/I6I/cxeU
F3w9AqvWJy9kspxCENL2iVwqR836e317LPHui/pcd/pUpGXVDt+BwaVlnGVHoN8D
9/0O6yP+FoqPIRWQOXpyaUj1anFzCRPI/89jxBZRVezahHNxywpVtkPzE7pG+EjA
EyCadV+k75JkRcWpA/nEMmbE8ILBOLmdVzMhwpiUlVFtgJSJf7G2HxfZuubw1EjV
`protect end_protected
