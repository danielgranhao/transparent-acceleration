-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
IibLyH2Jc1lPm6/wJSH9ypecrj+2EQdl4lOgH7FuOL6NSMq4bSgq2sFxuDUtUiHt
857WC3p+ZxJ9dZwuF3Msrwpbr+6Mxuwx92Ab+I19S9pHgez1MbS0bE/9zE14hvL/
i1Gpv4JUUXOoxGC7L6djicNGKoVeXPh9lOiUvnQ87/9koEXHztT5eA==
--pragma protect end_key_block
--pragma protect digest_block
BSqVEpaLpXaYE4VtHayTbQbw6b4=
--pragma protect end_digest_block
--pragma protect data_block
aibz+t/L+bMl7yW5Tv6jiQXC5oKoSH37OvXiyRm9t5sN8zlgnu+W/T2UbAWaoH4B
QSRXGJ0dz5jfnPtMLHDfJ8lyjbB/yd2FWSH+eXHGC3DvXrhm9kHVIuC4C6JAarzg
JdCMonaPoc86J1WfFPvxorC6mNNKO+ps4NbVVNvQjRcvYCDEOsoNxi1JhEfcI4om
NmmFwI/jrF9tYQ9U9O+fqaViwpdwQG1Cd+FK6KrEQyXrssT2sRptqTuoDHhm+k3i
MlmnnkSP2VFx4Z3+GrFpNbyFY4N6GZcMiVhcXnmERzF7GnBvynXpyCngTZ/+8GOy
/2M5LUge1PRABD/7Hh6eCGfEpdicU6Z8hh2SpnM5CiAd8KNzJOtVejcrdazldeoy
kA3DUbeXqzffqBJ7N6PgK6ooDc4ZMQcQmvw3HIPin6MDKZ5cJz6iHdemM1ZAvgSh
BfJyY95qBsQfv61AlexSDJEoO9oqpTn8rqquWbr7VRm5S81S7NeTkfNoNNkUsf4V
2vimvs8w5ehJPgbrPK2JuxWM2WCytu9WquS5+X3vZ6x4pWWVHQhHTDRLENYc38/3
AJcHUwLPXFEsV3gfjj1QED7/Uv1ltIsqxgMQ7Jdvdw6Ek9MF78wjZL8WIiKg2Ko6
8XaUCWaJAmqIorLtMkxmJpROKcfN8cH3tczswyLANOYl0BU0cD57549dOP/EiLHo
cu+3drQ9DCnP7me2TXPAJ9MNB8wl06P8gTXPZvA95nLM3IoaQehdwLIN882/o+EA
FK65ouhupfor+bSyzC4w4OIXRVdMKpJg9Y4htB4gpQGLeg+kWx8RN0d49nxPwIix
+C6AoBEsmKS3GbQnwrsj24M2M+lLuAzQ570kZyyFTRJsQzjK3lRaOR0e5jV1gMPV
yaYo2IPEyi1b47nMhLddvgnEm2Q//vHFv/EjwR+p9BM8we00UDrbprHxrS9q/wpC
TfXmZX046cocTJi+k0lMi8wMedJwKuO0eYRxTX2HOpnPAIXeWN+lIqovNxkahJ0c
kwETL8nxRG7ochW4bDaOAa3x84NFUhftUKZcIxWmJBfVL0F3vvXU2t1WeyAepMwh
Zj8Kdj6rohUyNaI6HF32KrUU8pCLtE5mImEAcCAc2jAEvdcl5Jk2iAC1JiHNTY2E
OZerpMQ1QPr70GnNGfAfsT3t8XzP18VlJWgF8yF8YrhrO5vMKsYfQpuf7AR7AxLI
5dYU0qg2zdddJlf2ibwD4jMrx7QfJGsMhVK9WSVbfVCzZjeWGOu3d9ROpnVyOVWq
YBmzc5koiHFzn6nJLXEzBXHYz/InQoNNwRH52qlogyMWXRlMetTOZ4kTwcCmcpt+
TQQiP5saLysCA2uEoM4kg3FqIG7wwXSrDZmHFNE7MQAoyt3WTp/faVL9mVFfy7pk
gExXq9W9CBSbqjLD84oED1ocVH1gOG9+x8Pyzo64Y6bcw4AEAJ5ajmekdYbVbOGp
ZrFMQB3ydWqt/G8jml2XEKJymQf7N1QpGHjzxwmCGma0sZ0hNUIwYeirNphM7DWz
+9e5+BfTtfK3q2XyYMtUx+YgZWXGXBvNT9j1gQdSPalNAiEMv3RzdFjkW3AWKpg2
rH9Dn/Oqkxrj/ULlGMv0xATpuDmVLrm2EqvujEyDizfLWuh7lHzE4ecek6ctQHZF
MOrUO//SajueFghcn15Ki3JHMY4tFAmUa1PhXfDNIsEsYZ76ItuE7QbMCDfWk2Vn
BZG4HCFxG4KKjSKqkUNzc5QDsX2xfkG098TSzRrfJuTOa1fJfCYKZWybDSc+hYb0
w4CJzBIs8CCDGtiuyQpwbeAkjnP46HfFPQ+1ujUvny8NKKeFFBmEjKAdK3Y5ifP2
BKYrsOre4BFh0BD4k80pug50csC9J6Y9gex1iQIstkUa+c480sGcvFe9od/F1NsE
P2R9cZ+QSGwMihV5QyD1ZQlLslyHpL5HMMyBRjVAJ/tGmiVbGqtLu6HkhFs/aZXD
4DbqAO1bGun7JIZq8BeANFKaHUmWVKiQ8V1HUSC8wE5qlXnwKSy+wpSIs5wljciW
fky1lbHmVxEdNvw546AGRBxuzgaLRQ1Gucw9LD0onSEr6AHgraBTr1HCEfqh5vP6
GZ08Lxf4KGvTHCjP0PWJ4AsoVSVil/CWL1u0185Cw27wau4xgwQzkb6JuUadlvNi
TtHEuBupOiOp7qSckWJgvdQ73hPmmmFNWH5+VP43XPA9C9H4AaQoGQjGzOAAsUo7
1G/YG4PGXMr8JefirFsDbEv4SQMsuWAx1+OTu/Yuzby3ew1L6qBfSfsV8drqGldu
G245E8clicGIGsRIUvAztFNjP8tPKp1HOL8322Fj29JQN4tujMuYnOEeIoAuv4Lh
OSFsetYWoPA6KKpzTtPzis3tKUDFs4UiXMDpE4W4WdzWGwPr1uuC5HH08yyjhFiQ
3zzxhAWOsBaTQk3vsdyraL1o3gU1bTxk67lQhHfcalvthEgIwxbVLa1kNck3lmXu
ahI6fBBtIkrvtEIqn1ilBd6RueVAMBSx2MXHPY6uLq7f0YWW0SwIZzzG6gehAZPW
9b1Q3CJqktW6NZhYTOt3oPVEg9i7kg/vOZf4vXacMxKHuZhIxjVwvm+gNAkYxBEP
REyJ8TY073e7S9iN9a5M2lmj+zWk1klEFg0ArX7bAdbVwm3WA1EiOQntopii6pBI
r4zUcvfwKX2dEo9B8aOzVD5eKjJyHCMzqu7XHNigkxSp+Ve9YXKXCtE2pTWhU4QQ
DGI8FbNM/gx2tH48aOYLwo7VSlTd9kXaf2AB6POzATOW75Jp5UHkiEaRq+rYcDo0
QCy/jFBHKadmi4sRbbHZJh4oFqW3gq9y7WIQS9nUy2L5gDgncTImTFcGSJjisFeZ
+sFCQfwulV+Z1qcSVVueaTHMNKIwUbrY/EKeRo7iRTvAp5hZaCgYWcbzO31ZQDZY
zPQswD3S1Gua6YddRCpy2gX6piwsnTJnbatJKXZ5wEDXO0A9sumHaSN5pAfOVuBQ
y0ShnOn+f/jvkNoleiHTcrrYnDzIYwdvWylPcDcgSkNLgmQhHHDoaOHKVThW0E2f
tY4QS6e//xFDK0zvRagS8mRJiqrgu4g2dVUQbpNlVE4kAT2eLKGMlHGW8JONJ6J4
21CrFIGzTbT90jd7qEOxsqbASDwtWYLCX6GimFxyvyVjyces7zkFZEVjXpi+s1mH
dkbu2aGG63kkfbVXNmAD0UqnuQnV58YJVcK/T/Zxd4jZtiXKgbTOduU9n5kZMaMF
7q5XqkJ/l5L/BkNOtsZz3TBF4Pqf7EXR1mVf0E0QXIBlGMkLS+vtOmfPwTaF2LDE
wZwMaqPk0I7HmSE0ix0CHLCzNsfYAqEaSu5A2+ZfybWDYU5qEtyELcNcKXdAKr5C
UZ/2xZXNfTpv2x2+BpZj4qNec49sK7aaQa7oYfDnbNmeXg8ZlY7aTj+E/8/yONuA
T39/diFCUkTFWceaylI9NiivQF2FdGquRw8VUsrVLWxFti2h8/PwjQki+LgqlqQU
86rQIV6jhuvSgq3taZtQ08QvfrUzZd8hpQLJAf2hBOO8KszzfxpcuboK0f/ZL9sd
10H7hwmjdywVvSFdhNWTW0TvhMNOz0QeSNwlupl4+xJBGyLep3Zgyr7ZHhzMaERq
u60w6JuigcmBS/7DGhVGzjj7nToLFlzgwQo674uxmfdK4ZQ/L+Oqe1scMV1EjXxf
MGxSY4VDlYw79Qaa4BYre+M9GhXO06Ed0U3wQuTc+e/GUMBkpUeHhLspqTGNvGvO
obegnM8xI0D1b3qf4txImX3xqlZhqhbNFN6PikahfpSc/Tf+9qgBIBlWKlP0FB/n
D2TXxhfwAozvrTQrMcF+Cl5j0hKMiXAL6r/QXYUHbPlU0AI4wxueeE1d058NwW/J
WNjMCSpmEIb+trQrTEHL9GmVjT+nUZWh80bipb3M36uOfP9s4D18NPVUO54f+CDi
S3dIutVt5S0e7mUWH5nZ6oqvGn0xmBoAuttbET08qmxtYZ761zgFZXHpqJHUir0Y
3YFlLTi0n0TyTQq59nC9fRIqKwDOf70GAAOpe8WAI4ftf63NQphnthDtNQPsC753
x6BAIT6g6donhlK+iqGt3qMTOhX+zdDW+KnmzbN35Rsbm82NU/VMs6p5AHe0Bw8m
brKm3O8Jw7R+si6Q/rnka+Nd9To5CFcFLk5hAhnTzOFtsw78wlvTEGuOSrL/yp+e
3csNv9mVlP2ywwWLdKrzjkRKb1T280fJm0UA8khQ+4gVi5i4YnO8+L7SlGnpWyz4
8zcf4tOu0Hh8CWEOKJbilBpVWfPOioqODoi/d5M+TWa8lyfOqLnajCiQh2gVr4L/
ac16IHmo58v0Kxc4ZM5SqZxQjLN5DPIIaJYpR7Qz28cdTxjvxP4HO5gjylrkzx3g
XTaSDwIvQfKVePEkxzodJdeHZXliprIpNyDy6SMNtZ00tp8D1yOGJWA9DACnVfGx
j6NvLG3PhKL/HW2wqEGMEN8xAiv/amz1bpBRaVLdf5kLIq1p2PpsFggi5NYT9Aur
0bNFjctYjK1MeWvrDE7CHo47+NlaEKTLJmHWdkI2ZGJyhevqH8JIMkbppdm9fRuX
wPa1+oYe2nJRzUM2ht94t2FGZiPYSkHSMWqzZUMQDdJUNGhffUsAgUTfzrxJEvFi
0fg4NPfzaPtaLJyXgWw7dozz0irV0YhRDrQrhGEz2ggWJd8zUzT+RJSsj3tlIlhC
lkFAukghVEMbAaI2gdwJAstLI2SxMeeAgpQOsR9JVTjOuu7EY++3PRnTuMolE78G
SL3ExwBaXgo9SquTxphEqGTtPMcOvebDl96ZxFRHwT7W1ACqQ2njwg4hg8sDVpHn
XsZpU60dFwbVEOmzp3wmzNTCn0+9KZnUeftOVu3W2Cdhj/pzk0ukbdIwK/nOfUOb
W+tcw4vX/e0jBsJywMd4KFKz4paatkyDe1xwreIcCNEV1VFITEqVFQ/h+CwDqwCG
zA+GVYVBIdhU2XmN6K1yw5Z8ebBLBsnFN72bo9PDLQcs2ahcgQBWCNhQfFvCLQHi
vmnt1u9rhoLHnLjY0HkOTXLinEg8bD71/70wL3fTVGJw2VVHYY7TLcW/5sP4L4jA
wxAdr2biwQGOa7jmqt3/1LcWsUQOB6GddAPKRbAzyiBRXxulH/iCiA3jn8flDlrU
agaket7KSG5NbQ309MRt7JLzX3zLzCa5YV7+B2PSYzp1xm/RpBJxsj0CoUemuUDA
dWxjq3ZFNqod7BULhAeW1MKa6WFcJwl/7Zoii4w4fnscUc+igBtIh2HtkSiZeXKo
+xWoWulmgHhcRu7UB3Ci5R5WAHHLpgfVqaGZFMge984tOmLJRnrebXyNqUf2QS+2
fxmoHhwyelSzA2uLvib0vTEsbtyu+5kKnyQKqC7QIsAdlnXBf6GYZWVPOOA+wFb6
051M4/gg5JhV1/kNH+0YADnJI4BDwG8gHIqCB12aNK7q/3QcxnniF/jr8v9jU7Om
PAslhk8o8lTfh7lZcf62R/ryu0P6JYpmWhqz5PHPIBKbyMgGBHU8wJ/ULsSdv3rQ
8Ufqnj4HhHCJe6Ve0KVDYTx9D02GOfylduUaYzQoVD6dbWiuenRT/adnOGY7YiEh
yzldQS2CPs+p0HVeI6iOPOU9RflrGO2PaxXNM5nUSLIn2xoheu8f6QA0jsv2UTaQ
0G7NOW3nWk7WN1b6Cvfyo+YmNmbP5bOSKCLsyY/re2OE87K/UlzNk1UJHcoiva5K
P+z7sbNs19daPpBv7o4r29N/AoPjsiW8M8NMs5r7IrOGlRZa+6cC3uVXHWTgBnpp
sc1Fa0/IdpTg9dbim7duTP0o+y4HRAUXrB2oQLJCFBvFFDLM1Y1FNbvM6EhTzdzk
23Kir8EJ+Qw0hbWPEyS10QJR1TYRjutTkluP+bv27WDhgUGRADMWjhHfSPtlFGf6
9JiOQki+UOnBS2KxBtTAglRAxKXmacMY+DfwfbniTSQYqQ3hwfCB81YStvL6/Prj
bGjw1yn+TZkgVBEX38EwdUfupx9k/8vR1GwLl9/prKhDeKs+uGJzuA8ilxPxrcDv
z5tYz7taCtBS9/t5njSyXMbB07d21Ru+MI7LvlifocRDMUjV0dsWgXUT7/YnCCDN
Zh9i8uapT9KDo9802sbSkmXPLN1UcfiG7YX5e0T/XBUbH4w0s1/Z6++GYd0Rh/jt
/2PPSFyx217QA9+wPJ4Zj1Rvi6X+QTgqBCbGfKybMKCydvH0dRCR+aCRCdfXPFU2
lcPs93pfZI3919XUoDJAsGWbpoyDRSUAgTazjtJNB4uSjgLxG1gQLpsTGF6quUt+
AqoSBVPtIXzxuyoiAUSHHDH6tVCiS8qXgbz/yIeUNfrD5Tni1Kf+XhMu3cAFku4O
hsp+8uWL7Xo9D1jwLweG07AvzmBboyt5jIN2WLL+NlTwL/msPb5I5xhtaAlnSIWu
1rtafYtIfJFx3W3hu551H0rg3n9Dhvuuglwt7KIyhHwgu0bOOCJsauBLpMroRuQc
mABlRS2PYq+j/5DIueleowfMMk4TJZUv14IgczEwniclTxGHHK1W0GG9B6IjNNji
CTPlkHP7HIZo4HH7SEkJlySpqpPyDZKN0VdbPxedlDC4Qo0CQox2gXQ2ZJzzTPOC
mqNbmzAyGypHvkrp+Pu78oE4mCleR+E7KnpbMAOi7AbdZG7fzYqz9kS3IFBrCOcV
2StZNsoArP1kE03RAwlJKkTgN/PdBjrEBfTWd2bWNVJfX0/6kyuPXHPX0PxinUSl
s3dOYbEePw4JKBy76MFIp9GPyiZsClJf9/lww48/A70msEr6+KGfhBS8N34bBmjd
BjME9T/QZF/JvzThbovEuOTIFdOLJX4mz8xAUnXbtb+YDZjkUlKsJ4nev77qfChF
+dqGVBQRpySgw7EFtQkajMaKNxoub7WCZkld3M8rV/MORycmKbWYnliZ704W6ke2
uQnxlnBFSyFZ5P0WJb/RLFK21nimYvADSIZrYZE2lTD9N6nJGjkd3F8mULoURrsd
uwnFY9uLtNbfVehCws/mqf4Y5DH8iDtWB5WwHDrr2zGfbGDQuPc1Y7AwebualMBq
fwG2FZcMVrajooBbCDbqSTtseCWdk83aOo66fjhg/QBfmHv34M/cq0kNlKPqI1/w
4NluEsdFVXa2pdf73UUhJurzl8j8O2BZikaKtbfsmEzJeH6V9swnvWF4gEZ4H8hK
abo9ZoOpD1wb5dpiPXy+MZfSrdTJdkchX0Jxtunlm72TKsztorWnVTjMEHIKIAUm
FO8vxRP2cDIdaJYQD7ItJAk4sC3pa1YHFuUXAEwjdVxkGAEfQYzs+Oc+7SFEfJHn
A0PHJw4YelNJlvB0uubk5MI0oYh+TU8erdeagkGwgL5SrFO2Pon7mM+xi5NCLbGQ
d4RBt3Znutc58gFy0C2dA42oqpsvs/rr9BOv8x4XY069r9WfvQdkhx3XL3ya8CHd
+2iOdf5pTnumMupbY4MfdnQvkH3pPI1BW2Fjr8/lVPXPyhSjbtGcPHrlKK+fh2Fi
XjHfnoaHBqJgzqDBPvQpugMpUFvQqnySfPfpR5BnF0YNGfT1tguS/4Y0AxzO1LIs
a8lexk1qUwcZK24ehSuf9A4tu7x5pjjznm87ZSi+Eeorha+/L+3v8QMzCXQl6e1c
8+dslYA/2KTbDKU8HYjM52M7+ApTuN7ChSiHBSf0FYvbgAhzC13k7R7Zv65TVq3V
hOPYjU5rekqABNQVjEpAaQ4GbBrP7kxg19n1KqynvPhDMCuO6VHngFa0qjtdYJ02
LQCQJPp2XGceBOdIp6ACwJ2AsXbpUNCKxtgN9LW7fhw3oOKTqmppHVTSTrJ8embK
cX1o7MqirKMmalSwiETQuK+pBL+0hofTy3Jt35Y5uTCENRhWbME8usP6L6/g1LWf
SLePTTXmF9cXZwSXpRmP7fIZTK/+42pV9vEGp92RCa7QZHUsrwnRtDpQNBD6zDkN
NfsuxAjZhxYpXEqBFfbdRrjSGAQKJ/NetmjdWYz5bVTKgh2cxuM9cmNgxUDM4n1c
lmggYN3zgAM84Ye62m0UkcD2dO24RR3IFqg19jm0VOTTDj8QdQZFGSixrpzYbuw1
b/ZyXr+5byl0AomRqRSYisbpdG1oCQUbE0YLhKSgBfiucWQ0SSF8CJVe2jSBYp6v
eeTid7GGBrrnKWvejU8dzUURa8LfxgMyGtKgjRPSmELQq9QWqjKPAXPM7lZiw9Tx
hcYZSnNbkRvB8Jf8eIPvVagm/Cb4KY6AANhlzY+MsuDxFFx123vY6usk3x90aqjM

--pragma protect end_data_block
--pragma protect digest_block
zLfGHjdXb80ijQ197FVsyvD8Qxg=
--pragma protect end_digest_block
--pragma protect end_protected
