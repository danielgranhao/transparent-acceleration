-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gZfQmvZjC21R/ea4kuVFFBAMc5H8zS5jkmyuNTNuWXWoH5rLfKLBSEOshnEnn/10
UFbCVGsuRlYP/Xc4Z1YlSQacCsvdNcytf3Y2kHtAMFefOTG9fBvCCCXnNj/OUmQx
km1mYZ20581h4gElPfjVRr0MlYrIGXOzOpI+6oPdgMI=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 4821)

`protect DATA_BLOCK
olbDsTh+gPIw+XdXT7h27qIPznjIsaafjGiUaRLVUmeiDjBYb2+pfVpcXa+GJtBt
C08S2iNQLy8/Apms6vf39Qj3IAlmQrRcwfA+8x3FAMZNsSVxpf++6JpwRS/ICpA8
dCjAc4bSLfU196sk/IC6Wj+IBX1p/RTg10Q48Gi/v6EVximGXSlycMUkgA7ldqav
1DqqoWYvDm+rNI6yeybW8jKucez76SIJYX0DUJbrbGkiz2PyGI2ra3IShVpY3hk9
KphtZLx4+7ewzaPbjKHVE6hTHR/rQdc2yzVicqOzpDz6Nz70p0WOOjHwLaOHPqVl
JFbQaeFPmJx9MiQIUxXyV+Pp9X4H62NOheE57gVQOGu7wZtzEmG8rAvPtcwpZK6j
QD4oxQpe2F7l7JV8yeonmGfbmR7wKto6Azx3v5p3nQ91VHfyxyc2fyAy+KU5O88n
F7acA6c82rqAEAIaE+eJxdspwv+gT71wdtADNbGj0J7/E8cv6x3ty23pMglHnrLK
FH5/fwkvXULr58PM6DHzAglNvuGJuxwaXY5zubKpy0DVeuSeLI8wBhTrHBYyNZVJ
FjZqSRNghMhjktuwJ0CNkuwdr31tZAfZiWp+l8J4Y2ygpTNhj7Fj3BJtGCWVy37/
6WqpCfFsdBOhuq/lHDX3Dqlww33Oarqr11L+i6hE51mOPHgmnTeWeJQ9PNbf6I9r
mlDXZnJcxyCvu+/OCGEY6uqPE9g35nKRtDSWR5ez+L1CxUZaCr/HMBsMy4uOBehf
K2AWqsy5+IWjQobpF1vytB4XomBkU6uXtzA8T/blqJW4CSGRDMyuYAaghtrrTJly
4OTbiINaHN0SVbLmjoxtM+BwDzhz5cAUcjySAzTtuVjLzPLQGWgqsW26W29zsQdS
5eBwyVNEJyGWD8XyXrc71kGeZQx4Vpz4f8kzPeYTsqZsE3n8Qg91IXXDxEcGcxpW
07UL4mWMV26hyrZB+17jQdRfSt8v5n4W891Sqc36woET0z7RqCUQbMKg+zLBMd7C
8MM9JNOKa11R2P2VcsBLsxnDokK+C7cXPZIjnpQ4l2oG2Uqg8Jen9xQA/YhED+MP
3RL+PfLpYm0OfJgxUcmVBKkYeYGrOymK2YWCHdgBHH3D6IHR+RSPtm5DUapB9wMX
QKTxSTctiUazWxYlovGN6z7VoevEETgSV7mVimDm0LvCly614EWLWYDAPKyKLX2u
Y5QmzYqy4ttZpp+s5vZX/iz18VdLfMsS5kz2fbunWXUT6LDGNvNIOxg8piksLXni
Cy9/pQcCTlx+D91uvCm0Tn1GwB9Z7LYizTIVZASQ2vCADJOVDTlihsv7YON9ET3J
1moVPjSs5IQKHSJ99dMiclM/sRENyBmyZkrxFDUq+yqmb8buFZYWU6ZSvZ0SWyYv
iPFZR1kKx+ZHkrg70Y3NYsBAoDSEAFVZc+nTeVIqqCWbE4ldPGm5ker72osMN34M
4SLQseZexJX1OMwMi6j0sZiRpUJMecChpdK7kAfb54Z48KMmjsZFYgtqiSzTV1RF
ft4dxGKrsBLFaTRR5agOYzAkRwX0IgMJVdInTNrhwgRGjfLwS596MPAi4MhRy3Zc
YZEuAgK+gflFLvAEIxc37b7Z1zgb5djoGF0nHBES1/WYY9pYFHrMTTWJr8wQpORq
LnrnReFNTWep7d41SpjQV5IhZ53l1ezbZZ1PKxMVXGH7LmsKMy5RfpgYouD5iOpy
89CvydsWAdj7409q3bRsIn7qcUnmFSXBchWdMzRhkouLRWNhdeyPbZJGxKu7cNux
uBPaPSnzLG+D9VoIUXezKM10kS1L118UE7MpogrmKmMXagKqJwb91I1lwb3HUZmH
MzcY/Nyhj3xi6TUVrkUQ2H77080vUtQAVKbPIzd0lLBwAn2N+PKSZXUX6zJzPsRg
IJ1KOJLYiFwV/7b+YrsNbzVXsPq2cKeMb5RJ7z5A58hBrZsejGxqpNcSWsoz9KTH
5fQyzFi12yO2wbhSI5aG+jqUK5O/bjh0vPDNMQDHdLCnboHJFeRy8cPJs4Iqku5G
wcmtGOhyIUStLuYoYlvNdOQ7bA4YfqpTjwTA+WVq8geBJE0EO0xcC9sxoTLOZlYh
s2m2cBdi7pvl9BG9x5sQHXIgi20tMx/GPp9fkxlSOFxaJ9dNt9/5Ck1tCNkWlzrG
orSzIcKoG7fW0G9CyqKu1Z4uglaOi2HMRP42S2E0S8mbnWdbY+jjYpagGPTTwg3v
uAfZP9JRhrsmfP0kRyutlw9g7wkOyJLSeTIpcKMmM+rC7Y5bBWNnBd6ObYhEJAVJ
Ccwm/zxjcyIkE7AGO+lShb0GB7aVelJ3DeehWKJo+voAbaYDhWCN/K7btE8m62xA
SCxO3MF93X9DSHjzWqiL4qhZ4qr3Q7GGgBDTNyaMy1NWIUfmCqxWKPsmbjUHDOsM
4EmGoZsXKf4mRt1QlgCI8GdECX1OlPLNjxt42WIia4J7r7Yitf99tMPlvqyapSXz
8mDJ/Uyr89xoZKoTPDHr2azBx+aoLbuJolwtVA4MR+LUZMe1w3Brbw8DWWIxeZmJ
0Vd31eeTpzW3z9FrPpJoF20v3gb5V3n1FIWQIfIopTA8lmhaAXfl39GSEagO/M4e
A1efXiwgYRQAZP+Y1aL8R6qMzMhyshu0E/KCtyF9uLWCaArObL7VitPWa4Ps51MS
9yRVM6h6L++VOF1HSxSuEL+54XMMjYr2BB71f3yizXPqeXPrOSfreb7sl7BxqPF2
fpJxV8lo9QkuRn0Mh1416Hz7KleymQ1xHT0SBXD6XJ0PSJZnawiKpLYUNmMZb+sC
eOaxx60YYg6KWFTHBYPkHRoI3Ig+wLpV1ZTUvu4DBrs43FBphXmCFLqF6YQBFq/0
NJRh8w2x7hucarpqoRjE77kRlLH18mebH7yuDANCJt12PaYxMGdG8BSzBA/CxyeK
iMpz3YDCXyU2gj+lOfRUQ7tS90n5cjVE0dNqyOO3IhfuSNWrkkAqq5kclnj3FrCw
qRICTCC/NrJtHE0XPzm3Qx1mOz39lu54okia8PHCm+cJPZTbre2ICfRSIM+Y0EGI
c9OSGKDx3yNCLL7T5C6J1ZiqG4/uDxAQbrK2gtE/ACgwjcaxPreFHv2X7Nu25u9x
1zGPf5utEeligFfLxOoD3G54uK4c5NZDmVjzcjiRW8y5IYNhfg0TrcEHTHYNc+Wj
77TEXVYOBjApAPqoOS+D0lZGt0trtWmmkcK4b6YWIoQ/d6e0ujdYpjf8NTI8lVz7
X9oLPE8pt6oMQIM1L3r4LYsomcy3l232QaTlxnLnyVUvaZnZ6fFlzn0aCwCZC/jh
K5ilyQzIohxI/ryxZ/YYD15i3YThEydeFuJGL0GBvfrXaxgaXbWu7uSPJodNc1oF
qE4chHaksVgoHN4nYTeXB77kO/DhRF0sECfRzCPYxoYVONokwfuUu5peI/NIH3dG
8q7xZY+ehbpnWXlnStyiHYll/rZdl+AaK3jnq+yirrDkfRLmuM5P1E2kkdzHA57s
165A4M3PvlHNcLZagQkioZTWad0vj5zUX3I0FM0/anQ8cHYeYU+U6YOzj+OSfFWY
isVCq/ZOCxThVaTGyfVvz94wlHMXGjBd869SatOlAb9cRWN1gZeIqQq3LLUJiBq6
Iw0CH5J1bprNfJSEWBYBlT2izEY/TnK1wyUlqtA4S1a4d5kFbzudz6PUSRgW9k4f
W+1UcDPMSAi5+jhrmMI7e1W+q1dAayMPoM6YKoH07LyU1ekXfPFd3+MrxRFnwwHq
hByEhtC8peTl1GQ5edRM42gEpQ3+QLrZ1byk+q3ZOBqpXFHzVE/aBV0gEc7Oy975
TMot+luE/ZgGXCai5mT5BvCFljNoLCk13/aH2fD8ESE8p3k06IDjWn7KKFg03T/E
/yX9ByY0xJ/OjoY1zlJi2xdb9frokelbymIQAKRCZw/r8t577muL6dQJt1eGfYUD
aCswoBOhwyNIbAOjT9XLdpkHqHG3vufcltEgkAn0EivjGmhwRwVxO94tnrKT+Sqj
OyPPivTOiiI2x3iowcDsX4X1fbtqRrkludOSSpiWdDd5R8AB/3X2fBF+N//vbX06
ZvT2J9dLWWZd9wYGzrx0P+z02LXCr7HnYt2Arco97RO6HPAeiTcLhh/Bom221oQn
rYuJSYokoBAFFnhmdw1IFlGYgnBHT71C2vfgJXc3uespOaMC0tbuymjbXjkqWx1H
mji6bi3f+5GKPqVGlyyZE95ugdfa6mEYLe2E4Eo/K+cqU/D/lgL1gXo3MEZ4/Y0+
Jd5xoLkHSWAex8CM1IkiFD7UMg9jpvHgXvF53iBJ4tvhAWTYYKs0MLVqlnfieZEX
YCb5PIZ/RRDb5EuH3JE/tY7OQrYOFhXP9f8iexazxzFOPSwBiI1qK6XM8nHRYUTC
xBJXou9t41Px49URi5ST03FIBRuz1CU2OorUwtGAVdvKUPyELfFa/qvws61E3Cg4
w2radjCdw8ZpphNAIQ+bM1oh3/LIv39gHvSFdJLsLeypFLzEzP2ZSlnK5gY+gLx5
5mGiyvbh/6gM66O1iIb1I9DQ6gxUv0GzMA4ygiREYOxNqORJhvIcSkH09naxmCrV
3bOysLAItBLELgHFKYueYVQ/30BDSzwnlXmx/PcTuAIdhnZrzXZI6fJiyBLFaPse
ADC3imHVQH0LPebz+4KHEslw09w2XwY8zbdZYZstv+Qw810bmQxOTteqwswgeGAc
4+msRbE6N9Xeu0byrTaiwSxZe0AGet/lv3MV+jdUCvacjpBYi4nEgIIGV73PygCK
BRzXY7SygnjMtNnYgLeQqwq26BWbTyBS8IGLbf86cbeyqnGNDu5Q84HRWR/2toXY
XOxWqLkGpXaSwPeJ6+HoIJMA/65jI92pVtBLnLz1580Iqd/WfnmzzEjOAI5ahXNu
EBor8G9ShDLjPXUgayCcyrM6tH0+ajBY+2NzHj2uYbSQyJAtCDvM/C56NlLozmaV
5VPFa4F1z1PVUcTAWz4qxL/4x0ov8aX3CPyA71vjKgz6diYydd0ZHyBlOjONNTWm
ABm1DTatb7hisfEV1FinadQMyMRIPI7JxjFDZVuc/pdOI5SGDdk6qJcAsrB6V4GP
9cv9V5Fvp71dvDGjyRHW0mGvcH4VyeZ9P+V4FfY6+hx2VFARGLy0iGuhtKOTLrVn
ck0HyCOvyPU4w3bVrXvcJ/hAQWT8Lhwm2mho+i9Tr+ZP5LEK47nQniMRSEHDTpVJ
MutvnNeUd2F23et5KtuwdYnxwFCQM1gSv9dp9A4jaevzHsSJF7oyk9Rp/0CcGsJX
npT/Yu6g2NH59a/Dh25GjQKUdJ+JhTazU77ljQb3vCOyP0mfJFa4vEt+ZeBMnvQP
E/C2l3SMQRbR+TLR1YFy43CuvJmGh5W6Ko9+DbP+Ee8mJdoVAYawdJiCLvRDyhXc
sZMhJgNLIrewLSVGNE2lNE5shS32X+cnWrWj5uGdv4bArFvegCu9Y9UxOQ2aEucq
+jIyXoM3OPcEbUiX158i6uVjHRToMfdez84uPdMb46sSL3LRwh5ixnIR/g84d/pb
xY7Oh1RWL7pRRASJ4OaojjFXVqnbf05Vycw9N5KeOzwRqxEXFrL0d4SwDLm20eyS
3LPyGV7RW0s5Ln0TMq4KCH09kz4T4dTA6B1/mC6Nziq87adwguUhjEcggOCgpfrx
beW61+YzVvg1zvVXla4K9eWkGIKtFq/SMpJXO4wTGIbAkxoho5AbYYy63WI2vBHf
ZLeJSzIr/ZlGws5YZg9EhJLeBihj8sy5NIkvXKkaj/YT4H/yrqgIGIKKOr+2aJ7G
bP25zMTxR3ZRkM8kwuiUdWWwfcDh49G+qZZoemJI1vJoswVRIRLXcO8Tbjr49DqV
KhyufqgYJcJOYT/b8uRpQgjAhlooPaFYVErKrtbXTko9AltuXoRGjPqKC8y96qlX
zjJPPn9vOle/o7yU/yimI2ABFR5Nn1CmcUPQ7+U9TxzcaZT6FZ5bH+xmPOPk3hud
TxaQ84APVZjc0ysrQBJzss39R93HYVMCZhSnOqH0XKfalpq+Ip3fkfMeB/a488go
kdncuKtsoHiuY0PBmlXJ9/sViYxLO1InnFF93TOxtaNtpNVqvYpp586tRQfBWW0/
NuuPmIrwc9qgGtdPSclsa6TPBMW51nJ4/7Lz5cgZ8j6198x+3A0LQxv4OWEQe0CX
OeyZ4YhWQd+HJOLKIID8aMXqCFouBNNVBeyKePFpXMEg7JFdeuRcQXonRdhximeM
TLTv0fvzOLmLB4yN5zrV373Dtwlgjqvxcp+T6JTAdeF1HXxcuqMn/o7meA1Omr9q
CQcyxhjZesS5GmaEUKfY+Ni4J+85Eaz/Jul/TGoRtzzHC2b42k6joltlFcmbnCBn
+D7gzHHlzjHKDRViAeyvvYHfaP00ijvalMjABDyETnDEu2hw9QO72zYMIk158xJz
`protect END_PROTECTED