-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
UxwBBrgkqRPWbeJ4TuqdYWTYCn3Kp5fz49be2FhWWistPvQe0mq9OQ4XZGD1R2kM
TxE9xzSCMPBHrNhLmVDtnXQROc03fwzIt3kr4/2WnkjHz5fWul4oaRvk/U6NqkFK
Xu7k1WOCr6r1ThdpgBDA1mXkbuoLY3MwbT/lLIED+f4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 9504)
`protect data_block
AJzy3dY17PIbCo37FAAWLszD4oQe5Wl/oKqAWVRcfpI0q+oHnZNWKh1UNicEsLs2
lnemLWEMD1LpSpDcaUAeWI6fmfrftbwbZh74cGzCx2m0ZYpuS8ly9QMzPULIL7bC
zYvRFyvlMRlAJGb0OtNr/cZi/a7M9QUczZ0DOxWWRORYNuNikhx7GzVRSiIvPhA3
d/64YeHg5tzSHvgGvIIzzTFApHsLpIRMGPorWYQ6do2ElOCsQ1F6alx2Svp7gMLh
O7ongGrT974zwLN2bxzoP7Mv0Cxa+yCzXVpvLeIMMn8gD+qrKhrfEuq+aR4W8D1E
skBPenNC4m9vHMDi/IalaRhlryxZn16at4/aexxSdDdlf5NqTI8n1mBLEtGjNGWz
yKW3zZWRvnOdl0VcS/xWoH+nm6EiAJTa4vfU0j6JGnb/v7gr+kd1Nbw8Il/OyODR
leS8Nfye5Sh2JpruVQuWLejBT/kje2GE+zFGiqeC1eyL/fphMFCQavW43P/n6rO6
yGGHng51t/BjrlAqadaLLx8eSCZI0LUz4Q3zd+p8WJtQJLoV45StyjGgBwKik8wp
hAJxrGC08pHkNCjAXbFcfogRb2lS8U17a831hYlHKwswWqb+FXBJyumUH9as4j1A
raVCqby0+b+JmFmN2R+JtSm0L1o6dclSjTsJN48LTdR52o05CDl/Imz4rUrYdtCh
Z5qpCQ1/gaSH8RkgivBSEoM+/B5gQjnShSPeUl119vLnhBDXCwndjBty4bJM9D8e
DrjHEwDYasBY0nHTtuaU1w8AcJQ3KZirP9T0HNxWsJOWGAImOkTz9jmVvOh/O9J7
dvADCbFzuIB0YZGcCid/iXw1G2SAx0jUuN0doJP//m9UfL5FLqC/tYOZS4Tt2eN0
mqXtbZHWd1yHbsmxnLDNMnIU/fRtBiRG58ed8ak2KvvlcX5yOT3MMva3P6PdmQiM
RBFz6HRimlJnoVzrOeXPmJL41rAZuga7RFw/Huswd9vNWuHpAhVZstwtGkjfWEBh
Q7+tcMKMDLYJwFlcrxO2oSXYHry5KLjNoviSZtttQrm6wzL9c7dUuaF1eOHwzt8E
JgDC89Hrje6wplRXkhPRDridip/Zdk/qKs+rboymL+042J+Uk3LPZOAZt6ytZYsn
RT5V8ihKZ/nyo62SSVgp0CzFlePOxs/O4JQSyvLDJBJZFI+z9FA3UZSAoj7Ip1fR
N9FsbFVf5rkRLIJKTRz1e/7t9TgFPX7vjjlrvoHoUWbErmWhEEidOUhVg4Yp45Kq
6DoKUoblwZ6mniIJSwqtz+SDHnCJZg+SqzT13al8AyX59pjgNdnLhDX0Y/ZSHmft
eAy0sJg9vnKddlFLM7c/+pKDJo6KdoTuevKokOko65vO4kkMLxLpKqYK99AJOqDt
xkL6wvRUTVcT8TZzaYvz18GxMoEVJQ+1l32V/0dfPewXKTZcqJJQ43obXhOrnUTS
StovEgGJD4jw94yG3GrbgNnBsKOtJPH6OLlCWz6m+jMBaHrjObqdIgBCLuj63vec
ZqMulhm1vPKyjIH4BNaqTOAolbP/J1rYy/39B2i7FdlAUqtmrAGNj2/TjkGd+ATy
9/KfXBD0N3D2rcluVRXsNGHu8Rrh5XQOzbpfDyb2rU5xGXPOYgzkEp4najcoDSxM
D958YHTADsjpOoMiKOT9tuXiw5vJsjQcJBNG/s9A0KRImeYBS5ds/JErrPLU/dya
Nbx0MQbAjmH3/tU/maGvbx9lvFLXBjihZaz7YVYlyDdGopzZXMlZJDq6MPitT4sw
jXGGi6uIC2YNzDHUryGV9A1Ff5jar6vFE9dT0CiVqJrQlSRCxmn4lvfLXCadne8H
ki1KKXr+7DTRNdozDAUoPyUcC4KYVK1AhBPkRnYk0X0LRTbZ/v2VpAthC/bwW4fW
VYllhxum6gTEVjxhG1r+fX8Pis4ZjhA/pKRbannwUnC40J637BAyHwc/syqFJ+Va
/B0RL1PgV5ymsfBYc8kE0FvCTFGl2Np6bC3xjs30d1lyOwptazLuaw7mOm0wSbDY
VVp9qcq4jxCNgxJdzkFovxBp6iUlAvY52CepLnK+S24yNnowm+v/XS/L1xBcpPO/
2z9URLA7Nk+6vyACjJgwDrpSM9G4ab/ZQaK6vHs4XI3j7CXaF2PPaVR8Rnbe5pH+
P0n4FeT2tGxpp053ZAjFMpluoBCn2YX4hHpRXCXK0PHteHSbIcoUrUzhxTh/Atui
bhUo5C5jz0Ev3Ye+noH3TYhKiYro80B3XwVYsc/ieGDVMIrYwd8cwNnbDLc2YL52
+ItlaAYZbrBfWKLZhiS55tPN97x3QZAeRCdKWkX4AN6MxzDSmNl3c05R8w/uuZba
sssfNq5kpC+FQQj0XRaDdoxyk55KeSxcP086o/1n+WIqLdGImVLVjPEph8J4r0KR
iftlEoeia/cZX45zptW6cFk9z5b9N4HJtifVCaXwICi1F9OO+xKvu+xoN332Y0t/
wALSwNkkuHkuqvZXMmVAPspLQBpooW8qJ7oUVTVExhnvW64reqdvODj0HoCjcCUN
9272VWnCHXLI7ISFZK8+ubOH7/OyXM2rTxMvSVdarUKybtCs6VG80Rw73NW36yCT
QuTEPiFj0MwTS76d5YL+HALU+2Vepvy+ljGHZ6txRB4oVV4FennN5BjXOB4XFfIN
d615qQULLxWMfq8jfdP+qvPBDvYO5eEIxva6ZGvac7nGmapTKI3g1ZHqTsqvXYqy
TRd/4z1GfB357tdVmGoxBccLiu6ksdP4T/SNw0AoYe+ShvL7My4fcuwLjCVX2aR5
O9vTk3a/sc67sbg/5MxFQsOXvSqKXpxJLkGfFJP6owHi/WUX9sgSEuKyh3tNPUYW
RHqdNBYrEMXSmRpYf+30mg5TWgbRhPkwDe9HlMeTIlcm75ZOc737Lc1TTDcjW3eW
yCs5uu/RqlbmkiP7T04Y6w0mIZ1czV+eV3s+JKM0sS9sOq3oPkM8egMbFG6tvFvj
9SY9Che/j64QkWdZmFkq5WAfNYX6O6gApI4V+R1uGKRi0nO5hHZbGTZc1yCyMtUq
vA0yBiLNj7VW9R+Ory/XJ0FnGjjQXhQm7t+rfsBVLPvwlTPNJhy8VS7oyCYfQcMZ
cWHaTwYhEhJloHR89KRfU2lS9QYGbY4HPwY1S0ZnFQDU5Q5xEjEZZLIbLviRi5KN
kvGyzb2unTcMYWazf59Al9mMUUuyZC+VSpCCr37ll8ZwhsxlX7M/fnBGpH2yK3JN
uoIZBsVBqiLTLRbhZTCoy+P7Aya6xH0zHOY/UmJKGxFVJwkXBIYq3U0zql1xzz8O
xenThOSnZuFBMntEg/n4nHDH4rx8w/gcpvOkUIb6MOOk7qabRv+6U0zg+xiBcsIw
Bu7u7M0LJZfGcKcX0hYG06AxdENWO6ob+6SM0pBNGRmalUF622HDnJ6VQFezLiEa
1NgZnqkBu7QNYn+ohPIsI9MnFTxcO8w1MBV/mEKf7S1UeC2I3pElCJvNK1noJfUc
3xgGapTSi9WdQvxWGvayBJwAzCwatfn2F1YtqGCyaDGWMlqSRS7He0Cr9mOHluGe
87TYzzVY4/SqOKEnQVzu7jvY3HlZHQJvSetzlJapQ+GQh92phr92znU6+oprtAH6
YFvC/354dTAmdkCaG9BsvxbfAXWXVJvFgT81kKMYm8D5bzckkVms5+9bxKCkgpQE
e5kkPQ/rT6rfqbGmjHPAG9TDbhU3Mh4o9CsjirB25wJSPrpV6cGC+cpMCdnm2yIJ
orxaEqicBhLk5kG7ugiHKryc5fjZBjFcnbxlBZLpjKReWUlGjkojAUFuRwnXmcAJ
vTtaLrd53oN79YeuppArW+wGMhoGGBG7rn6Swku5z+IpvS1UwvmDiM615WfY6dKj
nz+Y7D8T9LgllZnGEG+e0XScuNSkTvdgPIILXFSM2ZgY/jKFvfWdcY6AkyWKCdLw
o+XAh/1+X51pDmMqONa3uNsGcfi6oJOC/q2CY61AiE+tzsRu1CWV+bHo7JK8KdFK
dFZpNWR4Qm+ZOFKcIUHN/jj3LUaeqRQrvYTI62ZC/k3RxARn45dOJ65i/tda0SNQ
pBTJlJXOlst0Q74x/hoNBSk5HR4uSHmBB8n517IBnCDLRTDf+JlvTGVnq9jOF/Qu
du8TyB7fObWuedsMVDJ/kAwQkvYQNax4fs7WRQf/kvDU6s6zWQzEoOGwHsxyTdVU
dkRfS0OcepYXiBCexkQhTWWZbqb5WvD6EzTX4H8eLn5Z51jKQwlo1ERM+NZYJPfC
lNqWc3RYyojjHLuoijovGOCFVM60rI85X/0YwSc5IAg1ReNBhQiUK55JmXD1rrF4
b8bFGaAHciaOgHJWGIjAmw29OxhXgm/lNXuoxxIBzkCalGR79MP6mOSjkkmMpGjz
6PX5htLn223CECCvf78PKsuC2FnIxp30A+Dt15UiiJLzakHYFaOm/d8Ll5bYn0vk
fM60R+PRN3Nq0B/T2E219831w8dZaiQSGWwECzLf+/DkHdze5PD65/qHGnOpj316
E9/SW1HXHK5QudOmA733xZeQxucUdwlYVBk/qAIh08nJpDe8cMcpmEFz9cqnWBE3
1BN4n/jz0pVShrzpmU4u9Dq3C89J3fOqzhbyLlEAmfpUXdhyNzJIZydlRpK6n8nV
BnPaJ5Atr5F+4HrliHHyj14LAWKebmH9ALIj/gUcabVY+wYzBpd4NUd9YnL9lINc
i7eMLpGGsAtV/A04Y4Q0Mfqy9s5fHKdUpkX0DIBAiCpAHQBd9UshNBZ4/Hv4Nb4X
vgobY7xR83MJjAGUpi5Z1Bn0Ui20K+k2fp597U1Z1OAVoeqO8d6D9Uvx1foPjS0I
8V3r6tVZMaX6gQtAY8zt1QdhQvEJG4IVf+ueTOq2+zEC7bgBrcRVbk4HIDz8d1BY
p/fedAx+0ZhDDreOXIekhp1vk0/oxFnNBfTzuSttX2lJ+bbY2XTk5LbUHsO+etaJ
O7euBqdae1sOnp5JNqInHQvJzCxXeEIoGjYBaPNGjWZBfoE2J0Q18hT0k2QBrcT6
5ujR/pAd1VwAXPkXdO38+uh2R8SpQVhWAzDWqrzXRsvFlSq+fVqsg0LkolEs0M8H
wZr3tfStQEJxcsU5ZekV39ATgY163apKXe3bRxfAcKd8h/pjGhUlg+m01TGSkjSz
QVuuvx0N4kswJphl806vCSbx3PSKaTSHPX96dZZEueRNV+Eq+4nltqose/z3XHcm
aJoHC0PIneNkN5mTuKnN87AJEdZIJBd4Kc0LI/aYdzQ//DR4HLpyuZ7leYTcWRgb
hnN70LCulNwhSoR3W5YAMmJ/6k94324CF+hbr08ZLktRDI6SdyQ4jPWsAa9HP8Tm
m8HIlRkSKkC0fsAbn8uS4jCo5qd4yP/kP2IWeEPmJWE7dJWW3LIaWWbf2Zw6m5WP
VfdpINqzH1/ajjQyDCRKEeL20u6SUw2dEmb+ACTpmmb8+Pb1EI9b+BVkjSeG02dY
jsGLD6ZEWuBaOiGvaBTC35gAqOdNEL0cZXc8OUe5f+V/VbebREWEDayY/+VmC8C0
VyelAQB0OWuWn9FchhR9IuSvnVtMm0EuWrGOEt6zC+Y41RE2qrYZ3gJCv+MWrsXq
cuQci8Ya1ZJt5r0wnzIk5tFogYYqThZl0nOMycjBGX4jIO8G4n9bUlowcTOtKFh3
8jkCKwRT3jTHuf0s2c0W7cgJBKhUcborG2mga7A5xUh5hzEawQb5JzReUGOsDapb
joH/zabkJvHZ5h6+RabCwK2GIdkGPQEi77xXy0RDwHKB7U37o7yhDTnD3DQsTMlZ
5ujPmoid7z+GHgJ4QuMr1Zch0Vn01j+p5YuaI0WoJqskaK0nOKvIgIJhaf5ID8Mc
gzmOHeeb84qjPRvDqTbhCksdHibmk54vp9+rFI0OrWRh5qSmrxEIFMIefI+CeaQz
kt6hpq4EQ5lVmrY87aIZigYs7DphQXveE9ePWGPviz/lyyhq9H3Y0QoDw4NGxL1g
2hSuOU0UJE3KRAYkbEnt+V+LJv/53MDLrKyIt+CoPTzVRG/6qqPtn532eKnHdL9l
rVzfqsXIsQi2x/IA64SjRRHKtaRltcl1tBe4LiaQcQpX5jiUgBf+0eCexBKGsiGF
O6cuR4nUSwgtndXtAW7MO9BXYzV+XoJsNTq5tKIzVc+wKQVA0iAi7XdIwV5WzV5J
KCQhLy07GwR8WuO5eIOW/zNS56b5ytwnzQo1KFyuS41znW5EJ60kyFFu/CB6qEY3
u733TeI1wFpukpHVlYYayvCsEwg6Pon4B3Y3WqOy2pbmeXqdb/NVeEQ1dYAxVd6M
GOuWlUITXfDBWLeknxNA0RGW3ffWfW0lSbJOIIwv/uKZGHtlYq3MfycHSXAO/Z4/
U/S/1sCWJei7hcq/AWZsoKYAQAI+MGjO4l0pzjbbf59YRICl9FlAL4/HbIWN14SO
Ku5U9MnVYHznYdp+/DdCByEPHwCotoPcfFXCYaKiPo2rnkOqZymm1+BFGSNPwmu9
mz6+KQ8wW8UYXI9X7n7ZaAOgMbIfS/198lJeDReadr6LMv55/rwsXB4Fn8QjsrEu
u8Fc57Lw09io5bPUQzdhw/UAFUevPM29v58OtQS+7AQGsJmuEWp9S7iVMbBIhw4l
Bbg6jdCnW6v9S3gxL9c5URs7B3E7iaQ02M42iMzdumLWB2VjXIMq2gR8dH8po14H
FAl7Smv7kGa/b66dTgnaMUD+Ruowft7R9qeNNVaDEdxhzHVltdHHS7GSH2wqUhYH
mfvbdqDx7RMHxO7MwsSeJ0CZU4TexCaFHSxBJLF8pvXvEOrdWqSxHJTthVaYAGZQ
BWZk9BUcLPym6LlRmi9OFsaJW3FPYHS2hNVHdbZ2/HSUKxZJ3oLFRWOyEIJeBYko
iviwU1YCfPDkywqpIKbO+ayQMrcOTdzDUUzMvNxIOzrCTpkV1Tmf9VvqQoJr92c2
p7Dl0OXUSRq1rr5CyeM+4QSyufhsrN+q9Zhz3KZq/u20t6puZwWfZtxqQh9m2W5X
qGkfn3So/wwPTMJpxKomMKde4qtosIhPL53Tqm3WJwxBRs5enpDA8oa1RsKJ7Lse
O1OSp5OVvw7/d4IKvNZj2bV28LvaV52Rl/5fcl9MC99KTxxD6bIUw0NU+BSLGhcm
8r8D8lY8KDEM9/ulwgmZfIG7TY+HBKzbmmAFnB4IvQxxT0oxQWp/iClgn/5y1ZZd
PRYhufzsg4YaRrAAC+O3u3j0b2rF8SQB1ShxCV33BD5XpPR2v7or9PMmevjsQaxD
Nvusr7MY3ZkVyEvwumorUj/AgVMR5Y4J+UwY826/+Jh4ytPYH8k3ubwgILxaIlHB
mmwBzRDs3XkLTY7XeU77LBJsIgNtRBbfvaR4E/NmtC758ZvoiSCJ2JLyjK9OjWH/
DtX2fgVB4VTwx1Rcxa9S7a9nCdcK+K+3HZ9U6SxcL8Se0a033T+lSMyvjdVLX96+
glTpYW5F4ErTF6lrimMtRlAoE4/01IjyRyHmEbWBql02xdTj1DjjnYqnLNp5VDc6
1XkeuEoE2sPE0tOHb44jga+vuSb96VVKam1nkj27H4qQYf+Ff6+u0Spp3WcJLgsk
WbdMWlDHdk+pe+AZOUFOcWS3SQd78Y8GqHWi+MOcN+SWMKxV/bQzgIQUTxmdSLCs
O7KdRTNPWxSRJsi9jI8GAKI3X8LfDsp10EqKpOulzGwlRdAcY+I82jKnLj26Qkab
uqVb2CcxUs6GAo/9mJZGRR7JqKAIU7e83M2x1yNb/oMiV+hy3vrSS6IxnGUNGjYg
F9orGNGD2NP+r30E/JioUZYZKidDviDnhhfrJyTCQIHwpUO+mteZgraPiiCHyZN5
WZdeg53q/b7ojaEh8kHGs0IENrrLXjZu2M02wdDjbCxdydopQZUq+Y9LXLyDNrfU
+QBAyITopmncbDzU0siXrnrzykkru+hhRP7lE3LHMjE0sFamFF4UpoK1S+4vx25c
0QnKimbeRBbbvx51xWvc5dF1tzbI8PHXUhp1U0+EIDewgyYkKfk9hniPl4gTPzFR
kZQuLNs5pxCc1LG6bi1wh+iCK2TSePsGNlwzs2zEagSt2hQy1O+t56OImaFsIMoW
XaRKrkfkRcl7nIuHdVBAe6VqZe/HMTdHG2R8ALQVDyMyvnNm22xILH4D8t0FpDwY
0pNPRdx9xJcCiMQ3XdsiGoZbDE+oWarYvYtdZiDFJxj7dE47GzyQOG/wApG9/B/j
cdQkDGkM3l8Z9IJz/tsrdnd9dTnhN/gpLhmYwchfwzp+CwkZ/2iXeuhcauzzwMvq
EkSRyV9sgRMHaZ0Q9Ovpfp1kJ745x32tEbCv9eJDC5X+/JotG0tiOUgbDRvLzHUV
HLh8pSj58YGzwwhJHtnYhxtH3YLM63ssBb2XMlxHPuNYdPN0DxGfLWhxH8Xzkv+G
rV1Jzygm5swVngfrozBUgAdcpo6A3UZ+fESR6rMCXNnHfLpHRVi4XZmfEESeQUsG
sdP7ZvTK2hoBRgVV4hN0EaLWJ7AhjO5mLPH6D+QLpYngBdPUZ9XBRNVolsQcYqkl
KtkftimW8RGFABIAa5AtgQpnYPnoPZDeO6MtfZnHIlwbELv4Nv18FtCFiEAuGXoR
k34i6ScJRjyspFTGcyF72CwWnjBKnpnZbX9iXWPsFK1iQcCnMg+q1AJUyuabCN6k
5PDxoDLEkk6LJmV3uxIc4ur5AqNf3lYTXWT32BsIItETv26LSuaoG/mVliEGmuwp
YI1a2auhAhTtjhezmO5HvY8DRmxO3U6W08li3bEQUJ6e8jodQWISz9lEOAKsl9Dr
E4WO76j/NiDyZUfw64LM3Nz1XfZcParQSKhmHJaAC8G8pP+77zLmwGdMxcRNnAf2
jFOhIw5r0CtPN/KHy4M2zoTJ+Swnpu4/rJqSb47Tm41xYtkpgj7GySafSNYfN7jU
jMv86WohQ57ov8RyvzH7FhL5iqKl6PEpu1C73u7K7xqvVbgWlUvFWPP3D+jgiDjL
xRo9tYHXbjVw12Q4vA511RHOS6MWe6I0VCIqr4LsS3mX7nvZWyrXR2zG/mG7YSVX
PqM4C24QOsPDltYsiai/JvrZa6yBg3/k6Fn/4HS6FsCBrhy8IqUzojQhb4A5gngQ
zIM/41RB8XjPHOtbmBRcSWiPCwot7I1uT3TOjeMHcYkTzgaaQkeKXnLkqzn1q8+b
zCDn3EBgUtJ+o31LgeS3aMQpxfJe9244l20rSz9yXnMfMYtgM2iZkEZOX1ey8Kwy
6LVTskW7pl34MIU6/NVfdG0cvDthjsjDIHRaJmSPGRui2Q6nqD4kSpPE0xC+u/9S
Osx1E7lc3WzYBKv7xUBq++MBs0BAupZAV9CuBVrD/3H9sIaapvJyQss0KrHWmNS8
bC/wC3iYiiiPczKSse/NNZQEF9Kj8OpXSKXKJTQqjGhq/b4EpHgCNWcILXvmntjV
37GU/ldq2iqVDVXhuJP9P+TkfarMPZRojBgmKuDhz/ROiWddAXgiZ6h24brSAnvy
e04mK22tbfUXN4G3bxUIRuUZLJjo3vk1eaD0ZgnQRgPq+euyfjBczcCocznEjl1M
Pg9xk/DLAbyWtEjUF6DUdZCCPZ/fGvr2Mi28MrfMc+AGPPBlje3JRbKWuSp5N7H7
vaz4i8HgfuF7Y1niVc4AeyUyFfu+ZgpJ1m6pSU3QQfShW09wyzUczKtGFeNEUJxU
e2stS5PBRWhMiEFi+b/Zlu8Z3Sk1+Trh7bzPV5PWL98AimWEnp0Y9MgTGnt2S65Z
ISQlNwhcpK6q2Irj3sRxDgHNJkqC/ZNBR4kBY2OnvpO8m/FW2ne/JpgeB/vBePWr
SM6WiM96W7zxokxKIRQwqp9ts3AYNlREphnldpYVQBXbl9Bkp5xC/XiSlDSgQVWU
Kbae130InlundLCZr/PcMuxIofq04PRT/S8E3r/RZVOHBxZdMFO4GBv4yqq10KX8
H0FsmbAV4P46kUPUjL19r6gA2L5hZoLvOI3PXeK/WfkmPuMt9MvbKOpNkSlc3wkU
78wsMTtKmFkVkfwnpllBfIsxwHY1KllskayopGFvrgMvJtpG7U5RiykbnE9IWPvA
z3NA9/CfUGw6EUHtGzXX5FYl7WIUcQRlWn5v+RUi6rn6darYCq3x0tzfkBULEa9Y
+/CoSVlv7uGtm4RFeQP3oS/bgJ2C02oN1irsObTFnzen5DgY7g5KkDiGJkTegDKX
0uKLlb2qx6sdEvREslWPEIM7J3c2wEnVAcNDH6j7uknK+LYLMCDTvsVe6H8+A77D
+noxnAEGDmNlxV+Ap4yKpCwVhnHBLZwFjQqT0JE50r1DlL1Pju0peV1yaoy75mHJ
1D2u2C13iEN704ogpxsGeUE++YGSWxrYGU+vGi4igqK1y4L/4bwjB6cPyTowYj+B
M+fgDgDhFFouq1SDUSxMsYtiHOInr3Erxslt3nMyK50fk3ARBzh3pvtnUZzVTyse
wB647N92x4K3a9LbnJvBzKzf+4+4LatQyxkOkw5BLO+y0MSeaEpUiUaN8X1nVFgJ
dkUc09+KmZ7XToUY/KccsbH/VgVpjV87NC4Py9zSWTf8GQwgI2WXFFmT/opI2UHo
2KzibRTutGaWQy/S1GLw3IDq5uBXDg154lUn9gIs0SjhmOs3KcP/yz6fvDQrWsom
1DAp1YkiCTyS9IBZTFcM7G52LgNjEUQ/FTu+bGRbBkmdDPUqKt116F4y+9uG9egq
cjEatn94b5LqM8QyCHncbrc10i6Cro+m3SrZ58dWw0i/5qL912dPOuS5taZjnhiy
9ALdVQaJEtZuCYhNAkwVq+mIkF+EcolsPlRyYmLWl2Ay8Jr+fnr88attYY1Z0DrF
0h5u0RAsN8vd0LqMz7f07R4NDRHer2K/sMvzTF0ArnRwPYQaYH4Kbgjrw7heCw7Z
84fQul6l4yL5nCkOhSSTGG5OaxgO+nYKK4Wr5bxgJoH5BCLp0P98vO10D4iD0FYk
kkq2V9fxz5HqTujKIlGehbN8WUyFro6bm69EybSA2THQ8vrEdhFOe1z33eAZSciO
uFME0xx8MobC7CGtB0qVAzX/2qoEG2f6AHJ2Mw1snjCVP89jo97a4YEWKN8WYzfs
HNHiMRdxeMO1QpdJXPgR5yPYIVZ1t6OaLOzVYNTR4ZznlgSE0nXiBxvSOOkp3JVt
a77llsKPdqj2MqcLua9GFKoWxbD48Vv9UzKokZDsOGwaXJc4e2sDPjo1N2O1JoSb
HWDPDIJNODXKkgc4IWLTPvmqlIz0yy4WPj9CGlL2uI7wV7LN5KKRSHDnGQ+lCRpP
q3WV1U/NZUoBhnVTgF6L/kXQs6bkDRvegnwEZ8y1u4VY6lawsb7hC/K0ZSTOghVl
OQc9/qqtLGGbR60JkRLKU37w53TXLBblwbHdxdAeJP/VYsAMRCNinf5Rd7MGqUYM
sPZl8yJC0kVXfiliDMCHd6zKABKnegYBp2sFyaQQG9dWcsYeIrDDY+/dgt8l4CvA
AgY2RWKqr/WcZLy6LdEdgmMtPO5NgD5f41wTWYeF/YlgXkuqwnjkhmLaaIm4aUwc
4/GvBm0ncFbkkM4pnEPIdJF9pZiW1sxWmEsi/Z0PxsLzYumdKwgVB2vhrhoosiP9
jVSEIlot/Z2S54UXMs+thS6oj9I5Ra1eWNXZbtsLZSOOW66c8UWXFYzVabEYa7a+
8nPneZObmIC1LauWw1rSu745FmBCCKAvyJPEKZY2Ra/GPlWwIxVDo7X5b+xHPrU6
kxcpPC/HsGR9iOfOLIlkukCPsUXQMqTDJaZg13xYWTKwX+1Bgc5JYnfV6Zdv/8Qf
cbYVQ4AyDlqUp2juz0wczsKZHwTgIriS9FoEWj6VEc0YqNLTo8Dc4MTQLf6hp/Un
Vw2krFC2ShhYzFB1PtIay8/MX/Ga2wDbWKcJJlurHfsJEwgfp29ez7SL5KK3mCIT
/xgDww4mN7/eyWyk4EnS+vCuYBzA/x96pephPxLZEfO5xkOUjPrKpm5t8ax+RR33
Vh3u1TMilllkHXmuJYyP9IEu9TB7vAM91AMjF28PVoY3SYrDEKe2E/yIo5dnqsqA
GMZPUpuL1mfG8P3pz7UbqzEdFSikP37JUh44W0iSbsbuFcnxUJVrmHHiYCE5JXLZ
J7sSC8uHcMCQS1GyobY6+lvckl5LA3s0e/9UHwd9wXkJmfwR+v6HPzJHdjx7lTHn
OE8jkVRyNKjZKPo95ZyFouHC/2HEGk7bsrSAO0arMD92XyYjSCu9wzxKLgBId65/
YcMEd9pqOb+fK4xRTKY7Ibk8niqi7yEWhy2R1n3VX5mAZT3xcJj2VIULCGpgNAQh
oXpGsAyyHuo7RfTXkkOgRi6d/xF8i2jA7dL3+4w9kN+8PLtZ2Qr9BpYrQDMOfHuf
ABrCHq6kSMgYqR4yg1jlw7k02VvexfIoUpm9+NpQqeq96qOULOPARr3UP7IpRr9h
Bdg2XB/bxy3tVqhzUVIOjsqoWyzgL1u5Ahde/43rmdo0IEZIFoH2CB6tgTgKzKQP
1oqLIVVp6N78eQKRsCxfP0cup9R/M55AtapksxpYsYu6QrnLD/XjP0GsSbJIbXOn
FajaoPj+LVYCX+8lnvyUyIR0d2iHJZh3wdOLw4yJIyybeRsXwOZMQHVThgSDULBw
`protect end_protected
