-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
abiaGxTNtH2wIbmAcTF0+CbaucRNtG+hiwE3L/ztMFWAYY243AgSFVFkn1Q5e4Kv
mfyk5h8o1Ssp0ho0G8b5mnWYxWOzZXkKHq4u8SrFnvUp1CNNP041Xlgo9MYtxgvl
TZsfihcUtzT0u810LwbiW9WnrYXxu0fTZy/Ek0PVKGo=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 19728)
`protect data_block
ePvx3WMhRixqcxP7TAbGCJ9Z681dPhE9hABC5uvfUEJUpQ/AhrO2r13LfJLqpjzp
VopJGVgUH1NIUmHAK9stKpcNLbu46s7Q9nhKgXsppmgQlSHzVPBod6mq3eRXVYn2
VjybjCreWX7KDyWCEZhXuBv26Wek45qJ1EwSK3/S7sE4PSiy5Z/UtVfHa3LfF+CQ
IsVYQsrbBrP0ZMsspmE0EK8trXVKYtNt8wnRTfCqEKM+trmuhpnNJoSG1JkwxRqE
l0ViJ2frCawhNZENFWEeygI84y+E1IOyZtljDf2ldQv/Lrrq1KbgGUscXCcAZglw
nmJ1K4cZVm98BrmFE+xRMFwzbZ2zxXrP1sBAkwNQP6N/js5cEnLJh+ju9ZOH0BGd
TapwSSM3EM9OLs28/zEYKT/8HMBJ42K9l1qHqzH6eE1jWuHkLuw6DNB1E6zIO2a6
T+ZIo1UsR+apSoF1F/KYgJ42NGdzfTvQprKECa6PDTJ9G/CtkyA6xTlACcQ1vfOw
7tndjvlv+fLrz/+pbShtp99SnDH6McI4dgCRLfUNotuMoBkf5maPvJRVy4LMZ8jg
InXHWFf1ZSP1fcCf5YbqELHias8v8Sqk4hZwOhjuquRiIlkfmJjavM5jWfea0xve
NxfUqvG8a9c7baWEOZmXhZ5k1H7Rl2sIEenO5Hty0A9y/FCeRv6vstJLmFUDtoF3
6lcw6V7WCJeyY4Kd9ktkWR2lQLiYSPgC5uVpClcq/WCsB+FcJ4PmkCkIh7eSGKb5
LHqCpZR0caBhASyO6SkE0gNnHsAiy3Qw3AQfJ3Cg7ScWymmVoQeivBPhEheKu8sW
OV8mS0xc0hpIKyNHSiLYFrTZyn/900j8dFvuSKYQRhljb+B5h3G5d9Aq899vq7go
E/9QaY1jxfF5v6UR4jvMKQ1kQMlnWPKAYMIyEaE7S5EugE9jQi7ec35Ja66Sj+ky
CGMPhrwcOgvwdsWhqIFD26XSGa1VgPB0xKMKyWd9rlKa+XKsi0fkaRHfo3ZqbafS
iCF+pXBB38oa3dwSFCTiXY1D7nnXBBpLgwtckH7rtkhOJH3K4LXFOX7hCkEoQWBA
HsEKHT9dzKy34VwU6+fsT5UnIU+8gqMlAtsYvW8LPR4HYyPsqnEtY1VQORtlW6Q5
AVPA4uIIpNLNG6YxIx9dbTkdpKR/UZxPz2iVN7yqujV8Ur/8O4gY1gNLUaxnqbDQ
QM0FVBYHDk46k2SX/FQPZrf5o3EL5H/ZLVtwFbScf/1Kf+S8CX74/oXiLHbp3doz
7GoPmg4W50MbmcSz3ylWrbcY4GqJswRbyiPkyVrEE3x4dvY48jPnxQ0eecPNr5n7
n9wY3jXUIPb2z6JCrVVie4YkmCzcmfdbYOw7RivxgOlwxCOngXvNUiBa+7RdmADg
u6pKslQWtRmu0/quIM8NJMbHh1RrFnaBQ19qztF59/gwXo2oS81ErZ4/Lk/B+5XY
4BsHcOz9l9lT35Fyp1fT409tNNokpZWsosl9AYJ4pYfQb4l7UyEnYyCjyg6yqfY5
Orj5sIdwiP65pOtkhP1LD0prYJW9LI8mlc8NIYZoQf+aS6FOmv9mL44sMZjX9r2F
draTZqEpjLqZ7o/iYbKu3+CTLhHe+pP4HoLVy8ZTOujGnLeHDEDwYFMPb9nbqTuK
teJmvGefPVKJJEmnR/QGsfjRQIylaymND47Yg6yHHqk8d7GmqGJbi6o9cnBVO6x8
OQoy3q0jJWarL6yu+iX8FLsji37bauxOH6hnJksKdHS8BDaZexIHBojRl4W50bWa
5+7uTVerVXDMgMQAjzjlLEtON+L98UOJy3wAy50QFYz4Jsx5ZmY/FanDXkdiKlRq
lGOGvGFnA44wAKbgdJhY+ru+aTf+aN4vJyLIQbHyRxzSeVPdlckfsv/qn9ByKCDZ
4Cgzg57VN8NkVx9AD8tLPelCtsR1f2Fki+7RKIm1FCFYx/GAlSIgjrywH5AUuYCC
O9KyPV6CsmJS42s9b29hz+fKSi9zjorf5xx9SW00fGd8KKHE13xoIrNdz0krUU6t
sB0inuyeh95y0KMAxWcBrHeTiw0ZY2et5S4WF6Ex45TFsEc9FGgSnsTlFzHFFwHz
IBNUaJxdpfF34gNP8kr5Q/rjr2q5AxPEwjzghAa4HEoSRvZQuPZgXLlxGxcXOTUZ
1xRIb5EdK7FAZSB0pqCbnYiWatq4abzivSHOcOpP45cNivmL98wiH3ICT2Qor9Hg
o/TU7GwtXVA4CHR7+QCfiHzPvRVZhwLLN84rTbdpNFOAVJ8Ffcoj5/A9hh4eOUuu
nFPgP4kNhYnZN9770eYbrY2LmgkXbYFGngNKbsO3G80IgeeM3tl+hg+rHDMbAet6
feu7LA+5rb7RX2v5O2+TV1FADpwx7z0TXU+2pyripXrqipX3KJTuBM3r3538XZbq
CnoDvSqiLNW3yLlPxF+/tis+jjmXj6FRfxAmwH9TZ7RDMLiWeSmlZ5lqvArVEnxl
9xJNck9d30szQv9tmbBifhtcog3HhJ2r/YFIQDBpWHTuJZxrY16skmkA5oLRdJWG
vja9XtSzWOR6ZQJPGtzF/D82h2CvIjcgA/2/rR5pC221HBh79K1ivsB7KplYAJeY
iZ+A3dj0rDugAgO7VQrY4NweNd+preX8xXlOthWm/JTjrECDg9+/+KTKtGoXwCkr
egB0XsUE7Tb/XmHMx5CUOPr5v7guGfR4CX9DO5pLtrEugYMTQ/p+CbvKA5fNkeqD
YganuSSkiJWoVaWIFbEukvPE7eonaASuAWrQt5OL94bC3PLOi1F4l16SdseOrGJK
4/tHV9At78ViKyzvOLh0SkBhN3jxYVdvQlItBbEY2i2jn0cUC0mR9gErWb7wZKJj
wjDoObmFCA0znZzMB5k+1tGVIP9AaaRzgEf9flyZVV6uMajg8VCg+yTan750ai5O
f8/hn6J4WkqFe20ShVugSaYSu0V2zBBjyK1VzBhr6vV29Z8vuU7HTInIB85QkPtU
0KGf0w58pcNHy6ZPjk3/0cZZPtlO151jL7JIE/DMXqSiZ48a0UQki1WAi2aK+ENq
lsV931xU23Tx+EhBm8RGgUAhKp8JMQDefG+TXe1872qg7vs9fuItEtRGNJOU3o2y
345iQxH+tIZn2g9ysN8oUGnJ4IeeWiZUE7LTK9/U3qrpmHNk1XP4CCKeIj+iQ2iy
WMInZFDnlhUjj9J/G5XK4xLV2sMn4/6q2KlMj23fzzZ+HbRJSW/fpHSIXHHivoEJ
E8mlAVNJYwT7QljcKmK5eVeEZNLqcUxX/1mia/WVFW3GFw1/vcA7htyiKWhBSm4M
f9lYFgy+d7m6DBHC+Mx4JDq0+pXq7XG40C7kr4zQny51L2UTAWCsUZzbPvV/idvj
uS7ml1CRo43Uox/DOg+t7ZRS2dO8jFjc5wAokARlqkdnqjgsIr4m3YiMPGtFUytY
fRbqzaBpGqyORC6bnVMr9tl7hDJm7KZjYTSmyeFgfXkJ5oQGZ6nYwiL4Cq9LuOUz
/0z0/0uo702+OeDuAlcMxm64iem54Nh2woDetZfDONQlZUdgyQ4up5Lh2HwyTHIF
qBpzmEYErUsB3qBiDepwIB0hUfFvQkC126hi1i371t/mX3eiZ3sjFYPQYnwkXfYl
jkxlSehSg6GyW55ziEy/yFiAnyhrbpi9bYxB0Car2BjXhrQLDTi3Lu00u4GBDjHX
KhY6deomSjlivc0S/l0zrdExsaEx5mRrh7gUvOvoabhPO2kcvHZNktKvPryYiQE5
0dXZlt7ZOOMJRMcQbrtjYUvRC93VAz9hwGrutrziao4uyAVD3Tui4HPBbyQsAbjs
mPwN96YZrVWD4VW4DaCzCq+qX0tc7QjwepKfxRzAleD4On1ZCO6AKkx0pTGGakXu
FMUcLukbqhflH5DBc95csS/CtU9DT37Z2uU3zc1CKDq8Aag0+93q9XCzw65TtKqD
L12A0UERTXZyLVRXsnsY3H2L/KqXJBxd/IhgzJsKJLIC4wQPlHNAZ8K8j1GbQKdV
BOvQsHniFVDEx7+XGgzCNE829AU4TSUoHr/6ekr2iN7UsW6TpvWoHm9t9jIxhThP
LGSm7DPVznr6W0nL/EC4UBiJSekwWwpvQ2YEeF6j3Lotvhxj2/BJdWA0zlaroezv
sIAFhwJ5lKjA+DCdFKXns8qg8Kp4mTWtZwG/oARtDL3ZdMDzAGPdSmKK7FGPRgKI
9ZDsJetONQ9V0tnd2yer3wlA2N6LfBdvzjuqWswfGIu9mgxEod8eStqRmhAsotws
KJ7nWhwLj3FXQpYIRh/vI1ASlX8xjxluIgUMU3j2VzfFG8OMTuVkpmQIeiQZ+n1j
2nSneuts2TyebWj2srtyY8KVmaRGIxyaqDqW+/wWXqDhzPznFv9e9NMIK24E/7hl
nEZ1sGC5JYeMV9nIfZAKRLtH/ZUnWtNQrd7z+WgsZax4elnSj0oduYFaKoP5otNN
XQiL9MAt0+aOMp3scV6mZrztL1e3xKCuLdAXiNOWkfXWVfwR0RZ45ZQpmKFcTPnz
uskDcmarE2YuQDTlt+GkAx0ZTEz1X7XOUTtrH+VMhY99cINyVgsxr5q43xsIJQIT
CxmKo1vq3+Upy6XwOfZLFWjRXG2QcvvpMCHld6zaWR+qL8ObXFxnnu1ZokNkmxMS
p217eSVTwAiOPgTOxFLnltx1N0EKzhzckPA3BRtvyZg504X3RODeOOEBgNuY2WAU
1dSsFhdelvF3GLBLFKcVHUXNC0dxj9mIVzRxm8z3vQH3GNDDS4j5yOCd5JMwYECH
4JyeTkzGDXyoB1uYq4TfA7nIcaGPrqb3cBFivL3Ibp4Se2yDkf1JjugcZV6FXqJk
XHaMy/rsxDaoMYKe/jtkeRRD8Uh+zly0WW0XCJ7hSrEqGl+/QnTsF8fOdV/tjM9O
deehY5b7EMzr/dErm9i1z+5xaVbmXxxrmDUTKH6Gvku1egZqCagjpzyjVgzBtwUl
UDR4z2IPsFN+7dsxry977ZZ7IrADjYAa4elRiuH7wj2cG8KZHzDO6BoSmlC6cMnD
m64AWV3ZLGLoIUIMiOMKU+puI+DxP8nB8HadVrXFDXYre2MF8kvfcFH9L7HdzKOf
QlRDk+bcy7mumMZ/iMgTI19O+hsekWSy+E70mAfDQxfm8tCJ9j+yQD7cE7xYacXJ
ESi5KVJDsYzm8WfEbrENkzAh4ZhXgDZsDRONVZSdV8qF8sEcZBXAOW0p4/s7/t3D
2RR1KgOcMMefBl3RRCVZd31ITMA9vRf90n8dTIZsPKEy58oPZSi1hj3EXvBSxIbB
/geZCMJjZUDSag4qSO/zYsSHw8Rgmnzzpyggzeqg58iK/DBGiVJVSoXGKShhVWrv
EJ0ZELgFarHTN17tbUDHXELQrCs9aaZ8pgByIpjiZMEuU+qFxXOBrCEZ/KnYCinT
yqvp4XwTC+BO3a6Z63E14P/CCVRctpyYhm+SxW/kvGASQglIBS5b9PMmodkhM6u3
KzaZ9HxEI1TRCRnLvqm/kOpNAg2nfVgiYxpSN+962BEE4HHchkajREIxZaBvQB8Y
ylc5KdyCa1lnLyYd96ucbJ236ZJP3XbnGc91mCILobNIwTNOWJEJKuCGAtjj9Yw3
YWoIhRU/3k7lTbiWq8bVJ0z0WGLEWnAfZfVUs7a41T6Uz/aNeSml8VyVZoeQwW34
UjTV3cJh6JBU4Wt00ohtSGmbnjUMjlgu5CYTZpY4MGkszLTMXRGam3cP8YhYKWT1
CVbN55JENXH5J83Y25VFmUjxjhXxLcdu0avt+mlJyDlEyfvg/3xhO1qz5tn9ejhz
qumC5/TY19P6zSgfQzod7+bBSBMrFQUwYzC413jovBrL7QD07rgXm9Xde63THMML
nkE0vSO8fVkFzT1tT3afIQ8U/UqS6YbrUXgCJJ4410gLGmTSC8QS2P9xEfNBC3xE
sDAGJwkDjVLZnblYQSb4Ut3OXufbInZeo+7PIE+FFHHxFH4GqDYeGCvViib7AxYS
4NM+YpkoDFJuQawDLfhxVsQiD4Kbu1I+NOaAvv5mHkpqry88Yan4w2W1tbUAA2MA
yWD9b6WQkHPPQeTz25kZgpckJYXtTzyMma8XM5UkFqmBSHtZtl2HlPmQ17kiCd5J
7WuMUC4XfmWT/WTCDFtspgzCZTM3BsrbMhflucywEy751WBRYyCdqUoebuvIDi+N
r761Ye91Uw3kpz3LNHxR212s74tP7Bac+Phr7G/yET5PwYiRVFFgP4MZI9sSvByA
YY+Axxgf2/nGXzWrPKsmJUkTeVli5UOLjsi6wmhvMdvfu4fhYmn0f5zd87vEMdBj
V2YspBNsTqWO71k8cPZT6DLbhb79cSzgmfpDc+kAoXTvoC3MgZrh0PmX6fMe3d8m
FNry7lud9vadL6z0bg8aLJaw+xmAAyZIBXKPOXWc1NfqcrZBLtM1eboQ6EYdkAKw
FhybL9r4P1bBKjMaIcHhdeRhzjtKTUdLEa7E+qUa4F8zvopeq+yGuF0B7Sfrcsr7
NIj+o/eWCdmusF1KYLhmd61v8BBEfU6PUspK/ybcy75P4aTQ6iaNX6zgARU8b79N
usQHlOVvmX3HMeC5Lxc5TPK4UmrDRaOG6/XSIX++SztBUdvQLSO58JjHLo9WYYNd
9Ozk1pgPNzPxLQJ0a5M0qG1GlHmoqi/e9cJCZQI/g+j+PME0gI5y9ie6vcFEKm6E
9iqyTLDLVwVhvvOPZdHOJNKq1Siuv9GqXc1iEo2h6U5J3zKOqG0ZjmUxp7rTtnSf
/NvdcMNh39QhAuaznwFZNSlWHd6w2UURQ26rTKxI0RglyjIYJYuuwgUQoAY1ZT0X
BxB3I0rZntaSlyI3ldI6CT1Vgk2ZiMA2KcpSfheD/ipLIGo42Cq4ymfCAwB5v376
h3RnPxW6QBMoLbIElsbrHR4aQ6jwNNn8BlPe8klCBBp9VZFttpK/cBjLhOWK0YRd
Undc49r+lPmmwLbKrKz9i5lPFRCnXXFV4R+FX7JsMEJNZ2wk/aLlAgCQnE+IxZ2v
scAwYZC7KTHkT62bX57RB7ncJPIEKH37s7o2t2YLN9lERnFGRYY2ace8/3pZF4Km
jHn/4tmmisK17Oc3ox3U4D+bdMQDIfcPyrr6Q7pQiiFH/QY/emy3srhiHOD/75Ai
ojvNsff/eXnYaSrsYFSozxgwzX9ZLYZF1HVYKmhsN2AgSRVCdhqlOdJCLs8dCcVc
jOIOoz15spaVbpqoCgfORsyfJNHwRad+7kpMnSziCJnACdJHIPLhbVTgzT3boKPy
8UTqbVcUclsbYZdmm0ToKWW6ZfOwfkGcgJ/bTp20Qt7C/2o0i5rs5yewDg31FUET
L7n+cZp2j3EkxFk8/kdZ+e8SalnXqJXpI3DAkqr1eV2auZELhCExy+Fb/LGjwdCg
kCzZ+5UOFju5b223rhGbqZE2snSGJpZkAgsnCmrKTMBGQp2Di+/8d8xlo4+/kATG
LUaYlSf+ywU2QUGJzuwumac9oW8ueU+BrdRfBYFlfI16RSiPGpnCKbrMuPv+RSXx
6DIe+XSIy2fHtJdj4xHb3Mu9bXCrIe/KxAV9EWI9LCTF4IWIuEKmI+byRcs6jgdG
E6ROA2Gfp28df2ot5JXJcT8OimNSatE728w1uopAXw9WmW0jwcvJjpNbuB/bG3xi
mnt4U+hpcDT8nn88+cO18YSFf6z9BkEdSZW4eqYI3IxhYLt9jLafqBlsim1XW7KN
nAAXRyqeIl3FK2SuYhSBHrZm1oo/SjvUSrPFF2QQ+QDg68HnSrqAXKaO9Obxt3Jt
6rDngOKiNJzdRVGw0cuKJyLC4hF9+ynZw/AKFt9ps/8mHLCM8lxV0UDORvuv6XX9
tsnr08yt3GQx2PvkPS6G/4/zBPrSnm1rWFF+5eXK/AEMbnnJJqFxgIJGyOBqYeD8
JNkajGXhlinxRvuAPQbfBunV7KpYn6b853bCgOzJk3X1j6qNIVrKBHLwPqbRX6li
4tWR775UkkkTnyOC6sTzCzqIOWXrIWaQIFHsB9f5+hrFK4vr9gtVQAW5jtML+8SZ
J7w6eYfL9ubs+xoqYAEWdHqdTC0vnvf1+UFjChmz4HRYMPMquBY7+QV5JHRpCFuv
M3GusBnom4Ef7GWyngVsQSoz8YEFGO1kW6b0RJs7CalPfm22L9TvCBa8sqAghJAr
tLYJAMHb1cve3nKQoy4mlWAH8Z9NE6biQtZtDlStAhRLgHY7kjt8QXYESFvbnzdy
MmnUMr7fp/FcmJdGGFak9TQVRvfqjn2PpP2c24yIOECKhcvTTocRpQHV+n5yJhdj
UTJ91s+NY0A2C7m7z0jRzdVObp8U2Yt6qnUfyTYA1uKuN6142SAGCuH3VV9jZrlz
/D5/z3yMnLJsyRuC4i0hEDq1CltO1kJlGK+JqtJLFeDVDBUfLI6IBpQulwNmCuDF
fJzg7PdFb3MqRRP0BaM568sg3UJ9e2an5r0o5MY40500mhXhS2pk9eqsCbMg5JDs
05kfUteBjKXoc6ZxhgWb5o1cFmsgSZ2D445bKsHKCuFn8VzhI3Ji7tJynMwGLCCr
FbpUffsvM1ybWLgbL+7LrybTKBKgq3jQ3fY944IdYrbtDHxWHlER9QgXEq9BdJNK
FEHo9UTPBj6CfWqWYYC3ugLR7WqZWyKp3Fkfp/aexQ5xbGhcNGBtGeqZHcpXGJDu
7UOterx5Z4W5uSYtcvNUtXF6ATEOCW9e+Q2NTBNF8WCXtbl5szKnQrrD/5mW3r3R
hmHL/XrYehvNQ/dUgaIZMexy5JGU5bV09hmOxAsV6J5+KJ2rCV+Qr9ylaFV6xg5y
43fjj0/YlhyAfuMS3y1m6SKTHgNU9qv11dJhXOnNK8zO9exW2KukDmbuSm6Mf2g1
Fv0wZ1l1WoPQRXweRd/tq9oNDCQ4VmR5e5O8Is1NCKwPxMULE4nQ+7MQNpGARDaQ
Elre+00lhl2q6Epl2wOIBKABR4jK7HoRiu8NtYiBjL7Np4wegR38X9JzWmjePiEs
K87ZHppt0LYnzrU2pd9C2GNuDG0gxvXBDbOrVwqJG0vlh1TT0kICnLCV7ZEphiKl
zL+4Ed/vugBRkTFwMyFlz7KnktipGSzwB+XUaxHflUbQ37+S7xRZtW/lC/pqytBu
FY+icc/gCr2EuZxzG7OKoAGLsemTBHYK4bs2V45wlyne2+0ZBbiQrl1v0hcocYVb
/LMkQDLBKXmo96IGg2hGec9arrmTMAe92H1GnSiVjXzrIK4GvcSRvyPkPIZxa/NL
i4IPSU2cH4AsCDqmWEKhE3xB3XAtBgSuYhudmqOgpvZim4PtyGK+f39PZXzLDLVJ
768UXiQZWpHuoSQhEVVGg0JqvEk16r9QHL3IQ6SSctovi28aq5KbzEF4JOJc65fm
Jd7ll4EBjV3E7ITMX3f3hm9AA3q3LIgAaqrGjVgC84CorixFmZHAHM83acWz4I9m
9civT+rttgrghAqYvOrcKwvKAgZp2Cex1f79bN3n+GUxjN402gMttITRX2tuvVx6
v3H6UnCQplfXzzL0NpkCHdYdJKJgW/80ENW7eVJ/4WMsiR5Z3DfPik95rGaRhixG
sfEdYwLSFHOfgMe3/9gGzYOh8+G3cDGVvPxFufpN5stHHF/pkL0kblApji8IQpqE
8e43Oq8Y+piKBbZ7ypLgtcCLxKL3ok4IK1FXOYItQtXYHSWarFIUQl5S16/KfGef
PTR+pIJp7XFQe+4Lt2p8OzsabNiL3Lgufo9o7VQg+eHMaa4NKzRvbtjySTHOB/CG
KFYIovPMWg4diMrKK//GzbrAWdRmhxJVdDaOJxk1CMMB/fkHxvefhjN9V/iEO1pE
HXjpR/AVpT63uW8yxnFH6tLb5PtVDF+kIZ2vPesX96LuMlue8sbpe/aRVnHF7jB6
fSJsMU5P/7YLXr6Vdnj9NX22dUMDdViatBV6iFpqZe+FYWMmF336VwMDJCqNIDwj
p9fLjYR/p5oDIHRBTr9jUnwkuJZTFojtyyDhbEuNPHStMzRE4o1Gm5ga7gMWdC4z
zHS3+/0flwugiYJY5Hh9LgPXrJTzW4ICxJezpIY8fjM/jNoE0CePlVl7PQh915G5
F6z4zQi66jgo2ELxK029diiU/NXtaoFdc5LOtMlVHJkJ8eNgH72GV8uHAm5IsB2n
g2kNQ5uj9MPnQ2FME4Ao6jX6tpQ4x0xzjpjO/G1kEaW8bEzKXxAW5zDGpuRMC64A
HbTbXhTjNYqb6bG91Sf0WRw9yvpgMy+fcZtHxnqNKz0vXDOfv6EYRyAZqppVZOmS
hH7M2z4jgdGXoka7vLNysnsoNdKk0AaPuhwIhNlWIIK0iGApnQfEyPni2lPh451+
MGs7W7M0WAJP+1fskzgsMj8rYAKgeHJdV8lbo0t9Ofm3yDR5xup0G3SW8ONBcMcW
edEHedv0J6xPO9XXz5HemKMccPQyWHsHYebChZLvRSiSFJPdVqhBnYwbtHXJFma/
gQGZG4gadyv5ZNcFeOk3pryOBM/VhRiyykjRpceeyKtumbrOHBhuNRunVLlziSoE
3zrRScSOa4mU8LLQpOS3eMTXeCv98g1meRvrU9Np+e+3xskAnDm3Z9oGTSS7F9f9
R/6roNosaGKWLi59PO4luG9LCsL1CpjcvVjaTUou8Av1J59bhksawK4tr/Z7TOVt
z7rZn4aRr5PTNP0Clg2ixNcq7/ta+SPhxbT3xbkai9T8VYWmr/vSGhrVh5C5SHWV
iSM0pPapbD39sES9OKKqx+m2d7/2vGBTewZ/v80/uRpKaWoiC+NIS+Evv0hm1Bqq
GCxl7o+jIxHpTeb6UveY1uuudgUXJQOvAV2FIlSBdSLykeVS4+P78Z8Kjwe6j49d
+FOSRPd4r1O4kKjFImWvZu5jPS+KSFKsYRpYWTwbEQR6rRGXfjKMVyjvjY5AuEjJ
FRO42/pVUj9ZCS6/s/7qp5myi7n8d+ZDEY+zUqU+KH26NG1AeYQYl3M9uM/tYoPt
RsJywRfE29D6KETekwUwlZQuG/ih8541QxsW9zya/Zn2LGerqsKalCFDjzITVCqk
o5ojfRO6rhW3TbjVt5JIno6+A5pwQ9cbjEU1hLj6dvWsDdrbYVLBa1+MoSN4lhxE
JTsIxC9ba7PpwDNTY6fqcWg6uJll+MozPuZa+kJsBDk6mWALyogbX56XzplnMMBV
49WnMGcfLcRc3u60300uD0Ly+ujA620SQ+5M9phOXBToxgXJhPhCqjBYtRoBZTMR
l4EBLTbxFZFN9i8zfiD61ePZOagCv0QcpjLns3yHLhlFKvRJqifqfmFvwd9aAp08
M0Z2MiZA9ivDfONCE2gf7DMiMyUtUHLOqHm0JxtlKvIFKGmtknkmJs8dQk+GyDM0
G/IwN4TaKbwhUVjk96GNMDaMiSk1owT3ryUupoqF3uglowm9xyGrbCULi73KVrWw
keQOfJggfiiFbMl9k6q9Wg+iAMjIWrNmMcbqLtxOo0dk4sgMBaUeV1AOs2OOt4FT
9rzagqFqSAaRPBQU91imgosG0iKWTXshEsF5tQGRT/S/MorgxCRbkLlOkSco+/e/
63NtuYbCiQYTXdVR0RLkJPjJ1ea0/xWqxVGcHwwWOMw0K0NB6brdGdt7ve7fDjj9
LRijvqr+5QeSXwUEbiVe0pkMgGnZdiYg6YGBMZ31cmwc/Rp3VnYHLFJG/STnG2X9
KcaiLrkO6QXRX+gLXW80KU1nxHbCwysJiTrn/GcmnKfov+jWiYHXyAvsW56FbhMc
3YJaiK5HCAs1OaHYo4tFMmyDVPeU9Jys9zG1RB1oOMPfLOxo7hs1jsQ8RnBjcp8e
aWFUfwBf4oyPA1q7xLyacwlIA2B3BtvC51/dfOpLqs52LtXXYr88crN5VlLVt6Cy
yHLySyaIAHUYbpdWP5JMeIsRoaOvv4WmaACmVOQDrln4G0TruU6A/gVKk06teaMg
mrzKa8MXmoa6uDU5HDzp+cWpt5LAVly0oW/wsjEROWrEeiwGSYsrBO7Ga5+8Jl7h
ZsvMoW+ZTyQlqa2raghNcp7yta/pBcvESCS1Rxgjpu2gFDVzArXv1SxqMNLqv57g
ltFIkiiSMEXl4RU3WfwddeIg/Kn45buhv22SF7W0mgvmW2J7rqVeXjPf3FNkZrXr
NfCmNG5mb/aIZN5FEKbBNRNbSXtKyWC0dyc/D0a2R3R0JCd4YScY2WvK0tx1zQ8W
/yNMbxUinU2dUyIAT7A/SWzhHXaNduSbs8ETFacYcwW7FNICcUcjxY52xkGDEI6X
GlvxfVBlNBdFWwwhvY7GQtH5vCMAw0ToIgzae18qD/uDXzF7BCWuxhpPNh1q1Gmu
F16DJeG1MPEpBmSdRpIFG6V2Lk6C1mQZxhDg/ecMmhV45IRXeE0eoS4l75AhhemA
CH90rnCsrdNImpSQbswHQoUUQJ9uCbEtnRaoaWIivLpVaQ3LBLrg0W8W8Q+c7M4H
CCDfwYhrDM1lKTt9JdYpj/SlS8hsHvHTuumGulCqtfMRU/hjGxNWb+0/BLjbV+Qk
F+fqbRTzUrA/hWWMMjiuMNO7xhTrPT3i75jpdpvSOUSOE9zQ/IFDIDqIN9x2mIRA
/Rau0EqqtWv2lBuJ4+78pXwuz+Td6yG4ng8MDKuLclHDGirZSP/QDKBFuqqE45QR
uG9vsZRq9SrK/ojnKIhvA2GyR3V+N1W8mGfMjMh3SLbH/GR824xfoR9nsuIDouSx
E89z86WK6Dc+a8OipDBbiGQhCczYKBkqgtlCokvb5eNmTijJ+khTdTWdh8Simi3C
ZQeQpFXdfN5DvTpbLSQ64c9I9p2lzW2Y5a4DLt+kvLu7ucrXbXDoVoKPReLBNeeA
Yv83Bjhlgk69nHB2uyrWfR81OHvqDLq2SOKHBq4C+2W02blDcGC1QsEIU6tmjzbR
v1ztI+YOazWhfXvaa2YzYTYZEjZxH4qRBc/UDgCuxDqh/o5RZ1/+2ItcpzvgpnUj
sYtQLkYMN8S6abv4TDls0ddsYHNDdYRVc5GkgTk12VBfkDxpBTyfnQYLAsqbKMtW
s1EVhpJEjOBUZZXlbzTyeRJ2dz/NlvBih/YrL4l3iNf7rS4GMWGbs+tVd4zhKIz0
by/Xv6JEwerHyZthZWaruxfL60KNNh/ekmheSlCTxTp4FxkK1j5YT+iZOJeug1Yd
SShUK76y8mVoLb+P07iTZrw5f82dvymzoqwWFL2m3DZSL5zyzUxi3G+jVsmEjK+g
ejFugQ4S9rDGCQXKPWyrSuvZTD/67ItIvWH95GZgETWjSMA5oWGb04vKK8SgPxj0
ZuTIulX8RC4xL6+QB2dWz/u9H7P2qqoVFDQKfwzOKYs2hRidJ+0TGevtr3tTfkhr
cyyH45l6rjnSvOqBAQB5bZtaZixcD1c6wb2B5++kDqKUAFZbta3GYDazTj6h3c6F
++OjbwDtlxB//lfpc8IYZQaLuDyl0PmHBuf1SAwS+W9qmbTTF6l/q+83ywyfmTXC
8rkXRdo+0aVKr/x1TVzdCS51MVT19cnj12ZJyqWP4TCLpSzocigmQ1wl86YY49OH
+LRjZWTw4/YPzN/Q0ikBRngGKkFYluGCxHoU9CtLe8E4gkBp2SOPrR8U5gLtvzGM
hP73mknbY9uthHQnMG5PIL0OOQMnlaQqihE4UniGmhrdN0qNYCBsAmLkZ+VW1rlp
nsaCPia/vtmNem8kbi3JhK9cXFpVJP4tYoybdaTO9rYFHQYy29zkGTryUGW/KQ8L
QFHWsDmSnUkVl2fuD+o1zmNNDk/Te1osfBkrHGDU9SrOMmTFRff6VI4xLzznflSD
Jyb/uRotiWfh68vkgPQ1R392VBzkqtsF6w3M5IzTRkyjd67PEoM3EYu7jxKCXWc4
iKagi4wqZ7mUpYtaj1p67AYTL3ypZDrabxZrpMq52M+1h0s1/2v9QJw59hM+c14v
+4gH0YBKHwxQ0iD7CEZM9EPR41AXJ0bCIOpD1L4Nrpr7zGAxCqH4SKIWT+2TPJh8
7nCrrQG/X9JVmMQaMs97jzOEY4Ijxfjz3SefX2ZLti5D49h0ANbST0HhBJFwQZh0
nsV4SsE6yqJ3rZbiNIG2or4koFMOAN34GEHBuMgxuUqI4zBKxl1OYxiJw63HfyXC
d7/1Gag+o3ls0N+/nM4hWF5ckHkyLWDPTNTA8bqj6vJaygEu8p+w7vkakIpoKHrF
nCIGCyO+t7ANAJV9IwIjW8B8VTKdFftBfolp0a6iFSExpjrI9p9HlI2yNeCD+1Zz
Mb7+xyltgtC/BSIJOMMih8fGWIJHCdfShxVjG6JKsYsm2IgLmtXVno0E5YPLNFWI
lVOH09KvLi4glSevo9/cMM3r504yiXWbxJmerW2Lb59kbHFWvevG44ZUO5PEeeBH
BdE5HSVVhn0iU59EFTK48kusbQfY1m/JRslUHIILlaJp5mwkQyq2GV8NWScARfEO
wtDsNCy0Rmy+j2a47Casy1qyNppRJPzCMHXdbD+9IZEb0vv9cxB812fCCnIjJ+3g
x2fBcgovqJ8xLhKljYVbtIx9mBYMfDK9zLbvbRIWjsh0b1RrG8pGH1tGI/yoQI8F
qN45J1vlcLMv60925REUbjU+MSBNXuueLW7gf7f+0T3tYLMGaOOHOJ1EuKVgZw2F
6uEFQlAL4CVvkO76BEiKKk9rdwT56dXqri6cVog/Ks2XOAFpSOkbYjnEyn1Ns4lx
ryc60x9F1/yNvky/wP4ux6KiOgJdgQxVEu6kIXCUEdYOT98nTyTKdvzq3o8nFW8K
AEeGJO9PhoU6XKk0N3Vp7KOfebfKJ8BgvomJSkZxMU6cGOXeE16QQgzTwc0+s0Z0
7zyiWWQB0U+nSCo5EHLX2HpJCa3eZSCqgvYIuMw7WSNsPWHt3MIq9Mp/zXTSsUjw
8wD0fJWpgHm8lBYtckL1urLGIlvq7mr6ggaWEO/RACmjrgwp8MdI0Yq/26oRzmvI
gPr5m7IaJgoKKQ4g0h5yPBgfmjqHUvklaqilYed6dnymUUmwRlYJM47ywESgsrbr
q6XjyzQDb3yuqQrLzwZO8lMO3zMcRPwqcBEtkflEhtwKvQTMbGcY+bQaOoaq0O46
Z1jQkqBqKxCxZZ7eRgJwVV8BtvDzN8175a+/fXHxVkMxRN4q0diFqUo0FfPvqM8E
fTuMlK7EqtGh+RsoVPcHsBnnvarthUWqPXrbp7F+aBgc4GnRyFOeCuANoWkxiSPj
+jUw3NJlOrWcseTwz6E3lqDGV4XRjMn8O0pyB9TmNwlvVK3+GCF4tuAiXWXQ9fGs
j+ktbAbCucnjQYBN2ie4K7++U0CcZnU1BWB+GIu7CE9bII9EK/OPPds4XQaAYm/J
Q+r6R5hT0LySrj+hazto/BFFEDOJSj3L8vV/w01rO9CSa/NrDeFfwXdUWg6Ssyl+
PSZ9aXchCJ5QyLoeIcntVr90OlS/LgFMAI2k91oBmZjZpjdd4cuvxeWMyclLxd14
wsNAwJcn7b88dbc9g/rWZBMvm47h9rTCpYA+L+ChDDgetwU1yyaTWEFu6HCbTNMj
wCx9snyI/R1ULqphmFL4V+r0u+yP7P7edBb/ennZS18v4E35At+cgc8ljaAXdDDp
SpeKkSMrE7ribrmom/eHQerb8zMVdIeRvQGl/Elsnm7Fik4O0FO4IWwJcKAci39h
WmnplDhkGzovZGl+x4lzaJGpyHYBL/1hO1/Ee2YPDMgZcsrCtrkGU+lgIUOEMOe6
e3qCApptvaxWFt7R6UIZcIYBK1xLGMVF+elGqvCyqinS9CMPzNwE233PpbuuIGeh
6MY+oameVo/jghcnLMBfXoexZbXVgt4FaupqtkTq3db/xjcRnHJ1yjPFhKAmfmwU
lgwmHAIvVS+IzXvfaHVBT6fqcFWloZwZFuVJUtgaYlmYjjVskGer6dYg5FSblptW
HI7Vz2dyz5UGT0s8tTWqsmYtbcAqCITdzL0gFRL4dSgYzFpaxt80O6MBAfftiKdE
mQrYMt/Ebo/on/qIaujMDvf7nqFSHRAWB+Kj7gRlr8PAd5L/YbyeroLLczhazeH8
uti0rD83OVjrRhA20kYdsGR7RDHhbF4HCZ19MhN3daYoIfsuupkqwyImZppFhoei
nX9/K+zkm7I5OUPCrm2Wac2QLbLaJuWWPP/WUir1G1yFKp8uB+ZOVJaieox6qIAa
UxZLE/rN0tb07ElwfgfzBhVX5rHEEfkRaPg+8pEp6upajBHe1G3jAV0Wo2X4ZIt2
lBDMOyElES9ZSnbLwGDJT/YE6k2bjlnlzYo+MIoWzAWxJs4VfNtlD1Moy0w1pSvL
qqFYlxRiWM8iJJDSQnrJXrQPqzPQy2qVRLztWlACQVBxDz6MV5pH+cUjBdm3Cr8E
rm7T3T04TjhEQ4XaMRl690D0rJ7kwuPQjNXKjiQ856xFe3gP0OfNRSi7XX2zCOd7
u0F9OXFKG7BOHbjxZ9k4X4MIsMmEMDspODdI0W0hmvs5SU4CkVyVkWqCB26++PDZ
Y4YZVyTTRcxRZQ6qhr6aa8+P17q8bO9gvjNOl7U8CtY+P1mJ92CvrOAsNWyMdoDy
eE7n5Jf6RTm33KWb0p6Z8qulqe+F9hNJyawyt647FoGNPJjSP9yO2qtNDotKMXXQ
xyqT3hLh1ZCEHdIZffv4SuWtIX/bVgbdVO5mR29ft0OpvkNCOFE8m6aGx269E4B3
QPKFxkGhRJK9SP5sbT65R56Tv3VgvmuiU2Te3LjkE3rGrdInHgCtYekSYpbrN87s
KwJwhtlbCfI9pcj4BoFZzDrmkTYpLmYl5nS1eQ0Jh5Gau4P1GENZWPRT6HvWstm1
JcYsW5MSh+VfQe6D0DE8qTwzaW9JcUB89mfQPNXTDB3VPIVElk5ti1hcF7bUcEsO
5hNGEl3uf+7X5CO4lQjCHKyuzDUzieYCn8634am8ezhN4q5POMh+eOxae/tiH2nm
y7vlJdGdeGYIj2qFavzZMrnomY10/Xu6RhMcqYbraX5eZQ+T9C7UT14FdXkBpAYs
902Z3XFxLGlPZgRCvaE18OF0GiZOUMejtk8JjcSGhxKnf1BP6D/MCe3973nGHe0f
/7iKCbLM77wL94m41mdymveCcNHkcYgWQxH2f6472UvjMKcFBEF5Zfp9dlFqk9af
sJHALKIQgRDJl5/J/FbbNmnAVcSfIs9FPis9tBrvs/hUMRLCP8DYVVJcmwSYwsHd
kGmq79YsWLlvFUtbeYNdD3qqeMjWxoJT+ktDEPxUr63Fda3MVebgZVhgUwE7dp+2
eBQyLhxBr6G3zWsztRfEkFEzm63tjU4MAvQHjYiAZvpyutBWf8utHkz+4+vj55lh
AZl2B5ofxO2p73El/H9KoCFdaORofaamGhTB9ZnaVnzqVBgF1k9poGUkGsgmEUYn
8InPNxL24gJaImutROC1+q197GF7y9dFN2rXWeSKkzbZTW3kr5LHht9c/uxzJIcP
iy3oL9D7b4dzUuHlhMBg6jKX17cVzohd30m1P//pJOpjOa+ibAERYy9szOXXq9pV
wlNtANC9tw0GN8uhkBI7EqJJXA5m74mD/aGsvlRlc+caFjTAMNeAWMbFAV8BGrlO
4uBpa8/SlRXGQ8S1b/8t8rhXTf21icNmMvU6PVLTWkspoVDu3Ifx2IJOKhjRA6CL
8zxN6tbUt6l5Zu1W3hCIGA81Wq8lYmgICy9snsVN037+l0VSdPUrnX6veC8XCOgO
g0aW867WrIfvvHuiGHMWK3aNwYWW6xN/Qo/6ouezHt+vVZdJtCgvaJrkQkohwVaJ
Cs++Y25CYk+aJurh9oo/HpCDBuq2zQQH+fLXGtZOIqWobMKUm5VeBYUNPQRR2IvW
JzgjR3pv1XkshSaIvlnYPTYN4rQrBxo7wosnizw2nfgS99jOKlLHNUed0uWW0HtB
gHgTWeRm8zZTWqMOVaFOEg3LMdPxZwod9pCU1TXGEabpcJoApsMRkZ1562393DK6
aEkCfiddenkYNlypJu6lH/MbwBqthDObozsx0ylRMdX8+Hs67vvpNI8cUnH+UN7b
iUvQVM3KNlaUbAGw7uWFH1FIRmbEXd8oADuCht2JJUwePfa51MVV5zaCqR/12z4l
XlPd9XxYsT5XmoQFeTHKIBYAGhdnO0ogMXdJ4U4/XAj/uJlnBBQ4JMRIDy8zjEjG
gwMPk1WRi7qBuOQC392N0DI6WXExhJPpRKpX93B9A8wuWxL4Ycsk44cRfWDd4CBQ
ntTr+QyF7SQZUpAV+kZwIIBdzta3gYExxjHtxwPcvN6ZbwNQpowj4onR8GtN+o9C
iWl7nsQsv6g3KCbDDXwfsqANaqrDPMz4JFt57D84biuoOsBKjdAnyAwxT0RGVkwe
lY7ZvslqZSJ5kRoTa+pNalm0xp5g1PBvMccwo/ObsU/kW03wRYcrjT9I3K6qNRZC
0Z8r2hd/1UAX1UZzxOd9bVF7AgLX1GI4IDYWjKcJAex2+8sgJRwkJYwn8C/ns3Rm
7SXqHU82mNfBDDcbse9e4QUV3KHYcVUw8x8VKM8T62h3i8ppXSTc7cwwu3dRMwNn
VxAtF8rPBSKbmJfR29WtQMLpXcxJFOzeqOFAUUjsB0pmjnC//MprtoICkuUTmpzv
8HIQUyCDOQ4+vbimDEXWim/81ZhLWStiekkeXbD4T4jUsjYBXcSh06C4g0GFbsZO
06nToF2f/GRMq01HHSnwcFJePWD9eVQwNdiBLpmNVeZ69ReSwNxccU8JmayyhY4t
VITDPOerLn4EoeSxyMlxjgVvf2mQuq5m1FRhSIbscv8JNwY5zO8zQGQ5q+/2fgg7
3WpKlwoLyHJtbvTMYDHGq+Nr9O0GScUazusrR0mOi0BQMqdSh1NcvB+vAlDG5h19
HFeAbCAAFBnE66+BfGjwjOjoVb6WTmJ+2DzsAe0fNIyyCgwR1Tt09G73CGUsP+To
ZHhZnjAxbZbR+pHEelB+Oyk1ee6tsC3VGLTAaWa1ZGA6+8Z+Q+HScz1k4qX8uNFy
cSfEaOrSgcZwWklus6HrKzG12iCpiYGgyfWusQXphwA0kjuQ8sQYo8pSvSHWHPvu
AP6EgkFCasByv3V8AyP5o6nZPvJqSHTDYxhHMmb4MIcMiM1ceHDAuuCqi+rrKs98
5B1qTEcDeCLVUKqmcbRn0e7Swqhyk9uQeHsIsZsEzw2P+4CbijZE7jYhp5VQ+8ba
sYjHlaPSp+C/LtAgt7Obkm5O7MWWJlUf8uRmEt0k4piGOx/AHQ7dbbCr2RYD+YmQ
90kGAKc8DoO9xg04B6RX8P3a3Y/kSqjSZ/3AKKBZR0gDx6ss7IJZOCaPcxhnUznY
DMIxv79EekCrIR3e148KLDaOHgBac/5Hp73a84bXd6ds81JK3rik/uB3yVyAZyXD
oO9ODeFuhbXqh5Wfxzia60v80VboJkFsdPdu5nAVANTxEmN8XAYPsPAbNaI97E6d
gj0VKUsnk2yFD52dntAUaeolkPRnY6hH2MNM+DHGGrIlfHB2H1AS+vFEnHOTSte4
p5R383BqAtKpXJKsi1BasJ2eKQRUj0SIHGojAC+Woq7rkYk9qQW2SfS+RGlCTO5N
X3fXv1hZ6QHnY6hpf0KSE8CJ5zSi98Pr8nTX8OlY9aZKBYR0ns2kw3xIhX+JLF+v
9nk9D//CnLXIXMAL4SAfYYa6ORxDm5szHL9b0Nds871LaiXonsqGwdFqDBHOetsL
AYOOJXWwCWISszNG4+VcsgZ5ckydaSsISTomGcrQyJnbpwLcAszMmgUOmQiDBdCp
HBrrfkwBWQWxsloXveRj/lr1FqCMDIFZdTfVQxjlz+VVrxjoWl+zqibkJczcaOeS
ldl4q5gD3YFaOvUeJ8USRIG2+lFAe32DFGjyZaCegZT3x8S/bqFvAQ8qISJcJJzP
qmZpr+fZlY0l6Cx6zH/jCgqtTZtHX6ihIu7ac0ZIOB5lX2FRTCvsKses3mgTAPp7
qXZkVuSA+qBr6wRSoMhuoWjb+0mTp4+lQdco/cHVSu1fTLhqXuRfwN1msRoRt78j
GB47YX0zRP+A3ARnc3QAN9ObFR/Ek+w8+C9J8uHVLCKOZ712HnBrfBuxPe+JoS/L
9Yuzr4Afsps/Qo/Pr3fJvIHuQCpzYxYUu5es81F12AajsTIQ0pPFqnlMKP9Np8f6
p9kjXNs0FVrqJrY746hT0GPmkgiCSV3DTAF1J3yxel/YFPCDCY+7QdsrBjx0Ts+t
cMoq5QTv34hhrGZY9k9m3PNaKJ7eRGFpjkoAz3FJVksfcrdKOQzGnTcLLNTRahMq
gBEXSGl7YpEdupuVGphMGAVlaqH4/AXjLkb4xkN5l8GQ/nQ709p9/1hKSU7Bnlcb
qj2zKmGfkEUHE2offuyDk6BD/HqX0YvnCEL6td6PySEJcBmnQYF1Nt86PFQYbapF
jnHIleZWOAQX+k5FN4xqkN/5W5/xl6lmYLaKuJdzHgV3yIw0vWohsT2WEJjOEo4j
QgHUoY4Yn284TGpHQ1psPAXqrQkoqszACFIrjV3xcobCYTQB7VptDR3heD9hWtdE
1p900VPNq433uMMmd+KIlkDRC01mkdGGlhzsJwvV83fh0/adkhgOQZhV99QAe3ip
ZziOkh5y8o78HgglDKnl+XieEwADJuam2M88HN6tpFVGj1d3K+/qlDsvAvOcImYU
5+2kUDBbCZwFSuoih54N3McIetu7P6R5wRCZwKCmXfZxN/eVm1eOrqvi64ZmLz8g
aFyBaOZ17s9QfNugmUjFWIklu3NK4oxp901dNT6WmyrUSYlE6G1PFri4H4kffl5e
W5bBfJUMXhyzplRfN26LUmaQQHBKmjv/ydYuBflwqXiJDtsmjogoBBcJzX3nNoQ3
fagoIBGcdYP3dcCbQIXzojpOWuDpo/vbKy6NZmQtGtr8k59c6cHgIbRTwKyVJDVd
nPnMfNi9zGXqTdLPcnXk+gyFw1XdpfMRGNlzrydUFZrLAwGX02tyjI+Q8s59/lFz
KL9yHiY7tlvH/HvEI8VmaVUzuvqKMSHoqVIRV0MXi/zZwCDjgQy+qqp70FZupSay
LultkOt56+heSRz4MOxyP8NLSbn34sVR2EW6Nqbb15ksAhwEoulCiACwgr1avEEE
DzLRBz61+3ErtwvrsxExGFUEBZ5metZ2J8+WbXEE6dBCKx23c0XWQ/ZPiAHJQu6X
ngQPudu3WaLRAhDTtVX44Ysi4hcp4+u0CEqlfb7O8V1cXUFdlW818SJohhapW+gT
72+mRN6QAJXHzjdu/lULOOufLn/VJHVt2Co+gmX0mqrHvZlJG2ZhE87Lb2TvQ124
ufhHm7ZBNa1nxEkswPkaVfzgDgPx5u7i8GnGyFkH1XYXBxg2fsFPW0mTeFOjEBEQ
gfE6rJKxp7elx9u7csv0IjkOdsrJ0ASqbnBGKzkN0ASpts+BLEXG3tsKgOwOiekn
izpD3iI/JSLDED8WmG24sLSUTqcZBcsEdA+NPsJUQ+ssV2X1lQi2P9lnIua/+Uld
+tLJnOZHGldxAvDy+iBTh2tD64Az1tGDlzJxiOabv5Ida++Ib5MR05sM69f3nyYC
JDwD9MoJ7jcXg53rGh9KSZ3FAgFDeHMqJtSCjDIEayzoGGpaN80FfyZUhVVGmb2x
L/qr5O5a3kfTdO5JrW/IIcI5zPImYhWo4WYhIiv1QgCe/4Fp5gfv6TRc2LDS+QKo
2tqjJl+ir0oUNeX1TMe0WNzZDRtYPOhr25Xp7azrIMLqcRnbqJV0VmCLARGltQQP
g/NZguv6BHmso+UkcjQ3hh+tL7XZissX4n8v/4/BEnHC5G1lmaJURBc7mZfjUSig
ELt2g+n8WVvK4ByfZaJ7PBbiBAFGhBuITZJJCibhLKZ6jBAq4Qy0aCX7e62GwfHe
g7ue6xC102HrZYTjajJEtqgJc4HbtNhRFk2FFcCrA5VIOApvnlamvqD3hYSwXKjG
+FInpzBRPvRGI5026qQl9wnnhQawK4NiVNqYix4H9f9GNYg1Eeg2u4J0RPZDJjST
ixgealbLiS2pLwiHrRGNIdp1dQDyumeMtM0fBcnEClshTt6SGdQTqseP+ZhIoBFL
eKWcHu0GZ/e2ZJXawdpFm9yglitb56QTdZGsbMQpdYv+jflB9kz0MQsa2pWk4AWU
Js75XraDwH1MJXvdzzAGU+zJQCwUmezot5G/TswRJVbh8Ikj5Xs5wDNVqKy42w0h
eymeYVrNs7heueBzCqSH/RMzElvYqXbDEbrD2F9mIj0999WKXmrh5WVMSlilPFla
Au8hkCY/ss7pemx66uLsv7hJcbL1OIoAw9z26S9FGjW/jjdYpFlNrWKEXqBSXkVX
10MpQbRNE1NmlHeNPNYZYuelB7LLXGsLV69+K/4qpYf9db8mYZwIaA9lgH57Uqc2
GZ8hfAKupbAic3BZq4lOyDtAv2s2NWsozhINksZa5COpX4N7KWGXZazshTBvPNkL
77LnslIeofkmqZLbQvKXxArPuBoKsQSdLF+sUFiQQ5qlQ1/oLn9xWaK24iADJzHA
Cbq5/f5+csTvNIzX29n9/2audH9OKu7utp8vEkdv61MsHV+O/EO5fvRd6EvQEqNz
g3C+8y+P3sEhk+PzrycaDuUT58h5gI/tRmMzF0U8IAwk4tDFIn/dMhNNJN6RbjdA
iUjRZDGaQluNGrRJVrpeEOfATB/3e0QWfbnkgazZpmgIxJ55xMPF0t+gPiWi5nQ6
+iMrfwuJ/LESBd5ZDcPgPbqIWBe5WU1Jw0JADt3AYEYL/PDh0l4u9PtieRXgA/gr
6+1J20mH+2bkI5x2P/xkJA/X0/914HqOfG/3IE4qbCKX1GG2ktutWc+8ahdufzCk
Ch1bDyPelkTQoVSdMDaHN7l45Uab/DKT/e8ByVX4vTO+ajEt3Sjkf2YcghGjQtWq
a1tjvm2xAX7tUW1whemk5eGoBgtmcPvZu+r4Tnfqe3k7jbjkWaJQbXAcu45SVQVs
FVk1Eykll3kGRcKpHWmYoVPk4QWMdHmxhp3n0J3FEoVVlnT03r/hEGR21OdPz6l7
nmlXajPCmrI+qA5HhENsIw3VEqZnwoh3Z4DwcHyTaqEgMAkfxcd+9kcEeNlYePbQ
kaGKFjQu3NGwPTBVmqktxDOz/grEnpmkwMyLpvzcoh+5ZI0R+74xNYmgoaaeS6BX
UNk7ubZoIrjvI+ckC/IGbo11SL6HdeJ35ljXf+gq8VllVHumjIfPrkgPww1IcGZX
Hpa76th4bkrd3yh384nN/iWUTv08EPxVXLHz2VB3lvuZB7vEQKqiSk2Yo6Mt/7U3
AoWMjIf8birD4imvo6MtsazKHBA57DPE4h8Cx9+ykKVdq6ekOl5++j1shYdm9ZXg
VQkssW27Ig/aGEM59PN0n5B2eHlFZfxiYByXtBW7slFr6wvd3cQLyhXA/MLvcxQk
E71GQSK/BWtTuQ9K8ZXxR9aNkNNDbM8BHHGVlu9LDRFeTnaekCVv/0mmTyW88vzK
yujzM7tjUXJklhyVr8JRMHL08MEEdykkUmRJZeAcs1TmRcQzjk3UJznvmbWeyay5
1n7h9MiacVyRE0i09K3YHJ3Fu36TepyNWRQkoisO83kaU3e+moLcYp2LXS3eS5tw
Qn/i7Bi9ht14OWFJ8yjlhDWsGDlg/xMNmBHk3vLwXFfbj+VPSYLd5Mqqo4TWQGXJ
K3hBRUOWeCwcLQX/CuYNEyWZpTnh0QbybC36yaHi2zynpPCexAPPGcWxoBBAsu/B
0q8vMnkgguknUym4LgkDzw7jgCSfJfW2octRtYGa995q0gv8OqfX4u6WnG6NY+vk
wCUx/I2+dZRLv9M/dBKNeX56A8O5bHwyWMB+pHEaaRC0NZZNwk67OvRXB35ogzVS
5LrdS7qDZVrSEASNxolhvJDExhWgc7sDk4GcxwTgrZmK3o+7hEyzIjESHefQLQ2R
1t6r7hzUrFBKKjPxNbo5+bW2un69MaqD5+ZNbbedY1IACIAKH5Do+OWAbEdUFsFH
sYZnQRn/Qp/EiZlnqNldNmCL8TbMcRirkZFBTLTtrpspnn5sdAJEJ6FRSjKQbmtc
k3h9or96oQoPhuW9EdBgx4i+PJ+yIi2+ETzW1kUmNALzWQ61I7czud+3+BZXxX0v
+CzgWt58RCa3yZTwDEsLR2+weo77mAKHQLUCf87Z66wpk2Ulm2vuZg7cn2CAMBZR
YC0Xcqrv4uGCX8WC346qNUytW8sIR1Lmc6QEI222uycGF32LsjrrqpVM+3CFxAPT
ClA1qSAGE8iGagTZOMSY3raOyops+FFkpzSpP5TzOpQMlCJKo6uZi2Eetncs2RK7
4rd/fogDGOxDYu8aPNNeJFoSwoOEWvOoHz6LSZZPL/nhYdmv5WFgVLl5r33ows68
MazBMM4oXFaB8nqgbMq8aHmyIYaPpzg/LKEWq7tGG4Ua0SPyRZ+sMcqAkO4EqdwC
7/wNcIukpJsay3dFQPrIsbA94QLNvMowv4Ut01LXUjx5KFfwTSRcgTcQ/o+LINzj
+1Zp4pt5/YbI6SL4gz06mbyRi9UW3QnbbppjzWrOj4xpzwXc+baeLSn9hRJ2lKiw
+N8hR/LbYH+1aq7fkg15uRAsuXwXjX79xPa4DLxz2NmVhJOtY74OJa0Jgqkm5RC5
Cp6AdgygzI6YbaRX9doKJc83134fIncGtUszBgPGCLeGGVL14iyosjpjFCyH/9FM
EozyCqXdLmUKLDwK5LOhOTOivGIXx0Rma/7fLcl6CjOah8dzgb7u/QuFJrE9LwsZ
ug5C3jZHLvLOv/XTqoqCrvXLO071xgCxR4dgjmfzVhgTcUdwiEMj13CVn9XsNyPc
EknnbBDDokKuzBfcNrckvXz+umNPnl8AODxQi77fgXo42zr9lU1TGLHmRUcgrONU
II7bXNLx4qY+PiarnxtbHhh6lJ2TFsBZTXMFj6Gg8X0jR2fi/hjZMtnJo9nnEFQG
ltJfO8m0a40MPaGl8/PuTd9FODsaNFNtK1XbeDuMqiVB+LcrQ9vsRVQZtyTk9e1F
JQ6Xm3udgzJ14nITTOZUpwOy4RA2+LGqTRflZ/fCWkaDtAPxc5UafiGk4bLGj9yZ
MaxwdB95ha/RjBywUBUDZl8RMhGbelDrxS3ItXcOI/DFrPQF/s6LzIxvenL68r5w
4tu7Jr9mYr7Blg6Epb0lv4ZISyw1mEGg4Y4sgSk5a0RjtRt/+/Qih2K06OCjW+Y8
3dOswpse+uevFw0qwALl4+ox44peIrwTQ317irD+WfqzwIz7n9J0lnYfJ4O+VhSm
E7oplh0cc/eAvGU2zPjA4WRtHgwp/dKlmw8iBrA6duUqN+9ArpSep/+ov4Lmthhm
lvx3f4GYWllFqrf0E6FSH/l9rcd7iSSNCGr+wQ8+VF/9nYxDNb6spba1lwI65t9w
iQUrM4SjQAzfi2KtGFTv/orsZpoNKrTskSIqIeTFdC4iUuFF4Qn68TdTlPmtEJ61
2KF87r3X48C1ozS+q8MvcF3zYFjbKT8EuvnrZ4LwEBph7TwapXao3fhiOZcJG+mZ
24NVQb1vvB/2buZP+xZQ6m6GKXED8Sc9uzwif3/hBENsUtRnbgRmVwIWONPiBhP1
NvyYmPmtx8hFS9JamphJydRs0BZarqU5OdioIlao9p73hkkaLnMAYeND3jsm2huI
hrSoENxtvKlGVlTIRqTEYp4tiYOkRM8uCNfrAd0bmSKovLsJQnwY4zR5375kwmHN
SB3kM6Cy0+ZZOiZVlXq5CSfr/gxC+qhJf8B0gbWqQsYkTeGynLvRhdyGM+Rp+HhN
PzttpjSuxqWfar5zFyXKxl5Yg9NCqeT22Ch4u8yT89/s0y595h4wp0xQCdRCQrEK
5ExocOKjk4t4vaPZmGCGwdPUGH8jn5YaSklxS7Foek83B4Xovgu8czK2eNS8U4RB
raKBVpb9y3JnaBtLxx9Kuh36G237zhcdl10PnGQp+o82f1gC7q6HRilvg3W6mQHd
pwtL+VxEWv285O5txPn4kV6jRHnVCvIfrj5/EPiijxVTtNh0ap6Dq4j9npmFMV3H
Saqu3Yj3QBRrCvL6Ucj/L0+TYE1Ik8tcztEnJhJw6g1rjCSJjcRbi/tZN+NWbn5l
iqmbW69qf25nTSM/f/T5tFavxK4h4EwmRzB6RW8sEjDL0xl8hnbwyq5kseczq408
7bmsuA3W/5wkdxMxwI8QkfitKi90W1Y9KX6NkTSN2zdMnoXfIxtaf0NTu2uQNJiN
62VyJiU4IXXDej1n5ppbsXoDLFAzFzuBSmEV3qYrbSuM/IBbiralMYn1pmjdCoZs
`protect end_protected
