-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
sdU+wPCZd0dgjeuBq92gwPdmakxJghdFmtxM0femvsmQpgtkVESvWjfLVpgijjaQ
51wSpLCY1sf8nccwB4sEdu/jAb6W/aIYqU96rziXmT0ZYeNLTlx4X/3iHKz/+Ej0
1z7q83n9dmKhdAuGzIaLA/RaNlW98Yh9sw3JPNokDAlhFCQ8wkEEPg==
--pragma protect end_key_block
--pragma protect digest_block
WHpBkKWLUunjeTGBUFJL7UtoFZ4=
--pragma protect end_digest_block
--pragma protect data_block
40rgu6rnSdlrSBsV5s4/f/tkzb6Z5VDhe9NA2Bp1Yaw/af6pxLZH0g+PG5aRImyz
3Uswmo3gF0kiJEojLONDypJhCnB+b/bkgNjWw9fdwVA7zwTyrVELUhRgnJbGRO8j
LhuuzHgXZ1dZvelmQauzBvUpyPU9Uvfy6n19I6DIZ7NglrniBorG8GYwE3jJ12s8
9Dl1G1ZgxwahdCncnctGVhKIHBVSq6jeyBKbNEP8L3EPLEYgTOipgD0MGgs9SM/9
hTwlTTG17PRFy7z+yInrTkeH8U7g8S1CsNdLHKGRX2FoTE5ytbYCU+Wptm6BfE+C
xzIbr1GrN8cPYFz4ibAWtgDMkpleojoucG48NJSSQhMjQ/7LvjIrWHWwsNiFpqeD
BTgARiPi1SVUSmtRfxrGP1og2wvPMyvo6wNxwtmc4qR4TovEF++DnrEiyEfTKtc6
sMV/PLq707CFJTa5oCEJaaPOBSIQ7L5G/Ch+tIpNR8toXzOsoF1gejl/r8Bz6tEE
mHwSwkLvfqqgGaJowf8VT7jvZnf0o8pMvy6dg614m+dUmr85nbZYWCYPbP0jtuSW
9gg8Z0z9JOrAqoUXnJKUMznras8aPYwAgIIEU3mex46lhkQtwhLsV15AnBlgh5LX
ldsYzw2v5FYxbVFVck0CW7KycUEzQ1uvNqQfEh7bCm90vLEzvq2rCBIdf7Fs0Vdw
/OWqbDC6hKdhdhrSX42PrIIfuA2yI6OSxfNTWvI+KixY1kdf15s1YvA7bL6Z3lCI
Kxad+p2TCecnh1BtXkA1D6RiH8XQJJbHJH+3LSRmMEF/kNYcSOlGTmnHk6R6TaOb
+oi05LtqNKvvgRRQL58E50Lp0fKsUeykxHwsrcOWdm/G4LZbGCk0gcQX3k5vRFLt
kKxiLwfrlvggwtNSd9pPbkdiU2MU6QCfT7u7IFc0dGLapRJkD6JJmbzzFA6bF4U1
mupYX0i7WQ39ViDQXwTqi261xK/JLiiCVcMxeE/DbZGjFTyBgv8Amqk1sp8pEugp
ek4IgGQYvrHDp3z4HlxVyQ8QW88QJjdo1WFxoU04CrqBT7aT3OXOS855iahdqrU9
OIPvd3dtQriHa2xUhn4cPcodtgXQVcEg66OeByT+UuynGksD8M0mbmekDYJbWoqL
byyjJ+0yB/VcKJT5hksTxG+wPvFhRN1kyGfjUYgCx0KEZyUV3KfLxK2YlbEmx00l
kO67G8X7ZRWv3n4Fqnhn/mRFYEoeoWAm5wNGVmdJaTzjT/kinaSIGn0d/+CCh0lQ
7b5hnkF/qUEsXFg5rbvp5SE9svsG+G8CqFvqAqO3Q6mtOSc36pBu2Y6ue3xlDzkL
qhhbqhMYRLslv2oF2mUPrE5QO9zFQQUwQBOhvY/0jFOieVbW9Nfn3zEuXtPf4Rnd
Rxht5Tp8SCCsJCKKzzeTxgZDNpYPw+9xp1ORJDzla25mcNbZ3lSzN2davkfRhqrN
Y+4BWJHtSmvcbiin4CWMwggPyQeHGu1n5lOvvWrLv0hzOxpaMNJVBbJPWL8Wuqom
UsngcJESELP+2HuhmTW8iXgjZ4+7j+Po/VBXmjFqTkS7j6NU6mMANQEAufp52PyM
JkQPOcCJdR3GVWfHT6pcl6Dz1ozJFp+n+FybOJzUhoNk6H06aR5weay7ORZ93vqX
pmXrFWvqsz1g5MMGoajl71wfSdyESxYTYjnghqoVqLCw3Cqv94++MyacvJxGJ/Es
+qy21GkwQc6xPFGHND22eMyH3la0gIw7RB8fzDusMNmA4o2n8+DWIj8ca+cHefMB
+5WoyJiwd1l5lRKJ929fhYfqEONse4Vez+FQGuTpg+E3gxgtKNb8ujcaoBt3ry2p
Reba0/MII0rdcryGW1dyBewU4DZRIcmCe80FmPK6OCPvSrCaulEvUzwuDOMAg+X2
0VInmkmn9y6bFF6qPzniyPZaE6rB+g4v120YiFKCddh5jySXM/oKO6LchzmzpGkF
xjEtHpKMW6l6/jHUaYNkTweidfO7epxAQbpWQ2PFRRngisdSDoSarA4kw+dOmbKz
ZVSLxbb9MhlRGE3216L3gSDtfZ893ST1rQ2zLvZrtN1vKq6VEBLuyFMHxmzxoqyt
GUgneRdOllzEiMTIC+vle8VjLOeP9pnoddWGswqJW+ikpUAUjld4CX62Uii71pDj
PoPVjlNZdoRhBm64VR4TVne81V0ESWMJQDy0r1BC/52VL2nz3Jq7nzHxn+5BLsl7
WlgwSoaDei8emOPYdR5b7LhsPg4YOdNqQqOtfJ+SPLPJRufL9NbNb+etuL5/p6gq
/Ukgyr9rNXzzsZ5mD4fqKsltodXW37pbu6hdE/drtT8QIsbw2PbD2zBS2DSEXEL3
Jl+4xy3AtWdCAC+YqLUh6tVhge6K++6G2eibDZ9OTuNRm1K56G2Hy6iG3Xsz2AnC
fbt1vWsr53SFD2Vib6+U4Vsgd3pc3kS9EB/uaG/5CPBnqPyxBZpp3Za9xIk2XSKc
L7+G0QJI1fgdnjSKHp6vscK8vexfukjjdG49pAhvBzi4XjVZgyXMAyR057HA7Rwy
ulY61RI2WYvlX/Z+ThtcrVVnNk9AafazGbVdSKczqDP+Rz8jpjV0JovKHTcQOZvn
QpyCrLmUHZv2fWaO+GEyIIQMK7UACml4vIy7Plq0+mq1eJFMeckS9JewQdP+qv2Q
/xyy5+xjB8FocePVRRbbB1wUEfKgbhRgNWSMpO+uCSBnPn4vk7IU1ziQrcsAGuzM
tJOX84ogNjtsVDx5fmKeEzZ6FBhDNMG2xCUe5BwY0VXTUGBhProSGQgbpX8cvtyd
0YsOIwCIfWlgMg1x4PAucqBZi1ADTjKRUS/kY/j8Y0n59nDV8YCmzcqDjQm/QgD7
jF0c0IsEuYG4CMrIwKpTz4CEgwUfhSQN0OdPDD+oYjqeFDd9P2j7WECqBh+Qg8/M
kSkXSLKRXaDcVPxgn77+0SLl5jkA6afaHqUeRSndaHkf6nUdXEJbUt7SxPAR7jSp
ozPwCJe9XP0bf+LGNjaHKiy31LQ0/UzxmeS4/JW5bEcCzJ9WnaCkFy9bzNJBF1K4
7Wg+DwOD8jEAX4DmiLkFvS84sLcJDxx1WXYu/GNlAozmFrvOC5qBKZFviO/6cPNO
jl1WUvMUJoZXUUcAOqhsMt04L/sm6E8wDGuufMbEpKF1yRu6JuL1hUyjXUQpNhSF
KDMsGtPhZV+lSqqIAG0qbAIRgycGi9NiOLthJZ7yPjqM34b4rnw7Ctqlc9rbXVah
VU8QLIEqEYhUqRYE/GRFeNqAcp2BUV7rDuXfAdV/wIfhithkETR/kgt+FCDENyi5
GvL4mV5h/bNDm58j3i+zjv5jlEDHvhPLdlvxSZ2gwHzZLLlHHZvGZ/i0MYKR82SV
rF6qXsffyOC0FQ5KU3TKMs6KSzCHVZ2nB05I4nWCgACRZ+T9JZ9pJ/MdJ5OchisG
omY+pQlV5Lu+216hPteT8Mfs16+dXfzg9Nl+zjdv1NZNaCzljSOTCqBS8hTivBv3
YbGEFt3QFo7X5zwoscW75rFp5L1TZ/r3TaiorM+4vNCf63IqT+s3QoFPzRPnr9Jy
9C0sWrgntP3NglEgRgSVqzF1yKL+PczI6mCVjCyjri3XgCQpqj/MIXTDEc9bGRwP
ML/ZkkDSMxvVIWG/ZUCLTNSEUH7TZn6RhYsSnEqt1cfyUddKh3ncobGS8xzZ1bD1
8K7gEQ6cdNs4Z6MQA8C3VnyMDgmiQox+PudopzmGG69FpfZ8KTjvtXopap5tensh
RVINnjXkWtBClZGz/AEuywDLfcznw+BPqJkeUABOyBKqpOUQWBFAnc6J7laD/pJn
aTA7rK0FMgz1kRAm6zQsfvD3Kb/kAQnWeaWs7+Ac3WT+NyV25WPLUs4CGtWeTMpo
f7PjdYxZV7mz5qx7kehk4CAAcCSMFx+ffXlQIC0SbVasZr5hzAQw4Auo7c+k992l
n0aRSUs0oKvAWh5EkFglUjGIC4Ht5b+nTKOSlFP+sJcUZjBCiWnYpiNgonv/LGfB
keys2CtjjJYjWfWuY7uhS65zC76XYkCSsL1Y6Jr5Zv7uYBSqa98IIQQhcd0FB5p0
J/gljni+uWBgux0ThcicqdNCEcaoLhPYuPzziP4puChTzd0Ox6LZGpq8dqsYFIES
KKYVmS/LAbMUgb6z7pWNgvDbiR4TUPJuX1F7aoPXgXnYgBlGVZOTNqyfVFxPicMh
oYOTdXxobCg2U+inem5qIn0SoYgHpj2uAqO2lpMpT98hU5+FGIWJhCt1N+9VyHAa
e19zYz6T0+D9NJLshztTy9IL/KVjbKNj9WAaWYzQaSN/v6ZHRQmvm1mH5h5ouu7z
jxvTCcCXyLxxForBe5Tm+zDYm9biz3MUAbrKnrlsZvaV63P3AsPo0Eh5hnjlnSVV
2mI/PxfqBn3x9Yej66pYvtGUE5AN4bPd/E4w0Bd3n02AL2IhJDSAUY2m86FD4xu2
WJkycpAI1oF2QJ2bZjNb6/GigERW/mpl8ubPqbB3oxDSKC5hAFCGFYvBwTSnjjP4
7NmbHkxRXbcn7y/WdY4OuqjptoNabS1SUhHT0iMLOHqHrCOeke1DGTK95Ngfn/Jg
wYIuZcTzizwpd/EYpNNJ1OFXJNNPvKz0sOmdGFMbeveeRY/8kyQX5BTl77ODMKDN
gOOFt3Yo7pzoXEVN9/+4mmNPZhxHPDEwcgsP22Mb/Se6YlbSpOlUBXrTw+5bwHxu
zfUqc6JUkZp3f21GNiNqntvHGF37wcBAMDb8W3+2cyZIUrUe3dmHhGBDZQjHdSwf
sVEwpq1wAb4d0m6E9yFSJy6O+CWVztT2Q3MDgY/R2+/nVVjOTeW9pSK245jcVvEG
zFHGs064hOr5+TmKojNcN4CCOrLQXBuHAyr94HfhqzFg0ZCQnYH0um9HuAZynMVI
4zrK3meswjshrmD4W6xQYkOshiE2tVPy2U1Csy86Ly3P9bu4mXpeu7fCNHjlzeYH
GopykC8v2BQ8/BOWgXPrtCW/WXR+sMYsBCcpkmPr7+IrdqdyS6sLPB0qkjDncG8n
hBIB/ppFW2+F3dBnv4cGHcSNit1LE0mJR5YJ/9tF3hOVtz7EmMRViVA4j3emaDkV
fg0D7bcNqGIHk1EwAICB/2yTjq2vRDktrtHu9eMvv9/8SBodDAm5Mj5eaq70ceLz
dI5al+k7nH5Atw2uR7z1FYJN6J4qIywrAKHdKu0dyGq9iEP2PoQu9bsdRdMc+8ee
cHU3GgDsw2rm0xC/GOEQxqkLY/Tc9yGqY7vcUzhlbt8UDi8pX3rOLpCyyDR4psPt
f4zk2TyvqNK9o9T+Nkz0uWXvHNGfSROHNndnIiPmDZnVqJF3ndTl9H/kGsDc27rP
OV1XRgtwg9xi2zwbF3gxiKazZpUfXsl5SLV4NrqELrYrHKNpbrR+ogA+FweGjnG4
TZUFTiW9DjluTOvkxR1qDW5fqKKq2zcXx/LB+gOV8pW9m5ckn9t8vFvo8yGuM8Vx
DQ/cCLNoFSEEd16SupKCjU1o4t0eyCZFZw7APr2QnPObh0Rlp9gnJ43ZJjnl7ch8
4mVBaxf3U5iWWBmElxxOC+8KEDBG9w4teVD26uCQnVSOsWdVDOVd0MZPPrF4x2Hk
dAq0wpMMNwJuzFklnoxnU1doKSuDa68RGHeGs8whsMB7HB+HG04JfxZRkEtUq+DX
SCz2XlW4oRLJKIzHrjjcZGxoeyI1m9eR9+E3vYIV25xLmel9hFblbdulGejL3b2t
W5zVivlXb4XcXQ77F1xtRtdB0Ertm2zZx8rXZvOSaVTEugKAPQ2obNDWqS5/Xm5E
WNivjOAD2pf0Eg9PVx+K4blvE/DRvKuqPRVAGk0p1ACIWC6j37jYFjBWu09/uvqT
pATZT6YdqXTKYxMAJAdNUz6VKQky3t4Pguy9j8M0ytxfHIfDj0DcEA2pmn9RTskF
vB6jJeSjHT0YM4tipgkTpaV7w6kQ+LSOQ5Aq52+bHKEorl8oG6dOQgO6cpmibdDJ
NBkV1sxi29fqNh1gYHt961xtquygOnlrr2yROhfbS1BMR2ANkkbGyVOZ8BzGONUn
gD3nyGa8RQSS72ab2UpDWDunUv+8IfOXP5tmImv+5mb572YSCrs8HV+7z/WNSya3
t1mG9968fVeeKuqGkkPgyl5KtVvxN+GBNlnnMGN7TZn/+9GsWgyMxSUq5mf9zFCY
4yFSZW6EYXeCFCn5ZnO+h61lYKCDjLxtC6iHJdDFUsV1gdL4hebFmH/t5DCI7hPH
322PElzPIlMAxOcSP33kUZ2nWmgblHr2IrLIxlFJTNsemxdRY1E4ruhd8SCU37dr
G1waCOk5rZj1Lu/9xBcSM/cIOxMLMIIKTGbLqrcbo60FyR/exXDytumvIvO7Cz9X
BNNTNS3xEYBNJzJNQVtGM5kjd64DDuJHcBh60zS+M+RJ9UtWS+IT+AZ37QZbtpJO
bmbNTw8mQw1y7HSZwmmxlDtLujWgMrDxL/Zk6qP3aAiu3LNtSjTbgSqTjw2Uneal
JW27gbiHr08nSIOJ38KggoSsE8BwqUhj/xHqd7xbho0rRqmF+X5eBfSIanFqPZkF
HzA9nfL+V7mz1Y+9riW6uJE6I7iMCza+sVhBsxubu4p3dqo+rvp4cWElcCuBJ+w5
Ed4WY7eqdjt9utU3w+BugfOS9lYpbaA2ccJiOQwXbliDFl4jzwtgtVmnBEaKMFDV
gBBjYmoegyY5piNPe7HKa7ufbZbz3JA0qnohviVnDcKfTaKVGwfoMXtfCn2/7NrC
2xt2elQhsqub5D6wjegtEvYiYiwkb8Ki86uaaOoYnGtQmxy0fQo7XXhNypbeBUfm
tCAft0qh4bNYWtfog5j7sS6GhsHnonzDu0COhEJdLz7x5CmCRwMusJkJKoaS4h4n
rTnPDeN90qyMgpUD2J5KNx4bXXZncgpHTSPmmg4uPmi/2nfr0Uhuy1+eDVfNXiQb
A/cJl4bGkSJxbaLwwYstivqCOm9NyGk+KlN0VxSA+8rReLD75fSi/WfVda2cqxSQ
zZ9hC9uhWov9IP+yOEKClQPPnmPPHh/28aFbeUDS0nycNWapc8f44ql1YUHw5eMs
Llmqlc7Gz7B8Ak4o8vB0if/Y93q/R2h5xMs7AmBuLlC2vk+iqLhEXjLQFX0wLtqU
pxyEGOcGz/G7rxt2rX6uFPvVaYBas4k30L+U6iB+cGmkh49MMI/mT2pTxMlfiA5D
5vJZEfcsDGMAGtkxHMvkJi0dAEnbUEcovkuMoZvCXXO5P8freGfd+imCDo67WTkF
nMqA5YbotDtXdjgL+CeRIkiRH2Ti9UcGDIbm30Wwzx/b9GXN5cQwhJvCbm3m3xCR
uyEZFQnYHFiZW4Ak9BO418ygIqpDSYMsa067vQFenyajXCwJRKk/UY4stk4C6EMt
VdBGxfmTzRCVA5J0N4PKCbdhlwKAcPeEAlzra4W5JiLG+y2Sh3KPzIvsV2xqmXRu
kcTlB6dQYc1/BHj5FzRfA3Q/xO4g4sFX97KNqlZ5WkU=
--pragma protect end_data_block
--pragma protect digest_block
5izbfZMMYE1oxxq7lWveF7ocnwc=
--pragma protect end_digest_block
--pragma protect end_protected
