-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
1bgo5P+XK1VTXc04lOyhsMfocrENpclCU8aPISTQaASS1eEH3zihhtnCbVrCQJIe
FUsb/JYeE/h58hRs+oIz66bwyVShmdt6oqVt+pJSQswPpz7telQdmlUgVVBQbcHB
P+hV+fkNnrq9Ml4bGWTZf4LELklIKXaJlVAe22hHHJsKm30OHzEBbQ==
--pragma protect end_key_block
--pragma protect digest_block
uSQ0NHmKLKJuVmLzy/H7N1UIgGI=
--pragma protect end_digest_block
--pragma protect data_block
qPMgXD8SR+khyc/MZA8rjTeLESWliCH6o6sfinznpJx09NxPe5BVmbb+gl6fEzAW
Ax0oV+jASh7Ow10dq7/I6qT74iFPCXRWpfz5Tf/AA/1K4wPZgRW/sR4oxxveyMc2
xgx/aAdw/ns1SmDBKRxeAw8Ce3ebM00wC3WpCk5Yx0HkMfMFaR18+e5mMHVG2t3R
XMAun0eWiNapdx268XZPfpDav87vrfiMcog1ayERYUTfMGCcNux+77PIzfgL6OdF
FVi2S+RbhdtP6ItOAjp6bUjDn0OE0/NHxkTeuXPT2DfDIb6oYwZwJnbf6j5Jh8YT
8oRyECWguZ+eWV2+LQqOJXCMVKHIUi1T167bk8S9i3cZVRIq/vBNTzlMBQseEowT
T5zMs2Yevf9o82u6FWW41qXxrlKbOUYxzAic6BczUVQuQPsfn/9JpajSHgT9nH/j
4R62oCYHg/MKxUxdxDwtfkvmi7ywe5vXDFQnobEcEF93X7itW9ms+t5lMDmETJ8m
Db81kipq7Bm+Jbs4qfRiQJ/najeEG8pXsf7lv+ATWKhEhfD1lME1iEMgAWct9KAG
dWxyKH6+9U/7/7ZYjjS3v5ZZXZ3McTR8G/nFBYJbYJghbBZXFIrOfaRCiT1RL2Hn
5GjqQ/YP1wnmw95urTcqg3W9DPI3P6qTaaUygUjX6oFL5+lCdzh2nnWTQ+PEMWlc
2sDzr95Gv8tmJtae8U7HBJ6CW45KSpnD2d61NMCx+REjVO2hUNo0Hw1YLeJXZMn5
nSe+pmawzHI4zLSf67P9heaF1Mh/u/R2RPR+7NzhVC6aAC+Sp3tetWJuNRDOsgQa
gJcT/MerwY9FylwDfFvKhIepGlAxzypO303PrIAElJp3iuhXusPZwCyaBT2exPxa
LYk73j8UWzpOi6Q3aMRNV0WUWMPceORLqq7nEv8CRf329B8Yt7yD4O6neYRmGhBQ
crarsgsv6Yu/qHI+uKGDSvV98icTWvDQlAm/69KPQFwn+4IDgRhZyulZnh7zrsE7
GvwU9ejemwYnW5PioSTr1VCdQXnCWnB/6cY8OoKt98t4bpMqu1WhQiVyX9kcraCJ
u5Wsq3qZc/DMTifPCv8i3eg+Qiuoh7CTa9/UhB2R7LkwwrB+q++xuu/bPvEjSe1+
DhlHJdG/gpJICgKomP6hGJ1tTssjDNot5EB+iSs88OEtZep+NF/c/63t6A+jjV4S
8rvuDRLr5jhS3F5sbCi5UwbH1zyxEwe6asj2LgUC2yo800WeLVVraciobNEYoMfd
9V2G0+jK/YxZKdW9KSobZ0A/Th1YwMQcm9CsuxFgLzSaMAyUdTkXhgVa/E7kjG0X
JDN0HsTXjl/NsW3+t4xzEWr4v9Ycm9Z99so/NYDuWG0TyJ1WaA/p8ag7AER5tIuG
nt9vTLIGroYbU3XYR5f9jtX1spflxj805pWRNTUlaezVRRUVQJVHx0PxvZspW73R
oFP+ImceMDaAeGVJhoVJm2wMQ9pLnvLaT8MHrTR4HILdKD6OvOZvI79KlbTi1xbp
AKnjKHw516T6ej51C7K9kLhyQK3M1EljFAbgrsHOle6cFQqZZF4rtoWw8vzIjWvd
6LAahTm46EQTo1+mhtGG6IbV9pqr2/rNBL4xFg6l9cW/TJacm0uZMr82nSMp8TGY
xll5w8Zn6roklzjaOLbT46+2EkZ0HRGpDBfq29NPB6T0xnq9zF4hJO6LnUztibsE
t72qfZGpHGmPR0qByqSmj0ZCLzf9y7DRR7zh2URO8WIB8rloqvia8ZNPbbFaeSTy
f03eep8I9w3/HifQf++PHS1XrN8EC66pg1298tXaxo8nIXOWMBJKSMqP74EIKzLj
XZ/gCApGgntQFxEBU/9pwjjGJmM9/xwWVwRhFMY8JR6KcMmni1LU/72cEzLtTL1I
CyXksSwdaureb0uvdNMq+7ukZvsVbmBnVOLJIj9Uspl3dvi2fAfFRwGEHC03/J21
P7CZbJv3usUR/7TwnT/W3zVLHgzOWdWWH/tCe1cUeZFB3exFgWh0pQ3ao8Gzw4kL
vu17fHpeY87OZE+FUuuMIs8oXuyMNv/ZnQ9Y5yt6JVFNr8nx1hDrQxY7lpo066UL
fHPXMrSuOxGkdFxDoC7RODRVYAX8R7SJVSxgQv+Inp0Yb0VhX0uOsV0bLsV4AI/z
gsrvhPBLJGWXXlBH/mf5fC8IKKBJOoVZeeKAhFbcPKuUQGwFq5ecPMZlyf4hVMxz
9Ho+rdGQIyU9e4hnlIxS5tIB3yami9pNUPyH3qq0BlNtZrU16qba/YnnZV/a3nAe
DiSzVqKW7hnYQdZtmKHD+Jr8BY5kBZCDMM+Uuo8Dtq4KBfzbhu30/KhvsCDLUop1
TRmDiHjzRrt0tNFnMt7+wUzy8SaKIGbe7DGJtTd8QYuA783tdkgulbpyOWbAYF6S
UeRn2vPn0K8rM01L+jc/6vH1lEVgegm3DuS/gJEC7s1/IPdjWVTErvFM9gLrTRAB
IvYcJXqhxfPU1Rm/Cclu5qNQ3lkWLHMHfzfORLoSbjFjHOfeeHzt0Vm29trXnuXz
1+Nw2YbJJ8ldWXmJcPs+EXpBDSnYG5/wvppCjwXOvrnq6+Jl9F7+tqYajONruB7t
1Q6IC6TYaJ2KAaXReL6wJ3QFlb6z5OWTwKpZOYPaZNf5Sj3Q/xw3WcHacpG0Ed9P
Au5F2VbJQAeCze0BIhhpPju74VVo2IL7V7YefwC+nGot8NQVBOr7kzvwT3WQAOWH
q3HASMblsR0mplsgSF+JQ/pLoJjk31YyC2szR9qc/NWiyIguippg4ENmjQbTIGQc
WD+t/tIy3Vc+XGS0D+h9TCIIRXQwM1Dyad2TnxkKvAKT+TTQGyG1pFC2Osou/bUP
XmAg4bpv4DP77vyuftr4YPUb8pB38lTNRCwygRfO7dI9L6+EC50IJe4q/UnozjqZ
iwpU127modolh1HspPTGpLHTl5wyDU/og9lLtaJxJElkV6QzIpqT+Amm9emPWg5M
hM9osqKFvooz7xH2hLgit3ZqTrrrr2zfPM3jSuT885md3J//z1jUhpq9VgsRW/a7
qFp0ad1fMBv6g2AUJkEFVC+ppIIBvXLBeacjqRJxecM5LC+SNfgu9Xf8w7wVDNze
MTX0eYNUgGtjbNm3Cj0TYz1ejgyR9i+3fQdWQi9SJOCSMBXN0yajl+tyQQW0Ywoz
iyMLF76K0EZw9exzzx6v2w3sOKvvgohq81rOEixxApW4bamgaZPnyAimo1Am0Kjv
CFBYgYDVIkeaO8s/F1GHD9jzz1ctjAWay1w33Pkm+59/iEjbt677buw5gLDgQPLy
B8H8jO8kdtF5+0xT3HAux9kDh5L5ZT+jlB9h/5z2CYf/r0dCA8USnPc84SDusgGi
Jo4gRkBZ+Kjt97bUqkdCES70Ay5/TAq/uki9HdnSP9xZGJA+f8mxY7D5uGHa3FZc
iqFd1Q9VjA3DH2hUoJryf7gdZxOQwo0Kd/a55/rI43czI9HKIgr35FCytZgOEK/9
qnFSCBWVFbFcg6dBeZ5Rbm/PJ01kcp8pCHF16/YtH40YEhoLR5kmdMMjcQyEa8HE
GM2sK78nfR/WT3gdpI20Phmr/CucZTCZirjEts7y0Sga850e1WF6npWNIrxYzoiV
VO3jSM810Jydjuk2XLlHgVz5VYKo6vw1BxwcZr/TQVrrgks6p2mb5EVaCaoDCJZY
4+G96rOLb+CDs+t0ohD4Za4rVz+ZuPaa5ZS9ur1b/NZAKfEd0xIdgfhYhOLOESpT
GbwgYp7uwSbyOFrTggRjWbodvNuvzk6psvTICw3fOBfAoXxdBnOGLTmtyUsmDJcT
mJ/64y1QllnAjoKzIvuTdaenCrWwXit8aUSkDM2ytGFwvqpTFspL0w2ijEN+n3YN
+7KWP2Hr/y9BG3HcHCmapuXpz4CKqA2YkqxWmOUCx9m6apLyAau4MBGIYU/4i8BG
hC1P5zjLoMDBWnZr7bnF33dwbU3ez8uZpFC9cL1PK7qiGTYKkZfd5ErI5auOY+3p
BuIxUoSwts4sUHVUbotkvD7hQfMUWaeqNHyPSMYpVSLyDYV/suro75tbyyCD6tNS
C+AX7pWW9zOREqd+Q70eomX0eXuGyUH4CTi5KU9T86rYsiaiND7bkoFHS4hOqJnu
/TtO3oNi9bxzhO3vJUg2VDs0TbgCnoXrUcYX4OcDWKv0oMnG1+ejZihAB0KCbyUI
vTWj6jnbgbvDuY/me0/vTBNzupJeA8VYwUvePdSP25gsRQnk406l1jur/Vh4z+Mp
xy8lyTdPofuQwIcd1ZeEfQOnSR7y9k3ngRMDF/cB10Xkc2ukNk8l/k9eyKU5+rV7
L+tq54RNESMrxcdorgpNvtrmq8bg3+s9ZaBS2uCTPOBO1iIGo65zZapufv6Ii1q8
WE41969oHbajpFtfhhunZIDHk8tBcX1JPFsV0m/6TWwQiZkRmH9HIn5rhOpd9g7K
CT5xz3OsMUHLnuVJFtrLy+fSb4C1YOcT1IMaK6PFj9z6+BN6HwZgiMiCjbMXNe04
U4+XjW/aUJeOM/6UakpH5NhD2xg3RQ4gwOBIwTezdQYfpqg7W0GNZlBUiF/keX1M
14PeZuF4ZUMYxlE/Q76aSHT94t/jmNCr6gW+jOD6sQk7BKw4U7Mrz8OMMj170vRB
4iHKrwCRKmK8wtYAfJOQlLlgTajj+1OpGczOIyF/MRJ1Lc8Al+TZhg2q9r6beCei
fCu06YZkq9+oob4rBUvn/8f3bd6t2YJJlG0zXeGZFA8owG/JNYxDxLOIbetkVDBI
qOkQqEbc6fdNXRTkALgppBIadm1z783sTapp2qVXatLSUUhHzhwuOwYsh5j9i9KQ
990YpiFA0UCPyOhJimUBt8iExGnROBjfOmn3vTvYFVu0dl3N+9/2HXX8bVlAAijL
uCRgNHCpRXFP8f941ssUq+bEWSfLTAsb9L673wPL+XY5op+rXbDHKa1ltbk+gLrg
9da08udbazcMoKurmMxdb+3MEB/TIELvQNlJMEdJhTj+bk4n7Qxgzw6thBK6rlSm
P3YetKUDJd/85LxRpdBqaGqLbfD2Q0LibKn+Z4Rdrydg2TMWvnDpVT1OgkIqNfud
HdOcESIAIIjB8xwaTe6/hCaWq0NdgYoui2wNrb7F9KwY6+hHWHJrmGQhJEVK1uYG
JLPWwWbH5LtoaQQcsCDNR2Q/nZFAsTaM3fZU+3PFMKJ9t1b+LLQa4Zsa5hZ2D7iw
WQrhKE6MqxFkQmQHqMYcAX0LczsW+1f+QT+FQLuv4/goAnKui24TJf2jYkqgeIpf
0k5btAmK7wCYZlpY+3NOx1pDxfisXll8HLPL0k7kA6CwABzDMFXRaMgsPAgzir1h
S9ixmJOn3T23H4owsr/L5XaqtzYl+bDSq96DEUNN9DhTW9rOg6jncBj5nGhfKEkv
TNzvK9lgRY44NgELNI8L6pSRLlVb3OaVF/mnptefWSb/Rs7NGPbhROtJrpX4TBjF
r9o/gbOsdOeM/6fT1sGu5wAFY6QjWw/rTHAfg1tcmFykz5xVZHyVATHDdVsFwlm0
iTSUjL3EVHnqeQkW9tI/PnGe7dhJJnHZQ+30ylHby+2KJB98dRXP/aZf0vK8PGVD
aZzFHdqLKXqaGQ3Pl8ioQNnFryvuPdYoJ5Ea6wLewO55FPGRc+cTY1m9ZpEmyexn
kbApSqAb7njP6jicAkTa2yyJKvcW2uOp6+x0MNIIGY+QxhKKZeKJyDYmGECoteQ3
IsfdJYwwwJRcnwJL9j4Clgs8GVNJTqxP22jqq+UPTU0Xj21Aagip8ACOHLZRUkbe
dRsYu4TALnDagtww5Fgf9PML/qQSxfBCuyy6DsI8nzL1G6U7J7XNd8m2xXWzj+43
hWDV87Hoc1LR1MFk96/7r4XewFUQWL/TQYiq8hfrMUqTJL2QqUtNQGx0A0J4HfTk
fwKxAqaeosW7J+tpTcwGS3btiPljLTTsJf0krwOs81G8VewKvbfwaOa3XxQWQKcC
sxzQpPjX8SF5Z/aedNeHZYvpyh3bRseXytlDhT3jirGxcS5Y2N9FYhtyH1iCrF5x
B1NfZX4y0hxHtcb5sgtvBpKVxjSrh9byK/2t4tbYXWN3IjvHTvnyF7/wckhxSS8Z
WqWctmS7SFVBICoj2B4lFO53CIiBNp8fvmWGxmlOkish+W91OFeZYWfjQsG2Eh7J
l1/ykDOH9XLWYeJP6GPB/srSo6ATe+2Sp2DsesJ/rZfTeFa3FbwvGrlViTL7WVlV
bCwD3BnBkqYpQ3MU7lUNoPWYbVd7bQyfqZKG0W5X3OSrRLfQbrHw8AI6Kru3hbwl
3HCErbXx8cSI0HuKv5Ja+C1zt2XJTPbiIK8znEGHo3E9VEYqGHoVfk1z2tqTnx2r
phMvH5EkAzltP1buUUATvAVq5T9UVtV5aMflKvJwnTuFuGXOsWzUjigbd7Fa42l0
1fBikiyvOIymRMwDXztY+npvGJiRLWEfKbwGC+9DnuF6VsHOiL9nmSEcHJxJeZO7
HJEhZbmjR5An/PPtHyk4yXS5q4GsGAlBYEwAF0lX/8GrnVxv9s0bJyF6T2hyRcOn
hqFLAX1czWeUd7dga5PRX2IB8127/ERwRu5WbA3qjLOMJfNpMb2GnzOQFkkne3VL
y537mSsibPvBsPfNusuiGoAIl9Bk+V1O4rDEIku8V6L5y9ROk95yQgCAd77sCNlj
Uqjzq/v8xgF7HlRlnX04qxDaMSKP7XqSK4z8uVb9KCmDOGH+XUe6DgI02yXiDilt
BNu9AUSQLTvwBpfbcURfiGKea8A9/7KFXV7XdhkA7n1T452RfN0pQ8duij0bJu0x
rgVLrLwsvHvktc15gsfw/UaNlQL+gvNrzo00PVQn+tF8fAJuNchnQ0eRYjBsfk2P
2UnVP8iVF+pSqeC0hmfpVmbUXGLnysTpOwRRda+FVri960AVK9prlehfIIv7GHx7
/5Jd3R+ba75bgMKEJZdt64wQe4tidpXDCKwtbhsvJdGXuSdgQtP6foJY5BCiZFAI
3+w/vJy6yGqtdUcpu7gd9anS9tbQjwA4qea+E9oRp4i6rviF5I+D0wuELMt4IAku
BVVQJ/kYsJNbg3qf/IU6bkeabfllGyfwrMzBQxfJ4Ng0tw7V8g5DM2c7Wwyozhkt
5IERX5BIVwuXWE6ctz5Fs4F27pprXuLYKN34MWl2oOuHLL17AChL77P2y/Hvrfav
20vFfjllbbhF7/qnxARBsgkxvD3ntaSr3g4Gk4o4CY6jEt/G/Jxb4ev9v7IxuB5B
TRnSz7E4S6wPjMtL2fPaupn8W441KGiyWOlWXIdGbLWhvD5cjt9qslZwmE7yTp3p
HJ4855A/97jTrMsEUqY2zzLRXLICoVOZnQs1LECStJnQKjwwKeJJcly9X8A06fpx
cNTmRSBSU/HEiyywnMUcdjZ4bYMeBQKcjJqxvm4zc6goqnXVkSENFDDiVraO3y/P
TjsvUMx1raOWhKkO8dFtKnu4KhVlE4rNL3g1YzFkUQmdxLPwJESQbtQ+Bc9eXBdC
GHMBbLDTaRMlG9z82FvOBey0DjJPzClT1D17PCmAfAMBUADHFrQQzqgWGAZ96sKT
OPEwORR3QlDauV19lpH2wKAB7SqTeD0JOsOqDN/LTn/0dj8w1B+OB8kAurfrRMX6
8A4FIs8mJGku2u5MfIJ9TFWn0HQGdOZjG6uhtZTX+NFXo9uiOjkrzxz2mmcQBMib
Pp+o9YtjcK4AQqCDrNSrR3Ro5edbAYSDIIcJ6RZ8cTOq4jE3pDOg42Txxoe3HO/h
3lcPUV7SrvXeVlBCNgK2p32JGerRCX4kEtSCfK/h77AkOdTuuohbEx5g9zwYe0mO
tZmdu38To19+NPJDfMkCSAZIO82dUOrX3kDuauWHsRfb3Wm6E1XGwTOi9xhEjBps
9/QZyssEMxq8tfN3JpCME+AS/aqkFBV3rOPl+sw3Mpb8rb7Ph7nYJqZrrvIB4PSb
5B2IxlJXF16NiOEQ4cLPTlh9QfWeap+zkdOal9SV8qSKI9R83+8x4/95E/hKnJiv
iCi53UtZIaR7no3oE2W3t1JNO/2qB50x3VdP56eN3EKwX8Lt70IA0J0GcSv67jYz
QEp/y2C83T8Av6S8Vc30bekhZUZEENK3Jt2FcLHz5eMaHotIAdU6pfSPr4pIkbvg
Oj78omglhnK9gd989H8YGCWprtYEyFXnZY9yYY86B/s5iKWHt0qKoP/KpoEReymH
SF2m5h3bBWJSsSZLUawYP/NMsciwBdNkpIdgluvByqsJ3dUUY25/h9JKuz/9Y2k9
vT56QgercnSNrTv9HorsKeeUDtcscjVq3Cd26h97Ipl5nKNYzcW+7NfBAhbIs8V1
cQesBm5f5PawApRxkfjkx2bRZqeF1vu6UDdP/dcptK7F0XuHAJq7UyKt/ppnW7pO
EJddTJ1KsIXnlu09XKjsO6t56CIWWM/zfuJo6T4Wwg3xhIWxlsSQjfGL8kX40reM
isNqRLNbhV+wVfF2JHwV2sSrDwCuT0ymBNZePlqCvkBiKUyRUMaAb6HGJVP21R7/
SQsDCwIhXKWIVhuVdpmcsFr+6hEfZZCbJzgAv42sLaTxY9cabmPEp3dr3Y0x7foO
HAM+3BnDPPYeG4vPBUb+pgTkwwVgfdpMTIKxujl+4B7oo/kFQGATuwzmHpdh+jR7
r9lfWh5yzHODLSGc4TbFu1et0DzR6A++USTBIL9kecyab3L5eVJRFwAJsI6w0XKX
DPg7PcftCulwXhQP6m/1PxgxzcHa8scWbKezpk0axKwGg47idiMTcn1AQDekGWte
+uAz4l9eDmfqdfNrQcIDDmmF+7dsSuSlmlcukBDdr2Fj3PwxG4DaCYnhoZYjSXse
bQ15gJtVc+wY9ctl8mrpvhtLRypQBv7aKfxk4zITftVmNkLX1JiU0pvNcgLt4b/J
T/mRl5KZMFOcx16OA/BWX53qpwa1yZ4TMyBreZ626Zab9UD+Uec+6gTSF55KI6BH
gymAUYUm/PztiJPqbFDxb6I2b1xPxs5XJ1oWGqQBzDfv5PbCTZ0txLw3Ball2DAQ
fmmJ0NCeIvVi0T4tZTtrAWJyI8g4VOYrLbVwgr9+mOtU3dkIY62jv3nsaumwIR3G
Q8MVy3rLq3YkxnOzz433imnEAScpVOv8RsRrwXwWS/GZphppgXKDTF7UQvkdIuDZ
BjtAZzIOLhV64yOujaquKO5/95ckgU9yqLAUduLd6tS6Q/tcuF/W7mNXr7bVVP3v
hgVDzGerC4sYErO/njDacl/zt0/kasS4MS+hcwWd++IdA0vqt/zoHiQEEV7NFq3H
6FIBnZXhr0k0rPTWGcIomf414D7BPP50PtwSIgsyp7hyu7AaPNSh89pqN1ixTNO+
YoKhqn0ycgu3K9POTmPMLXAMHvMDoDdYPi9muYC4Uf6wdfbn3NTqwDVw0DTXZARS
ugAS9ZtwofmAGuJgK44Ldo3YtYpVWU65Iig8rO9y8567T+UJgAEhrkErWrVdwbkG
/dSZ7buISVJwgldD3V3WFmgGqdLmnx9yoG7xzxTdZcZ9Wv3lxkW0gx/oNrqn39wy
CYpuMUam3b2PIDr3rxerdETpdbMm1pkzTTc0ifPBK6KY7nR25ZNVr9tGiwHyChU3
2AbwkerJlEsGj12c9LBkGG32b1/5H9VSZVE6VLO0aAblBfOy9UXp+tS4kczxj/Ri
jvrvJBL/MGemFr+xFZE7FrCghCXaCIRVDCDDVPm4PZs/SBhsvH1+dqgYeFSYhArO
WAB86nrGNXKiREVYNjoPBTx525FCuhCpGiB3v0HkxmQAumAdwcQG9W+6wcP061C6
irbZ6JW4ED3Q6G/V+U40McN+O/NCegRwvXC8JcErd1A6WEmnR7ulMPMC4JLf1niM
vUlzI9Ua7Ee7ylhApi5aZmG5LLNKiNO7/0euxVcADt3aEQNfFa4PulhY0ugyLF7L
6J0nV/py2XlgNKThE3OO/yn3aqqJGeh81q32VZuuv8sixGbACreQgubnQMYOp/sx
Jra7YSzKOMaedZLryyXNxjb/YC0b0zI0gJy07J09qhUQHcko5pIH5ynomNQ6wxus
QmNliTX5tRuLjZi+mXmi9BME7hosne8Y/qZjkRny6acw5XLSg4+YPKUd6LBMmWHJ
/OzKVV3BLTFwm2pjbj/WAqjj6iaWUCOf8AlfNUFdQSW/IlsGtStrHs1O5pUQePfe
pkuAU1NOUi0bQkuaz4tR5LMa3MGbB0DHXRjbxYX1zTHSWgK/60vHogY5lm2JKGtO
ns8cVhNXEq/DuwpgQ696OogVF1N1FB0X4/KaLoMoAJ3/VLvT8SvNd31IB1jJHibn
D6L3zXUS4RyGmYlxzT8DaS6uTYh9YqJaegosemiVQ2GivoBhbP2J5xTPP36uFNE8
ay5yfJa02J7At0H89PPqkxpygyVH//yn2MNXGw5Eif5yYw1r4EwES2eleQYG3P4O
2w5hSqfi0QlPwNB5KDX5A/4uc3sM0v4GWs1DtxH9FKmFOSdqXhHOY6k96fFlHhVJ
idwtXcV1wAkCds78WzGvNknBz5GWWNdsaEJRD2qmv/43ZOpXn9kfrILgrOj8Vayo
3P9ejWGzMJ05uK7ZXdX1T3ApYzHWtNUKiYIG3MFadZciRShzkDNgvnmQFMW/+3gd
NMQubbuXod7K3pqKI0M5qRQSt46XwzVfoPpU2dUjEOVNdHXLea5IuOAXyXlD0Tqg
7sFlttR8myQzBzG/wt1UbfOQekU91ZWhY6vbXxv3K0U9+Xfr27vwqPwufADYOAB1
YI4s9dso+MgaC/yzNBaQhcLF0NxXxtNkWC+AXzAmxab724zFgmgCnQnnj3g75tOz
1PoMYuznH72BQ3xraLl5GzQi6+sJRP++CpQZOsfW7zLHyaLb+BWbMqxe1DgBKMcp
KSXuHJGx0t8D4Mp+8u73JfdxAfXdiwl7xOI54KzYSwwpZ0zhUUE7YviOH0lltRmt
gWEHPv6wWIOay1vieD0Mt6TCpeGoUEH0Bc+HZ5fIP3XWa37AlDlYBhQu74SSh/tp
V9wk8YaIjAtM3jOHL0L6j3ccjnLe4HOlTesp3BRMZ1gJogPOHwUmSzFNz/fVob0j
DuGJIU7PVYPJeJMamhb5shmYWudWScF3DjBGNwCe7z+rK8RtKBUkWg6UmeS4d8uV
1BdTozVqun8gEj1kx7TGoq4MqwOzeM1SeIp/x0a7CBeN+bFGdehH39sei/VASI0i
2IMryneegh9f592LL7s2SKYS0Es48VIjN9Hbk8vuJcQ3pK9i/VKoNSKBSivnHCfn
eW+9cFpzaqEzoyOuMEq0wFtWr39Ys+goviTZq4SMqjfg+TiEExOpnRKMhci/seOR
VP5yVgLBohauOJVy9kuUwqa8EriONF3DDQ1gs6UlLtsF+aCP4xuRaP3UrWiFDnSJ
GuW+hzHG+i9+niv/EA5DE/A//T93pisSNs5dcybRgdVNbyRY1uM1SovUJDvJJImH
jcBBqQmCVJT1Cf7QhiFTsI4i1prvDscnzySEQsZ6/8aj7ZrqM1RjLDm4pZ/5hJ4g
kEEB+683SPwMcw4z7eFxLJijlzJjfCxuSUcMPFpwgthEazFNR733F7PAV9iOkY7o
7QlrxO+c1f0/wvGIHVk8dcu9izQ8rRVdAEaQ1sXKU3Fht/kgXIpsHCl8AC9mSxXe
e5CZw4G5d6PFQ5C4Uyu2LJi2Q8eghnq+Gb4SB0RFrGYx+oTGQ2oCcUJvzKFrSZNV
R8WCw/igckGeMewxxJFRy38ObDMyPO3lRpGl4bk4qMBAbMHA9IhI6LKWq7iXjY3/
L6slf9wV9Z8vPQlY54XVjteB7DYll0FmrDdXfUQ7QgJPfjrRR5DBa6cFGOHS3fOe
WYpIUevyZB3WV3OpniKm4NXlNID8WSo2hJ5JKuEVrXh30IyrZvjZMLroGsgbdPf7
AThQR5xBmg2e7i2tuXvXSjyYw8uyxT4RwDKc25zW5jrbe2gVOTmYk4mDQSurHdDN
y8GP1beSRIZZ82XMy1Q8JW2tA7tbsLLBbdV7y6eFJGvADBZQsjay2nNiYSZl5xyI
5qbkCM9f+dPAJWps7Oh8iiKZGFF4URg5MtYnLojgpHY6H53QPv7FZl24BRE8qVms
AzLhyl5JyUvVhK+jK/US/tyMhq0bUXqWYzkpebP7Y80zB1gVfvLblVU+voPnurH3
S63ivmOHv1cHJvwn9zXbRBsR/wiiku001ki64k7A9Ti/PGPayWq8XbHx0kF8SY1X
QTo4VuTg7oB2QRrep/ocM8UB+Wg5sYNb3YxdsOBnDtOPvWQoUj4O6mdzw3IRV11B
KcWHNfTMvD1Ure5/OnSO5q+iKEwCwkILKMmp3Unnrz5VnOUY2VSNpEZqkekgok6E
XOuc2s2zdafHj9uNEjUhZmNKbb+gVn/Z53wwhDLE+Odd4o3CahghezZO8Bl2EwGy
EjXDLSMXIpLGm2CKxQiIkyf2tWU6jHMsp7e7AxKTkLiXwPo2A2stY5k3ErUK65Ql
zLV25rQzDztM+lVT1/yKivhpcRPvqg2+XlPlEKOPMH9sRxcyuFP1G+iQG4qZkw8q
wxhCA/5+jX4Exywl3i7GVN/kRRymAYKOMrmFluqZVuhKfPsdzWrV9JCeJfOsDJmt
9g9K/xsokExtbRGZ3P8fc7c+10svDLG/uhD+UeridGI3OQpSmGlnPlGLgYZMwlaT
Tb18RY5KogVzLkF9wmtD0r3Ul4DnfQDLztRgGov/yArgnS15vvNeguvKozqG2Z92
/khzhmDyHqeuW43ALjQXZuzAoMed8aOKpRbGdpoKvM+CMphRH3srcJk2R6fKHMQy
Hu7o2XRNEcnDuFSvNbngbLq9K1SAFKgB8QJXPBjhgj1tmpiSlVhuoosVbilu5/i3
3l5JfMdhomGtMflk6qi3IUNOZpD1cR1qY3eGzd/zNJiwkCfGAYul75W5AVIW3NOm
1U2fVZEcUpgO6OWJC5R2+iXJC0iP/pvjuCKMVD6M6r6hVe+tjfGHvxZxToXOO9ky
qplugticGoC1OZLECSt7m3bihDLpCKAqB7K6Q9nK2TdMTTBrcy37TFgvQRHpHOOO
fX+vxmPx3AUxFm5FUmWoeNdVFT5bIBgy+FPGuV4GReEIheu9XSj8qEcOarb/0h7n
6w7cTH43U0/P0OkHKNNiAFbqnOoZIfN9fP0XcxlI2wLvq35GknbAMfakw4lJ/YJM
j2q5EanItK0dkROeExTxuM5o76AvEI1YCfxxmnhF4vK+01ysyD47LScfyK3evNpe
6Le9wvtnIs5zMKHAz4FxWtIRFl3EMl6SaTrwfQtnEu7WkqeHY5CoC+b0Gh2HIvRl
+xoN18aLthBveHKt6VG0p5bpecILiDExU37RdscAumvLC1X92aFSCYFA5We3Z+b0
nx/snsZRp8f1dGdEFAKK6b3y1ibsn0gqAKR1Y0u1fSuTHARJx7LBXMs001sdljEF
/ipL3yHHE551gpFy0SERDJjChLbEUgR1hKzX/vW3trYYkupeXxKVsCP+rr/trx4a
frxr9pl2s1c/oWaZAGWvZeR1dEobtbjzr/14WQsxSsxhyPJYlNeVkJwTRA00FZDg
afute/XYcLERMIuRUuvQv4MI+NBRIKqbi+KzYcaMaCj4Zw8lr38iDy48y/E/jIg9
ZAi1+nCWlX8KN67oPLPHEVzPaP+h5AgUYkpPnEHs+CDxjFO5ELunif5wdFyyQTwP
MERHbqJk4EAd09gWdOnU6r1GtJj7HszagwjscqhRvOu0Yv15hCkD7CXPqFC747nT
SGbKzXSNYfD9p1KX1vwFUtjffSq/rM0YswBo5infYj9rZGS1uOgvGVt9Z4JeSaz+
mcUiuRq8B9xhipb/Yu1jUQA/GcpN/Ql1+zqwE9etbwOZPaZSKJD4uAQiZlleSaL+
mKTjXBSGe9zbANer9qqhvA1MfvX5WHFsH5MNfkPQlcemb0Op6NWjuCDEYdBUwd5p
sLM+bFEINJRBXtEZk5b4Fh9idyP+mSnH8Q/18SY4km3ty0RnPuFhcgbsItsqrXRK
rth4x/dOdwrbXVJFmIzUYCAXbaxHrRu0fyZ4m55XORSmZOJ1MSa7hr1Y5rEsQmJx
BCBZ2ozVSY8FweesS0aa9l2TQUQucCWwpisnwIh8io57MtIp0121gLTHWSXq3ox3
dFDtQF22uZUXT2rOl1FlmVS9lBs8my8nnjRd+5MdirWbHLRkPbaeO2qwT7VP+noL
hyS87GJtJHYqlgmpxyWnQdlTwLlBYjhoNJdWIfyiSf8e+TAJwEuHSldm7eWOC6fv
3ZMRmEhSh5V9X5wGx07RckIN2JYTX+IcLoaIsS5tn0U9B/nPNIiu09jDk0zAYZBt
oDG//zlQyqpxIqj6jGNl4AqhqBjjwBD5pOKr1ZYDatiiFUma/zhEm9P9KioasRNp
tNWa/9lL5kON+l16M+6Z1VLvQ8lTjSaaeLu/OiGVDiFLRyi1JgNGmQVSP9Kq+Gse
B7DQpUXkTQnNj5Y8TXV7YP4bVWHqf/SmzLiiYFiWXCwDUwOdKJnfskchEPYBWxe1
WjbhNaRHwcdEvkuLrVOmLqJzzQIQUnv0M+NHFeo6+B40SoH9AG2W9krHcGkAkONz
LAkhwvQbWK7TrsGhiwd1K5Sk69Yb5YOM7q56K4XIPjaPJgedoR+q3+36Fw1eI/4F
UPtNyO6vi0VvjeECWyqRG41pB45fMAfaRVV4ji2httlHqLjCdvrbF2DTcH7qFlWW
8k6h4W11zHW601EmEN/6p1z6OlDIs8sOKBUUhuEeY7SOR53Y0kcFJdsn9FMkXITO
gyeAE2/BB77i9H2FQGcx9t4mpEmlCsdQ6QNC8+ZGpoQzKtk8Kz0Ss7TMupwDbbwm
hclKrC73A1PraifCiaM/ISorBsSz7/8aL2dWsemrlhC9WlKk+OrOkpiVruZEeLLh
drNfAoR4TpB2WZfqaGizz3qSV2v6ZEJCQrtjNk9TsHegs1UKotLZBrojPpzlQS37
Or6DhVqLJFjeS/va7+uoQW5W/Q9Q9l9VEQrMAHNt3IxbvVhC2iNMR4KMLdlEl3Ku
pT+KQjndwRXs9FeqNTKoBqJF2rtZxT/bl/ZxA7fNxNoemTY9P6Xcp5IPr/zo5x9p
8CNzwLKhz5BfW++sGIjd2F9PVxKlpNJcmryebQMl+kDUP/XO1YeB+0PyV8TlLhWf
I2PWfRSIPU9w4+FCvz48fkBJT3UxSJed11p/vIViYLJECgY01kXPp08Ekbckp4y0
244sgFqYFbuVlWZtP+gR0lkNgIK58tqD+M/pvRQHLS2dtvvpmVosSpzRJlhsrSeq
GVzFrDjwcqOTCiUdqqQF8uksbhjqUsSXxZlLUzf9YcSBBufOEEvTiIY1Wgnf0+iq
J7asIPC7WEe1Wq/aIwCoxMixryA14u+7eiL4h/aGE6YyDFsHD7kyQ5Ax9mHW2gj3
MFGu/dCWzM1UZyh980JmiNUPWfjjt7WlQCE5g+1bQqemkEQzPNfxXjhowfCVxisV
8oqjIEYbvBX8Z1wa4mdJnaU++1phZRyyaLx1SHNOtcpxzX+GPdXepUT+pLFLizrQ
fETxMib4h2zLzZV2jFWY3baYPmyoe9RJ4AhR9a8gEYz3+S+WKfP4yCpiBDjk0+LI
fhG363b9xBB0U39YfIXAtoPdAXI/DXoTAAoQDAvQ3jUiBjISP1oROGbRjxXkdndl
xpdHer8aMr43h1wzrbTuoH61BcPmGG7LIwv0c6rIPfH/Kg1vXM2sM7/bnUGYhcup
GHsexkXZC3IqqGuUI4JeBjRgc38pJSWdBD5S/O+vLSZEwar6Q/fiH7k1uyNy1MIv
8r+An1joZirlBg4td/AIuI35M+0AcPAbMtWEHA+OZgPbRFfhPfEdzxyIxY4xlysJ
OkD2Hz43rhnxFHKdhW6dlfTPn95k/bRkTAjiljkf0dMs9vXNn0QKVEIMrPvkKyRY
bVbD6Z6qrIYvSn5zrF70/KBiYcXUm8qYujUNpP1fUgyGfdBeYg3WMujgjEC70kOJ
G7ZZqRphpPiekpLiPRkPP1gIf5yX5xWgksoDBuxbvWNdLAofTASz9pJ74JAyAp7E
5ib6dwj8LviFr2A7IQmo6Xd1CUrAOfhXYUEedyb2VjvI6SlIGlPjzWMiaovlvube
I19RpMgCxhgEXqyPcSB8J6b7gbIKgbJOolj98Z7qYRaptI+VumRTBpmz/v7IbElY
vfUHHFDydVzMqRbjvCECzexjgeh2AhL68aZTb03xpGewI9qnOSL4GRjY4E7pAkii
Le7EkzcQYiIWoSHC33Gm45V9IClC1N6c/OWf8Q7C8IS5+lbs44maCvsVqwgFCz91
VhbrsrPo6o/bF6D1suLO34Fb/rNKjp0gai3R7Sw1Cc3jAKWuagcIonwxXvcW6lii
TElMNoF7iuBdB5le9UFlOn7pz1VcHiPi0NCbN5e7nVkM2dThf65DejYAr166Dftx
aOVxYqcNfnFJ6eSYJD/JGHr0OAZlh+r4AsPbzVllpvfrZh1j1M6lFJ5KiHTg3Rhk
7tM9+/9GX3kdJ3sJ7Y3d83QrdVyQ7uHZn5NjBOlWHim72NRCr1FHnqdIHGyZHyjd
VRQe+53nPZdrxH9sTTVCusIl6NTw/OZ2r/J7dreafttQsEu5VZIg6IzJs4y6g41Y
pFn9EtkAGwnB5YpK9BBZF0T7Ih5JLJ3779zlrIdMu6x9wLRWP6xU7Py4nOuEMyfU
PT6A3dOTiPqAHgkfLUHyBxgJ2nv1lSJ7IUz8hfa1grhKvzdMADMvV5ylec6T9Ziq
oGYin9oJXN4kZyk8YpfaoNaYqGsR/qierfmw7ZNbpOISPTflRsnc7//A9BDe16cT
sKA+3N41ZaRRNKM+zz0AT7g+PFD0tzwR5JgsFYOOlLhelhBwm5K1t+7DRUvgAN6w
47YcKppQZc2ANKPELtiNs82Kmxc4VH1N3I5Ft7qI2imYZZvg4/TmMAb7bTrr0TAf
Z1LAh52uaQi/dltRKMLmxFv4k2m57Oxc4x9APXPDLM94M7xVPeD98i8P5X0pnUwA
RMAFGthGcXddrIArz0DUt0lSfHePSyuAapeWniWFMIgbWObT24PkCVR8zvCgQ4oh
1fHjinMQxqXKIXRSxhjOI1oLydeqslx/tvClBIT2pQArWgZkARbagi41o4G66DEQ
QOvHDulcIMeF33odTLxJJH4LhEVZJ0XwIfoN0Yz9QndAlw4O0CXA1WsEQAaKgqn1
aYI3u3QwuMZ7XYskuhD/MDJLkGDnWWl3zVFBo9nn9PQcrn7izVJoX/KYsqbiz++e
WSeLU3myFCNecEeBM7ukUGUN3Q+DANKKoXMSJNzxnzT9ypeAWgMO0cvHyK7EZHJa
tpiSS2IQj7UvC4KtU/2TeRn4002AcRE3bPsEzC3IA6I9wzKm+TC8gKDqFqR6I9Ec
mEuMwgobdr2N4RouKaMGYFFUmYaRDtdbfDjogDw7DjWEfZvUS/6wm2rYrK4OkLi1
HkD6nz+t0F8guK43DGe29d0cYhEB1MRjeLS0KldbP0f2fJIHFayXhGkKJECFuO2A
oMsos31fJ/1keNd6NwppqxoJ+Z2Qv9hIcrfQdXBsXprsJ96Qje+66jNA4TGl8U4F
Wqk8E0rOTlHuYgeWSI5UT/QuVmCQItp5eAAqyEMJgOuBCaC+EZIIx23JJkSGs+5W
/zquXfVi7QPNjDVoiGSUtMHGQZ6hElGfvMpIuAlTiRC9+AwhSIzuW0Xz39Vv/N6w
0CN5FH4bWYU1nDkw4D91sxuXGoaHzhzmzWxAPG3n49vyUHycSnlZzUEJUsAIcUcV
xBAjptraP4p7wqd5lqALRKMN3BERjUxBEka6qPt4GOCBXTQ+3d3d7GO/5PJqlxpX
w8QZxXCzoxrux97JryXxNvhZ25g/RfvO66Ka7tgqW0w=
--pragma protect end_data_block
--pragma protect digest_block
hjmKWennglAqaXn8WmI/ms0BP5k=
--pragma protect end_digest_block
--pragma protect end_protected
