-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
PilRUTubIl42bKB8sxO1H92EnflSSbZD/5vRNOst9D7lSttniEOoAy5As3oIxnOJ
9xB1Jcs0Lhcd7lQQJ/M5l1m3vATHxMm1ExoSyPUQGTfJyIgPEkYFPdAsBsCPAxpx
WRDE4B5azoWu56O00xUCOD2N4s4xf7+sf7f+HLRY8OE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 8827)

`protect DATA_BLOCK
uCEqDbm6Ea/YtLLsavXuyZlz1kmiV3PFreaWFW70e6Je+BE2TS2Fq921apOMc6bE
NqqSrEGoXEbuA1o8eeWOu8Z53qHSDy+eVq+qITO+RLQFcqkewhIiTmxDubSyRls+
JmeOGLl2SIzEHrVQ3wcBfbP4ew2/NcDzzXH3dRbWMFYVtGT7gIWXVyTLG12fT934
dYiEWQo9aNzgiPH9FiCR1InShTEiZIIylyhuD8k0YkN0HNCcMY9NMAS43pSq9yhP
tnpcnf84vicQljhVcLpRBCNCdyAFAbfn/CEI4tZALRy0vapIyTIEbJ0U5Te6SAiY
cLLYAxQVZXqOIHZXJRQwsxgrTMHb2exJ32YFw+7j269sSl7hbIEB8mwb4Widj7Tf
16j63IQpjtEaTOp93TQ8HwvMMQySO/L+nG+WwWnGNCKADJEwH+j9TDoEI21ZSfUe
fdr2VWn9lR6FUvZcJGweSGK9NrJxd6WiTSP+5fxp2r8/1npn8z5sD6+Cb31RCMkm
6CeXxyhlUPJjYYP5EUl5LtYWk9CY34U39QJPW2E3c0V69FZaDaCwlKUeF2cqILNG
2cBto6vBkPH/5MlXuTD7p4gwhsy6ZNNGqKjrCFVgkFVd4r4Jr7ceLLz6t8Aa8hxX
IkB/4b2kDx+6rhBZ2VZLbmTPsSjAG5TI8Q8PsLf1vGVQIO9VE2baLR44QTi8gvbF
UWoYV7zGJN8hcjtjvFscO+qy9eR3Koh7Dt2RtdTNB3uHbsbI1frPnmr65sdIKqZl
xDpyosXxAQyng7jwnYiGyjkvrLm1+NWre72+dxhrjNx9KDGmRNdb5ZycT7J/Zr5T
S+qRkRNUfYvH0be55sW1RrEItShcpGR1JG5DAOJyABkPH5L6oPgm6w5t18M8CWYz
bQGCYMrrtmWnQM4ihreK0RbNhx6qPSTN69ZNrgAGyZiUDgHpQKBv1K2wJAKZnqML
ZdmIyuJ9Y2kbDTYZhf5Kww+gDNQcpya/I7EsZi440WSKFJggJx+Q5M7F3D/VoarL
Xz7qKeT0NM3cakzTiclT268j2EpUmfdXMXHH/kajTEY1GHaTfnC62oxFNYr4pvne
cdAtjg6RZQ/2lSwVqPnd3ekhcgFnnj9Rdix6Du4vVhZJ3/R7BBYzL5eNMrqVCue6
RbyWgtmB6lyTMWPJddxKJQRpsKVYIRmrOMJL1sUBTXqOqxAv7xrgQMNKsZc/TZAC
Yei1mH9yiVv0oqEXdrROMxPynxjzFFP6EisR+MkN8WTnIsDFJoshKvuy25VAPsZD
nEftesh6EU03ZH1G6Mh9AdSe18s67Rf51KvJBUoDilg9IGrRGh8eZnXMxDWsWFsf
DwoiAYz+9Ss7RAxpNaRLp9k9C6Q3RODHpNWpfg0mg2NgiXsxubDr35dO1S+DIgZa
ikIHUMlO1wXvCuqKdilQ7Ak71Dcozbdu2pguEdLLRHM94VKhO0O3xuDdZhDrpDWi
oA0Kw1L3oyi6uBSCfu8Bsy/rx/yWI0INNx+0UXBl2Vg4+PT+y95l9RImDyO3yAh+
Z8LEvpJksXbiDFDVMifu/OPOtzMvZfX4tFxEPwWbGAXTMHjP7/JfKrO0jqZduaru
1iF7CG5eAPfUImRFrkkxJsLK0mQJt1IWEfLH3kHk529/6WnDkCB5RBPULLTTUJok
Vm2oi09jk2Y+ToDpAlVy80VMpDYPG7udnBTGOlqZXsqtgawjcErL2WfuIQYIwiUG
G0pEptl8cV+fLB4TyRM4Vt2a4I7xDNn6EZq54oCtO6Rz904ydXqjBHfXnoC4Uk52
ZhmeYw22uENH8zyaqyZ/mf3fp6yXGRccY3S6Q0VSShO0ex7EAslz16QWhkGIz5ws
HuYJH5NpwTTibtvcktyAdTiDgDbI8i9F9oIxBzYUkGimMLaCItiwX4H6twYlns38
6MeZPMt0jnD0Ok6soZTyujJD3XNgRkw4Z8ocLGszBbLmonS6kBjbbBioEiubwaml
hU6h+w7vFvT50iKBzG+XpGi5zjQqdsi2s4cnUV8nvok8SVNRsAL6HuF7Dg699ffh
8BHr/BxqxC8WFN5k+bo+H0PjKnxcuHchm27jMzk+tG6G03FC5jBI/WW+Claq1DP6
kW2TyWYJ6ssJ1s2CruYI7Ja5WWYxRHqCgTHWWvZy9ivgFaV8XNw+bWSdHW/Pjy+t
CTyz97CWeGgRH1POkSNXGfdSWz4SFYZkfa/3w43uGWmN6BkV6nTnSrUlPli6HUfx
E8yO4g9eMQ2D9yjG3i1LGoVvRfP2oGsZJO1h5ZFhTApunOmAntlRHRKfcRs81j9L
yTopmW3nQipdRT9ucJydMUz7DRCFXLRWetm6Z/ie1DxP9jywBY6MqzGE/vspA6Vi
OvlqByAJFbfZVs2Jsh8xkshlF8/L0djvJMl+MNribHnyiBkXihCPgdSZUIaFDy+n
FGNPIfu6QuOf3Q9UrWAVl6CNhkNFbu0VvD8laQSWYrpXMg3F3zgF45qLLT8ytlHx
XHcWYOYs2Vvp/UCvrYBTgwqmr34+Nw5LBdtYSzzNPHRXlbpIyyUUsbLCx709o/VP
nUmexBec0C0n9mt2eE/HH4jYMC5SAMFlKlFWm571j5XCD4LCnuQYzR+yN+lsNKZw
fYPcbUF7qrEx2gZJnUjtvyIlLDJmgHX4onu/fWUuZ4wDXJJ+6DLZNR4n6asQ0GKQ
nB8ZGiAQ7POFGSpCKs3kcuQdTg2hwledcYURRQxi0MAaWTM2F2AkpMaR81NzqbXr
HLNOAGCEyZYgLO7C+aXqHdUsl8JEWQ8I/+P/+nenq4P03glAu7ZDjRjgnwJ7qMNn
4fkKwLTBBE4jHakbtsSO6VatHyP8gjukrrdX92fuYK9SNZ81+3wOo6odn5PhhFHA
4OFzIbZOQm9F7AHW5xXWuR2Zm3utoVNs0a4YEIYv6dgaM57E8Uqy5vYKO5DAqXIB
L4RncYLw40aYHPHnC5UtZKK7VdPNu/bGPtJKcP8vpNAEyDZp/Fis8epzj4ns9eAc
GbOPeGWcmKXpWnEq3E/XO1qSSSIegR45TohbnSMCAX06Cxi3AD8Z8G1/+oQtR7TZ
Fp6DJTJG30/g9r61TevTb4+uPE+8D1c1AGzpwMBRDhVGqUV1FRrvVnBTLaCJsmZ8
3uNIJ5txw4+4RozFa+I6DzYdcCg/XTW3S0LVMscjid+/VZYFbGWA24+b2FU+/R9N
GPPDujqUDreND8DkjjJHAaSNJu0a52bXE9M2UyXOItJEzoF/lHA55V8AE3CmVFWn
WVWcp7tQItkiLq6yYbzKpGO4hrBWw2DfcC2JzUFigVnXJfGUeUOeLZlYnTzF6c7C
OzDpCelhNB1I14Y3OrAmqo+11clqJUa8R1kARZiophPr1sWpkYfQFnoJy86g5LyB
pXHV9wSPJOoraya7exatuWtnExEgDDfvafkwyK4kxg5gP8aKLSrBRYXy2CzdBJ7d
A8fsR2NSKiLQcUu6F46sDXDsRqLZeSyM0O08Ey6qfHytY/oWnuMkodS5CGEWNK1E
MVK7esPmwy+4phT5WjTrDpHEN9ZUUUgiBLCOSwbqxMnsrazes5wkIaUvKC9Gty87
CpfY+MvDoPz4LeMHkROsXUHuMAacR4++p+law3/6NNTsnbVU5mqXzzPp9mUoCNuJ
I82dqsbV1Xaes+Tz7IL1pIdmOKS/6kDpnIWgpzl3bL2qZwrA/wnoU3/6oFgbes/9
4L++H3mFIbZJOdE/Vzk5P+9AYtTX1iwyJJlCNlfnpzgwuV+5VEmpXzVZcIh2gWjP
/PO2pZYSGPVMTbASV3LbCnR0+I3zswaXgJBEcE+KXzUHEealrodXdSprHU60zFJX
PoZ0pm8hjGbzjExIu4ZB40/lZIy/i/DuVyvIkAOnlSkAi9JndUw7u60oBYRnY7P4
1+9dkPD00F9evsxk1tNJR3UU+rHPPKhwjN6e0I90H7FxIBGsNy6emR+S0gtOsIUw
sHg5RzBFxmF74EkTmluRxgkN8YVX3ApsuSvndVkb4Iq3R2KuQ44Iqja97f8ej7Ck
L+Bum0JHvKpzVX+ge/9r55zcMux/9nfwHPFrPblRppi8XRrHo9vN75hYkFsUkhph
FXATwQMcZRbZYTbs44G346aEsS8z7UJ16arqKbGzjYFqSsBrPumB3JWWY/+EKpay
fBGYOSF6yzPmGGsxti5Zqzf2QgdynTH228H60s5zrKNgw2sCTLB0wmzpQAuYBMDG
HxykfANXBGsMK539OPgDoAQl7oXPk8No6sXcbj9VmZAGzvJsYNSMv6EH137+sZd9
4/tmPs/nbVHJiW9qs6NDIfKUEEtA8EVnqCkjmxLbPgfRTWSspAIfGkvszqh37ymz
nzKVw2JZqID6hvSyE09A/ZA2O4sya0wwVTbwrWvf832rr5PKr6O6+xKMt2LYzW7s
tkqlzUPQUaKQ6jplcrln1HPMdrRy197URD9G+4IcuCtPYypK7KKiiAagy3vU1vAX
UCV/PqMOzk3NvbGQGqUz9vI7E1sQO4ggA43TdZnPQQDYwYABH4jHSMVFahBypjfb
ynUpWREg+hg6TIjglJfX19ViFl5DTcAk1/xUjEEojnBtLw0dwxwOchFVrCYx/Rv9
889JVNoCPC7vl/ZXGy32qDtnQjzlvxzhP38EcMXm0mpoRYv4QBOT9frU2yuYv0S8
bFAjLIyCnIN0bNWuvwWykDKZtb+rCbFVOWkw6OaC0tr+bizpyA2P1a0OdfTfjlDh
znV9LF99BEenstrg4mxunMtjVELGRH11AtSIh8l1kgRMMgAn0+TF3Z//42gr1GJ9
K6eKWnTX7Rjr516EXHJhA424LCBHnmpGITl0jKjgayef8sIhkQ4VmK/nM+b6VJOX
CJPMuldo98qMoVayOE6Cusk48PizUINtsPQLGLbENyHAQ9uMxZvVeU/WnzuiR5F2
WutcoZFHHRLqmxgKufLRhajO1VpfV2NZ0b3FsMf5DylBECHg6LVotj6azDgwKHlA
Dbj08lr4E/MpUz0CF2uXzMnGny2TquPM+osk22CKzYZKx4XVOBV8t+n4zFukp+Oe
HCxMlYrbdGvTUQlpOkOWl2IBoend356rYqxl0EjNgwtE4HLk/bHDf8K9WHmm9NZ+
ItduSn6HdOr1lb7xG4pwDglck1+HNrDtQl7en9r6mzMJVCSCDiHFvMnHWDbf1m/N
+GeuCdzSVMtMCrf+VnnGh2CPh2yr4YhJD/LTYZb9u7oHtalvV3IXbqjR3yfrrBxt
r/+VbCp+RuHKHPDjvahG2ELsc5boMW7w3kNVb034MBClFmPvJ9+htpBnMrIbsJPf
mrzoY+Ey0Gbjq9C7KZ3mgBo4JE/oaUOr8FKcMzk54i5UFYCDN8/k8pqxIo5WSFxL
8hMoPgSEYD+LMcJgkqsc8mLUqlGRmj9m+PjV2eJWDclngtqag9T1SL4ySe/xCM8B
TDpt+EhnYwVpzxqx4+R6kmAzCbLe+fO6tES1Wl14rHwxcNxt92HjJKOw2IAsd+gY
jNtR4VvX5yS8/Lc/gcR+9Yfo2Mxz2btkD8ehQY5H9IQx1V38++MiZJN6vV1KhG03
NZFP9wsPkHOXWnvY3pl5o6qW/zfT3oqLcxmexsFhkmo0/0gsknRka6e9IOpNK/Ax
odKSY2Z65V1Sk0+oqgNWr/NlohOos9eYhyFHoRGcFEtwSK2UT6WGNPeNEyEcpMGB
BUhV+9QEJ7izZVfdDd+rOIXzcgmSU60DFEhdVDGRQmXgtW6T4AY8MpuHjoHqdoBV
rMxz8UuoM56lGX6psuUfyczpb9/M6Vpb1VkdNwcPNcBgWVrgClegJyvhLBbSbiTm
YiPfkQ1upkG7oAfOFLRh0h86m38x6TEe1f365HLcdFZelcGPo3p+EA/nRJFI4QKi
bj2TL6gmB1zn8E231Eg0iY5ou5VINQZAaR2l+nFWNA+c1haZOIpiMasZroag3QNC
EchMY2Boy5TqsroTMrENUT1jkVqOotOYyb0oW9CVb3V8QcIhw81SBW8to67JHHo4
Ee2VM+Ety3uupApoyHnvdqPXoXaQjYgJMochQGHWa1bggBmEozijElWjB8rpeUGq
XtA6ed8ixXypFlFSO/fZIJI9ujdiUipC0Qu3oHMsroaoH42CAdEIJLdY3QzCYAX8
/RXvoynUKyOaFnVzNm30KwtdUIV7Thxp9iW/Eby3MAgF/wdZ+JzSwGRpSdEEpc2h
vNViOsEpe4NPKwmxi2p5V8WpxzleIdljaMRDTbvQQNqOiMCkCeXylCDRfMZ4GEow
F6wXIOa89uwNrJ2AFm8xGhMWp2XATcVeBSd+dMBXx9fzh6ZvDFnTVTXZL9lvT3zb
1o7pYogQ8rFCeYSc7Fvmf6WrdHReCoCc/NTs17tkpsgWk7hUx3fQHMblIkfqtTBq
bw0uyNpyGzy5eTGMrXDvxXEkGHeanjIBrfOGzeQ5XQeyl/7EgkmwmyAJPsbWxBEd
iDsuVGebTamY4l4qcTfKp4kQE3SuXoHJQwNf9hJHSp2njEFF+k4MiqEJN/ORVdJb
C3jbwkC744/vhJT2/anVu/br73g9JtOm6RNxrnh7L+ZPc25bCg2b/gwLnWM95s3d
OtYht5Nxe19f1hZ1hTrLR5MaWYuPegQ9pAZ2FM977Ao3QsaVOI7ZjXKlGryJuX7F
S3rt0N2K7dsycwWdxewyJpr5r1wkLqJYIkYV33g+ChW4kShwHRZU2d7qK003J89T
W2IkZniBE8czHAyfUXlvzmc4a7C0g/SS+tcBJ914IElEfwPgAXXT/iFop/4KEThQ
+tw2RD4WcPYjOBjVeswKbalLvK5z4EDvVgJ+yWhrSuGuhW46BGU111nhrZCElHOw
0sEBEFcDYXrMn4hYAveSK8yq5WOOCDPW0ELDB131vu6JnvWIGzuCVrlOj4bp8MfI
+XBfcXsj9eC6KuLpIsLV9PiPh5OoosXC3DYQWiPjWpH89UGNxw/tFadJNCKJBXCQ
Z91nx/pHU8/+MgNMBQHimTC9bWiLQi+iLqMpf4hQh09nUKPzfdtHi/viaRLubHuJ
wwlbaKUhdW5ay9Pky0qh1ioAyGIR1z6BaaSYPBGni6/q62CJvM8LwPfIbAFslHDS
E4FZRFvpNAQoqN7k35hbPpsX6WaveF/4YdNiVr+FwYIN8+QGKgQUfg8hgq3NDbhz
KlJel+oGJqRcxGsYQpWOFubnRBRrBOXTxdpvw5+bTizLxaT82ldpnRPyuTTiL6Vg
bWSDefmIo8LPRP8YqFlnwNn88asTNsAymQuXWTSyxwZiOuFOwgE1CS2V2yLU3Gx4
Iz8EA2Vi2VMWeDnEozZiPgsdBa5soaX/eLBZdMzhj0GIMmTSF+Xl2wd6tP98k+jn
pWuEcodStrYeY/jz5U6UmjtpUHxPbFV8Ed0fpYCkueJVFSuAXLZ6nlvcVT92sk15
cJxLXkNV6cLUM20x75BtxZndqw4Tz/zOWqQmjiRP3WUGLupxquj4UTE8TjbIqWsB
YS9VFeR1/6YFu3pyibq8SFwsQvJ+3grNPhM+tZSizTmVCZ+lHx4dkNkRQQ2kvfUq
sQy4QjZh4QEfdCZJXu/sirxFuFzUHgS0tQnV0dvjH679I+6M7iEwlBl+fRVpjEhT
7oq4XqI96sh6WzvuC3Lqi0uV0d7WcCG/D+hz3aljbldvVWQWC1zT/kTs29/17cyu
FAbAeVJWciytDz4Yy2i6DZayCmxQA8ZSzpXb/AiHsSSRi9jWAquUNRFIyB+pcvRT
nawwEA2Tj0b/tqsc7Xg8ToWMOKlUesm1jEt7L/tuAfmpn8AKNyB68krFkhmVR2WO
Y2q+NU7Yb/m+PrBUFp43o2rIYNv4S66kFPdP2upYEu1zBVgpAHSZomHGxwSQLNJ1
74SWk6sIqiBhHd6GaTkfSpQC+RPgvpLrr3YCzPocpUMuVZMtAsZSc7MfT4v1wMhN
bTqtjHhVKxyX4ZoE6P/Qto1w3UaMinKpwcoJShOZWeRSfPhr3Gm+1QJQvvNOU4KG
MGl5SD0X9Jr6Hb7fK5FVnUuskJ0MiTVi8LZ99QeAVYgKz/27vS7PLY4REe22y4WE
QQzbQ3K5YqPml1HR9uq+92c2x8jbnYAXDPGqsjAXebW8gUQsJyTYIFE/T8y0Fh09
v4wn8Sqtr5eqNfNV0WHeJkx26erlPFtMLcJt6rddHnsQwQL5fvDaHOyS19jD0gY+
ArNOu6lfubZWQ7vxdsuE8AYRmtXUbZbFSuH+00RNxDsfKXJ8hVlfEUfg25ThvKzj
oHvBUyL1QV4GfMAGE452AEcAjz+SEn92ArgKPAW4qybq02SstPDQAoCEfkLLldm9
K8qN4EYo9N5dWF8CwZzyUcwybNj+C1HcYOSxTqiphTBa07VlIz3jKKaWCHb6soLa
pDsmn8ULnI8f8nH6rCAtYoEioobdo6dBwQBbDVXZ6VlTLJT3TcjycmQdTppgmKVY
7kHKCm4J4H9h9hmyO6Qy/FLryRidFwnCqRShGBj41pctvUv7ypDbLSwcA5ioG7pM
sfgwZpzhUQsZJRAv2Smlyi7mW03SCIYa8zjYvNBac0/RyS+NzIYDBv2W0v3ZFfOp
aWJsHa1jNjfHwRXZNSgMvg02HtW5BOm7GjM1Zh5925rerppFxDaYH9k9TiYhODTw
EcAfVbRVL3x0sG9nSgTCAwqmax4vS+vGwVNomiJ2YNKn9pdWmL53z01Q923UPBF1
N2TQv6zq/4pSsGRYXyqgnqvInUjym0sFW3tPBZVQVSRlgFM75UcOwB4XhFImroJx
XGklU5+D7dY8x3fI4DDwOjvySkt2EU9LI5JFjFwMZsLKIy/E39nHK8/NQF/NZjYQ
1J5KJizCpqUKrLKzrYn/Kjd5kSwVvLvIKN4czTp2UjI31w5UlsrTt4l0b6jad9zw
uXwuSSOK3+sSFds0LswAnSDajW/buKWccmEQ9dVZMHQYWz20I2Tm0jW05sGpEygH
WgrCnvhVZcVQAIhQwlub4n5D/qWs6HVOfAXoi+x4Q4emCF/a2L7F7hcAisawxmoW
GfreKDRuGzm/eETjFyc6Q4ZNJjeX/PbEjxtCULLpPkEYrzEripFpAm5kcQUtwnpc
FbFT5DA+ZDeczV66UdD+w53K5NEXrcbAO4IHQnc8b1r8m0mDjGG1c3i8h3KhbVww
DPDcFtjospg3OrLMempQcAJulGKl5qMU2L+2xViOBD6FDVwaEw6zO8TfThxx2u6z
b9q40edENqn9uLPfn80YofNjTt+hoWhJc1v5xvUwFwoWKVa/cl1m26qIwQ7cp/Ag
uZU5Rm//WPwZk8zz23N4wrkxQ4wfVciIYd6DOh5kTV3ao2rE4K1UZc17i8vmIY7V
L64wUjBY+mI4CIERs1Sj7MmOgTYZshvjqxoRBf3CdGUe8+hrWNOU1A5UBHfqtVXp
gb2yUcQVda8V6KgSqUhC39KoWDFbELGyhANol2SaNlol8+LgAErq76G5RTuxaDie
g/nUrkacqB7GaQLcvbxje1IR9TgPubV0xgjNEAhY5lF77cpimilrqQk9MFn9fioy
QS7iAnEwtM4Xa265I40C6sQKgZqytVBH/ABnIYWG3C+rZjG6ScVypaf0qTcez05u
3hEFbMQ8K+IG0sf/k1wnXNW42Dc47tJNYv+o3Sf77yhxaURApeZxxCH36fiBa+aK
i70X0QolC3BkykN375wvHzfPZFRu37b78AZIhhJ51GE7qqOWttXx+YDUW6XgX2/f
cGQz9R10Xuefy+j2NdTYN4t05UAS3pD3ykfmuJ/kXaAAMxHZD2DQH2MPXwtT0ySe
tH6s9XrqdRsiiCFDsnjkERX4v2zk1Pdhrnp05lzedr3EK5A3CznXyjIqiOkEVipQ
JAUfPNDwxTatfB6X/WBh/qbG6a2axG2WFqJ0Fss/AbH7RBEnxw5pjm7n0d2tJiBf
BYTvvEm47I6Xa+oOLuYfNqnJGaZ1oHG1Eu4Yv5GWuiVr717Q9CNNrQoZgMwQVEPw
wKS2RYvX7VSQyGWZedaNTV3EuabLe2p+YZwNu44p3LTkHJOchGoUjYdJauKgEtq2
3BddfHe/zB5hEOCfNBDXqJLV4TSzbaNC7vFKf26W0p6DDCqDWBjqu6tKJgkitQ0/
eyKNNAVPuXlp1LC3QYSIxa3BvfRC4N4MI6Ppzj6xczrwXrbAo4TAZO4/suBaXpEt
x6bsmoezXyVh3RgfcSfowH4nvUURc0gx4klvCaBUOOKZ8UbriOlwsQnB3FW+K1CA
ZW0q6ZEZ8GxknWTkRllvX4UvMsuWnXBBpFuODxc833YXymktnj9gaCbbvuM9DSrj
UYVpYt8eDakZ759tZs78sE0ICZ5Y54I64zKmn+R+PghhZBLqYErjc9zMScwtkXS6
mmq54prVFbLxc/VOPj3gc5JILkf1ovN2J4M+JjlAf9ld7Xw+dDARzZ+J64udoSBq
/DuiXGagKOCZRGEaW6V3tbk30BvQbsJeXZkKGR1vX1BFIt2IhStXsv/3L0MTWq/2
3xaovt7S8TobFRo9Vdfp3vQh8ZqoT/7UK90+jx/Nx85+i9LEA5Vz1aiIDzpSqAHP
7PkEg3M9RxDGqqjNAkG4VjBoT9VYAnUoloT1eqWK3DHkb+gQtDr+YoI6PI8LddyY
n2Tz5bql+goBuDTqLLujB0j2tJgZHF3SWrIyUGO/0ijvaEpIzxd0zgtkFZDaz8t6
nlq12CqiOXvJfLMqstw/+EId+KlgYxP79CWAqPoyj3oiZ2DqOZTA7+y2zg2gIwJK
Ope9lqAomveNVFwqc3SgOYXfQ54qeID3iNON4qD6D6nFYUAGxgMPDxMZJT5C+hwV
ZmF+vkBGP8yLG0/nsVvVYrP98bhR/pEr94f0L6E4qWvN8kIM6IpK3JncSwqPbBI+
GSqWkyl0YJ7Go0TfkOguzvCwH2+NL0XE1G2zDDmm6I/GsptSmHUYwSLNNNAg8NLT
0ikmMFUDgd6MLplCy7Q7rH7WQj02256z7CoAoxFxTi6TqPfaJxnCnnWR0HAIZ9jW
dU2Mx5E78zq5a3588pXMdr3KrXIlF3hppfCUOUt2+tocMyWjYPnNM6+5DljN4BFZ
lbpEYiAAtzziUdSUKLgtPnQNDq/xDufcuYLul8DwGhTNTVNkAGR7J+mWtgnYNFQX
f9tt10N9PVVl1v8PPAg9LiOgAu18nY3sXopSrHuVVJGJThyD6356g1foMhtcPYFi
MvHD+oUOObuNcsbaSq/4RxRH1/SZL836S07veAcCTtidiI0MO2ZHFOOSCFcw86UD
TRFLP435hhfcYkQRhBRNCvPOxNqHAY4w2WAbrOFI5r0OWjbZqZITkKAahOoZpLRy
boj+m+JeadRoltUVsePe6AlMeCnJwch+KYvvkZyTVedyZLIz+1L6+hF7IXfbmYTN
4QfvFzrkIXWWmDs8FJnqCAShA7cJu64ydBsuAHn+NgvrOaZneYd+R4SPNi3XDfNC
G8BWXaAtA3fYry+td+V0PX4TCLavV4Cw5SJaVantQUiAlKf20g6QxkRQt4C05k9n
AKX98BsNwZ1ndaxUQCj1Hlgi5DIRgWxihRFK1AvXPaz6kCfKjHWMzQ+3VTPaU5Xr
5FJJYEpkQIESy+rh2AUO6hMzW+E6OvmhBnOGHK3y97Yibg9pMtJCk/XAGMfUadiv
knLEP/TGyInVUkSoREZuP5HR4j0YsQO7iwO1F0KIo8JMplLIy0RuGjhesRrxXg+D
Bok/cXZDyoxJmlW8c0S8tPe2JvU3vyXk7YLv/MbvvhuFvcbE9Kbl9kUXhjFxGLGF
q4y+sTnPGtXsGY1PifQ1bg==
`protect END_PROTECTED