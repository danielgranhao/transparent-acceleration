-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
iAD8P6tX7HacCld5f4TsepozHEPDL7rlqIX+mYkAt9wuky074VaRFbs2klYXKO43
CizopGjKPDxRr8vW05ycxTsgqBnPZquFbqynENdmJJQmBbubwzUIOQryiucv+3rh
/L6dSiotTvLEZpR6P3uPIUJkjMjHeE4EX/VsNB2NRb8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5694)

`protect DATA_BLOCK
z6cvF2JAP7BwR4mP3QuPL95pEh24fUKind6BxPVNOrMdpdXnIIgCflmC9Ix7iGPo
b/hpKjpNTYElbz3TkPCCAexDY4i+AvHjX7Psh8wg2BjDcowqXoa3NoLPqrYKcZRw
9dFdAUqNJ6kV8wTxwB19SuSTfHCJTah8RrbkvVRbNNmEFeiDT2baawtJZw3cMfsm
LTBFfS2Cuzjl7M7Z4r6ChIxupm7AXQWEZBddi8GD56nwUw507metoo6LZlPRQvRG
kxqHRXfR1lB0Zm+jiMcyrjEGfk6VOGhCZQGANqvmcwXbdbMnouMUPyOoj/OCuItx
0bfM0m5hEW8e3UFjIfaOX99L5vICnEo4YnEIhF1I7GqXMynPb6PDodkeD75LIL0Y
OP6QUfd5FMi/vUfm9CQHwVXrVsx+3vCNO+bcSwDdGyFSevvlti2QCBvLspDmLDCm
oR9xp3l2tJC6WHtFViG+o4YT/oEh/56tuhIhK/shPLzf/s5NUEWAUclsQt0/JIIn
9CEHweiyIpwssBRnluD+YT1AjHMZrPqBLwjeZ2uco4Dw60RXWNw12NuH794cgZ77
5elq8czgVanHpqVAPkj6kCO+Q0ttDUoJfBYa/7WwQN9d70IVuj47/fEXVFxI3UX/
BhzuNoz7vvCe1131EC8WdTbcRHPcyrzcAeJ0fWkDn4wOgMHftwIOfhao/pTe6ANR
9QUDI24IkIu0dJvFaEsfTaRcCrLn4nk2jEn8mKKWvCzxuIdTf10cM/ndW5RzZUzC
uNAobEkjlqEqHhpjSF/H37Hu0EieaQKMPQHPz6jXjnrQz/S2I/YR7zZzIgz28HwH
x04EbhJSSmccwGouVzw7hQrIyztSxb+tlXHDG1F9oWVDv7Kttt/0OTtnTd8osGBc
fzYVP3gw17dYue4Ih1dgGFX77n3PDQZ7C26QaEUpBiJZ2TEiUsVmr3NjbMxC9ru2
d6WjGtL6qvYtJnkT94OSdjd6xy88VP0urX+AFt5zF3nZUJhl7S8+GAudvR9ASYrf
muibnj/81Muo7L3slXFsRDf5Nsv1rQoZOODbuOmYPdQLFp1OsfTN30oygcyJ9KMv
P8MI/kjhwYUdiGfMWV3mkTEOHMUr/5N+rLvjSzY6rfavDyqD7nuLGLtH9R6/GyJO
dOO+Bjcr/7kH/uBjBg/HjVSbwChLPZeYK5XcHWIUHVQAeiwwP4iaupZGtU/Hu+2D
eQDt+QFKFuwFzi5bDSoWk62fLHog6chI0b0lL2f0VgJY/Pj/u0iWDp+1qUzvjEFl
P+jJgUKVwh82yk8uvgwnpD11AhamhVyA1HBs4Ua9RxC2QpDODRWlA8KLS8o1HH3d
LxukEYw+3Qp8JZ5/+dRZyTjq5Z8SoVz1aLwoopJwatvTTIbQQnXNTMOXqnxEwIM1
ofKqomaAbswS9WlFwrBF0qiBleAEjjIyUkRJY5XecttS03fSoOl5msXK4hOMNBp7
4MQzp+TELzv60EVpeT8qud33rzGYgG9iojldEtw4xEJ+v53g6uqfR8+OjTW6Taea
pNMtvMqJwXMGaegjMADXowwzDGzgI9dRHU+oxIWn5dm1XNOcmfcmJbapBiocJ8ex
aJbAPdCg/L17Iy2Z4ka2aiXGU+Ff/BO0JpCoGYZ8xrPrG+KvK1NwMqFT/jWJ25cf
B8VhzcGFfPXnabXIRvcz92ClLQl3PvhGFfWqx4YXmHO7VEzL5awIMzJRDtDDh8Xq
veE2GyU0ms5rxILcI7J5vDFT9+rVRvRVENT3m8D6VAqSysYAtOtQ3VpUGbZCRzww
co5ftWBx1ti3l8foE4gmeg0CN7o8zc2mh/DQYmeNJ2YwxBk1KqdEt7+89AUg4g+K
Y+Ag63ZhG2ak2R4Ho9uhPJ/v8eIeVTXRzXbMKrjbBIqeL/9CrqPXnNiy7KBCx+h+
DPeVUBtno2mDZ/9UM2zgJl7EBg2xT6CaeR6D3zBlj9PWNqnThs+cuPzbBBcpk2It
SA1J/qb4Ee7RoBTrCpEUTGYcgWkSODn88aKF262K9hePXE9t3fxdMoxlhuk8es+d
roRoCT5Uu7kZBNSXdYmuG+P4SeZGU7ktRWOzuabeulExQIyTEOc+5Mm8VMP0WBv7
bWgJYwfIbbhrWQCozYKdZW7dI7QUXObMRSiqan6aaZyfLdlWyKx2/wIYO/yw/FwT
MLf1eogWQCD59O6Zh0gjogXBIGkK/JHj6QXh3vbG9k3hHHR+Y2s+wLnHMaiheSW+
l6FQejvPGGL89MTw/xA61qNEPnAhdq/k8nAbPZfO3E0+SZrjs/NME3JFR0l8V8c0
kaUXTdlaC4uk4DbWWqUOo6XCHS2Ygw07KM34ZugMvgXjgruk8Rin3zpbp4ffLlFi
tJPezSDwKL+imUr5yXHIC9+M6CvQla5CjK64vKeU9RYmvCUVUDcFZqMb+zxC9LwQ
TV080HSnVldvttJyuIKbjv6KJNc/dskS5ibc/fFm59GQ9i90qTKbdnoDt3E/udNJ
HNB1csv8w2ObM1jMXDSOjcBfFzROjvbWZIB2CRjOYcWSva+NVj2gIlF2tdEgLRB8
eSEoEaae3gHCy1HRbtN3k01wcZLXfLEedK66SvkZKv1Ci2cNMi3vmqiX1WdCPm+O
SI4Ny3MBro3Y1xRMvk2OXe2/0hEpNzmxcOMkv3b26sbelFz/sQMl2kx9AmaF1g13
UB50bheJSH76zXNhPtU/E71bg5dcxo8FDnAHmEHRTnJWsZTE9whLTnxWI7iDeZHZ
dhFh+xVRCkKjNrczxHWKk6rDTlq+s070yuBqiLTCglEg7kuh8UxZy3rs70kSEr9j
3XD+S1MdGKwVg+Mp46rdY51yXj/hKSLtu1tj6pbnqZTlEzMVl1JSwkf+w6yGj3Y6
6ewGk9mkQ76s01Bo79ygUg7zG8/1MT/y0wvo/WDCJoA21k4K27dI3JHaXPq6tZqm
zpVCeQKSc83wRj4Quoi452RimPuwQYm4rHFghV3kAqr2BnPRPFK727urFGqI26of
zrrpVEoHv1tn2urNiTj0BT0GDL/eK0tzgZoddAOYJ/l8YjnrWW1Ci54hc1rEwfyB
Wk3av1KvwUw8CsRscp/KJ2bDrzQUjmJYLjHy8cAO+a+DYuZpKpppiehbmd2fvuL6
Pz5em0BbY9NqLeAambqf63e5fvdwrzZ9ct/5EHdz1MBEMpSiq6/2YKsiTVeatIrg
oq6jvFrE/km46icwuvm1AzcGuw9nlntZl/GJ6bT3p7qZWnmpjIDeC//sVGMjt5y3
YdE6ZMc4Hq02fA2QEAQTVxutxpqIFLy5LcnIQaGgEnuhvr21CNvmWbK4bhujWsrr
7c178uy6+uMaVjDi3GVlUg95Ug1iPUhaAb640eXx9mFpoChy4i6tkU5JLVeseFXC
OChG7nSMhlhC8UqPyVAXo2OEpaZA/wNZaE1r1MSGBXevecgejafBhXnZ1H937Z04
ABwGz5M3nsX9P0Lm4BGxoNnNT9oXrKR7yhbIfEKLJ1oO3j6+pARduxh1kran5xMi
xivdFb8zTyaYR5QQ0wL5ca6q+XqosxjnDhbUecS4B7PH2m31OMHSVh3ItBhQTGCP
+n3ISHTM7m/5yCTaoTopIUhCKZJXyhS9v+GsqFhOeBAKrJIOHMZKu4fjVYsXs9Xx
HnzydBWsHiP6X6+GgJFiEpUdpn8NVZnD59jrv9yjyO63RYPIvqsYxRjqw30dKyyW
j5gkd/q6fZhL9YslUtrQcswr8ACSI8e1Zui+cZGBZagvsqGtMSe8f1tzBRAA9BU1
T7uzwqFSAQIylltntg32fJBuxuKAxPQ5XO28yD70xSO8Rb8s6QiFB0AqNA0AFfhq
jYm/NoUMWh9dND12caI83RWAYlJuNUrvyMsZ1AqQR1rgU+tdCMxqrdxQC9Qyn24Q
l7k28dDSRlqv9C3k2ahgi3c/YaeApu4H+Dk/icuuXWqZbb8zoWMrez648qqkH+8r
5GVecnWvRIPFpLXGFXl8lz+/9aLrzgIiWQhHrOWCLKZFRVtJey1Tacop2iLb05yf
PpPGajrEVcq3jH46cc9a2CL7BjOxvG5ZWDyc9Rwkm8/MjOdBQ1YmwW6pA0bWSM5d
M/oNIlhTnrJuyiwqpdAReXTJdqUPB6kzuVG09utULUb9YFaUFqX53Rgk9fS9aR/R
MCCup0akwVJgZBduJgZEz9bb9JYf0vw7qI4oK4BQ1XC8k6vPQFzOWjYl6RzTX/SW
xml5fPnwgBFmXxOZpPQ731JYVptP7H590nx5H0Jaxr4JZ2mNLi4Fiv90tf/PTg5q
ezvAiC9f1FV0/6ld8E6ayUYJdtXoyifed0ZATHlldchkHSFJ/uZ/bwxY4AWgjLCZ
RF6sUyCPjWHwwpkELLGBo6FUKBR5+2jFWfBUnvhlEgDRzK+73bKw/GWm+I5Uiv1d
4jJttdA7Jw5emMyPpfhxEf42Sc1wGo0qciSQ9e1x0K7gPe2OgZ+x+rv8YRz0afag
aMZ1DCOnkJUtJxkwoJyHFbUCDfKna95wXcoqka6B/PtYsXHC3bf2947EHP8p++8p
nPUqy8WLI54boiK9sOj4hpayqBdFZT4YTzbnFjcL2dzoiD7Cbnn4gnoEgPdAolc0
E4nkcrL1abUCowXpblwiEIfHS815RnLwr9/JSfQiQhRbVmsnrfz3/4b82Xq0nbEA
9Svx5rsN3/wkD9gQ00b62636ZFAYlq5Mc2DGQQjwY7sYlXhf/FZWgl5BLdrN0MlR
HlEqJc2ZvsvamTWjWZb+vKpSS7/z4swTCJ8ID4NMkhYOgtheQ5DME5p8OJQqWbQZ
i1I8+uRPcTh4HWtqPkffUIIvl8IQvAJ45Smqha7R1iacU98R/4FWD+PDYEEwmQ0Z
8eICf6PZ6eBEzD5kpym1zRWRJ59TfdEApDQBnrStphv6+e78c2BKg093nAXUBVIS
bGw+xWDZkK1712BaRI0fsIN8Paad8rGmBcuVCmMiaM/vBPeUb8e+EbOsYQFLbU0x
tPNVJPNOxV/8ObC2P02rM9l/1HdZgWj/vilUs2v26lbUpP5VibgtH5l0yCPN+mQt
ku/BvgKaQ3yqIhNCRpHJG0eusT4Nj7HO5vMQdiXyaesFYeokPw9tlyn2Nn6Yx9FX
Yg+VXbbq0aFydnr7Iohvm6Oeck5WViDVmUc8a/Uing4/xXji9NXSY/8gaWuS9h9i
20z4lrvc0OVIgAH9zHXjIknpQBqetibZWArtOjiFHEDgSrtprT0OmD+nvLXdxfrs
K98IOHTXocZOrgNDFbjVAeYISLB8qoz/F7NhBNj4IulPz4hN9drjUEzWj4CoaP9h
Pef4ZutpWaV/h9IdgvDzknXwCMILp5UsnOIdyGL07YhHwgHrfG+w+GFEe8YCh4Vh
VFdExbLW2KUmTV3PolhTv7eYyevHPMZW6KMZDZEaKc+gL/rpYWo18tpNSgxlSV/9
zaO8j92KF3TThqBRlOoiEAEgm0EyFhowbiZInG64+TDv0t9wQSYtLa5QsI1yyPr8
Bxtxizyd8en+Sw60wD8m7KQ+zuOnqwO7FtStdxEyjX80b7vkVJtvqbCwDXQpgAI+
T7Ypo4CRY8CWzCCFqLfHIltCTZr5f2plrQwDKk1YzuMcuhiXN/IxaXCE9Oe8MDoo
XO8LhIyyTM34yvkQ4DSdwlmzhmCrw//qYGQ/mjqM17HTP8id/3onL8dIgLXHgG5t
mMATcHuCa6Fz+SogM28eGXMy6iZQB44Y00Ax5hAHFi1+yPN4fjxAUsY4jLJOnwEW
9scvDm8dJrcfR3dO9Emxccagikaae3hpxdgkC9ivuTjiDOxKowZ7Ju1p9KC+D0k7
FRsezqz3gt9vH6zCzwHv67fWTEhfer8PaDsUj83EApRyaHHujOUGr3X8rCKiCvN7
wA+3tbGDC2M7xCkCcINb8eeQFR6WEV4z8PQN91z+E01Wn+s4KO64qBSIBgbphC9R
D+cQJ/R29Sk8Lfp/yjyoDVnp0lhldrAXTU2QPmGZS2WVEiEpHtB1zvPJ8nt4Z9Z7
VOyaq8diN+1GZutW2h4+Mvl6AtmccU+5iBI7aGUJ8snoLsjW9J4GwOQ+xV8yYLOc
NwrYSQaLbX/hXI9XuUuKXGMmaEML5uesNiQ2s4u8G94BO3GHeuWnSf8glOEzal8W
ZGVbtKCEHtcegZfc0y9swne4wqqofqUPjmJhWztvdndrF8lsJ44q2jTNo9YpBZtM
VPwV+NgUCGn6dj15QG7Sp4F0owpBTmAd5w5WPUl0h92TPQ2PqDh2Zadz+lWs+WMN
tGVSbFDflVPW6xi38LCYkg0sXQuIKGCBg5BxRhZoBdeoIjol0fdMt80K00GNMx3O
7JZoK/5bLh/rC0BFAkZPwDwV+UlHpPov7AayN1nflUFVH4kCtzEkrwYn0vyAD0wy
vXxndEauVpFDhGnc1KuQFQ1HYvwUuzVXBhPgR6S7W0iOkHQUR0eX1oe70loKuQ5v
28Fx6GucjyzgA71vPk4IajlE2+X9BEcqXxk9I0nvfTi3fkV/evnmhjg69tTxTSV4
cvsfT8r4BM4PMfgR6omfqZy5D7mlA+tqmzcjmKGADOr68SOSWCBDcEymo/DQQ2wM
p7kjwJvVzUHx7CdY2RqdVUAHJyTgTr9SsBZ1vpXpQYhsYOe8rkwSEJ9785tVENfL
XIklYIr0ODBLhkZ3WDf34P/FYdpm8Kd3DW0PLaW3nKvlhe/XwyI1ZeAmhW6fC7Jq
24T5+wJxlEY+YKw5zBOrBPE99WKHWu6utXI9ccMjPBZzd+kvRWcPSiLFCHq1flGO
FY8Fy9BG3imR5d/aU20gXvlf/VzmGESBjFukVxQWXk/P2S17wono/5lb8/6PtMq+
cO/Mn0wTgsas7CpVbgz9IHd1kFjeDUx6sz+lj1UkYAb7YePSTd2/CkcMKfejtKHA
iMcG+rKDUKMIbDVzhcxH8+dDzfNHrUunYwbPkLr3lKA4ho5JBjziyTBTTQ1MO20x
QA3F3tLNft4jofReDuIpw7CrO3JTZ8kqk6KiT1bmhnt2S3d47sRPBLPE6LSMk7MQ
uJyCxExZy8PC6/JeXlN7NrG6betfdP4KSnOUIj44GZ5kPTBFXmVh+IX94YQCWRCh
JqX4rd6xpuiyQwxFCuJQ9jJN/LOy+wfeK9AMyOdpd5JxON2np4SlxC8b8K7PUqDK
5LW+/OQVCwAkrX+KT/ufiLX3s9OWUM+89DxZkhhEEunaEANuNBbl/UYv07Phj3mY
V65TCwyaK/f7jA59814969bnQcNlWh5SyrLe0NdfBIQIcOtFvLc8Wt19Dhzw5iZQ
chZ1MeQwksP0lSdEbjVCNQFIZBSvvdMwPnJVAW3PCVaZJj20Ux5h4inu06vjbYk3
qAlxf3VsN3DtR6gsTMbrhaN0wJ3WRnvNbpLK0CLOBhR0VOKfLy1uEBwV2qyXaW1L
rnKXkQfoPjfOVGCdsYB0uoA6lDNOjVZuiy+4A/aY+BBumLtc+WqLysdOFy5cBm2i
7ay3Z/N6Ju7jYs69wMXBDaSUcvMZd0k2XkhUOt0wC0aPAvbIsWICS73ATLtTnn1q
Ic9tu4C9Wf6DxUj0bCMnsVKvDWfdtrbm8nM7eHacjYpG18cSzA+qZxsPmcYZ7y+r
`protect END_PROTECTED