-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ke3kBgVCpk4oGPO/PAnDnfSp+NS5Q0Gv4ZgS56+7Wgbh1YY1IqL7uP76gc9IFTdA
rgmOrgPzrbcmVxfQAK68tSwq1G4pTycR6KRI82wS/OlnumrZJjy9x2/oOvi0bCIc
wy6ELNOuaqJwo8qYVplUx77CLyk+ZqqReOXNsmKznvLC43xuGZ3oFA==
--pragma protect end_key_block
--pragma protect digest_block
1x9qeo4QwsTPxgy9U2vsIK7jzGI=
--pragma protect end_digest_block
--pragma protect data_block
i4l38M1syJoIPESCHi4wijbnUe8SXGlPj9+vEeQtB46yUJb8CKHtbmKsXv+rLGCX
v0rmDycqssbi48vpykURwV4dXVmmHWPl+MDid+A1k+cN6OEMXZfdWNBLBjIP/S/c
leEmhHt8IxvTYUwySVwMw8ZCHJRvULh4aQWBI7oN2U1gfXgjpp607LrSyBKUrrAK
W4XN3oeHla7qV4Q+tZFzB00pyjYovL1NqZyNxwwm4MEsv4nJZmtiL0iHaMuk9OnV
EKg+Q8zX+XnrOxn4KTzqssbM/VAST3V8zkuCrj2g/Ckp39wiydUSsW8Wf5z6ZAZg
UhQ8Klhd4rknr7TPF+dfhzvA2jox27wQBOz+B+pej94oucEQDNLB/KlXQcnQ0C76
FDAW3247ngzAQ9NZahhazyen5R5YNPgSRmAc47BwbnXVcldoS88Tk87+yMWxFIkg
XaD/jlxNBeaxxZm/7IDZZUb3DfDw/eTOJdqxA2hHJ/36TpC5LRB6v/5CrZBRE41H
OyFf2+gFGXlCpfkk4Xd0dW5/4OgP0zmGmeM7zdvJrrlPxfBm8EtzqkVAsky9+ZGH
HeK0iOJgg8weCISR4CeA/Lx5yfBIbYBeJKuuohdkua/DkiduaXkN1Sn+y13eWO/z
K0HbsatUx+JDMtLZOBxIIZ5JaEdqLrTh4HvrxfJkY32THpiI0MHZA4XgWPR5PZ8e
PQQVam59Rv87TjPD136VLxcyAvxqsLZ/YGGYjKjsKy1TyUL4FZFJDRawtZ1eCfFZ
nLM8nXWwOeHzGJDFfusKSDk8Ty2IAvrH6hrNL5rkd3ROWoL0XYzi7J6UCH1EJhef
Ul2k6+XjYQ91cFoJwEjVLZCUScjiurVmH7Dd7KKShAXFUG3yHEWcDGeP+R5AYQhz
wUCN3Y0FYR8NXFO7V9sCPGcfLCUG+Q26VJO5YfEh7mCyfGw07irkPxJZsr08Nuul
vKga9BPaVuNuJw8uMt+CWxxarKmc+8NFK0G2bvi8CGbudyNYPbevKNDduRRPDgfU
otex3uU8d9FMYPD3YOGTKGVJRlQHzXSbBYC7rORk/j2xmvxKGmDscfFprNBezOT3
2MzUwqCSzQamM/nSsXjWlg4q2C4VHNwmiz7uhpXu2MUIdvWkSV+lSGI90edjDixH
JT7rtP5gJJGRbxePtvV53Hw8NNSUXxPJdg0+sEB7kSBVm2I39xhatvKgPms6X/8z
DZLcb//e+pCVBRvUslGwkjzaScWu7lGT2jZn+4IZB8AVb2z/Qv5GxGCjIlIGdoZF
dZyq9UQtt0mvL3qI3IyLvgksVFHFqk4SRHT/BKyvceCczKoPEF/LftG4XcrnOyKD
LAigK+zMBR1EGc9VDbtYHooGPYU+YG1B4NhMfM0VH/SdVLH/NjACGZo/bq7dmqDr
QiYlJSDSo5wbeDe7Dsoc4aD9qQ78zRr6/5W/OU7QkaZlZnO0HoxmU35ymixJ3LLw
ogrNTwIrTj1+H5xf8YqPpsFU4laHnhR70KoprU5YVLvU5OJkHQAAXF/o9jLhn7wT
+VxF3ikTIaVPFnCD7IZw/bdYRbJ9Rn42RZAqF9orJQsp+dPlyCTGhw2o5ZCSQGRn
cLd80FDIPJtzgsKGb7S3OZ2K5nZhhQjONm5zXWO7Zx3Zh1bglwJbc15/b2BguEuo
n11MNvlbRUdjObG6+O2umHbjqSjSfGYsiZLgn6fevu9P70Hd3nUj2GFogU6sMunH
8WOJvUHVg66M5V+yE9DpKf0W+XTROhblk7jAHWMV0q0+F2R3xTl0UdUbyTNF6pMP
rOFg2BKqHV2xjA7mCcxUGgH/d7H8DlLPiIJlCfXl4WeZ24e/BpUrysxC+jwHegdH
UXLq7VoqsQ2nbuJyzowtZJ0LWGB6p4V4tjgH9OZpm1TiQvXsVrVqPFptYoOR+azW
AqC2f+KUwV+KHpnogTpwpCTDgdj4x9ov5vKYN5rZ88ZcMnGMRWC01msTp750SwJk
DU5mzc9h/8GDwx+IaU8HSeVMzzmJO7WPDXW8Y/BkBY8Dvcf+w49UCm1SpsPTuUrX
AJeGI1ocj+b9FXAYSRLYv/uiy1N9uILylkuA6MD8UsjOhEMhxi/umM/9o3L/zDSf
vvxi+e2AZKzI/G5G3e6G9q/uhyFmrAuK+dC5q05DUtnALajAn2FdfwVvOylxcajR
P7q/XcaIitc9VMvchwPVENElPFqfH6GziA+HFzAI0HwploLkFCKxMKARxWg5zhOc
nK+GyQCJlrMXCZ/Nt5cwTonJsz3bYgyZioPddfUjMq7EPDyCu1uebyZm7mdWz5ZL
zuCD8/s58NdiAufNTTuVFAkNEh0Ki2YDvHJNwR3/o74l9ShWeAnUI1V0TcQcAMjV
5I0p9pBXUaEffwbGtwXloG6PE4QyKJiei+nmj72LN5hAl9fl2CteJeXG/1nVs47e
1KTf4keqwgtAR5QyDWf4W3tIXEaKeoq0rZvqNaJQbCPFGuIoVUHSbOeoe1Kw91e0
LWFFrSnnNIvU3BuYHVDR8OaqKOSFIYgEQY1VMhRFzvJuTIFiAXCndU+se2wVeZBS
9kKUya9qJM8YD6gzxtnv/nq5E53GkezBIUXtGrzYeNNQc/NHspmyD8Q0/MuKoGAK
t1PdBcIC/IsM65netXIkFmhRElYPAUWDhSQ98DUZgnWxAiPQ8Vul2SEAiPBRbbIg
snUDCTYQgWw9YTaoFXT/Zp+yZYPbQpfSAunzZAxnwPMLxxKEctdgDTRcWVu0odYP
pEKXFYQhyhzXL3sO57yIYryWtn8WXHw9cMfXnph0+3ir3qJyH6AyWN5z415WoQsQ
EX3QtAlR1wfnm85etOcKGxbjmX5ZwiWB9IP2v/jG4XwhLaxJ2CP7CBJ1zSbS+yKH
LPgw45xstEj0C6Ua+QZKEd9LEELhuNiFajBunTJdYKHH2HXwbG6K9tcqR0eFL+kz
XyPZnrOOrWXmuMbAmfD0TntlCajKP+sejiDnoiLGJsrI/xtIbdx6c/TAhe1Fno4u
K1Rd0IYxPLuTGBSKQcZilomyraRU85N5dQgcgAnc3Ncailfo2WJczIBQA0mQoWO4
xaSc3Wt5jC27nvPn+7eZZ8vVyKJY4UMDCu+M7lBQYMc5U71UXpkImUlal15mJOKN
Dc7fqQTV2qFbdl8o1LfxbK2+HcW+CmrojNPErQxlhc+Nw045hsClgR7QmApmzevT
WjxowKmYuAtQqUUnAjBHKd7SzQztF168IvLUaI4xHO2rtNWmbjliVP0y/vR57+4v
9bSxCHXR9pS0aS0BB/65Pxqgyou9NRP4r5C+NQqM6nwRPEN9c3tFj+9TyOESgtoW
QvNTXHIJoYmEgbJysnIWn2OkCKzItA3mNxAayBELy27WHQb5HXWf/FqL0BcOnm57
WHLWUWmr4iC6D1486n/p8SEl+1jx2ThfAf9Di9B5oLDNC+kkUdV06wj0SR1uIBCL
hYvw3uEn68OjsOmrPtVsO9NrA6cFrjXopV+jM0mDxFA1AxqW3EbvHe2SopKFY/AQ
ci0Uu6lae1YQcUvZo0nQ8xB4Zu/mIdWgEknWaySfVxOTSuGuWlPS/ztGDK2bcFOr
Sg+/PbndD+3ClkAYjteJEZsaOzaX63t9u9ZReKiHKMPXUIJJcrcNkutDQVopg05j
lWfVlOsnRpekeqLhAkKijfKCoaHqqTckg3wqZjiiJHGGfSCgOQwPwOI/qV90iZlj
PcUNtOgwCVQhYzYvP39q/+uaL6zKa+VJ6E3yxFdb7QG+DY4cbUCoO/67sfVA/1fy
s3Wy1irOKkFQwalGwSj7FSwkKgqDFMX3NzIILr/UmfMrFotE55MWhus2dFEp8YdW
BnnrcBdWchO5JdPPa3nN4Z3ixKPQ/7x8Ec9kPAySBpzcfa76tSDqsmHAbqOOFiZ0
WxMUveDnDBq8oYYBVPimyBvEMLy3RqfOsU3Nf8cfSVQBJpsP1OvH+l3i7/WRGPj6
q66csitAdXVCrvzydqG4SXSbhdpe/DTMnREbUfzTmfgv1ALicBPIqtsKqfyzbptj
3laCnx/ve3h+sZ8XBNy/2pnRBcJVfdbg2tIn7389r30heyIauWYERcAPsX9vP6Gz
Zg9p8XVKlhA6RRrApoLitNE3xoYyt1cwueS5BWBhahTjr8Y/OzvYuAoEgjNHjGfc
sSEvZTBbmXguqXEN193lwdFbhYHeRgCfVKYGYNpT/oshLm25KN4+hOsTW+AHeVm0
HPrt/rh1DbyJMrrvu+G/w5Q/D7y8974gUqS5y2qSBXRE0kDvFRCmg1VOZodl8y3T
Q6COcwfGtCWcTimVXG2yVVBjk3Nw+0ZcIKmAkJi3ELXHZ7uo+QpkNslftQtIH0dd
jvq8IL8icvUjdIQ7jsx6xqGrGNMhRq2Vlvjo/ni14X+7UgO3UR7h27Pd6HI8g1Pl
Lo7zqyiTyUSlEJmoEOkd/3JJclWnqzL6Yr/aW6tjQIVwOS5qg2jqenTm8omvPtSl
/tGH/NFPc05YMxplAU+R1VMEUVOe2xV3JN4eZ4NWONauHP3oqqwNjsxFY0mjwDB5
f6FuvH9bDF+nwkk5j2BjRMGC0mfXZCfMrfvPMm0QiPppHeubBIn/KwMvCrgMFNCq
R9TCKWG8WAkrWSOzBjpBDfNTR0S2kFQvGbOUeNb7IRRKIkjEJCP32YIM1EleASup
xJDaedkx7Xa0EPsAL/UUD3eigCkdZ2kU0fxRGVEd5ALkg/yBTimOcMWQqv8ZqE/o
Re58yiOPNXvnwDyf83+eLDwqeutlADWj6tpxpbz5XB8I2GGtOnPhHiX0PHBO1ZjU
uPe2iMa3xwXtyl0lGN4sobbxmUAOGhm7+wdCPUaEajUe3WHTWhvGXQbX+BIJXoNL
Z3IRCDy+QFNNcUqVsLNaFXkEoYbr9MyD2nNbIw50A8LAB/0LlT8DQgHIhGgXcl1G
YTs6ZbDWYo9A6X6ZO9yu8g9LY0QV9G/sYhtGeATZuazRLUlrTXjQw8KKrefiX5lF
YJJ9yLAVdg4mh4S6mUdnWYcQfW6zUwLgq2NVAc/Un8EwbPIWi9JAeibh4MRFCYAZ
oizQV3rGwrR4h0INRdSIwpYK67i1OR6N4VTEXs4Dc3CEdAHwqn5tHmgkQf6a5MSQ
qoZ+Gi5Do6kkK+OvgPT0xjRTzFGk2N4KpOX/0NezC6Cy/IWSyz1XnFwevxU7YPEJ
ITkC4O2ulxTfAUZ3c3+iBtvKImn/NoIz8swsrHbHF7/pqL0Q2fFJGYt4Mf4cn4OL
cCOvCoULD+XzPIJNsmVhLEKk0TZ1wrg+ZC9eIsaQvGe4Szi9gOPAzy/JPs2rQxwl
7A/Ivv2XBtQaMavMvLyF4mj74MLKkQKbmwl3BYKVWg1IwrLNi4kPXUPkSiWgcSfN
1lU52YK6/OcDJHoz1iX/f7r6ypRQ4m9USKltCwr9KRJIs2Xa1aqYO4S7b8MsJZB0
cWArNgdvGpg8N/Gn7z5/SD/xF+YKfCJpNkc+K3mQk48Ph1FYW+toAmFpPZBVajgB
JfPls83IVGpMU7FTiR7Lr2dkJFNEvFCjYTZgYlnN4xm/e6Gt5F73bGtoj0bF55kO
KEYSskWbSqf6oTfE6pHDleYaqdjIjMCYt+q1BMD60MRkgQL1n011Q5h14XuJiuYS
LJuqB2ZT/6rdqmuZX/2GiNNrd/jUJAC5nMcFAWZgsfkV7ZKcPjPoH0sNikTnycFk
iMnnzPOzUToQ09Eb9H9SvSDb6MLjfZNyPSG7+MQgu5IQR6VB9PVit2nDCgNWf8X3
00x6kT/0yu5OjK6ZeL/v3g==
--pragma protect end_data_block
--pragma protect digest_block
TqNNFsrGw/Rx0tdIAuZTjHq09/8=
--pragma protect end_digest_block
--pragma protect end_protected
