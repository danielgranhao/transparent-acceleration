-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
k2Q48IG8gmtdIxM5rcHV65NKa2PQSOKKZkr9W3BJ2AHh5C8tkETrxgtl+OC4tojg
eQ9igy/9zOwr5cbzBS/A/05+9LMdy99RT9uM58fCKcmUq5bACdC5JWpoeS/grff0
VVAuo7vrJnV1fs4N8eR+08dI+DDkmVHKeWzgApMmfsE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13600)
`protect data_block
rxcxE58WILqlul/oaIXew/MaikufI+KXn77SOG5qhyVqQnwEzR7B6xMwBhDX2TIN
t9m40wPuCJ0g32WJqVhLDiXoCjIj6cFhTK6GSMDULjX7Phr++qf70fgzEB2PDBwo
dsXAVmF1T23vfJdA2QW95Fnlra0PN8tl4CBub4DqkafGyQuUHPUeBDdcZYnqGDDM
WMYKeX1rSzqYAMrARyvsALCvlAYrPmWBdI97laNk0Nc0kk0/TyURW1hrq1W/zGZt
l4jdZUfcvRRG5Aw9RM1rX8psM+I5dz03Za3cWReRG2COUQTo9QqmAUk1/YqeFT4n
kLumA8WODVLhExHOAeIW32mRRCfBni8zRSSNqkUJN/A3x1KDsze0uKkrIOY8e0ps
ZNSmnTmMkPr8vC6R7sGC0PXcJF7F8+BRLSbSLOpPjANZuB8eTXwrAwmqTAFULpFt
wOjx6ih2hK9UfMlQjL/a0Y8LSio+WxsLNJGn4dnvNfAV51hst/soYR3fYTqZNph3
skH2AjVATa79MHsegzyYQo4VbjILODBxq1AeqpGf54EuHrMC9ibhzj+XcUXH+00j
cvd0t8lSeAymQbNlM5XAVSOYakbGXKhhmfN19rfJpE2Fs7gOhelluHdg9rzoQn1r
JVSOj/fo1uPC7qI7+ctoVxQuhu87kgqYVyXZ99+6uK2l2m6Ql028D/O1k4xgtbch
55FQZkRuF9q7rOZgb4Il9asxiWEEMC4QJjsdh/a9zd9/OShI6pfblQm1J+5qJv+s
5F3ycqXVkVRIpbGeWWRP/C+b3B+QzI2vV/PklwJTNa5fkCdCaIjrWZuUCRvcgvoA
awoCU3Tu2XeGwc7PVqBfOb0GqWxnst+WPgDqzdY9x0Dn6I/ntukWt1to4GU9T3jk
9/bXjjyFmmqjbw91uapzZ5PEn3yU7o6C7GyzGrK9DoHoJ4hg4m0Rv73zeydk/pk5
VI3F4nBTJLcKq19uVBj+dSrPe9AiKUlaMGayc5nC7S5FjH+Iuzwk6Cs45PL7M2BG
c7F5oX1r6DCOiu1UiLWFVn6tKaj/ulthMYbRWqCwMpwwREJkqEWJsuQ61+UFzl5b
WbxAuXsGwkfKD1el56BHevwEs8lAUvRGWUVMibAA5CKguHiCt0hd/+Ajv+uvVyvp
HfgoJVUCvFpxQ4gKKpr3pYK3HPfoNpSsu3VvjKjXzYWWA1gBGYRBn203yXXckFtV
WoLJ+Uj2VGJO6DBYT1/pIsNV4y0Up2t8u9oQV9r8W5zhZlnSh3+37ww0ujBAdWnv
iDhythKioFPtfdnM5tNsVq0jX51j66+4dsN5vWaqq+yGXBGpYyr0CqlkTrc4Njfj
ohfAudsU1bBjelqipxdOoz1s6wk2xLbCwbnQaK/tilp2Z6nCvDhA8KZIX+KN+Yp2
HgJcqV5kmn1SC74VnsEscz0dc3toEJrxli14IXFib1gWijXwgvl8Nrqaq+X0rnm1
WxkncmUsSdaygephXL2Kjwl/6i2sCRB8LqrS7yRtxs+q6wNOrgR4ZwyIgttrmhnt
mzF3C9zRgfaOto/TLpZxEJ3vIObCv9+fum3+gILFGwW0Q6jy+QyzPylfu+oxKrR6
zzsW1r8s2i+pJaE9wpWsfClM4xyIlhaxh/TE5IRCmfFLHpsRKPjrXiTQcX/IeeMf
LKpdiAzY1RrukLHqCNlhiqwbf1xFwExOsHblu9frQ8lWnj+FdFq2U29zVHT5Pu/s
5v9o263O+zhFKNBzLucBvxvfIYyn4qfaG/dt32pwrU/rzhqPdQ5/3eUthNGd9wG4
dUjKvruC6fl07+SzjCxFuKYcYi8WLRwkybLejRBx9ifLLYTvyytS49jivV884Z/x
z35E9oQrsCidU4EczswZvDkgOOWsqVXVWQ+Xe06KXugGvagAxTvNoruMFa1xZFg0
+8vZmpMt33jnY+NTO/UE/J29puiuCShwhbb2hmutxaUjyFO+GUYtl9iZI1MgWapS
Mdp9FH4siavHbTkbcdtyjmZYQNbCc3sYcCbKP4+yWTj/t2hUt5aL+xL0t7gkxrrP
1telcR9z0j+DrFO/KQTTgLdpblogQEomphHvV9m/bWq1xawJP/X7MqA/7UHOOVoa
GJYJaDB+G6bj1tJzaNF7BsuV9dnDstRH3DTS1xCKG19Zzu1c5jcx/NXbJxLcRIDe
TBd1vzuPq4f3dCbi+lCDdd4Bd8Wo8qUiorb7huXuPxDoL0mYBpCZg4QxRHDzgf7o
hX6MMpioPm2kDZFk4SOAPUloRiJN5fJuxT+DXJCjp2vuX29X/hkhWcxlIeDMoQLw
7oSZp4a7w7c1LRex0YwCRPDsM6rf4KGo0DEIIKujpypjZ44LIezjVM79Oinl3I93
etnaLu2wepXWl6E1kBN+RNgfnpr1NkyOy7q2J9ANrQxdLhtEcu/30SZgr9vXDPuf
opNJeKXJsH8SkiguzLiriNxSmDzhAHqSGcdvBttYlkDQPZLrqa/RSes96OPHpgXl
5deqyUw7VQIxH3+hsXLI1SOHuTwPFrIYO4s+3x++ShpH4bnCTNKIaACvRAzKtUYq
YrV2yH5P1GNRQkZg/jUnRuKBAJoNR68qxY3bm0R1rXmVbHvii/8RjDH+Z1kHt0Sf
ad6pgjXB6h3IAYl1yhhWGiucsFIvqUvYk/8BlE4SLXhsbyDjT6npFpZf2TlzFdq/
7CcDBT3tAXLtzANLxNYID8g6WoAn4oIoHd7PLSPwSeed8GoZ/20RDALP2jwwuiOC
nn0od8AJaEP+PFNY2+hBUWtpRCJSO0de9UGPkNz5DyBLl9ZYxde3Hur01ctxtP7/
PJt9TpmB/doHCxiZK/jeIqf1ePy/CaKW8ZQH9ZEWGUqpVwq4Sj2JY9lal47/8rRI
0nIVzDl1+EpCQm2UKBr3U/nNJHK5BvPyoT6f0duBYh6piQuhYa+B0Mk9p1GM5hMW
uEBC/zy8if/9t2s3dYE6FH8KrPY3QXz3b7zw9WQT2QW+GOIcwOH9oniCddolksGz
BnrawJVirxuBaR3Kp4JiJTvZV778Qnmvg582OvT6nNXd1z5CGIZ3defzxaHFcFUz
ysXvt63AbbXeaZ261+1NdbausF8gv0x12x/64x4S/SvzEE8M/DjzbbY+cUXE9xHU
rAbTJHCv/OeBcvoZmUji2UD0fUziSaO0iTXvk5nCU+CRgqWaG7QOiY2IldixT3Vw
cnYV/IVoVqQYdq8cvchyWwJwSp8lwxVM2Vgc/KDHIUpMmqlW9kr9g36+0+3da3yT
R0pH0J+z21PVk6eBXW62J7E7kzUlBDfmiCRRlxOLQLA6uzY6/k/D8sijJuHnhcCh
jy74EGNqTB9xBGin/qSTb4EACrC0SmQYnZQ/stw8soshuOdvbn6PcSE3e3AY8Ljk
2k5c4GehhGCOruO108jl/o/+UXfyGQ0ZhidJRsCbhUiw+yzP3EolUxv6ulRm1Y/+
pWSgulRZDzBZXrWMWzTpCVakevJz1OFFM0VnAUDKuvrz3HnAYSQK6FWbCIh1Iseo
Vsj3q+/o81MweIo6wmw7FhzVn5ru/uuDEeUTxYbEFDafB3kbI9BZ3MWF2rAujQ2P
AP2M77CDidYuAO4umbcV4dyvCdCvqY5LtcKD908epzxSnlPS8RR3IGZz0D9SEX15
weYICgxpeX3DwRZNm1DoCPNDeIzc6zz1cgOmIq7J0DEZq2wUIjU8eARy/rHyQG3U
9Lu99IpndAjTGkEajjpGiHhrsBb/NwSTd4QcVjlAolY1PY2vKAGvGUhezpKuJnHd
Uki7roTUa97MHZhsLX1pD1gyUmB0UHls6Emavd4fYN5FjzBgnLI6MzzRVF9nXQAc
JbqlS/1kYHVNki07NCps1r3V9tEEKWJ/4+mct6GYjBqsBETCxLs0BBlob0cdbCUC
TrsfsJ4sf+4CLlVa72EMA+dUhNT1NoDO/RzOxVCTdb9N39h3qSy/IDi9ieXhITHW
NvepIQHtLv3rl1kRZemteWeNDrRit/s80uHjQn9QkdXxmZmcxCxjmOoLClRy0AXC
aUC3lJQD8fiW1H5QcGXEF6uf62ec19HADzKnXdtRCTj2VqsveJPGuwkvxTs8tlsv
xa3jdkZh55jfMbeYgwigyrt0PrRgi+wi0oceGQq7jXYRiVGs4KKx3UgqGkgvNLId
rOKkPWQcTTmDI5cWw2CmRGzId4AKgPBxXLVkZBecBG32+pwi29n8lyMx14U0qn0k
aijnzyeknbfJcxwWoCWhN64P+jvtcTGM64dS81wu7syYTlDrH3Pn3P9m7fyvikas
qZR5EZH0kdifsMbc1rCqWw/vbHzpwGH9Ckvpd0ly/K9/odSNkhFTauaFM5VKM+QW
RwxBXMuZUCtVTF1mYWu4f++tZJ5IH2zjqS6wEYS6DIdIDzQc5m94FpTp+Mr2mj+Q
342oSaYMFgx+fnkhWtPWL1KJwCODrd+ky1suj/2iPEEWPBEfADCGBuepCsvEHcuk
VrYM3VdQjb/dDgR0dGj7c9bhnKSUo2XWH7j+3JVjwCQSpSX8WtZYfCwIJDmlZ0jh
uufUJNd9BqBhXzqgE8O4Dx6F0GCXNnUpoq7/4s8dbhGdpxRq2YZVWaixJoZb2ZJX
5qQMYd8ws8YkcpabjQq17ck13AxWML0VENT3pvxX6VYFXF9R5JuMRIQIWAEvM4BJ
vSDwSbxVH09i4R3AoJ20ivtFKKIknOAskJrJIZ/yB7j5Li6bqqA77PNGdtXmvVyM
IwvbWbJQ0j3p27UprVPM9Uh7XPm4Lo5VE52Vloe4wh3/Q3aWXJWUBvyHweo4ka6R
3asQNpYEniNNZDj52Tcj2exGTi/5gtXtaFCbrlrzPkkVYf9xc2/wZ/a4ht75DP8b
Dz5QMrEUyLSSv82Pl4EFFIpTK6KM1QSKpkwvLY1IfYaTzhy5hMUSYFMG4SCXCcYn
wNuaJC3NbdI81Y7NkvQmWuyZIoDwEsnaaU8O87HXgXjrXAqfuKljmXERRxVi6Wu/
okNonrJGK7vLvX9FSWf3LUuMDfU/a11XxXN7awp+UJJD+RW4vZnyU8hyZH3irXka
lFhpl7iiKwzhi3or2jYgQouY+DfTeK+C4l2PdxPi/hdt2yMFf3s3tdPaIPuy5DdU
F53t2Sh601HGcrswjYwejfnIsRz/Z3sr5iiQBGymhRT7aJQU64/RnZNMmO1OkasK
UzIlmvL73/Kt+pnslTgcFqqLDsaalMSqJwFbyUfFfLUtIWd1kiOyHUZ5+Bzux493
pOhzSaDcbZPk4bLe8zK93QTPSt6v/vuHViHqFFdq4Kdguh8gQkCwj42a+Lms5lni
4FCRZ4q43aLcA2fU0TGQE7ErPVVpfogzJWldp0T0rwATQ8hFWu4B6aARxIZAgxGn
JIqW9ZZ7+DK+Wc1dqAtCEJnO5NJuSzVGbteiQZeuxt/ZL+JqpgOQi19StvUKK481
RQZZKBppsfqykIfjZi68eT76io4hhytadU3/FkHp8Fpaf1M9qZlhvihAK4fXtNYP
eDFt5t3ThcvaKeTRvxEfs3rl6MmtiAiZNjXoFTLQ1zzRX343lylPv8Cous6GooTz
DilzRTHodog6EZ94CYgqvKGQXGPRSsSHxG/eocIglfopA57ThBJDHSqtstnxaiNx
iOSOL5vOjS3clktj2OdTSmHSIHEbeLa5XejW4mSerxkwZODpub4Jzay1QcWArP8x
favkGZ/6oW8sDvTsbAO8wI0T9vm52zrmbC3H84StqryiU47I8lOtmBAYU+oaLEkQ
fiSCdBuoRWM6ViLqLMyWS6eigrBY/NLxeZ2CzShxPSBWSXp5yX8Bdk+qdrB79+gq
OByoQDKS2PscIYVuv+65eqAaJuWOPW38hBn9+vup19NobZ3RXPy2z6V8ajy61NEU
GV1uwdoyw7wze22BJN5mYpOIIIZfoXSrEetkvrTSuSAlcVS0Xi+udiMBgE0+qENE
i6x8yV266LAAGL4cGDOBIC5O9FS9VKyR1/2Xh9fkEgBw42IYqvzDAWsd4fOtgTFp
ZZGj8sncGNz/CHPp5Dc4QZAw7HNKKlbEzRjUIi9UHmptsI3SOotph30V4KzIjRBr
ry6c5gclusBROoB5HT+feu/NcJsGOi3k8iiUEUy/AARboYd1mHP16fDwZD0GqnZ1
ycGnRf3KPjLDVl51ehuXhrSDw8Adl3t3qKwyqZL0reRj69W8Re7kDdIZmoJoMwcg
WpeDWJkDIyqEt8BY2VbyxgMqH+W93HD19Dgvqc0dxjaaVHQbXCBNoK8fyEutCNwl
6APUfHITkipEYRpzbRPc7M8hariJp2ozpgVrodUgZnSr6ambi367KLpfbO/cKBVI
xOMSzNd/A+y1/imgtW2zQBeQ/SQmvk0Tf7H+TfRdeymIztcAJpB2dt5auBXmpcYT
vIrVIMNDquNYSTbsQuSaTt4iI3YHmpj+i9USyKavVdG4F1msdfe4dd4cq0Um0c8X
fhEOPDgJaVN2UKJ4I2BaOKXgTSApcgO7OWx97pCaOTfCGUqiYc2Ob8QBpXUdRG+x
8+twSIv5W6h1nM2hMrocb26tc0k46nh4ZrHJPw9HkFp+somQinB04YOzrKhkOvkS
gLxqGqkmHs75heTm78vUX3QJv+yfj3ToQNVHADrzSAsndZlhCQHEc8e1TfQ+qD//
/MBfYwWOq2l0UeT95bptO8ZgOhkr4JijiSQgVGSYEyNV5/3cx+qUq1AkD9aG3WNM
Se9/4DqWMSLDNUs06g4up2MfHD46a2hjcfDoYjcJZFSCY8AxUOT5T0LUpZ5kX5R+
JoxEhZ/oPsjzddmgsbwJW291KzgI1AO3lZZ5IkLptLZV0Gzfo/s/6wjOGmgEcNqo
/lMBEq9K7p0Cz63Gc6stPOTiWkVdpaM+X9JvbejaIacevJ51Qqx4BUT+dJo0a22g
beAbtuviEmGqTwg40MB6T2h82qpUeGXC3EMuvWrf4JwUA8flt/6gWP3c3VJxJG7p
jUq5xoAWns8lqbpIpGNk298HBODPLk5/gs8ECIcYRO8GnwS7x6rAr1PZ/ymLsoCH
1DJ/E8mms9wkt1XRr3KI96KiSvzs/aHAtGXXyNV8Ih7kOhen9rnTgZjIGXWgJjzQ
9AdXmtTEP1Jc9O1pKnZ0dUSiTbAoNdHK3YHwzyoBPRtARcS3G2TCUw3dKjjdNuHn
ZCjBeAsvaTef76vl4rWVIvRATqAKyQDNko1rABdq9CdIwJ6QNN7sfBwG7/CQkDIu
3uaCvCYsG8OX+1+6n9mpMfAiIg1VFrewn9pS+bFKteo2amX6FfPAN8bP5LwQw7Mr
dvB0DzgqpfMWYKD9p4jOYFAB2HvYSf0bZtjcV/sBYJ1I9ni7H+5HejSTw68z7eij
NI4hl41+q0UcvJSC2cbnqKAtiJtdPUtVeF722eqxBkHtf7oYqtge8xJmIGEVxyaN
oGW6+wOcywNg3jLKJTqANCPte2GE+T7SThmidrVErHx9cT/iaT0/0pNjhWm6yMXO
fYfEnJ2Fxr3JZ4PovorIJCRaIrO0qV7Lb9w54aQelUYCCX5elNAuHKpN+d+MK3Lu
RcAduoSGNa9AO9R4SgA0I2a9LHYCyjFNbF1Y0I5NFnNREaP65Kwfnsbo/CVTKsBg
bSA/8UiVh4NzvW+UBm+7896bqD6qc4JtY5ctUhXJYQuGJnDRItCEROMGItx9GKM4
JGjGQ3ojvDpjK/nHr6Yzx5D8ZlmheDixy6eAK+VnwA++aw4b33csS5ZohRsIm8Z/
I+1Uf/WEWImOx+9DUnU0OxbO+pwGXU/eJumFjSjiCoHgTu0v5yX0yqsWnqfuxh+C
on6EMjjaHkZwTRlxPyq2TX/HdEpfr3p/CjDV2FKhtpv325gClmI0gks2sc+j81VQ
6gMdzswysKuLvkzCE/L1P/yHFiApbyqQ0mws976kTN7tWXOiNqTaylPovT+ODkN0
PSFe4ATv1QyNJbV2AN7UnStGbXPQOv/YT7LwfFMcJ+MHp9QmkM6BSVuw/wQw5nrq
Fu0D8EvamZsjh2hMKo2bIaz0Bl2qmRF4zj5SL44pcWgPBBwnoSEwSIyCIlkg0CLv
WCgL/007XZy0bfGoZ/sgGmbkRFViwfy6XD9rq0IFJFyykZpi+hEyRRf3LX8N430P
NfT4r77uFKFj2CcBrfwghcNfNcCLk9M0wF3lm7OpiUbqPdh7lQlOk2XTArXrIcvY
Kt2vLV4p3jyFxVyiQiGPVYTNJkRGTngPYqwZs50fD0Vwq0Z8mE75TG1sxKi1N3Ba
byWFdimdmfTMZhEwc5cukDZa6EzL5FtmURNRQ/d8AyyJtW/jLOJi1wnblYQ/haSl
shHOmlMVo1r+kVrFhO0xo4cSbsgYt4KqzSurgnDgBnTIp1gDP9mY5qz/HW4clLX+
9d1TUg1aqbFWv1BeuWd8MpVC69VvZuHks5c1nxqyBl0v6tc5sNiDzN1noaEnXOrV
RaO76QRqeXOfb5nVloBGSPjL2r0UUoVg8LBrYajyU7pNtBlnw3eE/Vn7b3BvbBiI
oxMlnSJgy8u4VwEJApJ7oYA2ALsWagcnvc1SukP2ZnRxUFSO/T1W+aEapMbXFzPp
CMhjELreC9nx43TcaH11MxWWa7X8JlGJ9a/8WNmVXViG6n6Ow6Qka73Tqfy4zalq
RGxJpB9RzmDBjmL2sNXWj+pGRc4lO06r4p+4AUlxQTRMSoy8sg+lF9NA1EI4+vQG
zeV5p04snyXiJYyz7nw4kR9AZiLxJC/owYwLyVsvX8iAKyMS+F/HDJGEDTKro7QX
XWE5uquMXvrUyL03w0Sb+mh42w2ItHlNUEZ3DWHckGwDeO7igFi9Wol6Yv8yjYvi
CWmXOgU8ZDZybTjF1hxHKEXxnADLu2i9i4tWsmcsRxL0hkgs18m/13gfg9fgLoL/
p+2totCPEF+jK6wGwAbA0nf63ikEyduuLOG3CstN8iRpuA4WnBZI6AYGc7cdH5qQ
H0TZo+fDQ8mMqwvlqluSq1BKZhnoTFjb8pxZEofRpZkLy++f5Cx9dvw/s/9PGBNy
YT3cL4NNitx5D9feFZpbkxDJevQZGw6jKcjfMft3vYj8m299VequGJUZHGpZusAu
Q4/obbvVFUUykfEJ99ZjLhJbWc5cTUcXV+TL/2X05T8MBemj1lkYingaIln8Mu2s
DPWgTdFmnHsIYPYGaPjhjd28yR7LouAmIVLJrzOL7MygFou1un9cTD9AVZ4ZsETy
nQQ1V28Wrr7DTG8fw8XUSo4g/CGn6tG7GQ3/I8vmhrtoU3f+yNCDvFROq8MB4yK8
5/lW9fBODfBpDsp+cOBB3n/ZN4oPsfAOalzX/sTit1+i6daJIlt6wShr4NlL6RXo
FkuupxhYFzJhvKsFRdBgu7pGVWtat6CvrYMedcfTg8aL+duED017WnBLVpZeU6zP
yUyHlCA9De763hCbn2Z0Rx/S8p/JktlzGfv4snOG3R/yQEbAg7o/jvEF6hKNs+fo
FJtXTsGbFp1HLeqOKNrGT1G3FBlelUTg+0cU8QvK/fL++Z2GHfaBGsS310pNxIXu
59IyjRPj+odIvjrX8hVLCHs0ZZNJl98K9T4UMelUaJNYSs74o4+IPrrdlGXmdPOf
B0aBEmZ5nGUZC3orFl8wq2yIo3rzqGCNFDulWiqCFQdrcWJXkSYIDeNG9BBv/+YX
yW6Qa3TrXUvuh5D8p0iPws9UZ8no8OCWAS/VujRfoancv7pG2cXHFxNmYTAzvAFu
KeiWeZULY9QTR0ew/DPF+qifOoyB3QVM0xay5mGvYSL/GMT94RpgiOdqpWQpcKuj
P6vgltFi656QEbTY1KdebYvrmnGZHr4edf3lUblV7XmYbr2h5nQyWSmUe22iJ/0e
N0DQQjs+4jhk5HC+NNgzlyjwaYnQM3UpUkEudUIISrGb7AZOEX9J13KB0OaeyljE
KZ/Mq7auviv30cxowV88cibBPt5ILwEPDd3kKNWp7A6xW/zbS4IQYj3S5Zn+Fzwg
rp8Q+WnBp4HHzwrB425IYrf+RGPBL+IbLDzj/HCj0ofI94Ed7gY8ECpxG9XLqMCh
hMxiYnKQNYIyP48kAXQ9sGInvYi/NCa8jNx9WEsfJ7DK/K/PrJeV1/UXiFMg4QIm
uRNToQ5yW1pz0PZ5w9molgTwhURy9RQG86+gifEV2rWn/pDFJNqNUHyqOw78+lyo
lpxOBKq3SzblrP76T6GKC4xWqWH6ZUEQtKNohHJUFDpGBJt/YmeJ6tRP304WeBkI
OkFsbkEtejS5ZypSgvI5kzSp++O2BenhshvtbDUARYvbQ8iWEFqd8EOZJUYCAuZk
VrZnVWnwSIys3+X2+BPzx6Hdj5GE1gownTZ9SUYkchAr1zFDONSW2EnVKziTuF12
jvfSu++QT5NAxf/FkL9wGflNfTQbJSMnjwzY4M/ysREjLct4Wcuok2ZZ7jXcVUX5
Qybx/3+oGQvRXK1pP7jg3mWx3+HnaXKV4IRG6NY5Jw+2QRrggZ4fZiy+qcT5SAMv
8278+T2SGx2kUbMPkqTbkNVDGHUQFtNMlR0CYFBX2YWozD1ROGqTmoy0qRswIiEd
iAaJKefg45DqerTP9Jd68rllw1BeiqmI9OjNcwyAdoBjOvSbuyLjxz0HpP1nFCs7
a77r+T09Eyj45CYap+nA9olDvOE+/DqDEIptZS2JShO3SjzdMOgllcuYvXiUHdyV
RLGKWD2rLRDgGIzuWJi1Co9cilCf4eTTB9JxgpR/ROuJpBjFU8iomDheZD70SGrY
jrTLFzo1hFaLcOi5hH1jUOgvQpBCUVG1K4n06BtgYbXOSuXp9meuE9PAcKrt4IbN
BNffRFvSTWaj7l+RNsVFMM6/eDB0Eb66Z75Q1aM8maGMGjRjJke0VEFa8CYaCUX4
ilcC7UUA4N9s/kCNZrPghkXDBvnFcjEisSxl1ij0rzUxUPyFBkwlEEXbZ2kdkOal
CaezIeA2kgKxywNg5pCUFj0NErTlYDRomEg11b3TKZNjX8t3J3M6zXjxLIhhWhGi
D4yXUT1KT18Zn8pzJ2KEphc9wFhjh73zMh48UDTY7dFkObGXRmMX3JfgeOGWpqfT
puU+CJdszPt2zySkqu3VhCVWFWoHld7qp8AOIbUVcasV/1U+LlNmg34eU+cVsgiK
3LZZq7iBieE3j4fjgbahEUUt2nv5EGuyXjgodP6qRB78UBWw5d4aBd05dkYhMYA/
RMNOPezPMMtM4gIUUR2ARxzawdZBYOl48BG2EJrLnGyXjxNHmKjUuUqPHL6HH5nL
LmyOh5R1MxTdY87waPMQeG7XKpFYkqrR+xcj6qTR91y8KnCBB97u4WUgE6Te6Av9
55TRpo0E6cdUzivq5nyTwIXRDtwqSmgHvURV6pVf5Qk537TCVzxr49bV9K7UepyZ
iCm6qKHtCsIQMc3omN7VsPWNl+Xod1DNbm0TWU6QdITLtoQCQOkV7EYjwGtE/2Va
IpKKFnvZ4t4GQsfixMsAqlGOKuObCV2uu+hvyZzDdhwjG5JFG6xKuKklUUDnQMIa
bLvOkOUszSHJmCCd8OMRNN/uJNmre48zUARzB99/NFUkxmhmyu+mVlZ2YK520Y8/
RdrnB//cLQh7TXGPbqESbtsXivo+vEW8mxRb2DEG7B5XuggOyTXRLoTSYJySD6n+
q+1+c8FjeAkkA3QVi5yaFyo0GixPhuB9b4phowiBWkyLVKvfUoXkGC5K/9uBeSvf
AhC0xcfEKVi+H8jABYMDwBhs8AFWRNwf2QOZO7fVBGy89GOxlQPJ4CdRa0gG4h8o
ZPMki0D7fvhq/T/BhbOBpnUrgwbuTH8pWRmCyWWcJbSV+dG+dlytAisSAfRSMcAc
X8yFdZpScCuYDJDPiYR5fkT7VSgeIoQ/t8IFs2LItHm19EkUMejpiL+H2/hQvWX7
XkJ25RZncKuJfLxNn0gxYkQyqeDzuhQzSjHCH0OTTgiX4ffkv9p+95tS8KbCvNCj
fEFOOCt7QUhsfaohe+VZGEvk+S+STVrPKh69sfxksqPKD+OjSfuXmTvUKpdYoGdP
sDOSzg/oAVS2EBz/gl3xkNRA+8fhJ8Qc4H3r/x1iC6dW8LholCiSrDzwfvu2zG/f
85MvhNUj9yzwXEPGqDZcZfwz+5ED383IleVmUGAv8gseIEENneb6+g9pF5BCpCJF
KVf9Xu9zJ53qvfq45rHuV+6CGwnzNOeDTepRqs2itdLZEefev5XZi1VM6lMp78h7
5J9uT8AGOUCZx4F76CQ4NK6AmsJjtSOTODMr4BCP2N4lLVQp8SMuq2mulYCeBu9D
8gMINpIHo5DU2/kbC9F2Xq87RAhl7/XqXBAAnMlYRClVecDuM0WUmPIQR1VoYrcO
A0E+2eR91SxHvDCRsHILX6/+CUXPtaQEU2lDX7/ks7DT01uLTXRa66J4/FH0gE7Q
WEpT5yYvNkTn4ipX/UCvBryakWLEZCNsFQQsInuUUqKqtPwsiapL+/Mpuj2xZHiF
p5bHSZ2K9apfJMElGZYw+LxIrqu1Y6+dEL90MTKhiPn4FsG6Wkb7EtnAElzyogth
qZO35viz0o1u1UKXOst9WuI7+afJwx57aP4X5lG9J5FWAHoF2ZWRN+PxDuXQyEic
vSP2A+EVU1zzKYuvChrepIZVrFlrSgFE9upLsVDgR3sYsIaFZxgMgMwp4aqPqDJl
mtdncYCRGYDySpnwPofEprKW0zw0aGzT1RhjDxMR3HWg+DNszcX3qSZNekGb4JDc
nzk6hu17ndRpIrgZ4sRbroPDwIKTJ32PisWgzUpnB3qwmMiRMFoCrPrB2o6CZ5qg
lNbraaELZtrqUenCcQkV5joqpfQX5PVcZ2Zu8u6z3zTGfaEUW6yDtlKysNel9CMA
yLlmGvZWuplEEvzbmmyx4u1Va67YCqMkgF4HK1TNauJsN7mVx4uqksEjUO0HV7x4
BdG3keA3+K6D7XWQMwNvvybvt2niREfan1aRwdZdb+NJyr2e/fLKvXN0ITz/BiWg
99KuqtttIHUsTWLhYrIwkaiONoqdQZv8uwtZGTsn0gTRWFkroVMSWxxfA8Tcsakg
0zdYUGMz9YRYudGxwrc2tAi6RoT2FomWO78Ksg3liWZnrhE2xSpo0jzdcZw4+8/X
Fx5gxtOrYPdYbH8E0Mp/hBBeVVB35qHhbikCWdcnOLf4WdX85twIdc5nNtFy1LVf
j0demoumVhI19mfbx42eboTQ+dpQI845TmjxnRvZVaxDY2C3nVE/v0mWAnQLQ3eS
SkX8TJGu8sVKKIghCqNQPYnnKa3tzclluT1dc1v+TUZSIBYd4LvrCVusWasbqfyw
D6LjHX7Xt3P24hG2d1Zenql1qDjbbyemUVJH7NuIT6S7ZGtJf7o4FFeXO28RaSq8
qX/VUbl3FpZUy+HV+g/ofJlj3YFnSSmUxGr1kmBDO/z3q0A67AdxaKkZKz6fhIfm
N9V345o0o2fzVRZ4QWa4w508Ip+sa1cFWBpimrFX4T9IUHZ7S58JyaxdbaEwypQ+
rY65tvsNfeqDKJC8qXYTOO7qDQoAkVG48DMLOTZ2JrXmuTY4FKRmQO1J2Zugt8Dp
PZVkVhvkeDiJV+udgNWqUCVQINPagUckOURivb4tELLQX+1+w/NvyLpPh9nA+ODt
cQKlFimLp3hJ+xkdp6loMPQ5iyxlFZf4Y0ArvwPd8o8QN2gSnUDkFFShzfT05GSL
yhn7So3aDXqbRUlzoz8Rd5/RMVqmKcfZMHKEEZ5CaafINVZnB6/0DA7bsc7LcUH0
HUNhmUisPvqz9n+OrqwfkibjkERQ8sI2Y9HkUuwpaMRccNWnRmEzuvNUXTMPxPWy
RqajpEUTs+0fvD0QRtRDgmSeJl9y9n6XVTExBwqeeT6P5xlSMAEsuCcFF3lW6Dz+
zzJaZvmrQK7kISxFHoU8ZjTKOtYakxci5543kQS9VC15D3nukNdamfYQIbz8bb/T
Q5LT4C82yyHZlTvEfA5RN41K1RCuaLXTE9NQGjUHy5Yg0+CS328CWPFGcF53cj/C
kx5wh+spz/A1+khkUpgpD8minI+fvzkdKqMmq1sJq7FDNNpk6nDCkxEN+B+awzGx
v72BSd7Rf2GPuEZyNE0Fz603F76n+d3Taea/cbWZ2QFy/n3SNGTPib8x7WeobjXw
kkygX6lcWxYwDZbIoiG53qHF1KGNbpIJBtRZ4LGVAFpqWMicgbfWCBgZh8slZN0w
e7bAn5lN+PFmngU5gPyx/GgtiDEUQSn1QEIDrTPqc8gSdBb2UxMNH4L072FbYVda
132IKDcwwd7wLGcgcJIzcNr85W9cjLAeaWIY6wOHpTyDBl1PMTRQWjlT2MidaAI4
nv6i1aTdtCc83hRZDPzX2KIYAglvAGy5huFEjEDve+ckVLtU4/lGY/uWo0fmJVAI
2PXCaQKEMss/KprMzAMPHVLb3jdoVZaMuiUhMFfETH/mLhXdJhp52XYd4sWEirkS
UFkN5vpZEc8ky64oLns2mXvY7ZMP4w7Ar3Siw0boZ4uhh2WEJO6lTiUR0SrAsv2V
K/5/UPTeKDX09ETky1hXp0ca8HVjzX1kaQIwymkOIZI90J9t9clB6CO/nKRfqYSu
rs+YDWkB8VfM4DA62ih6hdJD+v2GKVvSDjOBP2oJ9zddIlN2/rZhRvZJkoCTZvNl
nWOgbx/JeoaPk9n+efwpW2mlsG5dnQ6wHGL1dOvo0CwOv2yo27PQEBAACE85yQ+y
fJoquZBF0fwfcW3T70d8HKEJApC1dpuZpO7TpZFNm/EavhThXB8ycYW3PSD6VT/6
TTlTAnxXrljmrYLfuhNDZYDx5lxxRhBdtH1NtVGz6wSMnKG7uxhdgf9kvR/vqHA3
YCGI8EKJuLbhUe01VB8MrUBt+qt2KVOlvZ1OS/eOCzYxNisfPYbEpBSOP/Msrm0G
RQ4/EJHaME4ObFn72VTZhO100QmVS6kSLw6zto3CXSu+BV1qAVIm+RwwgoYb9Kxq
yk7QMOry6wR+EcFQa+tD2MarwyXitE5aVTMksSg3d+aPFKRZWunmxafVCpTT4ZqK
L0Xj20CTUtEU3/UXII/FE/j2jq3gZ2NVRf/kzM6R7ZSCBe27YYe4KQRAWUkaYPZO
RpDji+JXLbyMiykHUf7m7lrjy0REet84YqBSZELI+THN/kfnH/hJZMrrVy6zF/sd
gR4eqSNGyXmXKFxHral2D3853uFQCxeSM6RFzIHN7IZOCVSQ1xjGrXT6v7RJG1mb
KD4KKL9hCq1865YJrLNAQJtxgfyiQMCX+kE0OKtHEdl+t05RnQwy2e7Ul7x1l6aL
R+Kd0Ky7Bi9eXjeXl9R7Q+D6vR1StRjkLlKg8yfK7AzlcuLuVHVxNakXFa+p5qUM
5gCkFGu0qtONXWnCKvFIV4KCHrZN3K1Tyhh6FLk90W9rpmRLWtKRNZDtQZFnz8l8
Mena2iJQxlw2EIq2EP05D+JHtlM6JLNTlVvpGAS0VplXsSf6c75flkGqH/kILsdl
oNZrWuk2FLHqmQzjMeSPZJzpu5ZonJm6QZifyw/0xjLFHNjTICjic3ciZddc1y/v
pf85XZdEaxlEiDWXA3gYscjZs9aD30dYza7L69o01tA2I4dLA+M+ucp33+emjh5z
cmRceHgTVLLoZAuTEBXcXQC5aCsfGvxmQRRBaAKhN/Z0IBqFDtipCaxJPKvWmqFt
C06RP7uC1wX9m77NqKnfNYwOZXDhIGHAwxEaBhbv8vhf333qFhbIdEqn1097M8Ax
qDV+e4MNgoDi2EGn0Pc5iGrEph95FrmAmVnbDhwTmq730RRsozQU4voG3dB1LrA3
wiFUt/+SlVmLMJfPYu/U8AlsvzlEKQMS7GYsM69wZR70HxRoqn2H9TixfOzDIK8g
yXzfIiorr9Ed3bhWQ/bJda4u37Zc11KBnOcaMfNiurmV6JDQI4o7+21ldsgF5HP+
Bz8eP8N7IjnN2PwVsN4J6GBtm8jdx+XPNCAffFrAEVEN2dXzBHNVC5lX+3Nc3nxA
c951TDqbeVbiQxZkBy+1Tc2M3JI8V5MvzZdQBK9yG978hNLvs7UQyNAFbFlZS5+v
r2URB5wY1TNdPceMoeAyiJEmWnrpIMM4Xa2L6ZKbcJsuWbDDE4fjz/1uyQgHrU95
5MUUZTcKPmfVQfuU3BKzFt4/SJRAU0oK2HRdf0oAzKcJcY53AIgjyYSly/0OmXj1
OHuWLjLivub9SU2eV5Hn/7wLTRUTdY1eQv4GmPIwefxduk8mbSsGAewdFUkC7g0w
Z8uw3pDiNs4r4hEZ4duXDW0d+JLMw0tEwh+yCdLCnVoHEJccD6gO2Q8aj0Y4Sb/o
6YJJ8BIL+Od8BV89mf88shnpkERDN/8LU0yy7iACFLQIdMJytZNIEWpcBW4NFFUk
gZSS6rOCTWnMv9CMzbcpI/pIi9JE6MYRAqBsPuL+dHlTIBchfXpF8xYKzX6rXZ5B
Fyt+K0P2hhHoLO7MX94XVy3tHEEXiPnPIDf1A7x0poMARLWjexEWB73XuQM6kz4T
8a/ERJyUj4BzdJL9PAPSr0HfEWUkyWwHEGbwiQenZeojWH3ahnnscjjMM/s1ICa4
AR9P4Kr5Wx109+IZirI/zNdeeQI8sh0cxK/kirAJ4OqcDg7bTGQTJaIeee5Ymm6U
OjoFaxBVOeRLTcoAomtKAoJqdQokjCICCXONWRgt/8ZU4KmiNyFBOmw3MIpgF/Lt
stZZEAQkslHdvXnr9Zdi0568IACIAcwu6UKY5HoS6HAcRQ4ELU3TRctjY+AhggbC
GzNQ+V6TFNDl1ZEMrQNYUB2F9icfblHuMwixh1i8UJEVvg18rz918+VXJ36PUBhx
X4lDvfNF3IZ/7BUgZZxUzxeaXfCsBFjBBAxPczqdC15MnrH2gCPFerOZXzvRqwIj
6rexM0TpdafQrFzIyoAaS8dB8uIvRvpNXw1Y2ybls2ZxalWIb3Q3SrO/pzDf/56B
PyPUXdy4Cnxb3yXdNaS/5kIUOLzPslm8Oz+djQkL79iVPuyowFiYi4/wPlaECy91
JBEN9MsoRdUex8EpKzV90KONKpHgxHuSKT1e5gXlcl5dUREq52qnyAmCabVrme3z
rF5VUi2k7AVPbbYi8E8C8fAKOdCN1vycs0uBzM7/I0ADZ1c9Q83mQAU1nS2RPKwr
+F6NscKJ/mzlAkrsgv5U8onzLWFUjuw8leouLs5nQf7iadedixYnzg89bblsr4oI
F6wS4PYx7skHOjX5Yjgj4eUq/0sBjx/Aypm2xEf3URfgZpkz1DfBj/geEVtDOwWN
RKSBndgt5VgOjYpE/g1BQUyUnpTgZie4YOFmCt9TadmUk1emBPieoyEhL7Uaam5e
cE0VABOLZBRlZHAvz1XXwBpt0RT2ePw9OpYppjTolTS0OXweD9+Rme3wjYCY927o
+jtN5a9pHCjx12yOSGuucG1SZo1xHKYAjjmEMWzMcj3zr5XiP+EcViVphL6rhNMy
oW2bH5GttZbUKCC7DRopJ3mBgYZqHRF477VbqPk1URtbH/7HbG90CadkqV/9wbu2
SXboJVBL+ffD3PPCesMbPVxIZHot+0210pZuMWnkZWxKhs+OLcxEwgvUGFwl7qPT
Gn3xjCxM80a5E3Kj+TANVc4NL7nF40nMUBWb+m0n/HIfmo8kYIXez1lhmw97wtw+
b2DpfjLVW8w11OlROXcl5516BTtdughui4iJjHmr9ZtvkXrUtqWhC1stvxxGbgfO
Y5hO/0CmuWtNzDWy/qGDEQNbv6vj4gfysXrHAFYPkJVkW2ymmD3F6hibJ81z3kRx
lknUvjfxM+50jSyTsKJQR3rT10dkStGlvHNOQw6pKVL9yZ4TNujqgt7ep3/JuqnK
UU5Xmodx7JKrf4KCUAVJksnC0QoXBU77poYe3B5iyvbMY+0QuJczPSweT5jLMN0F
JrY7bF+hhyDrz+CfXqbZ+Fy7Yyg+I0ZF5xWN0Wk0WLb5oLOdiuVx8I4VnCv+k2fA
FDrlVJtMKvCQAXEU6iIPaWy2xD/KajaSiXR03C/dyKycarqwYwV7ray3/lz7QuZH
Sh4YvCEH8bTLmX+fYoFNdcRJz+Kp6wJdnmlr7iiV9Bl1q5i7BGnsY/wR5K720Rpz
KAlOS01c0rNcnngRAv5BfQ==
`protect end_protected
