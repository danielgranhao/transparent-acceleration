-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
Q3kL2nVeTjgZitj+58cqtpDUydQeFHnltilUQ+BLgNDfTvD+DgSW3xHF/rO9uR2p
DZ4lBHh8aBE1Ax3az7JdZjv4/01nUgzTlLF2uHTNjdYF8LqnSKsBqdyMw80hYqya
CjyEQ4DCCO2Q7yZgyLZQcJx9ZrHAHoCBCncbtQQfkgc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 12601)

`protect DATA_BLOCK
WPxElX5aVeGDf/6epuXkKqojsSY3/3wCUm0/fxfp2b7XwQgzDSImUdqvY1XD4Y4/
QkKm79Zeb2MYYHUlofiRbtNiV9wegPYsip6BUG3MwSVamuvngjNW8qbmZPPpQZdR
DL8tI+EKgD1ZZ2TYW2N5pWxtKu8FE6BA6hQChf0HwuICheOiPC1K3Nusx2Nu8vhF
Q7FGX7tokc/EIONntLhVxP2EA4cmPuKIswPnEQOPjvvaHS2NPECvGh0lqs08+Zo5
OGOPheNe6rCLxWUb/DdvPhQAr3yRihb3g1+CsOOW9bnxpTlye6GKik/BmoR7hjvy
YWom/IgeSdlO2k/CMBGMH0hC/vnk5X8wm52htNYEGTW9zfX+bPrCUvw0N6pEgcoT
HjKjH+9A/uByvnDBdHBKtIp9LG+jux3+T32H9CdIZhy7UV4xmfN+mHJ+bLMn7f56
xhxCE9+udyWdSEIoVvzK7J1cPT3A/euM+42IZE/sVIxlcWujR+2dSGTRoEwUndnY
W9cGzUKJcRuKU2Ji8zGUO1Fw9z5/h88U+NyhZPIzIpuXqOugVRAoon5UjqXMl8Tp
7cCKhXMSGr6qXgnJGCqs9dE2sjB+ZXx76LP4t5mimFijhEFTw/zBgOxg988WocpT
Y9q/4rDP8AWhyq4eDObXSFSteATvV+JJTcZMkhkjHS1c3GrQFrdNw/58B2BvlqR9
H1q7gASn5wWb/XhueE6dQMwAnCbQBlVjxeNjIj/ZBJ9Laud3ecJcgjY0VGVghrd1
vJ6R6HDqNLz3VwFKwCXS9nLZx3IFMM/zVCK1odRrmqQ9YiNhsNTKQuk5NW3MSE8y
mpE1hPTyf3mYmtersP7r25pFWlYCWnlgsh05XghFp8vkDJwvHRRbPunMoEvOaHQg
HjFMaG0AwFDvJxM+usBBCTgg5E/9DZ/lNPTcXDyfCwf9+ZlVHydT1FVxPIzzehaa
iBSMkkiaZCfbX8HCVvrTHQi1uPEP0EhW10mm6zdqiUv62U5jgc6CBi94Nby3UmT/
e21h5EiGjUNjjq/9aFTPbVM41XxC3phyjzEcgczEwcLoTosBV8DST3rbeVCZ87Zg
pRtaAZ1nX+TojOd85oNZuMuA4/N+dlE89F3hrG0eVXMHbzhh4x30Oo/eoFjq0G9V
PehzTWdUrzxkARSv8bP3mxWAzgK1G6h61OSpK/nYo1wxC+8CG//aALee015gxBgd
yfHPcIV8TdxuEfqSCJJyjmerYQ0jYyilychivsGbC3xkZVhzab1yM4LRjGG0OIUP
4EH2kGYDSdRYTwVT1hnIEWbGICY1L94JIiYIU3Ujook3bnDSE9Vi8jD6kRYrh6/3
N9zAUz9jgOIzNHkRVMX1jJ/7wmRgkkxR05KW2DRSB8itORzVrkma9LI8yFfMe4tu
uXHsAtG/l/9xAp/Ck7cuKcCWjy8fD/dCXf1XxTf3MHX+24kMZHCzwZm8texgzSP8
/YPpU6/aG8mcQEQ4tJKpnEBou+reA9lYtyK8LfP2VAYBqHmQEEVkov65CdkjH3N3
k2R/nyDBCQumu0zvu1+tt4abdZZDWM+6vAOiGm96zdbaSIQcOw9OuadiCr0Y34zl
JcV9eh52yk8zjCsM718AtL3xytBUPoJvVCAf3BzFtR/n9V9jCDFYOMKgIX0ei+el
yNC9Mp2Gd+A39hbcO02ukTGUIxFlky8uZzKS7h+ltVGQ3jjFuXnb3I3KlPZb/zoL
QO3r3baAOxJHyb7DIHzFpmSVLUACBWKwfO0lF65MfxNenalgP/JZpqFJ9tnZZxWv
hpKMWV6lhABR+O01RjWHfl8a50WMkmrkTm+wKbweyuhKiVrDMNNWHxoCW7nK0bJI
CpYE9FGtLoTBxB2OBW2q5I4hNOiu2REeFS/JGqGcKjlH3gMYR+D5GymTyUp5q5+S
O6gg8/MaaOjdn1TjlDThdh8yAZqX/oTX43wXOXn5QWq0bStfNs0G/rDJZ9Nj1xSd
LR3eg5CjW/TqFAYZ5lGwo3uqQi/rT3JmDT9ZePa25bDuPUT4fAPZ0SxcFulLzYEb
JtjVa9l7Wy20lFlOBTf7c9th1iZpZQ7pvjrqwkzV5AGcuOKpE5hfvqA3y+ul6Bk+
AFivXVzEJbx61x87B1Au1GIJPRsQvxb1+LPEeku0bV7kX5iScLrsXh2DHdNEMjiT
YgWPdxVn6aE9CzyRlGA/gp8nfjyXN3mlvvwXjmQEuIpcmKpsOMckqLNnVvWytCDt
rsY5j3euvP+Bd9MxkP7g7JWY+m6v7M2HtXBPIKAGFOU/UPsnfJ0FLLQF3Qj27Lgp
Gkzq8+1A+J7RT6V8Mkn7Ls4sR38IMnk92NSntiPdmvS0SHM/KtXNCFXqzMv1i1Hh
YItv6hThwFomCWOsHYQ3oxDZR07m6QRDGGRPhr4Ebw0++D5cTkG4+c3fqGCAktJ5
fMdMB5YMhxveqe+1fGBEkyZdsunDo+rkodygy4Uhp0KRZ1r6+FMmnOiRGSZ/LTra
JpY6IGgRJ0YdMWlmoRS5FBVAoJgvswuNiZKsTndPdRECv2pHWThr2EHNpkIgioIZ
bXJOwi2HO0YR1cA0MTjpe2hqEOpoqPqut39xecJ+db4/SsZx7I01c8i8V7c+oiop
R43VsVV7iM9/ZLiZeWPmo8Zwj6ijMswZSqphYyxsd7yRSjIgG2SgmrPVKK6d1nQr
GOt+FZH+LLlV4KXKL7iXYdkM5nCqXfK2GM8ZkbYNJC+fGbva+6jdo9dhbiUEXjp5
eXo9c3ZqkhJOwIm1goD/DVHdn9WoWkQDvOFO6gImzyCm7uominkca/pBTeqNSZ9B
d6HkTMQ0uc1XvWb6CGjirrHGkmcy2Ybg8Rv/zCwqcikexPHMD2GJ+mQn6s1zIdNH
dQozWSFORDKAJmGvT7CXrab8vLft3dFcl7SgdvC/E5bLTTRCib+v7vL1Q3HT9pdW
z21NiOrWOFyq0lz4YpygMstpncOgd6VdK+t9dlXqGcrcx2C78HXqoXFYiS9jR+tw
esZAkjSUgEYMvYIjkfaoTRXMWvEWePtLTW9cH/EaXhXwUlOupAunDj3oQNJSSqP9
03CDK5qYWiDgw7GZhxSdMckZb4uEGNBGupPK0yFksdmM0rHt5O6zAAAtuEYz6/I1
E6Y2DEEBQsZsqGw2leWFASBKms7zd5KYdJQBMC+DRerfM7eNA4VyO7qNp020qmzB
e610p0i3hzXf+6sqBHn328uIycPaXTif86vZwOrI5tB4Kt2MNeal1hEUEPwez12l
sdAIwvJ+TRSp41wGQclMamspuhcF6gdhziaHE0qzfkXx8YU443oxy2WP8j/F7BUC
XOhL8VCUKXkmt/yOxZLoIutMzCMD3+g1dB9iWACzV+QKXZLCFi6mys6WycbF7fut
iHPOPc+fJxqdHJhuKB9vjqy+vlgr5ljOl492Z9w/V043NFx6BLTh8tUSXcPCxxHy
KawHiManSnYk32bffeAR1x1Wu4qpOEW1yIyQpNiedLYii4I6Ou8WIk+PGi3wyo5o
Qkp0pm9zvtJdlrB/u3uWkxETjDWaq4L4Sdrmxs2CiE08UN7VlqazUkt5Uiez0DiP
J2+zsX3SrJkN3f0hdwQ1oGwzGYz9qXs3qtvnZn2MkqeWumAaGmvECLiaBEF9WSTN
YLyVA+XCl26ZaY3kVpnVRR+5RCA3YdSBtn4536GpwGRcQ3MoNVhMfu1W32St4SKD
C9asnyliQuordShdw/iXCyYfNDYajyZUQq6Rxo+nFSxMRkQW7baO1IBXBVp8boa/
n6u0jon4ZuNVpCTq7nGDAJ1HB/O825QeMttFKCg6HcH05Ip+acHIw8gz3KM5Jh8C
cWR4hUy9F2DI3oM0MzwdVIS/kuoO9pqD6xt54/2Hd5J9SvSl4Tkg/kcDKUWx0zsJ
BZ8X+u4Zf6QH8FodDNuSGKBZ2FjCYbpZUDQIs/TYqvz1vrmBho2kDtqQ/jOM0FbC
cCeqb8pcr5d8HpElTH4BoWipL+uzfpghs3A07NQLBoWipv2xTflrO53R9TMhF68D
/aw1JKNvS/y/LRZJltf78T8jsEz6SBv205P3arHHgz08sqD+vhmXegoZ9iXXVED9
sjiMzEWoZV7BzrohMgRrsjUWnk+e9FcYnZNL9KBzqlZy/00lrBQZ8mvnSCVJb6HK
SQ1hXSUSp0NgFUrvZ81fTw0Se7yQPWEve467gtydm7Mxs1wePll/C+phWRpFrhJ1
CUXLKDXpVm5F7C2VgfLend4wBW3NOLv6uO122mDqZaCKchL3x3FIbmcoFLvsRl2K
E+pnGcA8t0Fh8n0YKZYL/mUPzrHmBseLNYdWDyL1fmQcG4lkKDMXc6kN5l48xPhl
as2gfTycOR84ToNkVuhfsHLAHw8nvMVk76bTrRo9ENbqQdRiuMlSan9QgOafLzOl
s0ww0vA4bM9RQTqgJnL/adSkVd6sIjoNhlgHsQxPpF4RvNzaxSblxQcdkK6iZSw5
UTjozIzEkI37qZriyTgRHhxaLaJKTUiElnEhHb638VV6BtLZlxwSOUCpowXuseSv
WwDzZkqEZ9kEHo+8KkEOnAQVekMr3bNl4aSqEJO5buRnNB7O2fzZnli/7Z5S2fEa
ukhVbu+/f2xL4rkxRfHUIj2Js459d0xaGVPdn1ah3m7rwPELX5qDJr/yRQ2YK01j
28DgZihWum2qDSgGbC0VDv4pQ50SFIVydcV71V4J/8p9Mm1Qw2bMMgwS5Ffhvkix
cHowA3mPdEsKq1c00V/WmGN2I35s+t8+UcAyDpCsCW6kptccg8EyHaW1rtYo+2eZ
6R6dcZX2i3c56E2H7nOa6w3PYbs66sXubv/17HQKGsRZAzIr33QfMOwYjcEBaF5D
udNW7XWcZBvrHq069drIVqdAH6vVmP23jL0uEWP9SlXakeQ6Bk+fpA89+l1vh7S3
Pqw2KOV0BP11+OKu+SSRgqX0c/ShWSjbVmMm6syXGlcm4BAqKowOKJy/qRGXCt8c
w/2weRFUABS8/8yxf+aDv7pD/2W8n6GdjFl1WPvaIVKuBk2CI60xgjaNzA0KcJDw
KK5yGC3o556b/tsAn/2b+IZPSEfdUXd7R6qkPwRdDfxfS3TEcGRJB2hOFHeTWPoE
7yZ+vXETgGUM79BYSZ9hLFHhmk+sYpRu0bCKJ8EIWTQrp6OHEgRorqiMQdK1Isxa
Ty7OkeINiDqP9CrMZn49J2I6y1fMIZQfGwdjeTzw9msdTaY+RxpoCngvt9mUBqLf
3LjkiKz8YSzCTI28NFULbdjoPkY6xpQa0L5qeeteXq4IdYCXLqS93SqDc8yEpOXB
2u+sP3dIDUoy9jwu1P4uiFHC6KlgQneb/P88GnErEBX5s5n7b64AUiq9CX37Ubv4
hJ3xVg+UxundE0DnAxMk2Sp1ycAiv83XfRSl349HRVLubHp8ZqX4jM3RtFYmCpb6
ezWbHAPC8OLDLIeQNM0SqonAO1edilpRXOrltfd3xjVL9Zn9QsUScfRZsMdng2eu
jRQ4DV8mnLn0kedP6ihk0ZxUsN+Kdsl5hsVJoOCHC8UgG8F0EbQ23RDuFekOR3h0
11/spfpD04snSR9PfIBvhuyuhWG9cK/cg/p4S2JsdJYzW1+hQLTvvDsB9vkzqjM0
XHjnH+2ylylbCXRDhxs5hKdjHeSDvqxbrHbApHvjPWayrzhsR0WAXTsUSrQwnFSH
oQI0ScbHxRt7aj7/ioaiirwgKGND1ekvOx/dR1TJcLJtljaGFKyJOkHCyXl/SdEh
PJRAeO33BkOUqcDyBz9n29rX/Y7k7vugkI/IOWuE4oMR+pU6IBMa7G6DHyZSUCK8
s0ZPqZgCeRO2F6BaLM6KiHOrb22vvS8+wt0Quw8n4YZJiMrjxsphRjo8YeECzAOs
txMoRizgfeesXgsoJEkdYxUBt4CNjvM2heCppEiVcnkbpQpdjXkcfIshZQcJlRof
mNwoqPHd70KPPOm8WWFcxQxNkcmkc+NVoRnM9z1WcueRVF7Nh323WRvimXNE7wdr
wBxK0xnWrkNQpS15birYDWRJuU0zJM0RYxg5GoY5d8FwCObvcs7kTCZFsIHcQYv5
JOo2jbZd2XBcydwKjjyQ9Aw2AL7MIDYZtdVEFx3mHCoLPM9lvFpzZKOqj3+aEany
dr+xM7PL1hSRJ1I352wGLM2oU3OMCWPAD3ikFT9DJRvD1nU7vd0vWk248hqAhecx
kMBiJT6RFQC/2sBRApCqybVmM8y07BOCplOEEYG2YHoZauwdeCK5/whTXtBDF3fn
YpR05PYGTznA931Jsh2r0xS78g0CMvBNTyRQLwAVlpOPEJ9+13AEwzgKUnjbdeYe
VW4A1K9KPCUtObMH1aIaznT4k735kx+U1suC3gzFH4uvqxjefh1hHWiEKram7wgE
qXXBx47YOkom6v5ruzXXAKZbYBw6zrAnm2F3YcT0A3uSoRNW1Mz16sR0QF5mMKxq
L2A/p5qekw0eihMi5Y35orDQlHY6gOK0lUnorRygDRhNnazH4N+TR3YF6GkSbawP
kDCe/dz2y9zJpif2osd9Uokiz3bAiaEORYHe4V+lyD/pXOMcx+xmK539xIFgpnoE
hHGtH+d5Tg327trb9/fqnupWHk3bknTNvDOtvwdbOjx+QSVK+gwjAJYliFV6GkgR
RvcpI3OlWMacxEPdThG3zeBZeZZ9T3+LeWVDb4Xc8vvWcQQWbJFUwuVRUu5C1WI7
PHV/MybnSRfp+A6jWz/+5wXELu9NVymoXN+h2uscJqwms1dLNaLHaf60/XWiK5cn
1U6KpqLEzcTPtTLQ6PKat6S0Tup5996dTOf3wg/ovNvtsHixMK+DDtPnTT3n0GJv
shIkP/hmg6XAyYAOpVTKs8nx1tRwLum1HMztyOPgcb81ioapAuveZo/0HbBwWrno
ynSavw3uOAB5uob70rMUyqzqDM9xPkPftk3jbjV74qegesIZUEJ9h2TmuL5/XSSG
xg7SYgjHEZkSvAoxq7Qfs0kpj20PO+ESXd5cnJzRBcTcoW/g3Tt27g/o88Jgz8L4
z8rXmdDWQqWEuzkj+uLKrHlJiMjqjh5l1ydlNUWj9SmDOtTgdId6laVk6Tav8bES
Y4jWcD6UA5UrP7AX+L+MgwbbVOxGGYFVCRyZmL9r0XVHJdvRyojrV0IklnHgLoKT
60fyC//T+cf1Mf0NOZz7S/lsgzTaJ7iyHbEuxwa/RyRZ2r7adsmkEBUZJDA0qJOD
k17SppewY16Fr1SZo0sUoPemcyd/4Jd4cfEh0ygokYQiPw34dKu1jYW1NV2EaAD5
0264V6MO+AB+TFGU+s2y740q68XKavOjysv/7emrkVjEugyGdPz7A042BaBecdLK
dxMjk+IP6uyjWbkxXxPstZoMVmMZ+wfUszFsVEQsAPaXDamSDFcdC6XaVTfQ8knH
WZPRVkbtSHOfLneS44QJuls536uR4Tk5UyX5nDgaNIcuWEUztL4fm8k1AIZNs2k3
73CINX8vn31u+SkJXsyIcYmkXdoe+Oy4XiIxLoD1H+WSz71jGbj5Wv5+qZVVw3wl
kUKDoxhfsekzb0Cms3T7WD5TEp8bty2nfcSLSOZLeuajWqvmR2BxzqHt0C27VjWw
HaaqLH0vfp9sOplIpVzzfRTh61Is9njd/+GlrqhMRRIRrzYb0gsadTYVA81n84KC
Aq2qk/Z1+4CR45wekRc74zZeIJOk/FT6xJ4hJpsSr0NpA2+++EmGNSMZEDHv1JIN
Bp82Rylnu756GwRzhsc9Q84oxQgWsPgvIVPavuPuCE48V4Jlwcc3jdvpqQhp6fYu
K2ODRs6JAysleAtb2THw2JXYEFQvu/tl6zDixyJgJL6zhQR/vNqjPbNM2b7utAO0
/ipMra1cSs4G2nkCUWE+bo02NCsPCIc1k3EblGQ8wCnsrWZVrqKwNGIVVCUs3U6n
X34rkmDhyxhdi69WOZA5xzcY/oODqE9OI0UF7m6n91whBXs69BgIR6P6Y6hdrxnM
rCqusU+FHfCT/RUAaUbF+d7PfDRgyUm9lzL1sq8CKzEmt4jj3fJLon8J2qV8o1cU
zKrH4P7/zy99Lkdqzt7V5gtfHgYZ0K2M+Pea2wcbJIDXnzgNe1jq/eRHgN5jhfwL
LDeq6daQtXXxep+HC7rKD5Ow/Sk/8EB2UkbqBd4iHYc91u1os41BZnTm21OEG6vO
Ex37/fMqUhuc5lALUVWKhDDVDV+7nK+fQBWNtKqCBn97NTF++Xon5vH/6RmM1jjz
jvolfBV4c9hI70kMAAzi9mIbty3oqwEqIZGlRLj6yf/VNOH6REng1w0neJ3GGjv9
a2vAj1EYUi0pf3BEclhZFyvpO9zyCDDYvcKkTkxThr86mmL1W9uDTgWvCiPVJlaO
X0X2bVla0u7dO/PbSKuZ692FiAbmxVPd9Mpx5yd3W5PuWDKddfT92jLkbaq6lIeA
9SP6SJA4D72ye2JPkgBNDdSXLQPZ3to1AVIdVdTjZO/ZEwEC737WFHgeMAHP33Td
4/3U33tUOJLYiVL9qC1uRkTY57/bCIoCXFIoWeDeh+U01pEgpUJSWqNu0UcwY8hv
dcWoNKO9l0+4/bNG9BKiVMO7iA0MrXPhHdbdWDYTFdL1JAdtftZleu/v2hLq/ebW
heGzyQ9tIG+kYlsRtxGEL9F4IuRkaUp4UaVyShbjtEdgjXjaPT9FKoPBBcHatsmX
wQipOWx+Kd+p3PJ66I/Sj4pulUlXXwHHGBm/GxzQHuP9Jm3w8Z0dHM1ysxAqj6H0
IemUJP0IoH8u7OVrCK5HTS9E+Atnnq17DizEQFgvhgiRtO1St6JHmemvSeK3t+kR
ENgfMpZNLr58hncHu2saYt1Pjb3DL6BncuZ/6GSB8KEXUipE2xAwZ4urq2urWd1D
45RX92F6C+NpvIbs/PLu9oygnAPrcr31BQ10Ra5Xi8kv9yTJ6EGFD1cBE92ekjxs
rQ6n+udah4aFOAIVWxoFbuD9oPE1GRGtodmOxJBpS4i9BNPeJ54rvRw+/Fa5u1U7
3hi8dQ9ZK/izB0tbVdHJI9Qg8f0TV2fYrBkUG8WVM1HN8QO/H4dUg7eX7YdRlwok
vXBDr5S9Bn8o9N2oIklc6/DZmnvtbfZ3s4NKlRuRoEec6Y4qwO4ECPw/kNqV0hCa
slfpa9dWnXY+kujuzMwnBy1fagNzmYM8EFYVOj152tPEPH+UVz8ywFqNC8J6ymUG
FeShrexQxwWLC4GaRhFL3kLLtD7uw3MtMZRGxnqchxD/y65dMjeS9c2ihf/HrDsd
Q+OTOWcgbSdLgFZADfJYsUlk2SB1o369zS/NSP9DYjHQ1n29rrhVmCbbQwcT1xt0
Q6Z+isZUCzMvbO/edY/9BNFTKCVjLGGOswZHF69t3Hf0vqBFyQVsMgiXDYBnmA7e
vJnWvbOX2IOqhyJL26S+f2dCpAeXhvj2G3ztDwVySW8MIU1SSi8/19bA9NFvxW7Z
HDfeoJiecNjxkLCg505sUuty/xByc7wusSBA8w9UyrWweGuHuc4QvrRDX5cbLGQG
WB51eHkCrIWGCnlS4G2tKxigi91CW/tgygo+YlOhKLZmfokUywuHI80OMdkEidcD
zhGwTuZAKezSq6dgFwDYLuuIYl0J+2VYWkG9nZXpvWUt1JPwrmyr8vsgNuifVb81
urLFd79GrVqzTLPXGAwsZhxXe1d9F9d/r7K9rGJ1xL52g78tD0WpiK8Pc1WbosUl
AEd0sAACllf5mt6sYi7wTfTPKdjRqV0rpRKk4i1IsJIqmafU62rLbECKx/TcM0na
/ezD6aos67a7wC2tIJ3V5B62mJO5LgeuK3bnh49GqaJG6504mLTranWK5/+Rwmyg
2bWKqcr+m4ShU1jScUeRA77xcgEA+dMzQJL9+ihPUIKy0o+LPON3/WYq2awqG+uG
U8/jUyD12djjVw411SNry1nm5ud81meo55Gd7Zxoig9vdNCVuAcCMgigUFOnFptg
9rIIzWzs5ZO/EGZ3XXE3uzlPFeeovG/B/8dzHCVBq0Tv8ak2bawzHSYmGtUlX8t+
ngdWIAmKpShaA+9SIilMg6sdGZNhy8EMeN8eULCG3kjw/RBUbZa4wUdSpB2TggEu
pKIeim3AwC86TWxfMaIFChvHyc039xXiMMLEjd0CDL7Vx5NTEfjbvIoyvfKwL2UT
m/WDMFktnZDhHwFR5G78kuPj5DjyPQHXJCr1QiF158wY0PxfP7pg4lxlUQ4i7fzX
4KCnSmnUocPA4ElwL54KvP8n8+eOb1eEdq3iSCFclpV7gHcjkLhGByyKPPszAZtk
iLsNd4qyVrKg2TVcdvLW8BkgMaA3ab/TZoyH8cTDOxDAcx2iXK+5WoaqKCCmerXh
GwftQq3tEBQ7dP9339VArQ2AYwvsjc+vwCB1+rrBGQW00iMDq9CbNoZ8LbPxIYyu
HynL+olZOhUIi4ieRxyXbPN0tCth2hv9xBHgrGdBvsFd50aSaKzpTOLz6sFSOY84
P7Faa/vAd0kbUNm6hSCcRMv7UC/qSxQCR8rrKB8rKy+0DCBVFlVrHWOP80bwAPPR
Zs65xpCbhEn0J9j90yEa93wGwE3mV+QFjYbfJaBdEBWu6KMNvlqqDR3zOrDpMght
bPRbsTg60v4vSb14obvWKyisnJYOEarR/gJGI7O0V493QX10vls/bqdWC/JsF+eB
0smXZEZ7vdc11lmMBWYvJM4xK1wBKpEopcJEGd5b8psg4dz3yBwuvTfW1pBnS2PH
h2m/HQu3ywACdlNeM1kH0dNX/DtQ71d/zoWoGC++RSbvWn3KHpKLiEqcLCZBBZNE
0s11mzQc76p2b6cTyje9TukW+4Y4f8HAzYnXqKWqL6/XSiKu9gS/gLKfjYBa4Jbl
23rugefVO+ZOIHyQI6Uej9ZOpfokeaOm4MiU3AYPb9D06fLs9JebXiO0RE08JAA4
DkshqOYHlUWAoXRXtNN7LoJfdn5eEAsxchNE4+zuAeOnQSl0wICxFDOvR8n05KGL
4SnJTpYelNeE/rFBMM86cPD5pezdEoaYJ6GBKmosJb65wtdLCl9IEWscG8FFHriF
coiUPTcET6E+tQa3ZX8yaEFlux3wCxihmxD45LNHOSuBj7GO9eAK9IKDD0NlhYSC
+l4nfKTaBiSS3cmhCfKmF41t0N62mKd/Z2zZ7YchmM6RIPNExkVJZ68iz4MoQ/Dt
mOmrx6CZtc5jPg3Eu8KlloxN0yRi458QUZS3wGLZQJIHPoniJl+2kFaKOfNyEjOn
NinaYD3GntduJ+NLmGhye2CKJq6JEzAYlQev4G49Wfm5WJiLTE/U451rf+moXy2Z
EOEhWm2yyxOKI1bd0GeGRrWotg62roU0HIM1FBYkEWPHzepl1scDzaYT5R0HY4wt
xfRZZn+wAmAJeme0YPUwlBoOonFpnhD6xGAJjExTwqZzBwjPZOalQ0TgBgwmSqRX
lB0+62NdUEUzvpLdnKLDhuwgE4q3LqeIpGW/Zm4RIPWm6DWGXQ+h5xDF0drQbn+4
adt5bVnJwJDHZPGbNSe9EsAn/dSN1QbJhkiUfwcPDJC/ahAg8bth81uirbc2d4Zh
Wxhqhm2GfdKSTsoZoLUcuzkDr6QIr1ATqxLxgA6KYXRMHo10SL3jNsqplGhAlB1W
LYZIKa5GrwZeZBzuFrV4Fj2DX3HlfoRHhgeklCv+54JjB8qu+rdJcFod1xBwEfUA
wXnTW/YCj+DEV7qjolGlJpypkCNiZuGJNOJgfpEJzDZxemGhGxdfyyAY0qTpkO+0
a6CWJeSoowBdl9iQm/xAknOy5Y9cxUmdJoC0p36AeAFFv0ugYxkVEk9h4f5ADZ4r
zIMFrBGyHW8cq5v3DVYGX58Pzyi6XSdRQ1E9vhwbdSlyXvZx0Gc6FhRBSKtP+lwB
i5fBZIdn7Pww8ufxNk/N+NfghGOgHil0SmkgmA2BU8om1qMHfR7OaaAXRGMc3COL
OQmgjeregES7LMnH+tOJ2SL8/J3emkT1RqCQv9n1odyGj+utfkAub0xjSQZOsXS3
Xuk3Jz7875Yx6jEo6lcN0YoR5lSjMSZ7C/9ZX2nxWx9UwWuvXut4PKsDCk8n2SaG
yT52BxLrMfC7f2LADWlawoebRhq1ZAFR9ZpS8k/mgyxcVYn5ZfIOHd1gOQgq/IFI
sJ1cC5sHeVjQHRlx8pkvmqQOjglXvgKuker+xtP3qO9d+t94W7OavUce4U+LMx+7
791xDwRDzgp8msclLO0fgKFn+SnhUf5x7a3KfnUxOEcXRGcwL1HDdv638qF5mn/V
iF0qfmaHXPIafEDYUuECnV+WzUXBedm/g8uuPb2bZaWXKfXsQOiSpNJr9AqF8XPb
pt4uMoej/WFqwWl8T0qU6lt18fTRGIexJt6ezRaXicrzdkET2qcxx/hohePXrJh4
dmROAhxbWC86IVbnwjM1Man4tqk3Y81Qj36CJbwC2o+SG6Oz4BYFXWi/ytySfp9t
tMn9KQv75aP+a8TYIR4nQioB+shPMl84TTe51iLuTogGLMKnvhzKJmdDqQss7S5k
6c6fWDrO5069GeybpLGJWgCl9spZjrybFfO4qE/da0Mu7JZxfw2VMnbhgZF49zna
8A2e58eUHnWe7AIJwUzoQ88xv6wHqs8sHmypabX9c4tYhNVy2Aub5wfQ5J/h94VU
k4lkPZEBeceL5idvDdMiRavBzhQPogR+tU29f4wO+TJ8Scwg9LhZ2f1hpYNdWWQH
VxeN9gxqLtFOFAvaRJ3+bDgXZj+BwxNU9A8z8rqs54MPGkZKRdroFzuBNuuOVUCb
2lEGRdaHbVh756EZbb6b5VYdy5OKecwQC9iFql6AFRjfdOGgQSEJTi61D7QTsuy5
1MwPj5uakM4DJlowH1BUmy1J8JFMNgqhapv8UvWmHyiApTn4KTXcQX38X59iiJl0
JY1pOkiRMCj4A7p+rGGwaNBbh+0/HI5M+doZIewiJ2mUZuOaEWdZIbraxdzkdwXx
mJEMTQtmetq57KJSEV3cncNjfeoh3fkmD8/l36ljXXVU13+J5Wxbdvggzvqv6UKq
/qFEOQRd1avOMOzsbIsjcgy7hHBjoj1eh90WhCXVBqujGSvoaMzDbZ7G3a/Ndm7r
rJZ0ujSZztzozB+8cEtiRb1iEJO6MQjXQrvZwr7HDmCjbm5r5K4CdYGeQ89Ex6CK
MHlloP4DiJdVB80+C+valgM1GxPNGw/oJ6KbE/bwT18pv5u2zwOj/fZXKVXuEkqd
f80MPEbmrDvbX6RwlpboKTYlE7+f7kvFv7fZgE0Wg/numMs8Y+EtLRKiJ3CGee2l
rklFcT3GpKC0CK1rm8Vcu7a3q4u0zS/Lg9m/ni2/es3x81ZyjOAI7eoE3GkPfR+7
xAP93WZ1M4+/vh2NwXY5ur1dudO1ExDoPbKYpDxIaQoFAJuMzv8rYQ6bc7OvEx9O
9Rs8UVktgpbT07gAJe/NTj36nA0ikg5XUyLDKJQs2v/dgyPR0m8cgRWk+H+eCwKf
A0sb2Q5X3eczJTiaaswSIWvBHMxKHfEfQ/cI2urgEqIhX8uXYUE3d4rbRUefkLzq
wnzY1ZDeDCOtKjNQBgy8zM7mVdrbSyDFYzPFjXvStUf7mt8aKzuUQloXImUATARi
DGhBPzqDkHW8GGnG7naDaZuw5B2IDELYZuAXs+DcMHqU58c0rZcdMZao3TOFsA0l
J7J19UhemM22LOZjLXLTppqlWrjDPnMKbZ0IEM0frtGwMp2l6g8BK1P0JZTdKLf7
0vLcwsLSRiuZWfL7ch+kr2uOkM1mXvIDFeysQIhs+whN3Tl+CtFK5h4Y1L3SAUtt
8kd6eCVX0BaJiXqZCHV8uzflLUWz9OGxZSjhGpHO/IAWDU3UFWvnSekVFMtn8maX
UYHgKrtnjB+R39d0hJg89tAuhUKY35HXtIv4gL1yJtZJ5SjFitYQ/Tle0S9r4Bn+
WFkVWV9rNtQnphdiNRC2BLVv8zQ9tXJB4BoIyE72OXAgmu8YRfqULqccjynDBSIk
5eR5quZ2S4xvF2ZOoutVe+LWmkGuRcLUAOrkyqLzlU66L1z1h/hkQiUwbbYn07Nk
ZAWveSVUkhdrEoHn/cNab/Ggu5LWJMFefQ91qozNmtw/smHDcLfgQpwIkbG7ACa/
i3XAmNsWYmovm1/FEsrfk+OqroqQx0s22aRFJpYlrdqyl7KCfwb2aCrGeJVwiRtM
Jo17j/9U7UOi9+B/ZOBV0T+TJAwB0LCp+PSAYQ/jYOm8tdCZCpJ63jGwjyTU29LR
LxeS1ITk7K6vQ9qKzNMk7gYKgtAQ8elj6uj3RPlKPP9kUUlYY/YV+fByGQgWvOEl
WPm5MR5H1i34AM6Oh/IlAE/rblZgzfmyROl4jyNgRqsGhF2YRud2lC/lFu+dJesA
cmy/FRin14M8UGnfYmZTZOBeaGPBcWuQgSm500B0BaTl249MuXly3VlmSy4Dpvkc
iW9l20AYTbhp8h1B7HZrTg2U+O5UDPcdUSSIUFl7URHJe7BEvWTafCle4ucMN7xu
R5QZ8Hd/Og7cGm+QzM2na9gUcBSjN81gWL4+0oXVifmBHZHJIGxuFDrUH3M55OcU
ytTafHc+tfE9xfRTBAHMHglurvm8r809QiKIMR/3j/OympnomCnk7v1Wqtu7K0jA
F3hPKtI2wzn0L8vLumh4nPllIHF02UlabqF1vR9WfIAPwoWUCINoJbBfJS3r2an9
3Xq2Ind84LLwMPV/KxbT5XcomC669/R/i7TjZjncBrBFf3EBP1ehokOG9BlIDJjw
jJo89m1guvKJwGCopO5HSmwmfWaiDHZwfnAWam19an5m/qDcDSGOdsOBjDcoV59t
3fIzauVR3NfPRZMtRSNqPtFQSPuF1K/l8018cW04oj3N+v26RtwuA/O9B4mDbCx8
sCXBV5L/eU+KHq96GngyK5OnBkGWvXIQbhblSBYdl8tGxEykoT0koD6wdrzOp+f5
CZP9k6uW6FFSy8M1ZuuP5q8EnuQPYSnxbX84BO0SsSBxuDQkp6SZhyIjVpb4x6XC
Wtx4u0duX8n7FocLm7/XtrgEs64RzWuXuZKwxx0PAf7d34v/E6jiAM7shzT4FVH0
aeCshsuBFPyCTykVZ+hKIjW0DQEeMRkBFs2qEDsHpyZ2jtRL97+6G8lUQ30Z9FF7
UEIeLftZkc6OnYGPWCBRU59pveDTeYR+damQeOJxHNfVbpvFhm2EqyV1a/Sb8xHk
aCG+tPEBL/zPcB6i296clT1gtF5RKK1qdNbCeln8/f8RhXg61p0cQrRB0YD6xpF3
f3eO6dBN12j9b1hWqJv6UG62a26G36FoZGZD+mN4hVzPwdxWy8mWZhZ71Uf9B7i0
aY1xIv/p+OHQMQ4go2yjI0fh+cX2ocp9vlk0Eknf8z52Zc3V7ji9ztvnjQSvQyia
IybbQ57V7/Js3aIyibRy59qqlxTxu+zW5z1GMwOZ0ZELPApaf3HK7opAy5N4ROIy
w6vZ8cDcxJr0ipbinT0mGrMP0o8SUz23QnUbww5QJCRjyTxakNbSmup5rnNDp07Q
HsC5Cpbi6BJGwX/r2X1pMuBqH0p8MDw5Wr3DfPnhoUDW9DwmXxVMkidHC8QT1Y0B
8slL1/BrPhJND9ZGJ7ISsktnxh4VyqK+9QQ9Y3AtjZa8sfweBE++mCRJiuR0EjgF
YOKY/2YxtxYayC63adImduz6NE94HP/xIC85vMVp/TK4QYtqStzo5KNDMaJBhS6D
ZqwmwhKQv+l63GJWEV1Xad9bHuWfxnmsZzqBgsdshG38FL1vTfvJWzXt/oc8cprU
5Swb3wtgDL1jtjlukQNr92r5bvlvb2A2IyLSNkxOBCHofwZT7C+0t2rNNs1o/xIC
hWYZq2Hl9KdthCpQkRhTa2LTEWpxWGoil9glAc79q4sbWGozrHYnjelCr0uNtVwY
KCS0/otipRIubxNHk2LG5du9jUGgqsPbDY7UzPCwUJh30hLq8PyIKiJ8iy/ghDYB
o8HzkIdK6a/QXrt6mb7QQqzSKlPsvHWndAx1BsdCRD8wZFEmr79u7OHklMU3/Eo9
LvKwDyjBG1zMoTxjBPTj0MfqDtGLmkiPYO9PFlGV4+19r4XvlllJhMzm6MpdAaO9
Y+08lJ/4hj8OUUAzIoe42/1BGBZosHBc0C32sDrH1eHMExFydH5PjWrYKyQfil7R
a2rvzKqN8xnBDtetSXV25H8znBH8CZI/ZohOFF0TKzbnOTIBD3IjHYQMgbJ346mI
t5FNxhVkXUT96T7ObrYBxM0K+f6WwG7qNPwzZ3WLrVzOVs2fv8xuRC61UPL5EdNW
0KgMvTxc6s5xe3PDt295Z8kKFf353gXq419ArkW0VeQ6PtH38r85cvTiB2Zufmz+
FKmk10sDIQI/8hexVEhj2bLPOOVGmmFL0SuNvsQlVtKWMU/ZXojynvUEMVyFMTX+
1jOlqzb1Ag7hekzBLmOxdNVUVAkVCX5QXD8HUcd3i0DLSMQPYxDuqIllxld5nhSL
5UNW0nOWwqDPt5AIa/imHZtpb334YH6eoCRT4IFMMI8LiD1kaYlLfnh6lkkdt3ZA
ByC+KzEKnGlctiIMck1n3LTOni5anZkb4rOanGx1pU6Fg66wg5ZDpWLbbN4/Rzfv
O4iaAiCR68cKdhiiUikoDJz0okM0lpc1PVsvNYzliCA7nZKVXoZRFvCNxJuKDLUW
tt+A0t9FskhCFrjwLXLTm/7MYOjFrpK6nW57Za6i0LrBDx5GcENNCDFxKhiM4EcK
gLs8ThMzFMayYY72RtyH3+3xpINn1pOurZmwWMdxG8xNm6cwUmecAMwAGvxpFjJC
`protect END_PROTECTED