-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
C9wIUuMaXKQsCfi3gxvxTkxl4m57WnumcpZETKqzPn0TAlpRwUZDZns4Prq61kSw
D1dNUR7oM2+OaRI7L09sw7IWLPMV+nWLmp91Kw32858NziXv776H3sECikX/UQJQ
zV2WwI5U2CPb/UXHwtP6YXV2T7d1pmW/YnfWxRlE2heZv4iS3XHLqQ==
--pragma protect end_key_block
--pragma protect digest_block
IFX96W+fDxhI80I38X5N86x1/ns=
--pragma protect end_digest_block
--pragma protect data_block
rqobFief3LR5wqlwPjswWGddEYcdETV//La3aqm92GbB8hsDl8TSLCwNzDzI+y/o
y7bkLRtLq2D3mqQCKF7w/iab/yP5wQ/ZyOiRwBFZwwLYaX/TbalAKN6LPZUzlv8H
2IlADuDIUPSdZc4NPnmmSlovGwM7DyPW2OoenkLyDhpN+O5JOFkLUGrMgYw08m4K
4O9YlzPvXqHXICnTawHCJHM4w0et5H+VGeDci1YcirWllpIABrUAG4hOhAxWEKBF
MD2fInRm88DjYdeOr3tzW4ZMwka1QqxA/OuAaMzg0DqsKoggxgSSenMJcGPpezVs
/iZD1MK+AMDCcL91XtkPpDfGQU85S038GeG8H9YTaaXUaq+/rCcEAbXbDZjQBf7a
eVNBfdRRtUcexSnjKeZ/NnND5f1HPMWFvOJesUrFWdIQhH+qs6gc9R6ISUjGDx2e
dDtDLx9CZtkr9hjFvNMVfB+XIlAKrQR19AI/g7y88HQcTxxwofYE30hRbLx08r48
lQ263bjWgfq3redWhOj5KAJ+aFAmZrHIThe337UctIBDG0IL3qbfB9ySvWDuXTEa
YkBmfYeRb8h6jmg72EvSg+VM8V668Z3Ec8+4XEch5y+gK4OUB0kK/3y8Eu0ZUmaH
yRubhuiSS97/x70/7LF9ZMLl6KryaEnTTi7hWcgc2SKvQ1SzIR26c803Mg/2zxg8
eOUSkx1XtiOQe2jtpivFwxKFJpxYW4CV+JP3CszjDL2WpT0Il2eUxb/8sY5PdKmZ
jNUMt2Ioj/FnFQIcwHyU8kp5vkzeuZHP1Poh1RCf7+ayFDu53EwUIX9Ej6z4Iv20
O7qedY9D3i2z1AAPuFKSn26Y1ATTkAhHl42yROLSDYgE9ET8XlO1BDHG4OUwoYIe
nAyOUQI3KQFn2y36uVu1M6Y+RgM/Ioatf44ZNFSwWbpjk3AJ7Mn/InE9v+k5TbYl
MMdajdJJ/3bykgSgXr3WAOEiFawkA6yW18eunT3Ew5VzxLJj73E3xOO4F2ZwNWOF
51hi2RCehSi3h/XMP3RcY1eENOF33AOax/mdbs52UKf1daE9By/06TLF10MsbdiG
wcNHZO27PcfLj/EX8V2m49kcGE6tjvx2oy9uupZpqGhHAhcxay/IdGPEeqmO0Pdx
Oh25h6SCG84dmpOa/IRFnj1gf+w2vVHb+E/A5yh6UWr5tFuiM8ds0rEGX9ffVcgz
51H8wHAg2TiW68kYKB1S0FUD53uTjtGr3Jc6dwMpqpnz9ApG5wQQ8jmis1XE5wkL
oFkucYWPvENG+R31aSdeqB4+JfAhPUC49NCpdidbrWYt4LxdSOj0VqPSpKqDPTLl
281AawbUIaAC2pwC38Y3eq8v30KtmVNzj0+Cr+AaZm6MvMzLoOoDo682hWM2aQcM
XXhu+K2YwPRs5LGRiYFBpPkUm6cRRaXd6/kmUU44tx15eEe0L0qFNbtTOKt8ZISf
g2Hs43soNZh+vz9aAMOZ7zrWpSom9mFRFahjnPAC6nvVh3xTVJdo82mia7ePELo3
Agqvv9KGA2iRJIvHH8gHV89WBlb8GuRuh2GwiqUyPMJ6Xc9Wri4BGqLaIzrTez1+
1KXdnh+0sFXelTy2jc1KeOxgIYqW0MvI009e8diTj8K18mMbKQth1c8GAmeKRuHY
YV679v7+Et7mpY2iUC5UbWYTYDMcsKC2+Fsuc7Qsvi6DSil/r+zCJEnRuI6MPeTB
jQejSPmoq5Uy9QZLo9SkyCK8gzclh6rHi7ljcHPf5MgT9p9Z0q4a5vpBEUEAmH0a
t8UErggBlLxYK7HAX5/mRcIi7wSAd6j/VKe5/misEWeJQ6zNK/fd2tkyCY3kURA9
9f+XIlR/e4ZxzuS3YoknEGXagfiB9tWyUp2dqq+awsMGAPxDR7Zvn91MEZWEO+PS
7I2uv2toT1z/Rd85aO3OddzY+e2wQZsI7lJs8xO+wBP7A/1lhPfxVI2THdLq9Uzx
/y54pBTdinQuVWX/9EvyGecMMokA9akmRcS1T4SABPZvBOCLkPFPWc6LXKu8Z0Nu
/RpW7vkZL6aKohWF/ASo4+IZxmlCooVTlYpBHdL60rq0iqaY5bM1Z+yf8Cbi+KZB
PMwEd3jRaWREGTI9dKuZJdeog6FFBF77DkOamcbD7DCDA+INmT8x0aU7B2hxKws8
DX0JS6NUpChhRHBqAPlECf2NN/pvZx9kxGMParP2u9Wy9qVsg85HYopOhK4AyDia
wR/WPS+SRmfH4eRNgaN7cOnAEi8y5xdAt8XOgTXUEMKl0iVrDy/uMMVsSnleeLay
0bfoD7pcnkIEZJR1K4nVcnuhSGnCg+Yi+WYpFyJYbgsWSlRAYBJiJObu3FrfIHS5
eGb1qw80DvrsGm/uM8/MZ+5jyJie7xUxa+Ai4hS+9tTiGAj6BTkTjq1ztlN6KvYK
8QgjEjb/n9dBIwrDDeu30v88ctP987lg/6A9Qm79uVcoZk3TtAiJSi366HQS6A3O
+LqJQa28Ogyx0HOaUXCcnlxGXsfye8axiVYBGeE8Kg+lV020b4CERxqsuUQVTFnZ
FvNWSVa83vja5TWT4l/RBus+F37UvJKYv2U3xW5mH7WX3c1h3UZKwBoJZdiA8Icd
zKDJbmNSlDW5ogrrxKuog3bBNHLHdN0nqam4w42uMCfszKUk0pZOA6vg9GYV3evk
C4J8P80xqMB9O74kHANvZeLWaPicg3i7/YimtqQA0+pXdLqrB0hE7u+qeheXQGbg
PFkEsSPnscDbiN0u/bpMQl7fnjKfQJVEpDksJeULaLXZ87tLTfn9WXT5d6QPTIuh
FU11xVhbusBRoP/rw4Domg3IGKLlkbPDqC1srXlKmMzCIVR8C2NKrgIw8D8lrlhY
f/TMye3Vp/hLRD4JpxB7jK+leCcKaqKjRKEg4A0Q3RqwFzgAcBrYhQOwYJfx0X3r
bl2lMm2RTOS33JoVx0bq0+bgAOrvqa7Ys1c20JPbROdqKsy28N8nOf4HUknAgR+u
OOgEcDXgn/VwotAqyix1XbN0OJBxhfKJGG+G0pVQiok1MOeaixQIZnLQXbn813v9
TL6S6AcYTn1yAHMJYwwMjsvz7ZHpP5bmIQiiddEDXm+vNnWa93zEZpQyZdDfbRwo
Vm59aDWoSdVqkY3MefBvJF+sXRvEHfV9XAWX/GaSrHx96t9NZlQqbYQZE0sBqbhT
gXc80idgr3DXrdwou1N+4WaV5/FSEHYQtR2ze0ulEcm7O3DGn91ExSmv58ZZHgpK
NaSEOXSbYPEsTXaLI5Q0Zxww/zwRG8Mnlx6gxvlqqQh18Ggeh96mrO8nQJk1Dpif
nwWoaAjw6sDdOtMOOAYENHw0UEqQOmMYuEyaaJg1S9pOuFpOoR0iBKsJlckHNs/1
Y6JVyqllMWt66Qa8K2gDWxaAgW6DZx4QAP2yCSkSrI4WFr/0ad1LL+QIPIlgLmPs
+aSIjJ9KXnhQgv5dyMVasrwHROpKXCMWrk1SPky1AQ7rxbA+zLG4+JQR/pOVVdhI
ttbXXm5Pgw5GXY7BB/GgYQvRniVBAKN9fYDDVW2v5ECuEaaDoYFtfe4w81bsRd7H
qzRtR97MQbNaUgUHRFgvwcycDi0d3He0diC/bUf/VeF6bOT9vkyJlD46RHfApKiw
6XmJfwYUkmsN4/UukZTfGLhSjgwOdV7RlIIT55QrbadaeZo3H+Hffs//QKR/Ofhh
kBph6rP4WWsSmoJrGj6z+2B3WbgfvuKBipadQxMC/YAJej++QrK6oziDNLeswiXN
mpRweq4+RESnddbOMJgftUETqVERYm83TLtRGwOkKb9lHu5TCWXYjpO/ezbY9r1w
NDqMafuXjrOOOVzT4oX0RsvO0CJkURSO+eOv++LbH6zKM0Aht4R9NagHdsUbyblb
GCb+CzMcwjuh/yitqF2j64Du4wTknIf2O6jYsq1QzPF3tXTL8iGjF5A5eU+8jRf8
5R/I7H2QNmy6aetQiHgrqjFnFCWQDfj4HF6XEPZrHaA/sulXtM8WpQphbv/HBDEf
RLxFad5UieErEY5ng3SGWhkjyK+OFfeGy7UgzgQLIQkHkTDzqjmKyb+37SObmu1k
yf/TIJG2ovCsZuNsMVBPlx9BYWoR4+FaKwx12MsJs2+6vAp0ffzf4eswZyZv/gvf
BJseF7aj+JBHgYgFavJH0cpGSOGBfz3Ky0AmHik4FwZg15ThQya1ALS9D453g6UI
feWQFdSWAPQE0xXu/3Adeq1/Vk7DrZREKgRDuoG5UlRzOKRs1CuT2CmZIeSh1v+G
5rpqdh9hGVEuh6VdToYpM7nVOrXw7U5IizEA46a7fPY/PJVFdXF8fbtMfpukOmQl
vSrwuqXXoATyz0QzBkeQJ6d/2KyR5WK6Gb2MmylKWpPeRQ3xPOj379A74YSNXdt3
Tyne7xO5XlruDLP/VMRSHhkpglQabOgswp/vvB6DQ5jcU5Mmo6pru9qfLONuDjvN
GcoUe00RQ85gllKeOkAh8KSQKPO1HREJRZlLmK5gDReOx4QfVtU72jNoVO3wV1Rl
taPmeCr3jaTG1i5yrw1EtSTXvrLFEP4SuzEK5NY4I1p0aDNAaPwwVGxWc0z91oez
k+34Ep0ldPqnRTaWsp7d4GqrZsfD5x2qv76IMUtgdrD9CPXMGFcRfinhpt+J16Dm
BsL4PDMZpL3/zJjM027HtLiDfTHwzBsKVlkwcdyx8uS8I6WIT0sXiyAE4a32bxrx
K7aAy+sIPjkDiMpuUyMtXKVVY7q967yHiWfdx/CNNMkGqB+oSlfUodm2X+Tn5uTp
+ixBWIuIlSeeLcQSkLWnDz0CnpnSaNGCNZOeDghX3yCKfzNv+LxgRkNTBk3UxoHa
b6pWUkOsgXgpZ2LaVNS56Vm1dAcg95oraBaN4yRK72wsZvyNWVz5k2h4PI87w9gp
X2Hk0JMH1GgfpieqS9NfYXnSN1PW0lFTXA9/rd6FQbq3THlkW+5CrOag9L5/8zLL
dgljQ6rBLwKRodAYsvLxUFDg8nOyLAp6waD/Vjf2hSrfOJgmg4zOau2fcHVrKosU
sWXKOb4fDxRY1P+fDDCs8jmiIwZVHVquEwhzRI5prpafNgQ5YRWEckXE/oCTog5J
fBRe3RQ4COVgnemQnSs5p3rR4JIKsbt4emENS0kWYEFYklQmaKAlrCSr1MV2hEsC
tIt81/b0UW+RvY5B3iHQqI7/f7vggLXBLQFmlyg/vX45Iw3CSRZtTOrUy2ZjHe2a
y3g98BDHiNLCpiAvrzuFlhesYKGArCgU5BuhvKsqliLPyhTf8uu7bHcHtC8JIsBy
YBitsHXA6/8ifdN2YTdDvwbFekvDXxjNkwzTchFQzmVqLEjS+tHK2Tp/m/GkDUJz
heMX9wO/aW2ecc9JzRkaza7kUj0FuF3rXM4/iubVG6nTRUw5+Bffu0W0CYws7omw
SMowesTuYSs1l47PW6M6oYyrlWB5xk2Da/HQSOzFlD+2+CdSFf7KNUhYA+Q62teO
UenDhWah8LCq+9gihfAftpm/lQh6xpolNwFRaMRmCp/sEZ8h+L9JBEQfT4HvDWWn
QbkB+sxDf13cIOX4JWx2FQdhh3eyaG3JOHFvcPYsdm1I92hw1RmK51MVHmDewrAC
lKiLaKmcFHJW7KCUSob3TnLvA36yBzBUDs5jlUuQbMOjYDnH1E7e7UNCGf0TjcJL
cj+nzMcvhGSyTrstgKz2gOAiy5ev7RoFjPHnUALHR1oONyP4ScvdSOQt5LdNEZHz
W7JiOfhC/UBAtI/Xsa17a/Ln7n3Eud6bj1tqhN5cD6Y7UCUQSczZayCa4W4kSrLQ
x4YLlpRcTPg7mC+q/8VCvnVFp4OYclABQ2F2Iq/YgDHChM/9WAade7tP3Fs3p4z9
RjD2gOTzGQuMjO3Ud6OtdSLjAHPnuVlH4VIEgqjMXMkVrYpUcd+E2nXrXu3rkR3x
phbUfnvDaxNVMBsOwR6+3OLjyEGDhVEdthe6VI6l6OcCfV6sPEhHUnGgWq4zwSkF
Dc1fTbCW1o0c2AsPxCLndnpiaQJGbLDLDaPfigbKYpYySUHOTKlAxQujZAxHeYGi
QIvdwrKsgJxUXczflu8uU7LaJ5Zun8ygO+qROA4LxO5VNRhcYxAyPhgTw+ql+Zkg
Ks30Ds26pL9CmHw9K628vsDsslbzwauVYHkUP6Pq3tX9VZ3srSiTwhiv1T43kBGl
f3eg46SJI0fUvCSE3tLJ+Ck71F9pSbO2RVYjKtDKD/MuCjru/prZMLOF6yIRriv7
7uQVb9rq+KWEQxy+q1ywyGRTm7yyIgf/mG05xLBNDN0dvw3RunxfMuERffaiFiP8
zERzr4U/Kak3HWxbIt0KI5kHj/jENGZMGvW4HuI34vF5MwAaDILe8CJDzcPZYXDY
K4AjmHeAKKq6LI97H/0HnYMLE5AulsFHGlXw/WSTGhd1087Zu7yzbIS6b7HpJ6Va
GfKkiz1XRoY8svIExQgubO9gy/kLfclCUk7UlTm5kwQpIP/1oEp/b1x01prwgQ5m
nsn4TaaHOhlbyb35Gj0ju519C/dfJJftf0we/0nqdJLKTjQe5gatmJyfz+iyTsL2
uWxfsHAScto0A8kkdylm4Wg5PdtAwV95I3BGmqZdina2HjfJClxYCPMr9akEytWv
GyyF72wedV8IGs5gGgBdE8LfXPsj7vsJHpEus3swBOtIKUHlqiut2bEvQLTqlXtN
+liGvWy0VO3OtVTc/C+7tprngrWX/H59nLo7J08ajwtDy190z4atLZJS03GWr2iS
w6k/Nyj2v+sgA5+qiBEEp//MMRizrdUvr38fUp4a3yc3ArkSsnXQRtmN6dRrr6gh
4faHPtuwOT5YuI0npphrC+On8wBJP1Kq6xfEyYZBbvDRJpDIont5oP0jekzWjWdw
c8iy6YM1HoTa4iNYw9MCOFFtRYGTBP5ytj47TVgEcjOwDPvyx5xbO852q81pVwWC
G9GcgKZSovmfZUzkkZbZ0+qfwLMIznYYKWME5pXHatDR81NLKxFQ4YeZgyakYt0G
rlSbUk/5CRtFgV2SAOKyexOPuENkAYUdAmofafOADIZyep2XFOPmHGrqG0xd7H9+
wfVX3RDZvsB/BY5eXXvOVMwEQaOo2frCVieV7jk60VOVK3uSJ0wPf2vy9PAwW+fw
7N2kyJNjXpEZXJxnQ5Ou7w3Ma/i2anF1fkFyXsN2u4h4QlYFGRMPYlWeQtPjHmSn
n3xY6ClBUnmhHnrRaMuRJ2n8prDeEdaqXzY5dunitsHIFXlKoM0Yb37HvNkhhauR
rDO5Q/6rr0qTXS89UlNU550sM4bvr+2z00v5Zg+i1YRT6EnW+AM+AzwwaYLTi9vN
GbjpUT5QgpyVWQ3teIsHzrWSJmvRDCUMLgppZSKGp/4DOKTvQ3oBvlUNkuc5Qwc8
9lWRPty4LyHx+ZZDFx3vY2XaU7sg6UZg3d73aHDOjG174pvMu17jWFf83ZiWXzkR
8rbYQLSw0zOKdFNkofDu7NrOuoIMtmLwPNVjz5T2x887rCX13fidx5+mJDEQb8sE
BEOX5t1t5WNgCjjXUoFAhcraZbKz4Kxv8eqfoZAg4bSNDFBMxu2wn9pN89Wu7daW
oestLFetiq/1BIlUbZyaxnKGRIOnljAHKt/qSJbljOa4okbfxz7QQqElEKB8yL9x
Zl7dKqs2FLVVcm/sVMq96+d5ch1s5aeeT8yeQaDC68BXQL2xz6xpB93Osrb10uxd
usR4SG5OXj6laQiC+XFowhUdEa91Q+VRatjHwUxBE2ejrdj/sCOAx1jjmANdi2yx
IDWmpL6owrhGWAH7CYHb7P2WP916aY6hIyZTrOThZlg2jT0MFzAtkR1S7Hxds7aN
OhcXmLt9UIqwowMUnecMOk8/ytm41ABkWUzceIPK90qgKc4Xb4nDDoq8ZDPdMH6B
xRvw60KMYaY5oSfqQhWngDnJZTHsE9LnYuQtL7Ou8mYxdVwjYEOIC/3XH6viD9AH
tHgmXXTGkAyrf2cIQKsabCM9w7/oz6qLa6xPANGj0dziXyLOFpA5pcvvJcHvO+Yl
74YEjwhi9NuZzxf3BNi/u49nkApo2XwL8VzHsTynwGSzcKXWI9DZM9jcLtMfqcGm
YVbEPoFPM7RpNTDPwAeLr1R02JFO68bHjThnKp3MqUPry1DH9FHILDffg/wvK4E8
a6ETAsqUhmMtJ8msMwZlc7Is7nOAQf/sdXx7olSeH9wtcP6qrt7bZyb4pxn1JQmw
VVprzlEwvgrg7P4ieXiggonL7d0tUz+cDaqu1v7l3hNN/9wEXzJMWg8IL4I0cxiI
ptNnKcMs8/IrJSD6lszsVPfS80KyvDwXOeGaFX8S36H+bnPi0ogJ6Z65nAX4Clia
lnE8FG++iytzh89nmX+L9qsLhW6vp0MeFi3bMX3oKDhvIOdRAprT0yVteoDo9IDD
mmDBm1YuRP12krzV243bJVZEstIKvxlQcDoEvpwkgiGNfDw+j8k9e05+Tkw/LvyT
PaG+vnuM8MzWA1USsZ50kJa/tY4PVhCbgeecryw10neMAyd0W69aSXpb0iFlUNIu
VI5MCH+shAA/xSWMdLujP1ZArqMLrLHA6HAcgO4bKKEKsyURXPl+a8I6ixqibt2r
OTOOBz+FBlK1CiicXRVlyUI7Ldy3Suy1jrEboOA7T5K4SF3Etkhw0SCooOrcZR4f
VLWMlrGA1+xzwARENhtoNX2dgODu3sUvv73g7fuMEou94T/NiP+OOpX+beh8Lfpd
XbtDDPWKo3wRZZPhLZ6KlV6+KJeAyxbLxF8HM7Usu22mPanBZt7/dccOG5ofwaxe
ZJwgPWEupmqtoHRIBJMeYqJp2zZWhaL+zMlWJWyDUmP1LPvnizcgAc7rk+ZDpAoV
ycRAMpORnbGPCXc4xiLJrC9GjuSLhaZZ0IFD88L9eMc0G3m+MCB2ppeyHfFm4Es6
maWPGvo9Td+aJCg0gr82uOhM/YVj0e3KlmwF1Eq0sEMS7zFgdIjxvoglf5Pejd8r
Tuaa8svBa0avVWLYCxh2iGzl29k/lLci9saYyNhghtLv5uYkdwCT1nSw5bacoOe7
IuodBghrwcYiNkFQcR0IH1sToGX0uSBvXZb/xP/jXvGbthfSl3wxufZGLQd2S2oJ
OuxreRktWRLVAFjac9zbOpHqdxPMxkKHczYSsgUzE1x/Y5/2S2c8Q8axktAoL8L+
FsOiGLLwq2YAoUT787vLADO05e83y5D8K9PgFRkIi6k64/yCLNqvvnd89O9YziyF
nJVMXePWZVRPFa+zCpy+akxk3L6GaEgE1hOXlcTvRiGsqdCC9uAdUa4phc4rUOGd
dIlgu70H6440uLdhlF+TkS+ZjXsEZezMuGbpMjudYNBpnd50gYGKPtIBZ2TMxAM+
qIDFQBGeMBu4RnmXc3sbVRmwTiHkVU0rPk9arguxQNnxhZctrAIGpmljy3yQ6GGF
88+7naZdyImQ++ONg2gfPqe3k2BSjBDtzOdEKQCEdUVMwLbvWCktXpZRoacaktbd
kCho+ttfa6Um/x+cUtqlSvSDsReAFFWfnApIaChoDkARRbWWRw7tut3i09Cuirrr
NyW2wsNrZna/8ANQWc3GfEfqglRH5Vl7Ow5IQk8NAqRYtM/eyhnKafDHGAIcF9S+
qyYcyULGrU0IX42YmIYwhnokymOZQfSATWJfmQD7mor3z2aDdDWh5RvHs4GzjVf3
//BKQJSSO/uwsXCzOUQLAWpkkUtobhPBMd9TR3dWbQ/4VCDg/xb9ngaaTxswvZVf
F869a2GA3BOEPp5ShOILeUsRk/3cqQVJd4KU7h9JxHMApV3XeHjASSyZlNMddRkI
lUl+YUuyf+apAWkXePf1eNdgyYmj9Zv26Ug2HYYnUElfCw8sB4IxDLkXQ7U/V/Rf
214NcmzDaVMVhP4a2TPPHh6zOatMl5QLmW9mHl7/Uyqj4bXYQzu+ZQTIJiEffs4R
W8KuAhY7xYkGm8zM2IXrj7hUFjL9P7xku31TJXIk4C+K5Mk4URoD3rPlnBbaoDlF
qDOJxaQaOloHM8LKeuXmRf3qObbDHsve6JsvOKuPhyzjkzCdL3MNhSPLnq0Br7Ft
DfCvR2abxpSnZk8uGrbOHC4wh08zDcP0+1hDiOe1/jFP3CnL8pSF+gLc6jKaW6Il
e6XRFGZiaoARzoqZi4nSY3x6srCSMdRFZpbCv6gyMvu5ohNoCEWd2FAruvlBnZ4+
pyN9UKNsB5CKtfe9V6iYLaazwkzXpclU2JVA/j2nOmtnbriAQNvC6D5RMZ39AXog
lLRasibaOCgT9YXXSNP9xJzuQ7e39rPOhnxpKtvaZgVNzL12c8dQhYG69v6JVy61
ygL59ZmcwlyXy30R57DlxxcrLDxZkPJdc8VnExp1dPZxJVv5IArKVIMn14cyuW7y
IrlorO9UN/xAHqmwfDf0TRKgVWCwn/MRpn4cu+hsPI5SuUcPoNQ3NgyV1jbg3MHg
M5CnGVgZaQkHaIxycYr7EVi09DlE5dqL5VeGQLboPB3AZ9pYZ9iXB4SjXUEOppKd
DHAMInW7bNhRrm1CuhJKoYFQfN+QByX01lkStcOdsOsPAoudCRef2NwUYKKejIQI
oAJzZrcR+TldqBigQes5GcohLTUYm127mY71+hgJG3eCtVTuX1TW3E74M4SsoZKO
CUx1DKx3PdV5LRgcypqD/HGNR2l+ffJEEnjUS1KLKVdttQuKzscUPNXjC9IR+6TC
FoclzuDlf/bQjP6s/M8gvG7oiBNQDk1ThERjV6L3DmRFFM/OahTfBmcD6pBcm/uk
7fSpGfXVA+SkUl8rD8yaNO9e+YtyB+dYDcEG2mik1Jvqgf+YDzFP2SxidxEnQLp9
delMKuSkGO3jSJNGsDRLSf85LjcOln0VcP//0kiMrobj7o+Co45XuypxlIHbIvHJ
ac2D6vaF4Lni8jhQojzuLapw3ZgjpMYOd1xSquEy4nJ8mBcOzsAkEDX9vQy1CIrA
nLZWlrOAcb6O5zmNeXQVOSp/43QLh3zdG6sWY7/k5b0C6km+O5z4+8o63r+E0TzV
vQeRk0fZAPIbakFGFVuYlz2s3WAVnBbF4mjcXylhnglh2awZz6JygCeMQrGLfNB5
O2lvt5DdYCqeK0awMYqe/dbexYrqLHP7Vn2aNk7kt66It/nVwRwfFA5p5Sn4DIpM
6l0ZrZPwRrA1/3wh/c/hnacYOjo3qCH6KIC1bbjOPDROZkLKF5rcMPXI6oiTHfOT
7LsNoI3ifQqegdU3XeWMzlS3olqXIp2c3deVn9iwgvCQU4yBX3h4EZapXSDblTTE
U2WNVW0WP34Ug6dmooiN6Vl9GYJ30lT83XfGl53BIu49t3m8Xw43jXmUzHKk7z+5
pFguEtc2kcc3PvGnTrsaFEgTyQhPfSNdoINynULuFo8caf7AP/W+lJf3yQmPbMDP
m56cRAKcaNeF86HknmBm5MqX3uYbOeNaeps9E6RZAy9/+8GsnrKX7KD2HUTV9Jsm
cjHIjD+OaC2K7ioWVwBblY+NGzd3QGiiUSZz7eDaWxHV4rCY1AL6LregvOXHnmXv
Qm8AMErHgnrlWw/O/qJaTf40q9p/hcCQ0j9QJWtNgyKcBijBaUkDr9AHZZ1/+yXe
q85gsK3TTXnYWAwQmhL7c4M3U9VPp90igC7SiDcH93fLQm3Au6lPMh5Ll2sODkHw
NRMm8ij8XBpPwla3UXnd6eCetCsjXW9oG1B8KcabimuwOLz6RhBbh+kAuXiC6dSG
noE7D4xY+aNLoQ+C1njhrXZ9L3fZyNRoBX9XLs2PsHDnRDqq0mp34wLaVUQZ4dsE
ZV0Yr4OV7VJLzhuTgdh5sM9FFeKR33OCs/R+L5QtpC/SLH7uaZx7nqIaB6sk1EgS
/fnbE/4PqkzZaO9s8wGPdgzP713YfgJFzY6dLmzLTzMRKYQcoZy2XtXNubsyPvij
lS5tJqeJ9K4y7VJrSw+6Rl4hwuOvZaV+g4lSdSR3jAIWEZffR5NqjYlW3Kr0U4zs
BJtt1aIvj9SZjPJasMTh7XI6iRRsXLfuOACFedCUQyaPtdWodGHIgtXSb2aqc7uG
syVkYfxxvJsZOufkTKBh3rXaBnnrmTo6Q9g1EtMCBXMIsDNjLut4HRV1+WxOy6lj
9oa77lP7uTvFRFLhcnCQVnCToK6ETsGn8DF8FenrP5qjNCmfq7M+y8ZW3kSEXMju
cH+/1qvMmRLa4n3aMJZd+72Uf//AzW43zY2kWgfzOuglINKiN/IhoDKQQuUUXKkY
XaoBJP18uSjSofrrED5mBAgpasMfRmXz6IcSPC2jsDELKlkM14r4JHiq6NbpETwp
aser61+Lg2zTqTQfPsOCKZRte/xnoecLwZ4XdM24B3naqgRkqWCD8ramCheEL1b3
UIke1DAQ8SSVcp9RPA0APnvMEKToqFNrpHsCWLQr8pqLAkIQb0GGTlYn3eDWCAn6
c28LwtTgobRGdtKGfalduTkqZsaleOQTVNdW28QtOdVJ10IlOxwFBXiAfU/WS4r5
t6tf5VOOEFVHIYOkKNvzfxmDQMqGHVvrFay3aqonDKZyh4ewctO6StJAIcxpn29b
WE3oGUL8EXyq1Dy09c03Sxllty+WusRQbZFOe5wSwl0V0kig/VJIwsBLJEyNQ4hf
vRxlBI3qk8C+YeFub/pzycoZXBU5juMF7+Dbp3rzIe31HGq2z3e1qEgnRGH/5Lkp
vN3kt8U0ALp761iihggrKFdgYNLyWWOs87+ztPSMaxf0kKIv1RuS4Xfv2+XOKZJq
7ZZLvK7uUKc8nTtYqeY98xhYqWvkY92cvOkxT1QLtirYc9Kqn7LR2u+WPMJ1EGUe
RYD8v4LTrStabYD4ySYFsVo2FWQgpKCCXU+PFUL7LNgbW5HY8h5SYmY9FR8xIOD7
ToEMsT6BCjGxtMT8eeHTQ67wgRgb3aju7n+IzK1iKhnMQ2+yngQTQP0ECP7KT+Ak
/CV3bUfeZU0VFpxzzaNkjZuShTRiVFJplQPodtZYxS9ycAIGFMOr+8vdmrcgJ/11
P9eqFoqcvqujEf4WEAmk+PE0LhnpE2o1Pw7UQlJUYHmMXOYTLq9hD84Tha1UxoUN
a/VnbXqBCOpnDA1KL9t4hQhEJ13yhPXwB4L5eBssqD43E9PPH482dZACsTi+xaAi
xgSoj6GyaXJ1RXyvrwwZxOfdDTiOeeGvfLlcq/uiXfXQKnZ2JfzNPSC2dOt+5XgW
LgRuaQbbjegGEME8hT8rsdloqPkTIXbmSOfY/G7b+CMUj9YloATPr7I/EBF2uLSD
4Bfi3ErB+3IN9I4g2+1T4/7VCkI23BIvjRTrpGC+DQD1DAMt4x0YH1WEtQ1PWQZC
Z8OWs5ij3MgmR7XyiiIX14EZcQW6rAVjaYWLqbLrnruuDUUBWUjVEAqGHBRWVg8s
24weKDk5sP2/ttBKpc2OXiaOnCvPURgVTv8+xMhPA+Ym9OkNubVLPkjDCU3GryKK
tYEfiqgNiCL+DMVYsnyqUimLGWzEf8c4z2bQYZinV3EPqbl+wIpXyN1O5gXpi6Hk
OmwHWFvadsSHAvWj1NIRv/1xCWSCuSmZr7R0kxRSc2pi4yjoJgdMt2OVMGCsg89d
QEw/obJu0j8QWGEpZSNjtjEDfptzZPEQEXaIsFKgqFe4fVDGXakXclSX0o3wy3UP
WsF6tTzoLtRkHBns21AVqVGSo2SOvmlC/C4WQOJKHRttuRCaUDRNafmFi1YPWUk/
a0oR7rKdjPwAfBIxg557R9H6SmK5XR3+3YkWBRgP6C8k7m8HMUTUMzD4W8TB/QCW
GrokGndTji+DwYD1bCf9C98OWItJPRV73AowNQRaL5506M2DpzrxmVsPxqiirgEl
XR2KE7sVF2AiyioSg54Qdtze5O8P8Wbem4iSuDt1uHTpyaDqtTzR2Dcs4bGF9KAr
tgrSy0awlKIsQN9XWALN+CAgcNbsMQaPpueKCY1p1tjLHDO+i+4uDpoJ3ZC/26p/
yMpoNGZSo/vZ9fedMFMvMVm6NOAJchQ6SgGcJBHuzfMXxBjEQ1ivWzWChyLykG/G
u6Ljqusr6sM9X/qwlgETTA9z2rhAO4Budefwaxj6QuSBWCKexUX1DtQHZW+xUjWd
kg3/vK0ykQ7129g4pC/DmxhSji1dxluf4+AGnOj8gjGX/Usu1dVnuCcikiWl8/9A
HsmUqDXwYo4dXC3X1OQM/lG3ebezZpadDtngJLco6iLMk8mvduoJMsVlD35gWfFY
RbQOZgpdxlWSk9NWq50ACaAKB5goKNtXDBXQkE3+1W8i9eFYglOjiYCtbLYtu/TT
R81MY1fFfPeVOHYd0hL51GCba874ATZKfmvzH1350UxmuYq0mtfqGJNQ0hLin2qC
mjk1KBk2MqVJUPpme/WZ/b7r62XCAh1yZIoQfIoqJ/PT0p0n3CZG7MK9I6ReE7fc
yI+APSKAI5HFipS4h47kE7JczaTwBlqBN66qC9XP5trvEO8FftzNq2J9Ds7oSF47
NuGa0xKGAk+H5L3BLZzsEG15m4nSv1yHf0YRoFeEwNW7FpPOuv1P/10rECCvWiqU
m5BniLJBZ9XZYvoOohZ5d7gGQhkb6Ag8EJgM7fWPktD3xmDK+LWhBclcxgivsd4U
/3DForMfZwTSyhYDu0Gfhc4s5Uha9S10UaSATUYOzA8fMn3uXTFZHlDyO69RE7+k
ZItRcleV3KRurvAkUNznpPYh+C6Mdl3Qt3kKS1IIvW2H20tP1Zc0c+B2z0PIb3p8
pPaNceaHlU24ac/Xj9ecE7k08lzh19/vk24rq2NLhIEIwqdvTS3GL0QC6eChPRJc
Z8EXK1l2XamJ20ya2XuvjR9+rJdcsOpDqdvxhag5+I9cNJ0t4f/LTDa7fzouKZwG
Oem0y8s9wMjBo4XEDIIygUdj2lxmI8VuVdRqLVcogWYICzx885d6cAEg+cE2XUPz
bF8y008l7S3300BWOzJaCsHSpUXzsxS/+b4rJqSyVfJR67+ajmMn3mrvFViu3NLS
YRHc13SGzkHrYul6674ZQ/JnxqoSL41gaytkHOZrBvA0d5pHK4PqPF5AVSxk62zt
3FOJfL/8Y3v4YBjIttLwObYoav3jOz8j1QVVP60axQbOGjPHy58cvKv4/K9wESmi
Pzn1LpmaNMTD7UlCPf/B0u8q/lmJUeyQNwFbMLI5B92tj3p/JAD65Z21w/SwQTew
ktTQF5yYEjK8k/rrl6Yu3/MBu2zIlubI+QLFwlFRoei1F+HQzzF5mk91gI8ukCk5
+5MjkJRJAh6W1yM/IfQyXBQFTKdEWhxbWWAD+N3ku0RhzTJ58fSbOefgiN620DSo
IS8eF3oEkKCI2yJZXtjfmgs8neLqDzs0F0taB7TaL1ikknhaqEdJcnr8O5m7JblF
b0QrAKqCOB9S3rnTo0M5efIelMS2MKclg1y12wwWumr3gQ2AYE0pPdqqFZlWOi7E
4jHkxVhEJY/hR+8GwUVUku0UBE9IRh8hWQcSzkwvYF4W1IU1nS4fXxbpocltLIbY
T1B7Nrlta7xWbkVQo/36PCT+STwi7Msi6RktOUDB3tQiTG9o8vuzCbQYO6XveMS0
PkVTKQge5UzkenPWJquz1ohCZrVyw8OpMSkEruXIfgl2144XgWon0gRq6YdahSIB
07uCPF0yU4aKkil2Arn87I6PxJiY113a+wEan/AqrbMiyUoCc94FBAPXsTAEhyQI
rOd+OMjKkjVB53QZMFXJQJMxy/AmAFXrF0P+gmDY8BBciPF73DcC26+gN/Eiq/BJ
SoBmmlrM2kV/J/7H5OsaSBM/UugwlS4tECeAOGUuVH6CamDqe39dgnATRROtqRr0
T690cLpEOLq5sJ41/V7e8iVPrrbO3v6V5XP4ZvMeWkrT9AZs7gm/jugRBSXo51Cm
uNb1wi8k5xb9M1pFOiwkyvWHxe1MI1xMi1mA8M3DGWqQt7pRUvHmuRtGLY/8LgzL
bpnMH0xRe9PR0p45hcHLclLVxK9E8zbpetFq61D2L+a0v0TXFvpoMM/fdjaWVcLt
WiX2540U1DheqzPCj+SXQiATd4iV2ZjQ8R4ZoyqOa7oT8k3b8RfljPvqlA8ciZuz
/zdsVW/zPFF764aCD0lP2x7zSb1meV2Yp7lydWUQhE9eJCSwyvMwnDEyYbT7+4bR
wl8FqiTW6JtBudQ0g/4LboEy0UEpTuvx/l1oTnzmsQb9E/O5ezVA0S04jHgfs1Ng
3VOsBqKawIyutAcRg7kZ3zko+uG7MVWp4OlyltPA+HCt+ycblfiOlf6eLHmnjTE2
oUAPHx5abYSy6Rq3mf2Y/WEw0F8nayRXIqoTUsj9LA5yGlkZyR4200YWDqc14UNg
gtM1c2ekoiJORFV6JUOyo/LfAnfUvSQKr4wcEXfZoONvHN776MBYw0AVu1xq32A4
pBN2Jy31LYpP1Sn7H4lc1AOPDFZ+0C0Jviy0TzAtMONZq6QDDqMUMLwXHPS9v7JT
h59nkDhNIxCrW1lVVne/Y8dTojVtAqWKz3CF4NK+NtEl42u+BilG+WEUeVEcLOSh
rLvbePWdfn9HLM3AiU39IOegVTxrc9szKluL+gc7XBdIJTZt3MXHupjOxADcPvuu
4sQthIxV4RYgf2LyXCLRN5y+xC5G+T4V6U8f7JTzocaIX003T+cBAhd2p/bdkOac
KzR5T2yMA/vFKMyMwbmxNaix2TOh4xP53gMGsvPK09tSN8xT3vAXo2cYJrsm8cto
Il/N3B6im1Ob+4ipODkxnkCnVkC93enPoDEOhZE4uogl1z0pEcrFabxCDdiqmweU
vBOc6Q0991fKksFmZUOVMK9glgQTjNp/n+MANEAKCpeZCnNMRigPVLpSgMppifRn
klViHdCqGXvRU/05yPjdmzqID+/Xa0vZ2S1McA6lNWJtu/l+YK5G+H/lW7DuE3jM
O0iqJhx7plCixh6nMXLTItw/gnhUq5AALDVOFU7442BoMIaIyakyR40+aXg5XLaU
uW60czdt0yujpFw0aslsvsZGMgJ4N/3cAUXfw4qj0au8aXq2XC47YjlGCEcTozYf
5rRw7x8cj0aQgMJVdbcA8tNKKxsB5G6ieWOEurtDOqoBICe+gD1lEzBaFXPl5lTX
u23hjebIdqR6CC+YUwt38jr1J3nsDnd9dQd+QOO4OUSLADsHWI4XmsPsNiKd4pNT
9S3j9fTRW45BToKNn+ebefLfJW/TfEvH7gfVTxjMnn8WO9fSAsOnSo/knIHYZ9W0
VIy89fMdC6nhHSsJNGpVDTeTqCeh4Vctrg0p413PCGmAHhsnM9/Fp8HS6fUaIEmC
vqHgFWo2xLfrbXhbxssE3fsBkrQV03PYyN7TaZkKbggcPjbed2mvrzTsVWoBjlbf
+3miN4CMdt1UdpA3aPCLRc1No/IRXx7o1a+aYXhpVhq3Xzc/9J8SlNSCNjXNGfCV
jt/kGxIdAyFvLubKuze+WiBM+PV/hHwFWrhZDZWF9Xe7yaRjnybFnlh0Mskd9yEN
LdoQscO4rBlZJ5l4daYQ3SXA9oArImDVKPxS6Iq/bUtFgGJtG2C2MsS0HgzvsWhA
4ouYXbygEmt02AZZqRmnPa87SBC+Hm4uUOpCxuQA+or6V/ywd35ThiInvH59BPuJ
FrGlA7mor38Qb0vcz8In4nu8PW/6+EXW16LkILZLf9uwH4iVg6QYd6drRWXpYSR5
y2BAPudQ56MqTGJc0+Tgn39tGUYbFHY6r9rboUs2q5sGzZ28O35p1J/ze3mvaeXE
PjHvMpAbhLMIGj9/XiHG2Q0KNphmbrwBY/K/XTnXTZZwfQ+6ULgQaMvTcsdLpcGN
H48rGymNl9EQgFUyxz8EsJ81DGDwuATyPBIW+5LfhPMoD7gvRY/jm7N8ASG5hmbn
XWBEb/fkSF5yj3uXT86X6x0iQxPcHeXtWSTEoNm0wuKMF8oigoXyFMTizdnyxHwL
lYqkkioGoKabVBlZq8zrzuhPsqa7VsQCVeWI4TlAcf7kucCmNN1haSnCnMB9xJ+9
lmKHfRrOfxFNBpspLtuJyrP7j3sqKf4ONn42AxKcsOHrZukWXz4pWUVmgIdRlVxu
fX7DCmFowRegRx6csdwMcTh2rXskwlNpXeQyAsTn2fitQWcxqKzuyjBL9sZPVwo4
ooF3wkr6b5dN80/ByGuyP619GRBKPtiLBG/iwZxvMDyyI/urn2tMpSdMZMjS+x9O
wD9oCB6ovwa/qOhheqwntQ+mwT2n2CPGcXNJmnHqvv6mh7u17ZzE0w9WI8QDmsAz
NTpxHgkGf3tTRzZgIphyBQz1G/5ul800TOIqX16F1jN4kjnnaF5VPPhZ0uOMqDHf
W+6l/myCZtmFLi6gKRT8U656Uu+8vrSZ06uDD4rk6zhelTyXgvKWjJaU202Cs8j5
iqEzyobRqhv50hz/EjTSEGuEzxZZlE756m9SBiaYEikKdPAe5CfP/huMPKi3RZ2Y
gWkz4XhQJwk42sy3AzrbcGYEq9VR3ehHK8sjJR/GUMYnJQi9A50mS/WDXv525SEX
IiIxPjukDfT5QhXLWODopuVVaNXCyNyuZjbO3WM9AzrusENzTLzFSTjYsMGC1faP
eSpjUgfsPMNNj+mz2Qqe6FuN6bjaMoKOxsg9rBWvVDZ9YJmMguI32Bsg1wu0vbvK
bZ0pZzRpN6yefLFOi1KkWqAAaQYeaUQzotyoqBMGJB931pVyZntQctZJ/istdpv7
0iVrZ/QeVdft6blEquA3xYF2FyTO4UgdKlsQ5NCLwYeTAmQL3zliZlauQ4PJtcCy
smmwwZKPnTMhx01kb5RlWSzQxNyIFPA3k5SD2RG7xC1NUPS5kIJn1nKP2wDK/yCp
WmF9PWY3OZcFVSbhyS05Uh2Pdst6vAcbka2vkcyM7HDKNVPLmecU4InmsB5MFMlV
RqPqwGDNAkBNJnx1Dja2SSMtoUrJ34BsuyAl/pk4tMxwJBW7cKNPTTtSwIDOYEhP
bdh2+hYYRHNXEyW58351tPj9wjvArGdESvZDd7su/CHaVxiRSMaY/rywRXWfH3Bm
l/RLSfPuvp++utXP+AgxtcQ3SsbEtQcUAQTcS92T9rsZ3bEXSBpYr9/0SuXMB7pF
/bcgUbgM4TJk/yPw6ixDIIroHsN+gH4Xjp4Yoigke57QL6zyMkms98cIjangEY9A
e4H51gdZoqh/m48nfC7s6UwI2NjSacpCLjatkSX167WmXD5mCWaUzsG2lMUls+A/
VVGF7I+9HXsaDYfH32E/qiPO0CXhBW4n9DIwoRaCDjhZk7mQKiS+SS01p8aOIaLV
woIYyEgfnRrRAuFmXzDs8andIX9WzvCUsyCfnVYGdaNzkdAvZ9m+w04nXZ9dpghE
xtpSqf2CwZeZFOKsbKMf8nBu9BJMKSRiwcCvnQ8NQ6b4eMIWnEFSQczgSI+06PEk
kPhyzmOIhC8xgS2m6rVuogDOkN+VwXUrIBwI4RPoLGv6RB/0ZKXj2LT3Bq243LQq
y/sivnlf+zKhml69J3IZH5oGVCRbd4GBJOIXbknqrtS5Fu/cx/ouI2S6oWxN+HW/
d3WvxDMThNj9Ldu5yytIHogIFZDjLH+CJRG/K7a/pUxxxKaJTXUIvBkZ+5/4UUaX
VtUpdtZj+7teiB6eONCAfSgz6gszmlQIY8na5tf7jf5d5i1el7KMmWZTYMJ4J2h5
E6X9AihjTNKSCJbH3zHGWTZ3yMgfsmn9HOD9Akep/HLUZruT4jmkq9zdjiXyFR65
EkHdfFcLqm3cVhvBH7eyojPFr060rv/Rk5al2LfyV+sOJeltftXfwmPQQe5LMDDn
oDv0BYNHL402lSbZK8EguaMU4IJGvvcLS2iYcBYj3z5gJcDEvoZIvxsuZQtBBqcZ
zYhLFXxuOgCApUfYBA8ZTf5uNaatAbFKryip0RfzkJZMy6u0OrMYugrW3DlcbLSl
M7hzo1Q1KpEruX1uKSUr3vhGHy0oBQQmIBwNxiB0Q7T9zny4wdl7ggH8l59bJctF
tEiGtUwWPwv6N4e1mGhQnb8EQvoj8GDSor+naD9r8Y3qt5aGxNW0kIVRjRnYTPbF
snxl9eeMl3k+h+FY6/WwlAkSDktKjw8IBvd+2O15NMBmHam1PUhXhJhT9uWhGcjO
qCOOU8EhOagwZ4sIX6MmwW2kngRWiiWp65ym1uNwoekCMHtoYV2KM/WcW+sWa+Sc
H8jdrhpc7il1OBI7sA/wEEAekNhA1GQisjY5gUSutkFhUi8fEJwmc4qzVyspP/9B
VBCgOgzf7MKdke7ecuqIw4/6w59r6DVFwQ2R1/cJz7psf2xeNt2glEISKv/nyM3f
rELT32ThkuJeC1O9y9oNO4Peyv++wtacvpsMTNBf9oRpL1EacWFQ/pjYp6zt1YE8
ZoNUqzWXkNKYuWxj3jmWvZzvFYUyqsZROWp3Z06ZI5VRxNyUJHY0KJuMRqHkNSPZ
90EqTux3orwCdanH+fOsUL/IHeoSjxVPr5eHHDfqkpOwGqqpEOo9VXV26Alt9TGr
6Y92OLkE2bBcbwxVi2mkHhyg+e6Tk1Io3Env8Q1DCPgOWZerzGMFCW7jKTgRh9K6
ccJjrnORA9DN03ePT0gNhaOIsluWgPRnsYWJ/yy6XH+189veJset9+ag1WIcxWcs
Lpwnl5yy4/YCr2GNwpbI57dYggjCnWCc9KICZOLdsb84OwF7GtSYfphzg/kzRgUh
oAGMCz3JgUGKQaruYs4bspPUk/Else3dL0Uo/gRQVHiz/GDA4/DoUOZKmVZP2/gy
w4XhfICbQsyjkh7zdNGlJTLTHsTKo2dZpoHebdsW443NbRtgoOoBv866bJyt1EMw
CUEGEZCHpG7nO61H201z+iNYyZ8/mcQ4+OJuRy+2eGcnwegytbdKyLGW4CggNkZQ
u6cQtOK0tMHLYrEqbNOoeq+YVEzC32S7DPybmsP05Ahaq2kFnaeyVksOqPLobejz
GuosBI9h0oTjIJspxY975X5yQV51XhjHYt9sIl4d0qq8U1X39yGLeBq+eMoGeir8
PjjrkXMeAQzGPj6WhuOfNQ2nltg26G8tj7OI757sGcQyuFfO4/4YPRSpJoL7VspE
ZQaTkrVeOKVqEcIx+lDWF/1aTJ011TGkzq0Z8cwgAJkHHbMiDqI4ZVpK2foC5miS
l/crE5GEHftac2wyfVMsvQn3M2M/5VJZCMg3JM6rWNZ+aPWhC23k/X78cUmxKp/n
oL/xKqrrHGhjVKqwYYNBBKiOLI3zOFr8yGbYR6W3hZUjHNaAgpzVF6VPz8jUPZsE
DPpgxziR4rm4uGVZZfMv6TSM0JoQt5bXCyy1RhCHELAHDW9olsDxueLb/zM0YSv2
oVNXfg3CxzDAuCDpVf9HoX5Emi/gqfqndNmQvjk5hqAuxTgnHxx3dlPpIPO36xSO
JCoE9O1HSBJ5DSxTA0hcYCLN1rjAHa0fGF5x97GfaZbUoCSXFK10oQ3nM8qkxsJ0
gO3NBQnX9x2DO/Q0f7htZ8XPuSrov/XYsIf4NP8lxpuOYOzRRiuLsl4efpsIEG3B
JNWUeOaS45XNz/weE2bCT6R+axqNhExuq1p+BObUy6HsYpb8TzFXNa9jVod/DW4p
s3/xJ3xZ/Kr1PXLkRSXKY5FETITZR9/AZ97QRx3E6eHh6z7nKBthcWpBSRWZ3KrA
Ky9Sy8zvEl4ug31g8poEoVtA/doEfv9jgrU8WexTYOqANsVxttNAnuszm9+TFsq1
EEoK74AAd17PcSHH2rPwz5/tbHj4aV5caZO9CoROifFX+Rx4rMxfTprY1vKRaAau
IiBNVmBHbsjQa640ClhIcjvsSyXsqqFHW+QndvNnr6V/8LrFEpNjD5rxPG3WO3HI
DyROeEcHSGOwsW8Sr3i8GpNOth4cO7tyWVEw1Z0Vh5qpcFYaIdvSWUSnEIidu7tl
BNKWE0O0Y+3yU6zWPzTNYFEaSsyvqe+lCfaVrWoTwiDuAzoRfInlk9ndjA/yGWzA
wVHgGwO294Ed24C6bqZF0f9KMfI4f4O7HCHzw19iopKg5ZW++K1yBm+DcpE3gCqG
FLB+x2350aupEMvU4JthfekoVnt/7FDAwzWXQSid7V7anh38EcB2bIsv3BXYWNjG
CLBv40IUbwWxiJ5bjkMvsWkCF1kFOT7D6dG9dHgOKhRlm0gXYJ/zn3uVAvqFNGPn
OFlwGA8i8Dd6rBwPN11olrunAxiRvwYPC8B3LkDTxL54n4gN8gNkr1H3NHZH3a/a
VHKa2yzWL/HMzPts55RVoUjoFfORSC9j1DFNnQhxi3qxOn3Mg13dUGDpxzTa0Ilb
mw4whO3euv5oqTzm6HVRljPeD4W3I64LNrLKhgcaPItTHBl9w4u47w4mScUokYIS
aESKybB8wuXcd7IQMbXKU2TQKtQ48U1v8lV85KPbvQOlAVc6UQnvpz7/+MCgVE1H
n66v3ALOpcA6hOabj0UGVjVkaUANljkQc2hQ4I/0ojTRs5s6FD8FR4++Qvgy5lf4
7WskeDFzxokv1+R06aVr7HksrWqi/pI1gHYlAr3qhtzB/LXq/rsLwWzksF8VTq/i
eqao/Rjm22Qv3WRsJ7BB3jZT0/VgL9zPOoZR+xCJWc/9RWtYusEk2fyTJJdMZzTj
dy4Hx7NS3RNG7jbYgYRagkHOrutM9Li1VJy6KuH4dIFwucrMCFQ5bRn/66vsMq+A
UJAQ6MoPNNviFqlMACO/qIqGafFF/Z7JvfSkRlCiQ63xPXjLf4M9Kmd0sEqOO47Q
N4SG6Noh8dq3XZCh4nkrl3CoXm3Gm7Pj1QuhOuScU0nWfDBei0H8pou+NPzbpoMA
LpXuv6lO/FEmP3nNRUzKhDTKNLdr1SVPdMZUuAGIQAbCCTqohY2tvFmcZBJE1cGT
JEJrAKKkDM7rgXP0XUoJ7EZjYoAM4UC5JxZjjbIK4CGSCBJcfIkG1AwgGaToVxY6
BHnMETL1ubQnM5pZPezzJSYHHrmi/utivZRlndJgKABs+2nlHyLU+nHJ2OzzRkn8
PaD6flDNkTnn82gdwB8eH+US1NtQJw3PEivEJ7dFHb/G2JQTeBCoevAybMbvCHNH
UzYXK9/Mb9NuMDvSQ8vWO7RYwzhnfk57REg8zfUwboaXOBfmsVABhR5TWfw6xzvE
xtUbVIygWwA7VGTF+zdI3PTZ7jKFp8Y56an4LF9nwPgsMckZR6rmBAdiHhyWa9H3
JQfwNWPJ3thRK84BmEPaBDAAw2R6vgrDhs7m2MSbz/WRHFLZ9W4tzSK+BQ8Jp8y7
fNRzwb4tbB86/EChljzgP4vwW/pTD+PvSASaJGGT7q89+DaRhEgOpmExiOZZMHxb
c7gYv+3NnPRGSqDAtgqj62wlOEsWCO41V0FMfoMC7YyKZLWGqKK27hOmUWeB6jRM
16i1gwgpGnUfEBBoo28cdo66Wh42dZHLORHpTygj8oGygUx0EqGMz5dO2lvIT2eR
9Crv1ITmPYEMWHIMYEKAPQtXsPdmG+PmydP+4K+0yAuC10pC+d0JDYj9aYUUosiy
9/ACrf6yNWuM/6upL5mhBi6n6Y4seZobYn+uEWxCembLV1hMQtCUKdZfK/yCEfsS
GQoy6pJDN/2P29asb6Yco9co2hYzsvA3/qlZhaaWYU+WI+hVYmQLq/YNnm+DtPqC
25NusW/LPJJxlG1W6NXsiBPP1ea8M5AZPsDPRUnNGAfW+42816LV8qjiAbaY6hMj
4Mkv01LtZGB3gef/rFAws1bg37RMtMUbskZl4QAPA4UJ2QLYJBeXNd8FBx8taW9e
/PZruLLKFCiRlCTl6WIduhuoJ4UzV16YbBSpaa3SJOOm3VS2aN15DvRl23yX4oUp
q/DN4jl8qvxijZvs9Fw2WMr0JRVr0S/wqDCybqt9KRZJ2D1v8x06vByg8PuWgYUK
GjsP4ILWh7ly4bKznAhZfF4hUKl0irOJtlIlb0zWXDxLccU544UUEa1SZ6Lhv1+8
2cMJmkVCb2A9mMp5T/gUMOGBXmxCT6tqN35WaQafdfRSclF7gcrvMRuJNs7R3xKH
PQxTCijK6zj53egWwnirn8W2YPM+lguTf7RWTzVjcPwrlHjRbaNs2Ev+CG/2uqZ4
sx4ux2pH1/mlUkeoC6KvOcLcQdTqgY+GnXFTyy3qpysrn0tEsOZz6JDyc2f8c5BB
V70IKSwGjj+i930IMlkSf04u1+U6YtT7cG4nD+8xHx7balDTvZC5ViulsOGRiXPj
Dv+kj0jBTSTQEfmcxhFtue39rcesgwPnP9O3HAaAaNZrULJvC0WI8Lon+4d/r0eD
2IGQxcqFAIqEjC2i6LUBB1dgXQFBcSLq7LrwHIUphTrlHgr5sv1wuKoaM3O2/gd2
hst1yx7Luqh/1kADRPXzM77KWaBz1YudoZMgMYZ8iQJESsItEI5Vgcu77hd9T8pB
jUtbmdQee3EqQR/qC3Oq1Y8nLI+4gIRMXYkwdG7QLCQ7zoOGJXjHALXgLFTtxSJW
vWUfa1r0/MRwOOCiuiRWBrQq0bkxfg8rCHLTz1/5xVJMZE5Wy38rBPPBIZLAizIE
MGPTuhcW6l/c6A00X8lNg7VlZf3qgMItAwPQTn/YdY/hImBEi/43F6/fvvWBQVM8
m2uJAN1gTkhtHl1DJ0Y2jWHn6SVELrg428yIHbhO6qyCv21s4gc+DnqCNCZ8ERGd
vT2R2UsCwdxbk+IJLo0nU41govpEKxmV/UbrT5juuKWxd3EhRuVUkWQSBCIg4t0L
+0YtzSXOQhV/Zfql93j7flVQ5gqPWV61XRyzQlQD/C4C50JCKNonTsmJJCgguKaZ
gD9YGP5i0QA7dLHDnMep2TmHKhZb3npTi86LDAX+a87R6YK0cTKXW1cJd3OwyTOu
OX6PGhFnQtT3rHk7EmZ9ibsNsuF/g0E3h/vXya+O5EbhvpfcPP9rSFOKmRXCZcXv
+Ae2eTNi0j0s7uyI9soHGjzCEFbLfsXX/2mAUOGW2qaWi8YfDOu5XSMOcfCXS8B0
YVCXKMriN9s9ciIzbRWlKznV9EDx2EqPXmbc+uRQrUE4LtRW0AeUiJtkPFCNxZYQ
sK3IYiV1Mxnu5Z2pDAD9BmUNiDXg5cEeqToCYMSJ0j9D8udA9NYppeD+XOF0KBoO
XUpQjz58nrEiaD1BsdRHRyax+hUtqWe0bcekB3K+96UFiTB5BUk02LVhJU5xJo3f
y8sYBMCh/A4cE4qE9Qd4/QFj5jKUdKlhRqQC4RGXNIa296ehASFZrLiY+y7BNOxc
0oIjoRPBzJKrnoMTDm0RF18JbeMbScf8VvN1h94ADnhly2LRJPgNJTPA5CLihs5+
EqNPfsKk+TU1TgAv3byG33/IKJFsSgNAR0CK5AWztIJcta3KoYTd+OUC11WTVU5k
jd41JL+gAIZAELfpLk1ZK1HDTOAmeXPJkCz21L53A+blot+m7BTsz8mNRVhR85Cn
yQQtr3BUCjA71r7RSiCKGn0KowOxMNO7gdpTEbhV9fZhtVN857MFfRSXChd8x+MQ
Hah0vUzxAISqpyOTq9B810tMFmF8YlJh9iLxV1SbLKQNi7oLx03NlAITqGL28sJY
M4FIKh2nrjoS8owgSCDGYpw5xQxrMFYjnMaguwwj7D85+c78WH80OtMaRPFo61VV
VFQQIIJMKgcuSe01GNFKZATihigcrE8heX0Gh4Cs/N8X6tUTtR6fPcHD55ms9Iba
/mQV79TidRuCkmoONOjFRoB9ZXtBCcAv+G7LxibEh+goe5Wh0yF/hnHLj0DqG9M7
QMur1ta4ea5HIsVzOXORWXEGlEMXS+doKHFvN33w5yZbVOh/fC7npcu0H+U43izt
2qzpXPmLX7PStZPboYXyvlljkHcjg+kzXbqEQflkLmQq17VYqF205APlpwRkPsol
M2EMLo/kveE6EgMmB+0YKXeirzyd1/npQ9/HHyub0wlJvbYyZbNsV+Pmp8hXQ1Oy
7NpiDjbDqlg9Qm4FnkQSlL/2xmg+hndry/d+GDN8mQlJNZ4eoztaif/6EvijgXeg
lFGhnMS5RszXbOXBFTcZ9AC//SgyubVn8XFEn/L7Lxao2oR48Owkz+XzG2CYWg1e
I6YgOoNHSBUJ3tgYK+cP5cYG4dYUsF2ctZO2vB9RZbEedKzGkMuF7mPUZs8FAMUv
t4dYFWkyePskG8Sgzk/3DnW0gz235wQt+xHa1PA7FSrYAAb45Dz490jT2MRIAcFY
uvv/PQHUIxzINd3DYZF3r2DEe9zwPZORH4jqmEgahuH0yB/bytEGKFq+5UtnYJge
/3kEbxEBJGGc/LdxZE6pF21ZbxQ9RlFalfMcr+s1Ppq34pGChBCQckSfvA2qHrAJ
NKSb4CSGRl5kTuKe85IZkmbPCvsnFXePgfZAn08s1nCvFqVqfwr8xjDIKE6TQC+M
lNlqkqLZbE0FanyhwAWgaSrM3q0+AG2vfC7JAdgTZsHH9qA8JoFaPDmoOshpdKR8
hYozGdkbyobUgzA3rcQ11+jd46uCW/Glm+QLdCPddWVPvxmos6yX4r3JjZUG4vBW
Gqx08i37C2IOsHnxue64TBEt39JXeQ9wQrgnixFkAeCBkVkPqJ53gPA/zrd2gMi6
oXEphEqsuU6crwKrKrf+z/GyOyk7q/Yb+w5f8RCtpi0z2X2G4kGgPDJafiZjY3GO
WDVLPS0NmGZVYwoH8+RbzGGzA+pHpbYyNSNCB8mcSyeE+/3AQ1XIhcYjbaMMrJwI
/7kYEYtWjr8i/wRFWRC1ySXAosca0ypp+1E7wGzlojg90RMJTRz3WNq2V3OYgiiv
vfUKYLoFWMMDYwYt3KPU+Rc/HkMYSve4zTijBzKwuQiaFM5Htc7rPvBPl0gFAoPn
0+4sxBcr0DMXfuwLDz2UorKX2EDi+Rb7rrXfJc82paxl7c/0uSS6w+2G3ECJmkTo
bmKzPcGg6sT2VCoYj7dmAHmsZ+gZESYwv94lhg95tiwuSsK0S2Br/c2xlJ++/NYZ
82TSd8eajOvcrGhkNnf4Qv9gTWNU8SQA/2pVaBFJ8VVVGscRtCqjG+6DwzbGi2yy
jR8EpAcjmcs2EJ1JS7Z5idCIbwF6MozCC+HbbpZCrbziL6r4DlxKE0tMBb0npJZs
vOYhtf4kn77BcLEl0b+5EZ5zw5flHLloH0mYTvIjBtoKJAaKASqpWGsj+TcgSV6J
zsPvXbvXYrAKphmoU9ScUOy2dlGkmnfQa4aPu1qPISr+KufCK1ByQgWqIh59AS4m
sI1GeIUR78sz6KpSqYBfApOYJ/sxXuxsHFMRmYtwsTD6M69MbXqHGeYHBP8OJ0gk
SIZHvMA7k+L7Aa4oXs1lMQn9yPDPJp0OnZBxToaCvgy8zm2UrnGB3b8UEyXpYcGh
stgb/obT0e42OXRfLoNqSZPhfX2QUb7cokTejiyCNRqQAWEgavhCF6bu3nhneSob
fD9dISmX833MsUuHN9t5iyOI8P8efX5xVpHDo9T9FNEOsyks6YWEpdrFAGJvpv95
ND3luiXmJ9X0dHU+DQKFgPGJ2a4A6XPQ95TSeYpG4nuR3Qs9JvTI0ludkNgYKXhM
6sJ0apKkzb5yfriYnEssbu/HUmcHR0MVt5015lGxtL5PzBVb7oVsC2F4B8eqfMOi
9MSy58fzn87tm/RB2E9rGnU9i2i4W0Ui7t6BVFDmSf6jlBMsqoCy0jvCbMu1l3D+
jOkgaS122yTT0GvETO/ybQ8HSsyJq1AL8DF1HE/UflByB58mPpPgMtvHXqaa/Y9Y

--pragma protect end_data_block
--pragma protect digest_block
VuEEPUDjd2e9fz3gZggCQQQHp4I=
--pragma protect end_digest_block
--pragma protect end_protected
