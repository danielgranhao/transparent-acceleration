-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Nw1bnRnSUklBYzJWy+XY4d8aM3aj9BkGUGpi8CwuZsXQXO3PbRvVFnEr6/Ztmw54
nVD7VRU9Lp4rI/vGH65Oed2i/OCdZjitAYb1d0AhKWoEkYyYCZfQiOKPNCfSjurV
3VT41ncS+rly/J6yegEgzIYnkZ/KUlP3y4Y1mLqA6XNVeZ0Y0HpfUw==
--pragma protect end_key_block
--pragma protect digest_block
am9gxd8jsJ76Llk6RUBXLZSGn6c=
--pragma protect end_digest_block
--pragma protect data_block
xyt4rpi1iW2+r8wbHm0/H1m5GyXE3Uy0l0boujl2WPOeI6FgX2kIyPGGgMC/3HCA
iXTPRgyGY34W3vrclOrqk8fPpcSrHxuv0b37oqn+G0MlJ83zTcImWyc8I8ENaQxF
bfc/slmpf7XiMgf/4DErJ5BRZxxLgd9yixtOc9pRC+hRgGYsAahxguddK+T9xR8K
WDFPL1lchfNJPasX8l6Psd+70pbxnDu6NWB98Osa8uOF+HsfnHr+mrhlSAj+kz24
paoHA3WNnjufZoozIWLhlBgqE6zzPuv7Fis4cWh+1W/BDba/aWNjRBRwKoWeX5f4
htapdMQsNv/WuXz+a7ebnnv3s3cigIgPZe6CWrTZAEPEqOs16KfDqIMusko2VzwB
eznSoVlH296Mfyk/Xup+bOIOWnic/OsP7Ls6iIrKgj9s0jf+Dwud/9OOZJ9QdGA5
rUtfuCXWmqZTnfPLviX411egXy7yawnlT9TA+MEMfdnrrbk6lcgl2s+J3vmW5wIl
zkwj9GTgvR1fHFz7pufKupxLMgvlDvED9Ls9eCvM+9H2W0TVzPQH1gIj6bIjT6eb
F2VdWYV9OAisOrCELm9YByyPfXWbkjmBaesf3yOAHYr3P3LioiIgE3dTp2zYEEGI
v1dRAlS6DyzGf9u1m3i5kg2ubyTZxu67k8tvzHwlCtqs6IcVD9LoDVaWMOCkU1+B
VV45s57NQKHtukhtV2ylG480uZkYGWK06Lm4Hw/YoWKMhu0X3geDm/8iBAVhQDWF
Q3Z3ZSFwEuf4+7++uGNNKNt+tkAOBjwD8QQIJWSvpQnt6W1wsRcfSKk5vBZrv4cN
s8+gsiLJ6jtDRnwlGhJ5CDOxPeZaV2WMwll1N3YyUPd1X+huGklnlgWgzfEulhs1
Gealpr6aiHgnqNtSZLh6ELWJs52X2PJLUkiuUFwZDyEZD661RP6PpiWMJkfaeZ9g
Jk57n1p+GjU3g4bkKhyfH+ZSBD2xIRdX3flG6B8ONKCmSPSwgE5BE5gaBI2M6u7B
PpbamWyMiQ/M5rKNsDbHJQy1JvuA6G5s5cKq115AToFoA1wQ846SSqFM//yDJDva
hHCUcUnebWJX1v9YbIudrQl0WC9LNEvh6zCNaFG7XW55tdv1r5Mavb0m3bXACywe
v+Onu/0i05QKTUbJyw/PwxZqvXhmofM3Q2VPC7rOzwDInL9yQqPlg9TbOGVc5ECG
ZQjb+I5yrCYic2/6p7PsirlRGnAAsO5OFDOsFipHchP8iB88YiP88acvKrPYjbU/
nUMgJbLkpIZcjFrjBQYks97v0fMmKNHAz7ASeZuYPlXyE9d6XNKzwbv1LD35/1m1
EA/C4fs+VV1ngmZt2/wz3dFjrSxN4OigmjWaOXNg78p89zolElMIOQdM+wJkv6Wr
QU4suMEgPyMCs+7n/P0TuIKGAzVvwSHdBMAcsVOv72fiWxXKRycLkEnxPtWH3BxD
Tp7hQKdAk1asmloE61QnH/y/hy57pTCFIUNQjP0+OlyoOZpSQpLuZ7dWA+piS5Tf
wiyQtt0PDfF+N+wGdkkzYTaUbGVimY61mCGMKnB2WcCYWzcHyHux3ybADvqYZ0rb
9moYeBlSHLHkTRVDlWIJkQS4B7Bnu7OQfeCOgf1DrHWlwXivwkLYNrUpTKfhWxIo
evjp3MQFHPakZOW4/3giTOSH2zrJdaN/KLPhibrDqUBKHYnt39to795wKxd/GBPO
O8ISi8iF9Vv7BTpCmeaLO5EDN0BNgQMrpzjiyh3gh+cm3OUfszNLVWQMW0yaIc+o
CP5RbR2yGD815uoiqC4YxscRSVW+il16DjhmfnOT9EZnoyQiyLtHOfLdxQBd+/X5
z4ZpMxJX9R8FyszFJ+DOqN2BYggogVI3lDyzM+QxLnIUi/2nDF4BZOKHY3Ycl8/q
t8SuCfU/r4IfweLvSPOOCki/dY6kSnCHlqzIxLIdqYhTSWGEBQ2MtU6JinMw6xKc
w6jYnEAIgIB+rj/+eeZlz8B2aljCrWV+qdr+yjKVm9UipiUv56B5TBuPnmnNqwpj
WcMfD4JQVww+M3xCx7nSMlBg1wGtWubg49Ov1h1sWWY82Im4OX+kYP7JNjsyqEdW
sV37v8vU24FmBUHvBJAPl/9PvaRe2UdEElIJEih/64YZEBCZSBwaJJvVU/ZAtWef
l3u8y0PV8yMmx+ruoKERZZ9T5x+t8t0AsdY8s6JFMDGTqVPYw9buZZv6rWoIPfq/
103GNwwO1fZW5oA5TZa4Dx8OI1DD+eSXXt7SMfMGhV41XzA0C5/Heji5M5L7Y/Z1
wt7ohysZIatUwD4srjaT2lcZ+v18snQd34XdYYGJB52XkRjGFFf97BkfIi3sXXWr
lEf8Mtb2YQo/63cii6Yof7ulRGIVAtxfQx8lEIsgkA74ZGaE6im+Xp7iICXmMQhu
is8aJ5GuEUxd15kDGE3s0imQUCBiaBBUaA/MfIXR2Zis2aJG2TBHfGzik4TIf3Fe
3T+/s/5mvqSD72kUpHVCzVi7JDw+b42jck1lCchqlfafVB7+eC3XkkK6RZ5EqPmU
huJyXom5N924Nxn48mIvFawNja04mB+WirswimcYany1yIdQV9pIbR9BwYJuLR36
eAdYj3pEU8uqXsT2CPNRNXqiCFL8uWV7fNd/lrtEb2Dsnc7EFneTsaFmEC45980j
hFeQ1M0wYYD+xO4+ZfDG7a1CPoeVq+gy4gG/Gav00zxsfAwh/BDcVRqQV2CU3TV5
s/ePQAeB4kLxf3vyS9vLQ4/iavgV2Zi1/wUmoZSpsvFVj065YU0I5OLq9vlPOJN6
AgOcJBEfgjI/w+Z/yL1/KXwpOLqdxW9UMvM6G5ARRqXMwn8u9spT9A9hAkAGs5Wx
TIbOhyTwg9u+DjAgNcq+EvqG5N9EOsccKMaJir0YBqwcKzgeDwIpksaElI8+D2Jw
t9gl+5iQRbbnfnbbWLnivklHlcMWMzsrLoBUcPbdKlcYU0yEIjc/5mjo9QF/Kivw
jO957BXK/W/8hpc1mPno3T8AqI2cpItJo8jhnbrgHG/bcXxuYzmFPPX04F1PpXRd
0ieIhvW2AnTIZyx1l59ypFqW1MVrzRPBAISjmeWF4bW924scNhJKU5xbjMVyZvRA
CWMI6kthUpuKIDyxopbP9VRk0iNdsMSHkKL8zMAZrzUcfzeKM4ZN8frusOyhrXHY
kC9l2jqn9dhHyGVNGowbBD6X/5O8HPWaw6bjP8gS/nmWpku9cUBDeJieYHXccB6O
VbkclzJqkzrZoEa5NOosEGIpJ2d7h7SEMKO0V/R42Q2+FEVQOY7KX/Oy547OpRm1
dU37kUrJSQclSOunbqoimcM/iz3z4hzWiMkU7xu4LPFVvkc9S5Qc6vDeHmPr11vx
Ma/kdo5xf6SKKuZ5RSwb1hSnCd9QZPmQs02/Y65uT6DWBOdGGPr//pr9pWEuw5MO
txYNMhFY5uV7UQJ/9O1pWK7dN6RaEyNBKgJSJSOFMh8Nb4mx1e4XeIi4wLDnQnEf
v428OwG0K+eAlE+osZC4jV8luCRejL+81G7zvNtug2Ygqo3gZI9xCNhMRzGDVMOS
kkoTqpUGO2romA4aumNk82LIusWxRrYKUhfGrGLCgialb0U+ckJgmhDyMWTCPkf7
YqGlGGvSBbYb9QjolSYX7NLifKD//efp0InknIPoZ+1akNSkrDSOumX3GL8+z9ao
gt9nDPfIGZL9gCde2y5xxVQtgDUcOwqwhxD9tEaYsjIYcxOj3P4a4DmqkJKczNVh
CcIHSRJe0vfvRlAdLGLzNAy60cdYuqhtFHCeD6TNF7XLQXd0C4LLRgwTst07f05j
gQnD0+0Q3G/pnX1mSsQ0X2wmydNu9AlhL4BqI9/xTb5dPrNFZ2u9BJGaIvwMW2qH
l1eZK2dGzS65gsbFTrHOaDflKZdJrzSNof92lpYNl0nEfHsu/E+rmLc0fiirKAwo
nrsjZhAUdBmJxnzsHuWMLduSpk42BC32g1hBLB9CMtF1y/eMqQIirU+4sQ35Tf1f
YnNuUyw3d6KEYdxsSnRAV2P44fazKgqN1ElSJSswf8ksU8Fh0mhaVedYrmSCx/+H
8FhctZwNCdFNNIj1PklhcTLgcT4tyzZDAd6hC2465T8aD39MDXfwMllqLvuutIai
dQmyCMt+RCXygP9Rpi/jyeUPmKzWmwtD855YsLhtru889UT/+kjk8isgLCeJOlVh
PS487x/+u3IpOHcBSTbmaIOOBVUGjBPdacl4lOjZRD0zOWm96ljCYOQ8CVTabp+8
re7rfA0WGJmpk15hbbe9zW8dcW6aqi1hBFRxJiN9uXKR2iLeBDabsN9/ab/naiD6
vsBzZOMOrI71E1eLCXOC8y/WsoSUhZiNGr7mCvQRS8pwHO6ieuf21ZP5/kmxLRiN
kJRzHhu3/YOL9Da4ydpkqepMVrmQMXGJLDyYIJb+0tCM4SDcjSoDOgmtfLmTxP5l
BJjEBFjqTkcGddCUsoUQv0JzO004a9OCAuvc9WOQi3CsuKlRgcx19iOth89u2kS3
11g7MeXJXYaCCR891SibNkj2R/xJXmWqD+4lWRqpyAYv7Cg+SQnlhUVFRJPKND3e
SF2Y+sXD4WKQZM4rNiotqZsEMxrEoKxp3FrxLKOhzdb7qGYUnhg0dTFYi8hkxUdI
pn8+4v+CaEBnemN/lOHFw6Bc16p3M2qs5m+daOE/kqmKY85LMo816awpymyfp3yy
f2teKAYmwHLmzZ9FdGOSQCWfs/ZH4rlUr1fVy44SHTPkdYYpvU4u+itkzfzG01cj
4Pn1PGRpBgTg1AZEnvsOFKP5AZpxTUDrEgJ9EMM9cczCEMpSYKr2Eky1kcx0dcnX
2MCdsHpTw+HNJRZwxYlKpdG1G1YQ3XBXpcvCGK9mgxKYNgoDvoqnbaGbC6pToPkm
nS9naD7zZ1M2pNMrlI3R/SICWDZlQge58WcvQnIQXOqiiJ3P70CJA90W4QmBoM9l
1Exdo+AXjUMi5vw+czAY1f+40jYAtdtdDoISn5ZTIy+fXBQngVIFkvqSUxXwRkXe
VLqFO3FHq0DyBSyOkJlwZt/yxU3kzPpu7HH5pPpmuujn3pr+ADlm1fixpVR6zAcc
uv8vMsRoKSNriKqI9PYdtQWutvZ+sJGx3u5HCbwqIuCP6bnV9dLnGxvs8GD5xUl0
OgON0Uf3LUGLFLISJpN32+MFsp70M9UBqcRe7mL2fRfg+jFdKFwJ7JxwgX1Jysib
L6EjoD+pKhVQauRirCW+fGdMkuz1QEWIQdAcxkrqbrWRONhpsHgMSnTUBRdwXy5t
VsuR7Pk3GacWs/7RQHHVjQGKMD1D7ZGSQeY2YnufefW3YXT3jlldPYjZ/e+eoAjG
V2X0Xq8KT1HBYkusUHfzIpbxUWcOB3/8JGrgvTrcfPOeDztZiAbNFVcic1eikq3g
K9jXo1aylxSNqvBizLFZlhdMl21iY4mRx3CCiu2JfBDLK4KyTnb1/ljTffTolDQA
weW8klbQ2/mlFWDK26LYHxyKT8oy8RRpQ2CsFHsI078lpxgFurzKUoBp15jvsycU
fJyJTKMUbY/CUxKZKrTb2wr8JM3drviv+yNNUoxAvSZsmiY54aglIAGyKq0wamUz
bDAF85yLHthaxiTQV0Ch58lXJ0cc/TuLxw+UH1Ef38uYm3ly9+OWmjsC/Xh8Z+vb
qcn16WT+9sd7hqGocoD2HEACNY2T4XXK57+giYWoEiuDuN/yRKRs60k5QMICt9px
KJsHgZYWL9l3xt9gSZi31sZEtbPF3KRQDbI/1Cc9zt8KcYXccr7ljkbjIIsTmKXx
IbLislGazrrte/qQSDT4aTH+Z58gWhwGoR+Q+6N6Qc0tEPDI8c9qv54+voZcGnC0
j51kfPHcq8QyUpAfkwmbO9NeSO2dW50Vsqb8l4a1h1HR49/r4OyQZl8BiMAGoTdJ
yJ2H2xX+oNFoqViFOKsRvORRqDUkvvOb3HrDcboI+Y0oXJpgpbI2Jmv80v222xBo
HFmPeSpkcCJlcdkewc+ODLPncpGhvBrAnU47m6cYwiOrdffSq9s5AiGYotcrUs0G
2tylXNdkNaFHNxPUErYtTPI2cfICoIbPrFLjsD5rsNuuG7bQRQwQpiSWg6gvMUaO
K4N7P39H2Sj7fVhpWZJbqG6ityN1RlmiN7jEcWmXoMn062BL1ld8TnGpkqsmUc/G
s98qeEPDny943vcKQQ5qBLgrbE3EonDS719LZKZqcW7b+FpLQryqL+V5CFA4Yafp
Q3Uv9LesMtl+UiIzhXfgUSeqdVjCLSou6OvKzcxxvCULnUe4XuAP/cPJSprK4rkZ
aYp3bKYEP7o81MaxrbFphb4HG8EFYtGrMLQcNxwvKik=
--pragma protect end_data_block
--pragma protect digest_block
/vFMzrqvUyU057eKpaRYJSAmp6Y=
--pragma protect end_digest_block
--pragma protect end_protected
