-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
pSV5Qn3AtIJBjo5mwOZjH5KxNWv/qJ9bnT3u4JBe5S0ixC1gmuckGpUjV0Fiv7/Xu/a1C66TTqiA
oMClMH11WsAIP/QbEoKGpkx6pOfaLe3GMzhBeeDcBPGDuwexleCiIoN4BhHEzC1Q+RZF0TeYXWzd
cH95wRuZo8x9weaAh1mwgJtJxwrBjVFEhRXnO0Q1CFv7YPiwUOF/u7UR6f3cGYq9nT8M3mv/WTR6
jyDHHjUvUIdGsS2r7U/Mz0QoAPsalnPXLOdwSFiYDa4gdAtxw8d1CpbcTfLxzVBsYwHBy68PUMX7
+/rWCfZ/KJ1FOBRBM7oTWVhd6/E5zad4GnBiIw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 21424)
`protect data_block
C+58/rl1OcsU+VrvML+eDRXNNuq6mjb0cBMNn0wzQOczbHM9HQE4SWf9URW4sjrSswAIsSXmUVCi
Q1qv//JS57fq5cPLftSOMa+ug0i7eJmXjqSz1coqDwAgDTHG9f/AJeA7wkCUL84GgYgU6hg+5L89
M9J100fDYPTvbhPLfoyc2ajCzyk6ANHgqdzkzTlvdMoZnCXA0IY+prGchrRy7yZfZpdjoKQIvTqI
3Jwa5Fcfs9zTTe74SKjVFo01qoYMFLnm+qtoh8Jq7MW8PTgJzhzzWs5ok3h6uj4OscNQSqqWH7T7
+vgmQsG7qKKJ/ZOJq+BwYdwhgJQZXfKocjBScYQY2JZoslILgTNr/03WVvORkPZQsKLmRnBg1Nm/
aLEFXbgYMJag4UVhgkDzXmsqopUAuOi1mBUjv7DUMwZbsXLWNxJwJ88SvdeNDnFmcezuihH0y4Rt
JPNbe3spCi5SXsbo1WK0vNFnqTwjk8mMxXRWvUPJwOsIu4jpjqu0gPYnIjyHzKEpRjIdZbEsJsD7
PJkKBe7xk66GJwOWKq9JZ6kPUuHP1sjvT9Zme3oxczm7aqOmAI+hSMM/FMfHNzPth6If+YGToCyY
5ohJDlRuySA3nJrQ//+0jzh6z2FSBWDj4DlISIPpeA34ZyCRtzXlzgZ/yBwMdBpCoWoLqwaPU8L7
Q8EkeyBh/YB2eMCAgpIHA6mmCu2zwNyBifWg9xqLDKBjqRvPGryQaZYfLUiZiD02OaNi5Ncin5PP
ONKsd6+6BXR5FJS6oEy/22JIe1LeuPgKZQeIUysOwXodwE6y70uTjZpXqPg5zGJPCfdij2RkOlFj
u/ydidBjAnJ8pxNg3rPq99gDa1adV4WHhmTwPQM7+vLyeLORCxh3lfk48cK9usCfu/yR7AOtfayQ
QhjKVfv/0BVyhdB/Zxz8iMkuFWfpeMuoesE+lQs6nFksfHlS9Rb4U2ER99qV+CQnmJ/6Ys6KrDcA
WEVe1QhC8ApWqJV+VQuYgRpZSzGJ0HeNmtZYk2wsGHPv84RuNIfQmqZZ7KsuCV2NbRUnCRdrvkgD
XLPPC9x9xGkhvIZDTbgQM5Qkx0mhx+XL5SzJi9+lAfvXqbEjUkKsJfYVirJTw4icRqoWkpymvOo9
56OTfnaHXUuzacKDEB4WGbcJWIW3N6BRVd9uCJiMNejLPkGgriajHFXEVMpT158kDD2UsCtbG6Pe
UuCIYGw8wOm3yCt1FZ+OQkiBTf+Bmdl3hkHmpRYfVOxSP6PCgbxx1bDSLZ7hSEvhbRdZ4GCqMPKY
l9xrJhkd5DWFBvlPKi3JEqkOWnjAluSJCDpTScFWB4YF6Cr39K+IJF90CKSsSQsM3FpIiyju9rjH
R239m+i81XI8+aE2fXvOY3ekrkfBrwN+GpP46OoZi9n8uUcingVVAQxhsjWjUMnlDAkr493oCfJ4
KwyYBu6V1ZLfg57Znw7Jl3ts4GRVwNyeWDJKfbCNqItIbu2MjKI5TME95IENLgb4JDKkve/xudqt
OLLIlipPudJusBOFM0COU1ekYx96DGEgceq87HZ/NVKuYGLkMjqHCCFCcEyevhGRXUM5UG3ctHkx
46BS6rrKlJuvdObkZDOryR7WGScwFSCYNGCdqCllqzKMuNyjpamT/5xE7gbueik+/GjbzvNd4Bcg
7kPXjiP6UraW/76FDbcnC1rrFVlMq7DU2YxQ4JZFtxGoxdGe4T9TbGC2r7xxptu4P3FMGA0uJU9+
0p+01otA5pfsetQ9S7oNXVLSASrT2ncqHOCcxZrpQUvkIXkcFFOXksgxrNFpXDq2QvJgPdegva5m
BADeugfUPGXPXI1iOSOIrmH1Wz1AUfTA6gN8yD/IdGkQ8TRdSHwIcr1fLI6f7E/ZN1AMM+5b+3mb
hVNtvH7swxRdfNd6OPUwkUbxLRoogHw8VxhpZeGYHvv+z1AVdAeDbbIXrtXEWuP5q9iTpRLQ8qaR
th+Jp7dgFkHXu+ErZoipK5N2+KRMaXKlKCXdaGa0R6ZPg04R7EFaz1btV9cXK1Hyro+Qd2gjZ58R
MAsOAjzDZ+YjxWstEA5cmdueokKWsLfTct9gynbNPm7f53qYWeV/LTmqwerRZHtOO8XDExU1fwuG
DydJF1m3eA0MDTfWf1k+5xPjj9c6iGGK8PabPCDGy+jGKXxVeEpqdADIqXfkvMfgrcpYa92gtmKq
W56fdw+UGpVkqKqQSwCyqRR1SUZ5r0yi9zHnyDMt2SnAZtkHkVTRJjNQsu25X1Is37+HTXRuqlBO
ky12HCoQAHxtkWoU3F+XMrls9ktNeacztS/vVgJ/rO6coq2qYffrGI2TqUEL0f/H+rM/ZCzgywC3
4uVajsx7Wn8CsnUbIIBss4gX7pWlCxAmWpP0cCPzXQZ0YVX8yyxTXK58bXxOKPcM32hGSN33OGW1
0Agfyj6xJGju/HfhBaZF6AxRNHYL9dmK+1uGG3/DKPc4QZ8p0Gl+ZEREOq+4McqKeV6qFJeCA7NV
rLbsFIeFu9f7m+lCoCIQG/ys5RvrNBf1Ank4CxHTYE9FvEjFlVbfZb7TDvxsvyN4JdHfR6A+GGmS
+1N6n1FGZd/elLNp4SuK3Vn6dPoOH88znKUGsbk2owXxCrPWXH6v4eVc92NlAxErtfNhL5Xq8S6C
ochgAIdLoyVXxeUd78B1LWo/+ilVRdBFrz76lBouaZ5/ZSV/5ZPsm7UWwDCUz9cOjgPIQ89mfhD0
exDJtEbj6CHXDwiSZSNLPcCmmihTPPmO/oN+K1/Ui7QuBy3hcJkVQiD22kW6J/lZ4nhJgiAlhQWA
KzxC5kFBjSRluoUNA8dS29SROr+kpVBsA1Hi5HLW5NmQc8TJbua2so45jUghgRFuOuUiEYL/nVtL
EBoq2WKeMxOsX7ecybaS0KHy238sUQHdwAoc+QCpYZE0b17Pos4GfAboocDe0h1KTfBrxq671zI6
T7otlxpv4NLcbISTvLRo0tPDPiV2Iazejw7e2dfBtBm59tQe16fYmoUYsjL/QmFcnAeN9RBbU4be
pG/NYsn7gMUqOo8O/z7HNcjf3fWzoYv/+b7jtg8PoKt/ZcQPBP2C57H3BsHZR+GNnCiAHfuGxGyw
PyFy1+9R582s+q0S2liIsM9cbM4Vs6Db6ZNUUSe/QU0wfCqcfNCHh+RoZ7d2W2KIPbyvLH/+DU4M
XtrP3jYkYwIG+7bIWqEKhJrfQUlZBxnsKLiFGqTM9ovjYL/6hBB/6K+2XfG/EXKJfLB5EpgVBE13
+DoFMBpLDC13azftR2/g/wMv/EHjCzumNu/ghKCefvj0PH/9NrRVV4QPh9EhxsdQu39SbR4exAWq
ksb703g0326lU+92WXn5EIobf0HAeE/muowlD7a6QPYTOqBndEH2k6ekd6CxpfVLdH8K7SeaZjeb
gsvFRRd9G6Cf7sqfU/cq2BFVSvR7A/gc8E4130+FdtAjzaZSe7ptAFk7AtNaOLJjq1dYZEwVrFTv
/O+NoHHDQjsxrVUiAHSUdxF2DUxqshLZRSFzPaMHIL0aAinqLMbMK4XRpezds/S4nnAlLsp8t8Gv
uLDigkAc/I7FS2Kp5NxHhSS77vv05Atxu/Kpmvn8KIP5hPiKiCET3H5r9gYR+QFf7u1t5tCF9QBg
TQWtDqyFLYLoK5Ji1UNbIPOzEIcnVvseBq1z3YJY289bOB19j3vAA0FriPiE/gIi8zHp33ZcrVO6
vQb+XlQ/yjCASsuZttL/t1gf6Tcn3Jv4dDLSMD19yjo4gwG/NxIwiIJdrpumiF5mPdZDruDa+i0E
LBJ8kJwsxb4TV7P71RoKblmXTy1zUst1lKBJx9/rv8leZlzsdpAyKqn2iA0nCqMU7lTgMAVSd3dG
j6Khi+pqVYdzGCp43LCa94LUxJOXtyIcLffGWI7C5KyG3LvRE/Bmt+s1H4XPcJxZXSynsGcR/0V2
dpIkCO7h4kpnpt7uR95jx+VLf5bkeTav+yXt4i9MTkiksiTEdZ5AdIDXUmWV3ie2g//dUy1JOXte
QhwOAubTSmZSGQ3YKKsO0S/sWfDZtxmUp3svKT4+DTTpi0CBmTzQrA467krVvBbkXlk8x3CR7SAy
p6a5HQPYDwEKn0XrT7aYeOWtjyAFn/ezHEBKk9gLqrAd6GWWzwIcZ2JmqQt2CcZz94jkLbedBCOj
hZGHX7u/RansR0so462dUBYv7KCG1W7/IbuXC0RcZLH7xgZIQawY1oIuXt3RIInb4V49k0J+UXq0
MTYJyI/sDGNHaC+4xayOiIsLp2+O35OOwlqYwsh3LbSOiJ7Tnt8FyD1sSs3MeQrSmn0YhziFPORb
V19yIUGBLCI4dZgMue+oHZx2ZqYkxd4bX3GUniojBu7DLbnxAAApjlqTQWLeyHjn7Xv7cy9kYkl6
WDs416Ja9UhpOiLFAC74jep+tPslNPG5bUhW3YZHtNDdaVvD/llct5zsQwe6/d+4DyP3GK3wxQ0T
w4Nc1zxrrL2M2pGtbCpDwnRIPmYzsnL3sDnj4yFxOJ0i1ZrdLIWxdhFshEMd1yvTYaUyzq8d6v1+
SMFsx7gT0EkxSifrMaKE6FvXgCx+lcmi+gVm0TXlTJa9b7foqCQf03NmU+3vL5DdlZ5gZstSxZww
7dt3MkPaH/kZGdZFLzwblT/fwntZKMDB8bJIxzQyuSnRSNY4uEmc9Y0TeHt4mbEJJBxiYfwLfaUx
pNobSHjmLfMCfdgVHYtOBYRi89rYdAEbqv9ZaBL5gWRBrAyAgEzUqyzHM3RwbIJWhmHrsmOCVRxk
BL3Z2MHbDIXCq1qGwNZE8cVsduHfGFb8AZKgm5SczjMtLj1NReFhb2PELJRmxTMJXFjCg/fqW/k7
LQ3USgsMzlhNMtBqBJ6J0ZbiWG39Mrx+d+HnP3+4szaZVOLf4hqn7xjDvR3CjUi+S9Wfq74Gc0Ma
QuH21xwU8w5pkB3cPKS8iLr4C0XmFbjmO3fFfMawiM70/MdFwT++iwgOxFO5O+y21pWhAPsu5Rhb
gsqGYUtrIBb0NcSdFzkpPht841AYjkHuWKoxQp+lgLS5CJreOY17QvaiJ+anG1TgfNq4LdV54m8b
89uIdtg5PLcg+4GpWMCD0Nj4+ps0uNUhTb00qweXNl1oboPSA27P8i0QjeFW/M4G58seTzSmwV/s
QwHm1SDmbc6ah0+KfjwJsoq6v6QWKxenGy2R5bXVQHnOYrcC5lh5BcflWNDSh9m/8TjvCqQf++Vn
z96HH14Y0Lggv1SiBdUGk6iLjz5jBtjlNANznyKoqS+bPPnlH4kKfvhtPLbbpkkHa4BCtzluDxzl
EBjfdlU7O9fl0yL8PKLJxQ4EF8iKr3dba+LA8YWXHF9KtJ5rkmZ0DqRUbhnrZOZm+gK59Mms+GU1
RIfsHG4Mnf57SehvMM26eHL1L7GoRaFnoFYYCG+c/ahHMAYOESVuTsui+YP/gbLzJWA4OXKFN2cq
miBdftIgdB11r45mcUzsSvsf035Sm9IMlxeHHLvrt0dgHQ2LLhOS4K21XjZqrlv9zx8OWtYvpyb0
KCeIIOF3J683mywzhVSWgJicIL3IoBB7vHCOfmjhOPbHiy5rbMKTetCppMgojCQEJOsnylihKNys
m3OqPbBfr/wNGk6otpRiYPSSIEh/M9ivR7saQynrcBW39Zi2J1xgNy8Gv2RvVYkwxLxHAtOxQjor
eOjqRyRmvFcBI+lFXgAMXNPDazB/PBXRe4Itn3lb8utK7Sxh703il5+CwC0uPxGfoYt+zWqkF33b
yhAYH90uwgSdLOdDJJU7NSzO3866xnhmtoCEgl4FxeXaV79nZlElLZ+RytmgsV4qnT43NXVH5LO2
IaOPIqgjiXPZjwkpP9ish0ynn449Z+6vS+CoC6HIaFDkDogtf2OD+aMygTj3nUPgO9BygNDBrPks
QEL4lgU8hUdQf61/sLunEc6Wl3G4sf0PPZjlaOAVrLyz0zH6I8OASWo/koObNXti/uK5BsT5oNWR
AAUvHFDjqrwejODvhaq/ykcPRQA/KTamYrld5Wl0DIiWL25TkhPQG9zfaQ3GnRhWa5Sl7v3eIY97
KNe4zzG/a73R/mtutS3TH/uFSpqtOhjiCBQ/Ao7ILpxxmCG8neQigPP2r/VQe8m2/EON5/iOcIJy
3UYNdq/C4wCDfVfDVYTBRgcqVymWZa9hlx7WSZIQUZkrYCpFzGhvLsWPd4qKX6b/WwEfIFiLHKb8
MbZts4DVw1kwrOBVyOw8BYqi7HGDRBmLxAv8IE4mKtBTgQ6NDI1x7Qc0USEJkcst7Kve1Ya5xolH
Doa6qF4Y8w9cgMcYBSS6lYylg8bWtGMnMALB53P6J/aq2vmfj01XAhNV0lP6qJZDEP8Px+IJnpZ6
PJeyWoRhRnFPEHoXGx7XwLnZceJ5yJPtfqXAtwUM+Jg+ZCW2RH1oNQj4VsmWS97cItjKrzPnkgdo
qFEpUQu2I4WTgWFzIty13ppvahNz79d0jj4XbSqjjexvMvemptpCWWv6kBo5tEJ1TqV2rAP8aS22
/hyjDyuumQKG7dbfQexW6f0azz/SrmxQN3UTeteQX+QVIve8sdOjsj+74P47GnY5CwvPZx+JlTgQ
m12C5NTduk6l0Y30m0JlZCg58oWQDawT37kTztNA339Ngdcf+Se9WoN4MRIO3aYWxP1SJkr1inbE
3hI7umImYmSOoymjzSrpn6FR8i/d10H/AfhvSnQJk3rGwh/4eAsvlW4y4aEPY3xS+A0o8rCNqbtf
WtB4NodOuJ2ElzHfTJJqSM0QO7xFfWmlqgbrI1zuaRnSAac2h4/9Jzoy1V3UeFD0puSPfaN3yWZA
MvL63rnEChHubWk33l168ttkjeuvlwgwtuDvW1zSh/diEr8nsIu6adoxRo51wip9POmi8qlXdQyA
ffDTUyQGB1p1ayxHk+xM8xKBJ1/s7HReHmraV3u0/ugdwj4Nhcyvxq5IouJTdFLx7gwPrrKhrzL0
atMinp5tQvnG/TgFQVVZTjWozsD4wEq2JTFAtoaPzv54zzQ7ACbAl6/DiMZJsUSylY8f09UKANsv
O4YU8GMRl6uAfVnZl2zNXv/b8sEgz7X7OpWmt0WagC0bzE1ooNShryR6+K0Efgbo73yRm0ZKFACt
fZwiuWWfTx0iF8nQSUi1D7lUC9VePskodpzgjWOQ9YPhnRwJK2usx1R1hXDhV2P5JrLisDcUCjjR
IJ6v/aCaQp+fRZox5hsAdJ5/aKqeGPuw35mCX6Xg3XI4n/Gri2KyCwbSPUWATpsWsZRzrrj7dq10
bfGPjOq6INUw9Iq152JvxDN9/7fLrcbdVSGVt6C/GGme+b8NsAaa2h0jpjc75hHjePrR3vsfj2N3
ukKOfcSL5pdE3CU0HY0kECGKYnkOHRubjST2kHEFYCNib8ceg+b/BJ62JEFVUwHcDdzEKriYI2yk
bwHpwhmZsGlNZY+ix+w64j7fHZfVOvVkIxB1FBmgeb9svLl2sU9pxvHMTT8JoL92k44uqTX1yOr7
2Vy/GyBEyX8jPgc+RtsYsP6sFtJuYGnpg5GMrUm6BfqFNM1xZSBYoUoraTEgs6aDgM3apr/36NKB
7i2zXRq75S0NI8H6L49pCpSr94SEW6aLZbIrdOCvzYLgRx/d0R33qnGNdylAL1lmbXQUGik0KCJD
UKT+qXhyyEjnDWqTR0Ce3zCkEMVbE4Drm2r6+YHrTqwP5Mn6F19AxNnB5X9GmtqxLrzkJcW+SDeJ
AYyo3gMtqboQkmHvp0aBv4WkXLFxDobfNTxk55DfVN7RbCJBIwsaENshqFxwZGACBT4iqBYvD7zx
1OG+9fB6LRDXHGpBkrj+X7p7MQQ8KoSPlcrbgOl3tPMDayErC5JObdhkMrtT1LYfWIhvM+10/ERN
TSiilrEv1f6K0LHsr3VvAaFLivz+NxGjspmDZx1D/9OXabI3BO4amD1A6MmfsLkqe/LapWvHf9Ty
N07xAzZOtHFF1ZNFGELXkRbvDeHUtj8RKY46XARJPVH++U03a47Bp4cu7pwnHum2OPCpOcOCsO2d
7h29fWxYMVMXW2Cd4XYLzA/T0YnxOi5f5Z1mZ4OaLWL7Kzl/AQfntEE2rPsHivz1uegspx7Rvz/I
yMJLfVbd+/tt6yoOzXzqUH6ShghLC/V+B5rUvhLyYfYv/S1qGLblVfZ6kedW+7bvmNjtp+Wd8JPr
utczbNLGQQ3Ew/uL/sXFsTZOBAMzJ7A+tOP5iS1+BAzK3x5WsxMT4Rlo4QPIswnwJSkKzK3ludqD
WI8PF0/NzszDtA9FZheK9xw54RsBnJ/vYFjdkxmXa8gkXs5TCalWyDjC7zhXmRm2DNFd6i0ChPTB
iA3pKeqm6GyDWtfsfBotRw9KkW3ssmo8xPDVZZL1mnhKJYEkHNmH+I0vHd06pLPOE5RBaNyo9lMG
OiwujGx/Cp+9CqFUyC0FNr9qoBunBNhKX25qdh+xJ8LIIh9NyyYfWAIJUernFfxBALGJWsXDzFoZ
HY2eelbQPxrtUAmE33hqCuPurVYNEkynxD3fuNLYpVpP3TXf5PFpOcrrBlLs1LuInji9vvyLI/FN
0AKFRYEKtVds2T01wqlNJB4EkBbSyQjC/OUkjxyZy6nYp6PUNn6SEbBWRDv6cQyCsZbru623HGld
bA8OQhRzMBGs0FIEGpPk9z4rzyqZ9c67sUb2g+SUJYZsty/h4gYyXphFtBRinurjHfsk08bAJzbd
t8FdT9MoJPD2dICGFoFhoABa/WZp9GwPtafHJ1rijYlyt4a7mkR2yTlQrDEK0GWz2/nv2Lrl0uc3
WF9qc3wJp29UlElPDb908lCd0X1FQBklawsGdyNqH4FCiOlu/qtnfPXVT2pFRaobQXPx42U/Nv/V
Sm7SjxVj8IyH7IMKrBCWweMOZzBEp27kY9wZxJCji1/6uGjzjtWYw/saURshih56u3AC10zKszk5
gka+OCKr6fUZ64vpq2lOECAq5Tt60fqo0eUVggB8/5Sn2yFeH/ZHCb0nYGY0JmpYACwMDYWq4sMl
xEa0X9Y8J9j+5HG9UId5WwHbj1bSJyC7IN+SxWH3lU2taILEq7tTcc+TGyNIh5/QkGYeZ4JH+5+u
6D5WpL9LVTkwsA9xX4R7gi6iQ5OWSd3lr2U2z6/ZeMs72/oPT8INzbG2bpBvXM5UAOUzadkk+c4J
gQ+LwPXbpULwQjqgdsGubsW5tXH9RErMwsqwQzX5UE3SswpBwnwLfwxQ/wiMbEzVzooht/kSoZGU
PRp4Fkhiw/oGD1KsWIeN45RR1LPiNnyikbq0wbs8gtCb6r7LWpd8l4rv4vRiFMAxEzFhoQNVOTTm
4d1zFJLJLtJb5K05ZsmLQ4U9GeDTwQTdOUl+6PKAJOA5j8nw01sV1CymB+tCUnOwu7O5cKZjiTLg
oewdN4DgAjPEYqHtf+m+caADHlkUUjqrjPczzkEzp3YyOXhp8WHC1BHxtGkvBQtKZw+PkoElLouQ
RGjzJpj8nmHZwh/o5LvGHVY1ilOxoO6f/qwjUUyQduGQIH5cj/a+6FlIyoX7vQNOr48vFVfo1BkV
+q4bEYeiEv4//pNC0yJJ3YzL8d1c/h8Oo5dMp1XDVomHoA2v40uCN5/jjaHLNuVlFTSAkLThw823
wRglJWl6FwOwclzOBTmXiA0t+XA61pl5vzdIVSX3ZSKDzLC+8C0nCwNO1Ktw0mFjcMua5ohUyFx/
nkbgZFRJu7bCA13mjyqG2C8Ja9Auks2mjSe7LEe2x8mTk0L+jHrpTId3Ll4KTRQZK0Yo7lWuoCZ4
QM1M8D5Gyd5YeuIUTxA5Y1Ic9u8Hxei4RGT43UEC8F0JgI/PKnkZ3U43YnpAEX6utRj3+orPFD19
9BMAWbKnLnxFgWkVvToA57KVYtTMfspyg41fwmETWY8OQs2xwv4NwVGcnzHa+qPZKavWcWXkBQ12
0L2Gq0S7sj/aZjfYWy9Wd27rLRLD4EJ7VVm1WyL+Fdg3qHd8YmwfNIXrIiurwUQqfzL1evgH7mDo
MobKM/bt2F5wAYsHkIBT4XaILdGqQLeHcNjFvtnkzoaaIhFnidAkq4fPtLzqx1pl23618YWKBg7b
k4MRSLJsC/cjtRGkosKamcxyNUoodLBrimvAIFgCDNrqJ2x9vFR+HaS6ya4d7VW5zMVB7rkZGVp3
rp1M7TxVxeL9R++6iSxDkuiXJ0vcic6FbgmW4ebBvYDhlePxIqrkXrlm8Ga8zVfVPBb0+WSSphZ1
4OeyXYER1gZD63ViigbRE3WLHsx4e0RrPBKFmcUMb1xBZEl1AR3oXL0og2oUS82mIkS3oXWMfjC5
wUK4slX5xHnDrMvWaHwdUeETYrWRwgqs/p90TTdm0fFiQHbqtLfLa0+RUxXD2JB/tZUhT/MqDCQv
uk73rNZJ3zuCrenCvVrhkFZHqHOuUnf8uy9VvzU7K9M0Be/gxVzMLzNAxSCn1yxAmJSO9FHcoSO5
TrPCDm7O8kdNyw29ASe/1F/NYXp6p+guvl1M9GpkbKOnYZL6SDP+sbXNy+A3GanEXdiXNlzlU3vU
epY79nsdyi0JYXa5GbSNw82BcXiKzv3LoPQmmhKNi0yFwV6bznGTZo4lHt/NO4WxV9pawHBnCT+D
2jII+UwXV+XVtK+oswB2A5qs5ug5NVvideg50D/W4MD9XZ47lwWDDHhQwIt5NxfSaGyVcAzvucs1
RSBxFV3AlMqg3lyPIxcPAZqOpYczF9APh+Malcq+PJNJ0f+zTbe5bvx/BwJKEhBi1kE0PG6vy/4s
1BJiiABpsojhWucJc74IpA7uf/8K1jS6jPyJakgrHFEqzaBtia3uceA4GmrOZ1yhJlgvFQSWmcOs
DVAHHrrejlYLKmPXzLNNYcnfbv00rMSyNJMDiZ4vDVnBfD3jcZ8kh0E+g9Xgd/Ng5zyHXuszP3Yi
YThRp5PaQCzTqouIot8UJ7cSiV+YCfCpdlg0+E84PP2p2gvS/7boMW4/WWCpfsNomyERbb0Y70mZ
FudPyyoOcEfEVFjhAfl4Y6sA7SH16uarpOW03p+ZRQZ8fLR0ajEU9Tdq7w9SPsdRBtUR57Raveuf
w2nSd7aplQGGwpYPBNYorDNU2Zvj8cvC+lQ1VXCnusDR705fZeLAhF8wBaEXphX25iByA5Wi4r6x
S4yfTRJGOwlF0lAt/7Q2b3CPgkaRNUHaFw3Cym+HRIFJg7jhNG7JxGiAbtzVCqJ8aPU5bawtJcux
/loSBsNWELztc8NrEXjzRMpx6Jfki6Zqvr7Q0I4fzPi3GTx6wRGUqQYZL+pInZMF7vnr05lzpNot
yCRZlYEnW7P5LDhJVJMfBs9HuBGuH8x7mpe6CsFvO9ABjy66M9/XH8YUGRZqxeOvSZyJ05O3toQj
NdVrNAAKTveFwfgWC8W/JIRWUS3fNHR3yxhhfLXV12LR5Wp7MAFZOY159exJB2NvpYnUTtZSbdSL
DmSmuGs/AcGCcqCSqDMZ7BqVJO1TigEq72c0uQj90rJvUYO2deP5fXd6NpBEJB8GiiFjhoBjnp3O
hPBAr2UolzJ60B2/kFcJ9lMMpYeqtdJnu27LTb7sdo5ePy8l7uEee8nCLx1mpPuyP5kc/DCCj36b
reQpr4m1NyA92AxpCj11ucTYEg0BgtV13WxGVqRlYKIGDo8YrVAy40xZgtf6iiuBKUI3oxkNU0Ya
jfMVX6Wa+C8Wh2It6UVJdE3uyVYyvf/lJ3HDh0wHsc+55tlbwJWtQjb4jf6SHLC3af8IxVVyk0IV
t6eXTBfzqK/Ng4BC77T/AP3Wf3KppaYXTwR9RWLM29yxHhBQeMRNNH/WwePjcLR/VoCv1RTaYjjV
3sBmBnH0H80azrzMWQBPZhoG5QsuDJYK8ATljSC3RPK2iHybe42DGj1l9JJGmux1A9vpKh/hHkJ0
qh+/IVzIAPl6t9uWB4xyMoRRR8/o31G/hQuDOPLMQJ9ODD0oxD4bfoW1CMfJo1D7JGk62n+V/C70
+mHmFlvocfahy9p9q3fgaAvfNDqTBSrg2LSb8tbSIl3ZGAavPd3cKYJLm1N6mTTAVVk3erDdtrzy
AfK9df063NWLzOtd8S/n62+GsYfHCefdM+oRrS4cEnWiJHUPhAA2qNbizN9h9n6r0ZCr+8GuoGOY
POueVYYp/N69mGlpd6gVB7AUa82jpomo2OwVHr2Amj2ot0XzByEir99Uqq5i8MuvB8d4ije6x10P
83AshWn/x/K+qC9KjoTxsU+bb5+ghcZzUILt5KKfI5sv1GY6wM5WfgXFIvNFLQI8QMqB5WtalszE
WHbww/Cx7Aj53bVpbBYpS4tev6X5PqepCUljKf0wzfzhtYYWNQ9wsftMCa+f8aTpxRKTbcIRkY5T
3yZquE80UI1znnZbe3Gvu1IkJUN98tqfbr5kDAtQK+e75C7IqyPOgErjE1Fz1Ye1cyaf7o0HujzC
FAWiLl6PRptIDC0WW6aeubIot/8GR/7gJ6XooJZhij11ssChkPPiCW9/Rp4kGyvzveoI8TYXbfKL
W7Ig2yo/3tFKfcpE9dciWfmBXIiX/k62TTK7yHWOL7+NcxbttGn2hLdDkjmdyX9QK3izTvQ8PkXT
rWXyNVlrXQzoFIKktKEF8nCOJpHdHZvU5e6oCy4y5MUvl/kZBIW52oAPBebYBO5Jcj88wvKBW36w
wNat/LYWmKtlEziNvfoHXPNylyhiqOLvTAdU59MYXyNh5JXZnVwuadSRIg9dcfiUhnSrZMmLIQwW
V7+kgJ91rFt6OEEDspwe/lY8deMqfkqy9GhUYOA8udiLySF/eLfn4pwg9kGfLKuL0nU2PcBkqPCR
7SNRPWXSY8Ki8byWDxKb7pV3ZPWCyYAYkVtfLMgT5ICCeoYyR1BTckpqOJ85/L4v2e835dEoXDlH
HnTZ3Dxqj5ZBWXSYj6LCIH9z++KZQauHv6KevWwuSAAtXIHS54kwjkZ9r1jwoKuLVimFoWi33CTJ
sDc+A4JW3a/7/Cy5zmDe+isAEaSxcjofP1vneeUfkrNuBTSc6PoYiewbJL07OJ44qzecMrTKuBOj
ZyP2sKxFWDwcJuo2VlklR2J/IhRJNNL6T2MnVTK/R7IEiQIaZ9IkkoVZ9M3PC9lWzxUil5bEhQWp
YbV443eBc1Hj8XELKqJEaB4NfKGXcAwV9VX2Pnd9pVgKN8djv5jVZsvG1XjFgc1Ldhr5scpsHbJ7
zubnzVvHhhU6M7q8hF2ZSdU2zeOKlbi4g/VtjBMCCyi8jmWvPmaQdpfKVNJABXIy9w2lXaEtTy0a
jv5rzesoaGExEBDxcgZRxNK7nGxICOoatFU84h2T6j+knLxyj3w6dGxi6da7bhD09xsLQSxvPmPx
cW02WkkTIO+pHbfH+0hPQLTOMnkXvfp/jJil9LXweI8T/nx1wIDXvBffy6s1B062AMoM3nnj3Gny
DBM2Apr4beBB8G0qoo3v1/N/RuRqKV2KuBrc32KfhIm9L4L9eEwZNBY5899T8PUfc6xT9F1YvRRn
uK7b74C4O4Rx69Q/6+yKolXR2PfGbDXHxETOTNfpbGjIHFCzYvY3DvFTww3ZPn+ab4jhp+wVu1EL
JemUPIkhOgdXI5g0j1Af1nHaQTLYMS2XGbL7cDKCmqWwfNY0d8srKBaCcmbELDQ++Z3mjUb0RzGM
2pEoOSGIcUVR0uL5vTIeSBSn2ii7G6KMvdSXllmhgAKR7CXI/4PQav3Rw/gxVgnHHGZnVtFFCGxQ
ljCuS1ii+1TKpAvjAZCjHBqHCRIkYCkdfeKAAnOAfQvxlpdKa+VKWPdE63wR2M+hcDKsP7lpVXZv
iJBcKGTlM2d+dLUsnQE3u/Kp7QiFgDPurUkV15sqYAQE5rv6V+wLJnUiy6jxX8xlgNSgBI1L9zDY
e/4U7GAumYi7s4HK51GItI8S7GDH9g43WV0AZjUhsHjtxJWTJSsAGXHhx2+31Rzk5a54O/Nv972y
0S3cXHLw7uczDeJq7u5e8KFIf9H0vUpLJBrj7pNN803evL9NgSkcJeSWTbi8IZ498hnMu+KmlaqB
jjQTPCRmV0HSWIyzUKsHcVGzAK6MdtJB6C7uRtlc0pPJ1VNLZd5pZhhUz77bTuUUix8NkodvOhZ9
pVtft4DMGzLFGnUS07TYwvtriXfNd5AQRve32qNPdzxMIxcfxgDaLrAm+/oBxIfBdpU9IfxD71k6
ADO2/VNAJOu0ILnC7MkxzsFHCf7xyznD6JJXAVCmgDYJw7i/0j+LG8J1iLs6ogLltq/PmsA5ekKM
SDq++/0L5alQrvtqbMz8iFIdCJ2IF0388jdA4ltioeQ7XNQ7Oig1MEDe43M0KHWZJJ9zyn1h56V3
UGYuG9vJl9anxZDwV9QP+JqicAGGfU2Ks7pqxKCJP8V2RFNWdKiyYuFSso0OHyZ8tBw0zgngxrSZ
Y1LggKn7A0SJu1PsSwuWuRn0flx3lGTfEVIVDe9ysE3xaDNEOkNYnQiAAXr7BFiM25AXicZtn/aT
y7czEV00HEEzyrN5NN2FjgBT3bJ5k99tZ4IxlKa7Q6m8L+TgMX3/r0Vs0fLcGq1+htCAocD93Qve
ob1zGj8RwHspwfV7it4CjSKYzbYIbG8IyApl+Kbornf9m4RDGFN/efv9NqkebRFMBJVw3s5E7/jR
G9oe1ZCZkaftXVL7VceIh8Q1nNrl4da47FOLry/D91IKInazcbq5stvsOz9jwEZBzluzCGKYg65P
0Jh3SFlsxNc5tXybptYc/nnVJNmAfXjkfyTJdpJm+5Lftm8qTy2X+yPXMNmIec+TtbcGXx0QtN1W
4VAebIEumR/sNVzh1CoYPM1k80sjs27FsPVEN4kCvivPG9Qma+P7QrIa+49HexxdC6a/1RShuHbz
oD07TzSm935fSeVCAsNn0BvZQtXlFQwCrcm+CqSiFcNp7yxhW0DAn6hsljcx3jNXuXblxh05A9Ex
9KE1uphj3LsEs5lz2c4jucgVAmA7kt/dL9A/Iz95IP9eIRohlPHxBmyYt7wdsQ7bpJA3k7UW1DZJ
Ymk8I3HPUg3DaYOLs5TaYXEiVNSxhRfbdOjLflDn1L9s0HxXAIVcH7OKfkbarBAICMEHSNWNMpPt
SdOdKF7sWYJoDYrL+No6nfHxl9bYNWaz6VB8h5GLvKnaSkLizLHqx5e+9MQOaeZGia29yx0DyDmP
gk917BU1O3Jee27YFWT5dT/b+Q2s0nnNN2Wr+dXEhTKP1BiUMVBhtB3SQ1whjU7WspVUaY4UZR6D
ggqJ4WOu37/SmiMRgyr6UI0a10OXFWQ2omrFoUCBwxp8nKJRbxcZgZqSpCI9UwejUmKxMxuYBzfq
OWT5kO73SeUpJ56nywV05Mu4m1POfJRkgrTd+hLRkZ0L7bQ2/kDB9LE7nGfpy0i4PccPU/qpcp6q
SjaFn47XlJxpdfK0aKwgpnQ9xYYTLx7vFnfAnVfW6eWeGeVIzvEm+6FYul4qOo4YOL2RaDEgAGN2
haYa7v1n/Km6RmtDz69Z2LUuCwKB7QghLJdRCrEpcDO6dqJ2+Rdr6OGuWQkouLy/7jivYyAvg1LB
NlMbN+3gT0hSGMtkIm3rj9s6is4lo5uHkhye6mA4Ch2ZhwI4UgkAyXaZPIdPYM+rAYcm3QhmlRlh
g2SiP4HFrrB6IIE122NizvHsQ0V5sGnt17CVLls/0yBGe1O2GR+4yJKN8909DL4nFpiFbePfPTb2
MUfM6sGMgVRAVAUWuRLf8h6gXXDyTdT8u5m+k/gVD6LQNRePMp8fLXC2AUmfghfhLIcs3dZVo14/
Z7Ws7ZBSbPMfoD4vpW1riHF0ncwBlxLVquRQYl2/HUH5Gl+iJ5qyVDkkpmZMoM3NRzlOBNdtB8RI
rOhGFy9Rtu7KEKfkm+nwWpzy9bSPNfqcMBgLMwnQauXLU/eYSAZlsAF3DSIQfX/wxRjiPOkEqtQG
lv58uC0E/T1gmHWX9gkVDvlKFTEB56tJNBNfJ8EV2nO0DVsJLovAdzvpWjdRA0+rIRpZvGHnFMAH
4fNty0XLYoEOJgiv3vdb9jaAFighq0wG/sHpfOqUEJikdaapbfgBk67JvBvT2OU4cvqRCuCgUvg3
SUIlQyMDBeruckFOkeVPfnFOaSOU5LxfHkgUdUnRHYBcgAs3663+deC0eBW1jvsw6YKsOSCCipuC
TDqKFJBNZFJvxrQW4PIMhIuckzwF9SLZcQ1F++l/L3PUrt1YdREX+7KshaZmx6oZJlqg8x2WPAgF
hohx6lYaPgmt7lQRlsioHo8XMBoKzmoPXM3OWQMs9qWDGPuaP5tn1Tkg6QG5BhnqP8kr7zfDp13S
M/MLD+obpAdHd4dgtN3Qlc4mXdx9FbFq3WvR3pSVoQQena/+AJhrAB+ZpC+KQxOraPU8OZGaziXi
L/er03Gh404F7GQPCWjVjWyxluOAKgM+d+Ag5u2NcXc20VKLZ4mcC3vJ/KyEF71oo+ovo0J0f4ys
314GZTI4NUNiVAaYFlAwKy5ZWRSXSG5U3HbAUnuhCw6x0atOYcrzB6Vi3fpm5iQywDsDTNHmX600
PNX6jEGavJztAtgEgt5yE4poeINSRHwwSW+BSZsNxZMtqGeIFspmqI3qlGXbtQHln1wCLJHlE2UL
xejNEv6jASmccUZUZrMl1auca69UJip31GDA0etMnIKX6Za1RkuZhPpB54TnHmRPqgJ7M29JYA5Z
Kz+/K7qWUMhzuMAOXo5ZRzFeetApNt0Dqgjz6bD1DkzaPXuNIr5fgva0hbYUM+8BQAleQAA2bWMH
E6lQSgE+B5pRBxl0N//5CcHv6RSDSBopEa65wgjbD93RE9qjq0MQWxYE5kQGDDYSOuD3PGpzQZgZ
l4cz3jJnk8sC6QNlgbSnPcaJwFeQW1hkGlsUp3ca0r2P6krAY0p5LYrrw98mTKGmXckOL62PI6Rk
9B1Ug+aYY6M1X9qiCuWlwoLOjvw7TzvTPygynmBRoqp0qysoB0xwcQDJ/MsaSmeQ7iYIumZbDdGD
PK2tAJiFGHjjzFyfQSCgjzpWs6/6zL1zucJj1jcQeCNM7U4cE1SClAOmElAzEI7zlpv5BhJ88aXN
0VwgIygZiJ6nKI8sNWd6XwPj1TdUHThxQEzJ8uRoTedEW7gnOGjAUpdrPzlHqgR9UntJO3pag3hF
DxvnvC867WfTNXRxK9xY/TZ5jREAgr6tncxc+uf1NXmVebbK3YrdVbDfVeDBx7GLQ9xqn4JXLLv4
kdqZmpAmksO1k64cWPEftJumFP2QV9z7VZWAEj6RnJ5cI9nxrbPiLJMYaVDTrmqHwH9JKjnVp53D
WObp8OuJ3Dx9KKFSlxOrU19kY6dUBYhNWlJ2hflvr6jaMIHz//2UmUlJNS+XasrRvrbwK6TCNXP0
Z65cuQNicNbx5DwpNJRc7oT1+TWb4ZXsw0Q6nHyE4O+8wf4GuyCV3TdqXyGHhROEdS5KUNrX5lT8
+SQfpCvejLWBd6yp5lnl3nG+sUqew6R9hYmw2Hxlgs0PuCWgVm/qIay4jG586EAY99EP9gDNGH50
MLomEAD2ytWvTA/yqN1gB9wejiJc0S0tJ/miIPYdGoEEQ8yDhULTaEwKjObxgYkzIahUekKuoXvG
g8TejO9AIx1OxfYl4e1Hz63rC0DoMUhZOZbn6fqoBJCswe0rzYR2vPYjK5J8RB3frbjbRgszz5sA
AG6HACmw7R00HHnYrVm/29nmeRZZrfr2tvME4blkVRB7CxfM6XgQeQdMcSXTVTctGIYG/JgaFrn9
7aWnc8rSKy4lfaF8JozsyhznRTOA0Z37c1ZmlbbgxmencavLYGNwH1O8rE1tAfFgDZVs4x3iW12+
K/CNsXtynws1f6pZTmrtYwGSvRd0/mvpMmp0EBwi37ZkKwOom7wokzsPI0oQo3rv9+ssDG0VxzaW
T0nB1rAKARvYFSqNMFi+buCpbgMzyBb4dUtKPUVoC6ygPX4G6pmqoEq/yNi4aQ9Q4yFGFAdd9rW+
wTHEjiEm9ULnPUyC0ZfdQImufplGiZdh/1Dv3DrlDyA73dsrhKZ2wJPID4eVrvmM/UdqRG48mwAt
p9XqhMvLF/ecQKHDXRHZp8v3aukWOA8wrUP8Xk2zSJmFWoWyHU2D7dovcELMPeBBEM7toi6kWN4V
rV/RccwORpP1OJWuOEERW+tHInwUBUJCqrjaVdGQn7p76NjJGJyBTEaK1HrwEv2i6XSdL5SKeSEz
iwN3yH79g51SrqL1lb/zXjCfb+Eix2b8SGNr2m9RFTE7ePHwAQN0KgGyNZgMloJUIqHLpiymlaCy
pTrESittpvY4SQ/+aC0Y5ULKnYeBRIpmGxhwDwZk5F1Sl0oDNnw7IiupXVpr8dnqZDh7XfGCtcJo
Yz/ZeNlGwjMPrBAjmdK7IPQXvj1Z0TAYXcJLWskzf0eEta4QULRaLKciIb2xwrxuy3XYl5vZuxwz
wt64CSxhg+tf2IP+qPYjtkNk7LPTh6kBK5/kSiIg83vp1ENtLoWmbzjG+lI6EmdIhtaqU5+JQKdD
imBxr8X9H2REL4oSCQgaDtbhMj+RbEJ7uVss1cLWlH80tWQWmI+yLwp5Oku+HE2hGJLHSoLEYP0z
NEK4ObZPwMKboXtMPi47xWqCQCcfa9X+H09wrvkkc/mROBdyClhlkP2xG1gCbcnNQzEDYY2GBEWy
WIoTcO3sshbzu1YHD0m+Y4jlpSmjKK8FJbrrOHtIZb9v04AH3RTOHaepY1niM1KvwXpjHD4c5XFn
8KwQmGxEAeOAu7D/tilUIUb/b0ERqxQPO3DonOtJOAdXK1NKgNU22xU+akOVV07Te/98BOCl2MlT
7tDBoGc7RG4qvnrctZMNWZNfwQHMJPvhsBZ3GOm5qxOU2CrDCm6U2raZP0y4gxs/Wii/7IZm5Nif
+UnCAyDDewpkLpDPYyiZs0+NHXp40oGeBNK+0ns/fLc4+Byi/rDNbuYOW6N9I+I7PHz/Vfk3twOV
VyKARv1YVdDx79icP4Y2VWvk6EvkWPpAPXEY/HDmgoiUvYpGP+J7iA8dir/dtng68dCYNgItfS/o
k/gZpkIKY/iut3HfYq1rutD9JQ/qD2HOSxmwaycQuaovCWhkW5wMlVMbwUu2Jh0AQg+OgdKBI+28
tM7aejqaB++6/7iyvAr+QG5Hlc9Qz5Ly5yq8DKUgrmB0perICzVRS+Xt5w9SPUmB2XNC7X6Fz4Dg
ryS9oYc/uk3IpBaYNMA1/JVD/NBq64F1set03d3VF7jIbL20lQjs+C44/atjMYDS+H1nsIK2eXVA
XgmWSUE6JjYVYs43PFaoS/DFIFDtbqGHMOjJda8dbM76YE/iOK2QH5lRBS65ktMfo48NCtmt552P
aJtxl/9qFnafF4X66cK4vHoKpLg8ZuY0XYc7eDRTICAVDUyB1TMPQ1utOQgSaF76+X653QC3Wa//
nBDTCSk4osE6bO/Nbaj6esZjtRKtzAVKtyTG3rgZJjSp6D4PZafQ6nVxc43XLxlwf3G7K+0goeCs
5IM9G5L/PV+Vf5GRj/OK92AL2nCIa5iy/8JSjCQXIXWopfE05b4ZffuBnHElcRVDBVel9V0DJzM1
d/U5rs3/gxH1YCOcAQS7gbfYaijC15J99fdtD/itwUXA1FZSHmoBsyi+1UOW8cEY48P6Zq/w6ZRE
AfvIQegsjVUKFSNGtxeJ0h0Rq5ji+RnWHSCv1PwOr0t3VBojyRPB1hkZTbCObxaWppj4e3tqgm40
EhhSc7kOvtzQzSQ/t2v+BChzToEOT5MUGzCkTSgVk532XtLMvkzI1ju4J21//nTSXkW5o+phcRLs
pDR7hyNRW6PEO6QBuaK/oUrD4+h2xjwjWDi59TpBGU4QTflrGG96hoSB/r4g6zJreppBU7HiBmAF
exraSumxuhvtgahkXWTABFWATiWIrPCa+G4HPyRyF9DnQv6d9EHd67E5t3bqDSMfbm+ki6I87RUz
RDltet0Sm863s/ME7/K5yPxpV1qrWRAL+zJ1lt4JM/AKnzhOj41d5uCmkqA+Nqw/stD+odRYYkyt
8/evN39D+CgaHkklxmGdYkKRyLr8dMDrCu54knfnNDW/wjxj0HFJpDyRsOe2PHOpmeWD8OE/IksU
ISha2yT5ZgBk9BnbmmVBYTH9WGBLVS1GKX+BPbueMlGpyq0Rm1qyrUq6+m/Or8lcV8S+CVzzyp/L
uLNpxHsfRHmjbMe1UG2b85MVWMwZBlad5vIS/gKqaa4p9NI/93AcEL3ORt8roSMrWd++mHadrF+R
QFhzY/nwNJmXDRufo+G7RN49GfFRUppd6PQJ0vuZ0QdMIXGY83JYzw/sPFzFcqYRYQoH/zvluLlA
hgvx/BDFcqmJuErZ6blNVLeIsKQCcZNElB3lh5Ml+3NuN25oViXSKQrhII/tNe6+BE8PhXU9rafS
a8oSm/84w3gJIk1IXp8SFE28IbYZHLr/W5jfmVxBJAYPmj8sCNNA9pW/tl19J/sVm4JUAU+vCy8K
qLqIg/RmprOJ15ffrxdMSOl5vi8U1W1xOyL0da22ixv9yy+m0W1grBJ55HEwBClkV7xSwA3PLlMA
KZ6l8LM/mtJooqmnL8bwtZ0AjT8lvhFyZD2vweZxpTuKM44Onh0vV6e90Paqklw0HZ22SMWPg3Nj
hVOSKB8jIGju9c9WsmcJhfBT6vaoe6VbXgOotuKlWw5UMXtr/wNbIHfvAjzhAJzatMVaSB5Lss5g
0QUcly7Ym2+tsAYN4wgNo5+4lckz9KJ13ClR108V0ZZHaNaBBTFjyVmiUMOL4g0IbSHnehskomCV
SnA4JZXeEAviVwYzV6Vib1XasmZ03yA4xAzZkfRoI7cIodor5yGBUiwJ43DTcbwwBbfT3wqT9Y+T
BjxBmrJfBFqfDUP2MpM/OVpmioJ+VgiL9DQSzFDbk8jzqFKj9rPw6MEhr4FTufnuTK6lardYc6X5
/otoQ3U7Xs+iWtSB46dF/A7mBeWLsnlNsHfNTEV+tiAcWJ3PDbQBg/EfgFu8NfgF5dH/VYPcNs9K
NF19y3xNuO2/hRV89VDzF/B3594Cj1IQnfJhRYGiny6P945ChrZfkavNCc8Ch3efNzGjgzXQEHn4
C0wV4PyjwW4NoOG74tWwqsJJ3D4OeFwvL8WqNzqLFUGAlhoxxknBJq+qbChBwlcARxWTBrdglV0C
zEmeeX4AcrvV3ZWrbgHzyghzxjGfKrgyz9dH1/8LBQ7I6lGOrtwfwk2dH7ujlzBgo6JRIyocq7Gu
mi0PARsIs8MRhAmnZbI2K6YhKI3ARiYnmVZ/mP8+HFr05fV7invyDMGiwoivmh/avudm7hnHDWR5
MmTb5QkBBkh8t9DOCQocwsiNSFSgP8XJCuqQolS7Sl3YSPP2lTZhI6GAB4GXSlTH3AFSx6r1ccLc
/x70bft/Z2uA0us7ERjC3f0Ii6g2Xiz9gQh5x4ZVikXbwRIzRfoEsQKZo857B/0OUrVqO8Np3cuW
pMLFqAHDfEla1D8CMhJ0NouCAcGEymEFRGATdY9Ucel9hMT1h4GKCWST/RHu0X1/7ktYa9syrgVM
5N0UmvWSuUhyIFu0kynSM0iU7lTW+amss8Gz/UODf1GmXGUQAalgsh+Wegw5i6t8bSLwcKDAVqgY
VB6up585SIz5AN8bVWTSovbVmZwg9vQYAfqbC29NuO5rn9urUTzPrbwy561F/D5ijhfCaH3BBCYu
0QNTHVOq+tuZ+65Gy8J0gQZv9fP4+nMDNMHqdZHjM7G3sUVTCp79OpANkRExX8blOsDKh2L69ZIU
PPVEKN+EClrfgEgccXYg+3hz0Uxr0ccawAuvb3oQIGcu2QGFzaBlbDDUXc/6ob7tvqKSpUaOhVQm
7Mb7+5cHPpRaBvND1l6QDiFNp3yvLX/XCDmlw4+DUV3MZKbM/DKcXERa0X2Ofb8YiN+OgoFUQqgR
FUZqt8uIoZDFGiu2hHqMcbzogxr+QylPVDPoEuNyld0flZW+HgFpO872C/xsOgazk+gkpARp6euU
Rp/wzOwvcwCkQBTzApJgBPn7ChrQcK1jqL9xzoWFLn0hcxuvr3uWZepcEdRkAlYLHTv9Op+pXDnK
qKYU2/MaXbybtNHsZr6nXdX7Sbn4S+zaTqSF7foCQScmg3gUhSh3XRvDBbTypq0RBr9TtOZsh0zd
g7NVsy/N4t89p5qUOfC4cjyu0Js/2xGVOpHtMPJ+69cntyq0zG/Ac7knphbxwJQa5DxWwUFT+8b+
kIf6smxEYp5h4Zf/DJUaweL3qIr5LECb+GLCooZwFLW+9tpCOdmOY1hoMhKh0hczrlia/XpwNpOk
y4VhrEQcxDIkAOsakhVGup54h4N0CbgB1saKrR7r2qUk1MAfOCTKIASM1K9r+WFqybYgpE8GTHn1
SMeeQROwuL/+89IcHyJ7UhInZioL0pJG9o2o6sozrXgA6b0c1jTKpY5dB7zxpVcgQT+DCLHKR36A
dJ7bobT81XVsF/PmwZynwulLcklmJx75sesjUA5/Ju1YHxBcNU0rFBJpKeZuGVlFEHcegIuN0uFv
i90ymamoixQkQea9czkoIQSUo7GHyGYZnT2lBE1UeDR7bGBdUc4h2+nRkaR4LYszHS/VLgq9sgHX
rzfbOql942uUY2voCfD5SRZ3shtNpHK/dT1Sj/5fw9OE7DKsllnbgRPXJ9Lt+AXEhtzwDW2DoT5K
jEAI4pSVN697Dujw62UQ3MskAfsNZEjsOU+y4l5ynp5TSCJbim3C2++iHd856KFvfvFxwVFelW3U
KnHRP5DFdEQjRrQi4kjTD3Fg2xy0N74lr7NJpbE4SJPQAk34ycwbYV7BfTFRSw608zzwXtJtjcXj
Q8pM2clL0RRQtInLAlTNRhLjmiT8ryh5G4Y9XQVLnADY73O9kyaD+OLaJM5U0dE85Lglc8kRvqNO
bNWIhdXu4xPRz7qGV1xh3PJt/AHY4htng6Ip24ipYtR37Bg3xJWM0MrsBhMJwzPoO06o7MhCV7MC
R3siup2qLTnedW+Mics0cVef0hoQjBGEWjhg1SusikYx7o2gaAQvh/NahfrnAFoJU9LDdNPp9K2V
qRZ/n1M6GALryWv4A0C3oSGlXlBCEdG9CvRYs/sFHU47/5JkKx3IwxeHyQsvBmSDU8gZODzEozKl
v+2SsJHee7U+vldZbAvUnZPh7q70WfWeYnsUIEGzoIqNFkZ12O58HlDG9Mu+uiKHiu8hZgNBqjVQ
+027kT1i6o/ruzbnfzFyDxkYm31Ld/yoId9POldBgjGSX8vOM8WoNg1+meMZUUUqLq1WGEpADzqr
HmlRR6HRmYeYGQ7o8fRgrol/e4lpiEM90FPrzh5pE9UBd9bggwiXuBzQ62DHIXfuJLwu9dDZ4zBl
RaX1Q28Pe/o7oS7TJXZoo7H5ka3hN/9nnv+k1l8BqTzSe0A6NChUTer4IYSyx3RSEhPo5sRhGHAy
zNxUstRtMTMIwiZnFEQRvb6dV8HanDb27vPbdIdpkaBrqdJgZZHurw39XXtQbnEBwHS4IAuaQpRP
2HoD7NFDxrJsuul9xnw2QdcWuj6c5sDVyyiGVqwFSUPzPpTN9NBSSwFD6w6p6quMULfCpeWx3lvj
0Rj91EpPjGkwFJCeWkP1QMsSsCQKqwdeazQb4rmuyKsGEd3DMnrCv8qNkrg8dSwwxB6xWS2+BFze
PK7mFEL4lsABQolwg9uPpk6vAFtiJ3ICTUV5czSWiLAn3hkkIgrsLPb2z2Tbw2UmrZB80ejJgJ7N
CZ+0USRQjOdWFfmUab+GJ0uDD/XO6kjQxnzSPxIoLBorx8JG1EYBbaH22VOj/F+qOPlODpvp1nVM
OigoStnqhXPKesRraWvo3/vWZAgrSVX/VB2nJbkXtq3C+e5j0qYuj7N1tEZKqDVmuv+I3UVkvbzw
g0GW2fbCJzjxtIuM3riHDeeUCoCgEnXn+IVl1c3vX0EAGcFZ+jhnVQjIkuw53et2UVfCWHN37Pp1
to6iQ2wAkaYlG1D5uHsbHWbiwWo9X3+pD35x7tfKGthxqR7tk8C0alL6HoAHo3hsNC73bMLB1C+K
BBoteX6oxAS2KmcHjOD+DmpRtEc2DBvkjzQ8qkUTbDKVikrElwCnXI8k+crazffXuBio+EJG+xSs
pD/NlZJhwCzo4RD/nTpd52KbixiSk6/SeMqtgGamNCEmc3EEVovMKB9oErz8VKUU3cAZBFhDFFa4
R4wYMjQF+x7EggTQTWJMS+JlEYOuMGJWCpnk5FDJzlYiG6uvDYtmK3pK1R3CiCKDZWqr+VFu06Vi
1ZPdqMR66ggs1Zaa6hV1b0ZWAEQoISfkEmwQcu+27F0CIkz5xt0V0i9QDl8Ts2zFU0agRqAfcDWc
OfvQC4nx6yx8nakVEmd6WhkAcnRDHi7ocqNtufrU9UUO5zFtk1kznMBnCNjsbusIkGGhtt6/OfjG
Y30XIx7WuRHexSGQ1SHH3mDF65RiaPHHJUPZEZ2bev1FbcFIYN/zD+9Bryc8dpsKEulvyBkvALDO
XjSMXPlaxHJoLTKKoI/U4nuY981+9RBcCXVDB/0VFUp98e2evY4NQwP56rfOWfkWA0GkYIwH3eCR
dTeLSOTo8NhvMVHGHH/Qoq7wKPoompfNQpSRbEcJnLclUhQBzMHRzC/T1d5Y/dxh6IG/YUsKM6R+
3a80KE6NHHrl7XqCz/zsUEnsnMYLDRib9JLeJUpqG2zq+bO5udSuGa9yMGOE4mICA8ty+RDZugTc
LWziVD25wKN4Q9xJBr0Yf2nEbbwlvuZ/VBn5FikognudvNMAM77KiEA5YkgIALfQ2OQwdffj0lcS
T//fiOyTd2t6Jeai83eRp0RIZ8Ks6hkcT8h0ZELALnMchhqJinaZjCK1REHAGQmfgu9Y7PuRWlAa
VvbJ0trzjC+2aPBN6c9EzDDg8K1I7Tll8F05oMHUCwEGx8j+gOVo59SKpY6AUbyR5X669v9VvMHU
xEltS/QhG77g4/wB2YSvFPhZqjmpnTspFd/eQspNKAq0vRFs9G8smeL8Nus7kdOWWPVUKotwrBNn
BrWqjr/NrAyaMBYYNYm2Jfx1dvlH1dL/WNVhnWQeLvXdz5YEs+0EntaDV0nxjb0oL3+06+AyMb9a
EGy0vaoxlL39GdLsQqHcYZLJ3CaGvb/df0kH/QmdYcNFpGCAyHz6y3Ws4q2Uxa4ptZ0EsGAt9alD
bFnplfLB4oH2RrI72iaUsqjrNm/KENsBiRdTPgvZuIJ0MjylorLwjbwUhrUWkVxDb2Mshkhw4Xfc
002aRULlJ5ogsZgbgv+7pj2CIW9B5tPaUmIlB+pKFl4qcaYwuwXwU5IWQnEyDyinJpLO3Ue789Ol
vOC5x1bk9Q/ISyPRuJT52+Se1hxDzFhNxzIStBinjCyHq8wZr+0Ifc/BHv5fUChMHwLhhUuWkgF1
mkq6A8M7UdOXE5flFq8xgjEzB586UZTNLlZLM35jkKuvhzG7tr1/Zuy03gPstGYANf06775P+ipq
hLn1zKI9+hrnpf7kkCfYGX5Z/5QsH0ybJwSTSfFGU//xrcYQT56H2kRR3WFDenMoXjTMJd7b9Sz7
Czr1kWbPO/pHk2NWsECLMJI48vMWMpDqzCruqritJjf/sc6KUXW0RlEj7pCbkDyDwnoLdfpCVheG
Xu3v8iXcPNS5tTvV3CQREVWjCxi0sVJ9inNcFUsv+AFhbo3KlMGXHiqvMWB3Nl332rJ7KWq1mw9n
Xm5vsm+Y5laK2goBVSV/DrKvnTS4nzVAmpwob9Q/KY7Gp3NlshlBVzGsFz8FsTRAqbFiUilQ7gCa
wYRs1mhw3bE9UjJRNqn5MrifnTz8k79SUDk8TaYnh9h+WUm+ok8xBnv+1zwZUdRhW2jiCqBgi8fi
3athGhV9TFQuIY1FkvDTzdXubcT/+C03bhsRSXqhwdgVgrfv4p2i2KkHX3oXpbPAyLIfXPbarZbe
ns8EWKnxOH9jxG5Jy5+DuDcavBdin86IExs4luT2k0cwoVmpO9hb/cXPffrT4NIrj8GIQBGXBmgI
cO++6ruKvkhwckKd1Z111DG6t8/47BNOB7I0zjkN0P7iAAiym0sh6BNSd1oM2nw8BlcgNZmPEcL1
rhw10eVI89H0nX/hqw3E1mN4ugS/JA3OttDFUT/RAPuii1dm+3y1V5zuClwEKwPQ0gQ7XuaOFo/5
Ym5SnY7ccyiuT21wkFNTF/2ZNy5VBDEdD0JOT0/2Pu2GOZe8+hBW7zmyupv7HdJPPwze4G6AlzYT
UR6J4sAGKK5+G49S9NzGpnMPWplDTIwE6UkE089nYnSYh0HMF1nO9YfAlrCcGnK1DjEgz1WLFuch
fvaC0UooNNSmCriTFgwq6+uQnZAR2Idz42uKDybO3a5MVB+G+7neQaRacbJ8QuVGcowY88GjqvZb
3NI8oc8EyP2Z6hgRwLP3gp2Zv2RlXbtzkbcMu41n9Mop7MWG1yTNwvApJkVUT8EIf/c2Z/PgKpHN
10q67CvnrJNP3FMobirDA1MhzAryYABW1aPzHzX86SpnSS9uF5U9fQ81GywdjbBZoE+w4/8MVPjb
2yv4NW0/plQY0q4BqAzg2nT/SKZsS9CuVtM73TEYtNcOOGbosaP62tnWDa278kvDRe9jSRNzykCk
1VKC9CWv3gpuKMQSJGQWG1dc54l/vGdA34ast5KB9PPZuXJmXZnOUY8fz8F2FCiI0PPKAatnx+mc
DsB3RPLaSKveoj6fFwvTlb4D6EwW9G7Z+78CGQfJLP5iLaMgm4YWTQUwitDV5kcwROBnYWJjZraI
iIM/tOeS5+qhipIjpNJRtkwIErXmdx0/NX8ziP3KcqNgyNHdry/1kjC0J3Q97/zolddYy7AblGi+
2Xl3KdYBc4JrQT2c1zpwRD/Rx9nq0cbpzMHbJKU6m+vRP94+5EK/gcmfrPseZm61fv2XDHbMgqNr
ufTHThyZ5Jh+3G2MLGdYTPTp8LBBLbFEZj/VgwnC1EHlUl4orPe3PEUwGUF4je4Fj2R/0dFCosf2
FGStYOBd08BYZahI29r7qO0VahUJDSuSfydTk+H8iB4ZEalYntUnwtTnM3BXPu8SJGra5qwWjTzH
F6L0ILn9A6BonH9SQIP0GEcHVe9OTMDxanRtsoV9TLaJ0ZGNMmjbtyWWFnU3hfYr0QeXVh9frXxc
Bu1uSc7yiwcXyLjmnhquPE6z6lFwyaiJ1pn6Hh3w+jGTlldkRatNZw2sE35hGCqfZLcmbm6us5Jt
F1ut/0k8lRzLyqvmfuTO3V0IFT6PKx9f0J1cZYgrb/DgIBXQH7+1abn0DiXUiVX3ei9M7+kQy7/f
cidQbWGywXQitfQdyJ+Rdd9cCkDC0l0WSeWOklafM4dkR43x0IoypbkbtEOumbHLwLf99ag7sOWZ
R9Sixmuv96LpImOfUwZ5Bi8e4ilav7fM/o3G7r3J4KlNPjkQqfvDOhrVR5PKBW+lk+4zgfD1s/il
FSYgpmTz/XuA3wEMhWrDx9+vRdU2xa6yPWjOBsKe3mMP4FM23UkEP+QTaEcaFQ2EztYL5FpJrHxp
cBqyb3RAj8L89cDOEORQStHPhpspMZxJsEChQlkTB+vHv8ouY7q9EEmCUdaGkQrz2bRhKqY14FwZ
OCsCQ89igm3z4i6w8xmc6rzgelmYaeDNLqqa209FYfGu40U6kuq8gpCYT4ahDsrKDuy6/4rmPaur
moy9oeXyyht2mJOtfKD+BeHK6LT9eJPDQO76l6Uclg+nRf/DcsBye3YVzeer9t7+vi9nUYlkYhm0
LwaU2H+MIKBRqR0wwm3HubPwJlAW9FK/huA9glgipuOYi7FE60hr/AW3LnVVRkocgWvpnyNDEynO
gbGRG6LcHcikgfhlncoRnkhjkphQEZMk20w2BCWlxvHLaXWJmrxK3KzUUZccWFBz3H7aDuUInVvk
DU6E6G4vONIfF/Zt7sbwd8YOdZ3eIVPcReG8AejX3stk9HO+aP2/+XmM0vn4Zg/eEoEeJmIsPuh6
AfJcFS9G2bIx4gikJ+rQ7oS+IG4tcslwBSVpIyn7DCkR5dADcVhM0XUtMdFwreMO1DKHyLJmCMya
dQOndvJ9Ivn+3TlN/q4uZ9am1cDgmHr0n0zr94KbU9RyH2bbEVIO/6etapWyvrjuNHWiGlq7YZLT
fRxXB3q3nWwuSs938edksOAoDI12nbgjipXALOv7PH1qr5ahUUo3+whuz+YCOzfM4EjWG8WEW2T8
+PezLuyfuBTlJzNJcdJD9Qk2Kf51L6tB33xQZRHKDyw3JIefjYhUAHe5umCC2cPIhc6OzQDQUkAs
y3iptcicsqDUVOYjAmChPkcZXCVPV0q/0Msd5gmFVwGlrgKHxqPA8WXf/bPcLQVvX6LO/T+cbjub
wWGA4LKuoMZCbzBCKWvpWIo4ry4RouZ0O2oJt85UBUmZ/vh2peFjYcix7L6Re/dfDyKtbvNT/2Rq
gJ+LwsuP58UpjN0fjQUku37ldgTSEW6uu+wIx5Su0enZgD5VgDzl3+eq/m7J01B4hw==
`protect end_protected
