-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
uFmm3uCxGmgcPgX2AeyJyH1X7h+iLaH5kFQT2ONJPAn9sXzHvL/YCbowNAyIZ8qHu2zvTbRc+1lF
54kqhVqMxpLDRen+Z9EYUqK8QiPBz77uHXD3xpnQEqCKci7ql3w1GYPhn66BMVowU+l1gD+e6vz1
zJdJoriS8dal1X07gVJx0nzyU2XXnJ6ObgzPm0wgnMTnKk4H6/Q9T/OYSuQw3wf00N/WPuuIqe77
Xik4lcyen//61GDR07cadQuwHXLwxbm806++aYRYrMqumGdWvRBJGmQkzN8fYDMjgmtFsm4CPSLB
WOX+rAfiQD3m+WeQ/dP/sXL6YBoYbk+ihbVX1Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 81712)
`protect data_block
a454b5dU2CuuWf+diYBgGC+hvsf5kRh29jxbhP9EYbjyWHcMQ664DhC9yESX/JrWy0PmSTItquHz
Hj3IODV1YH/CueEoJfwu5Sd1T88MX6BjDT8mc5pGeqeOulMM3YtMas2VcnQYwLw7g8Dgk1v7Qvza
S0zqkXy9Y9X3HWqgy8XDAuU4MicB2PYv+PmbEBUF/diqYwDDj9/MzTSGW91ACXQKHqe3rdnEL6wz
5BmJ3Y2Xqnmaum0+z6fNNlpwe6/MBjd3+o65dL0ZJE49TeSAqZzRxufRxD0MExO9GoJ+6u73Csc3
qtLgch++jgLWA+CKR89jWpXzn0j7zrLcKiOT14p09HC+kRZ1BQz/rYvUwH2jpWB4ygUFOxjYbI1o
EP2SIkP8pG+afS2hcjwrG6Il3OJDqpp8yfvmCuCPUmLnImNUK+bnZtTSvaQffXaxckLk3CvtukVE
kg9K+fyov0ZNQul/6iIU+xD/hOwSrUddedTORTQOtGZa+BkYc20BNkPdvWNJ3d8C60Ot5Etb3lFM
Me5AcqHSnXhrAqtvIYKZFdq97iu7VYcQCramczT6kydNzVadR/3QJX+hlOx5dWxYqVMIiWtPv6bO
mDtw2MtVPSxf0hXsZFaw0Eo/nblA0hSsP2DpiBBXK9HzC0LYUuKFV66jPI9w1gXunOXcSCKtDKCY
Rh3hR6deqOz8NHmkAw5TC5oA28I7Luj231bF2kT36thghtLXPUKjn4rjaG6uRxik51Oh8s6kh655
Qjf38+JhEqzriJb/Rv02kquqQ30qIqh7jHHDlKbxf6FU/vvrtXjgZsd0jBMvb0tIqfTrnvs/FluM
S/QuD0pvxikCG1HTuadkgLnordpuLHSWQSBW2oxrV55OleENk+r7yeIFlyFl8J4ZzVKFFBQQZ1BC
slsn6LgxNCDJVPggZGnrAoF4v0RPZwg3j6DkOf6jfDECqTdolGH1C6EVEWGwCKIo9hvhHD8Pj0hi
OOd38BIzInKk5hY2CIailMgp3sr85DX1tfC3P+NtnENalgEOKAbuiU0XqwigbbQVDcA6lgLVtJQJ
qo8VLQvtO/osKjcrmAmrxyW4fIu9xSE2QwcYTlqbrtnOBXhq/URF/0XQIcEps20GrkLjYMYkEMaL
1TTqkyi2A+fKXGy/lnYOJu9AbBuScog2g1D+TWPrCMjpe5/rIxFGkRXGXqhSpS8mqi72WxGf6ruy
t7amZBNw0TvfsE2oWoBH64iLu9ERABjbLPS3LVbdHJuq6BOG17zZmF9lLPcHgagFIuKY6YdBZ2Ze
AbrNDWP1WRHp7xZKYVEPsLMtRl38TGQeSY284KQVRz0dpghP5DWF8TCKnPqWiwv3SkPdzBOH3ijU
/KOqhjwham5MdyW1aXl3qn6lY5OgrWzWmL+5jLC0BCCIF+2AkQjkuiOxZAyszlgIJjVw+CCy1tPE
vVZixSmuu4Ag8c/1EeOtBvwgqmqQi9qLh1QHI3ZDORsWWjExPKOlOeh/R3FR6WWYN6NRakr1yVWB
Eqlh/UHg+OO6LFOSQAhfSyRiqgrz3oR6zfBaBnl71OoTO/UY7xpKuS4ucrF5jhLK781tjYBKFm/X
K7UD714qUSk50Vws81Ox9H4uIlgIhYkGRDngVnX9kshrruusfmV/E02lMdoBro6K+0Et6JZiTqXN
qNlmJk85mE+66F4fW/famFVwoFr4fnqZ+xUPs498xoU3n0i7RNlgNnXnrWvURwOBIB0+C8s5/qa/
n64zvG4xU3L7U8yrqRa1mwDhy5vG1T6c4UMuSGgk1msBHCp0ZYmHaXEctYUfoveRadGo8NKWAmUh
47u1FTSdCRcgTxSkg8k6m0Af3JQGslC8JXR3Cjj4mwzPnPpJ2GcAhBji8CS/bZKUX2AM2PJEEFsG
DkOUrDT0d9wAA/7z+MRgARq+K0fF38rFHzlDbvEUtzlbIXnSoU1kYP6HuUfB8onijemaA3qPzQRA
A/ScoVg/Jk/GoYu+UfTS8UMdPS0DUdn/aMQwup9Hb15RuQZobpx51OxI6fPAiZk7ytV/FTNkcWwW
Ca12BCzMMkqSSmQvAvpZU9MDyP+ghZHW/hbXiLVKS9Ov+iBoWDlj9b3rqH0tmlXI71yBNbTtk5z/
cl4j4RJ/E7wcrcxKaAkS0/ZpjGrr4zb+UoHtJWS7gXbXr7jc5Eab0P2FNgkItG5LbHQopN/08AHd
GT9ewOXWVJTPLnDlH7VnBOs2cYKUNFE+A/1HuMm0Qozpxl9nHBV7RLxuKitY33Fj1hft0Rp68NyC
sfJlWW8561b9vs5mPrtFkhzF8S2CCFOPdoTt/+uzuzWYbntKGHk4gznJyAu43FtLGXWw7oftPT7A
kFvpmP87gNa/44aS7A0ofX/z9v3emcBzjlJKk8W8b1XGhHBkoZ6dt6lNNevtrVdi07xXnPLv7W5T
GkVG0/bd7Jde/qePK+m+/h8C3a2gbFBuB0Acnh+FHO8xpDNA4FXmQudT+7ka6mcxsctmoVOMNU+u
+O0jzdRQZPHeWzaW9VmLNgofBAvFxaeZ6bN5ps3gRA1i1KFgOqMla4nJcNAVJIBIZ0AmcZf9ZXUp
XqwaDfrA4AWcVLgHE53fjxmgX57n1OTnlLmrKDtH9AE+S+hjkIV20PSVnEL9t0GDsDpgJD1GeMzK
JwXMTTyasrdyIqRHThSdlX0zY20qqXK/HcBe9ZnRCD0ZJgYykGM4zz2ca95Rmuonk6GjmdPEjZuv
97Do7uEFAfl7nRxcmDmWT7NvCcmy+a+3j2VBkOkquIIuYaFDqyXrMkM8U3tPEkleq2Gid3RcCII4
miEqnQHeQjyfFaZcvOJHZ19ajcokd0eXMfRik3TfmMww1yh2yv4o0GV/bu14i7V0XJmc+K/b3rok
XJQKGR9foTarA14vlniUm2nYV6phZMzq0iR6Tfvz+3BTcZtNB9IY7kNXl4e3+UbJyQDWpHA6f4rs
C8Ynu9syA9emcVtI7y9kjou8T2ZNy5NtRNYgK9cmBl1FJN7lxHB6pDazh8ywJSS53VhMJho7pnch
tP8C9gc98dfA5PY1TVnL4+3h6Hs1d7i8lvUq2JEXUvzYhRUinSMBiJhIecdFeVJ5+eTwrkY8GoDK
+/JuPrzCCULL7aluOTs1VpbkFuzHvX3gSrQC2azipElrmT6iJVMd4ke6COd7J26ceW+gT2WSLHZ+
9MXBcHOXvE7aEJQ8v97GMlXd9zscl8CmlsZINeEDGIVaX/YA+bpWzNac8ycbcG9XPtXytTz4L2DP
aEDhlU1KTdWH/dCVIpLcqWv7u1S9+n4oEhn8bsElf3QAeTGMeIZwZdC6sz/3fUkW8vV1t8OyqHLV
xZDArhlZGp1I2o9UDwQW760C+7Qn9Ds3a1vcHlC1z2nt0fuDx6qCjslUvJuh6l8rUprg67dtfuuo
ZtJYgcYjKzH4rInMshB6JzEzJL8SdtN7eilOhmT6HtGhM76F6JMc1OBNOtG31VPf90Faf9iRt6UG
/iBbb48/pyUOB7W6vXlhmsPvUkH6dn31KXXc0lxInd2hDDvhw9O1ulCa5nTP0uTpv4exZDrIxk4M
7wHZybNHomquVgG7g+6oMM9M3JsXPDKi+KHg1piiYHG9XTwheI3a1f0YvaVUnCbNCQvPmfo0HeCF
3ZGZHP3w2lPjJqkWjNod102QSKauITYpzDEiFammo1+h4oYwnsZCZKhLhvhjm4BbZ6A3ERhscyUn
ZT74nS2qGY/rD+fVmRm1f4jSxJTa84QAsQmV6Ls7EgJ8MGwLrvdHRMBj3frpMuNudyVfMVHLa8Oa
F8LqxBLDMgQVz9LTFFM51+Scc9yXsKfeoei5ExH5yWdBJ0zveOPZ3OzMY8n6Oa3/s1QUgihyh1j/
g+BSVp4QZEvJze3VxxQuT9dvjtIpmyaJCcOdU1TX2zavDhSRKkheyNRtrOM1UvMHQROsnHfDp4kk
xppuPsIKn/M5eq6nOO1HMi87DEUg6gtjgRdqQ4wXCROuWxEyRT15jzm7q/GDnYG+5Kz88fKm0WKn
W8miVoMxFfg/wLgOE/MTwVKGxKOsXUsEHc5UK7Q2msOlZU6yZNVjGc3JsQNjkSHaGuIss+37HRbk
VgREjkleEHhH99ionXExNNGcrRVZjQbnOe5tXYzmeiEuArM8VG9WaKCwZYTX4ZIwmTCHUmPl77+r
Pwjf2vRVk4UQHnhd0LJPvLipw4leJuqDu3TGP64p3p1oQxYxFkX+pniXlMukJ8BycVeuVrFyZXpm
LbUQ+WfjRd73ymjQ74s7MrKGTEW7HaomY/STTGk0NL5bbBBOPbIq5WddC67MI3GER8awqp8a7PDB
N2ZPMr8WHt6yu9cut+qsbGChdyzpC/AWS3ODRPFd+25KDdeRrpE8AIAYe2kjkjK5nVTaJIpN+81u
HVeIL3Os5WOCtUqNWFLz/XLVjKICDqmNVrjRZe1uA5BLDg6H8rwjsMZqLokgx4sU/tcz62yRjiz6
cpzbOO/4CNJdGfoPkKccPPce3E27D4KnC91KhsWqn9abvf6X4jzJWnopKIZeszBJOKnMDALvyTKy
tMJiade5HSMARDVqJPbH2Ru5hIAnHM8fx3hLsxQYO24yi2qdLgRhY3Vz09+hG1VHMBckBiARvgFM
/usENLgd545fDLa86MGpPs0GUT9DcFzg5x/0gpbkS53jO9vOALUwAQldaB5b+T0Mw0GE3sJwO8YR
IgXXOpMyeRoo4TuFqYsr3BVMf3/PMSeMOP2gV9fcIO3IFR7wWICVcfKC3mgZn6T0M+BPrHmjj1d1
S0f6kiWv/9nhTIdEmHGkne9NgRA8JFiF9d1Iq3gp4+yKEh/fO0Kq2KIroHm3h2wfXIwVGHOQH6Cr
Jf7QKYkyAFZwHLBAccw5WtAhC9Sr75vcdCQsNIsMKp+fBr2aW/nUd4ZNhey+nZBLbd8Otl7txdRS
kTvosI1MZHcKQSdAcBI8bouzk8GylRW7R7WyENCipYxROBJ8hyYm+hIO87TuQOOn64L9ezeuoZ7a
y4sVpoE0KLcVgXqQYucvffrTQvnmG4TqP0HUF+y4+wZEYSxOxOXpR1zdorRjuw+/9Lvtmv3acI2T
3e/G+JXHcQHDG/s2+C2SZHR1I4A8tp3gVxG+PatYXhHX4czeLa2sP+eXnt6DZNQEkYdU9v8bX00X
OolvFYOJlkkO1g7w7s4OKcnWxN49/9idYUUvxyCcGFR3tKmkl2j2f5+KdD6GLtSPUO5nr+I1tm0S
PFhU7D+e/6BxHs8cJqVHPzQt4BooiKQBLTy1ME/wGkSIf3n5GU8A+diMNQLdMchyXUJp2l7leYR8
auzetdYz4+tdXZevxLJaTg69ic/+V6/pTCKGCrDYZ53cPzzmJCkNB4lsllpgYFEkokJaGc3NOlB/
RwcuhRP2HzsjmtyCRsi9o4hRApu1KQKqN1K9KtMwxglTiiYudixqrvAAd1G2+1H1YnvAoecOOuF5
DXWsvhV68RMPqF18pd7vVULTC4lXzGncyfmaUn3zfMB4WMUoeZINhQXRvoRh7gOJ0v01PbAilKWj
UxSfuJNTvmA094Z11kDryEA6KsRsTUZPqsFRqxuQ2zdJIX7RlMWtuwjfiPCDwpi5uChLVIlajCMf
2lDE4NRrGgEn4kzxzEOfLARPcVTaVEJuxKsBDQe+DyPUWAFUvdhREqspxAjj4OWN1t6I9evIAdDQ
Rf3Z9NQGeNGCmB/SSQU/cK2aDt2OQFPTQArXo180KKXpulexLsyQn7pJyoruKVHobFQQnvgjem/V
7QUx9oxkTk4gNuFxL8BiClNR+wlpJ+tn6j5czLh/0WxUpdGmhuipLkj67DsWVfIy35D47TS1SMBF
ZO7u46m/9g//EaXdSe86agIOvD0I82vGMf7upbkY874HpmwlMcQ6fNzGhSNEzIgdk/nbBLE6vPdE
g9ghcqt0mbgi1EO26Wx+ZvQKCmICQA7mfY5jXgnL3cHcKf8Uk2fs8yoI7qHh8L63HPFE7r7EHnIX
UWdhTpSnNMFnkrv94jWORsithAWV8KaR0chjfjh7nIsNJEhLHQm8Az+C1sIWveioxvQGutHukvxt
iKPbCe2DsU0eOX6Qr6djzOKs8LvTNaUCYvhT+ZYgDVHdUPC0nDyKZTdOA9PBbC9V9OulU1Waxq4H
coK0bul3Q8aJRj3fGeNjjaTWS7halYdtAnS4zFuG8+avYr54lBew5pOL8f0tRld0abIFRgw8pzvD
a2CcxTnmR19iLZm8+iFrkKhYgXPUowy86yO3+e1xQSBmGq/bxXQlP9wMFTz9PwxbChAh3EEyDQy2
Q5dQbAIZ+8z19tEwsxH8dnFqkcDEVhM2mYA/hgyd+72r4RDng0H9Mp6mNw1oQA5vL93V4oETuUhk
xaEvhac9jq1Rw3DxeIJKnMPABY8u6dhJzrjE/2ZtmGdu0/GzjNj9DTJXIYgdqlArVkvJrNFwFfPx
XEf75yMAUNMVU72yvMRL56o73gi4/GSjqoeHylKeHZRVV19blWWJvvP/zjh/cCa9QWaVgCqMXnNl
pvHfAtPC+FwlbxT5sKHvcMSC6wI3CrgqHqF/jufuC/8C3WEYBQvCvd/5YrgqLRYjftA1qh0aB2Fm
rWIyqapOj4GCmYnqRCg5bUnwz+NJQclyv8uX2i9FYVeFA0QJ74AmFKa+nrPglvakodDuS6kjBtyz
ttcGz1xaKjV2hmhdKRoCNCx9vX6cWAVN8kFAhurxEPVOXSfaFlkpF0T2W3UJOQlob0k1+L846aUT
pl/5MSZTUcTA1/N4qZ0aQCpWC5c7O5qjkWTKSleWf6mAT0sz50t+L+uCDbZ9Cxk2ztR1TXZFJ/zr
xXNgeTaB8qvdq2d5IKXafz9hTPIQoLHYevT1Xsi8ohfN16mGps35EDIs3bEKc7Y2wctD7UeRdHvR
KBD/J1IEs7IHY1YEZf+hsrebqz1tfbGXlMI6QLXIswT2syrLRr3YDZ60VJshC0JUEoTMRKmRJAyo
daKOdP8Fz3MTDRydunJD7N170kYhuPeUgj0N66j3l2MhOChLbMGOUKis6SZcQquPC6q28vYQePg7
fabDQdVt2WfU2jgMRz4B63DT04N5aqEcRkGm28PyguYxO0leZ5VFEzql121NlzFQdszI/suGQhlB
CmlvcphUZS5F4TRprO1//656728W9jp0GtYHuvBZCPBKhAsdHskyCdizBDemOHgQepCxcJianG0P
XDrDSIiiVD6UyfAuWw3E8aG0EC+G+NdxOsKaO9LRIs/Mqs3lCGzn1s1WHCgHl0PvmEGi0CW1Pi6m
T4B1xpGQ1FSNrBbtYsXwQoQ4nXpBu5W3ZklK4PI4qjB0S8VVe/pA0UTi3FuWw4jOEoWGdqfsrS/O
fKgvmNOmxEwk17/gZ8IUE4RisgJbTzVWBtqyfJirGGNbm76wv/eYr+V80CocCX2OsM0Hcs/zH9i1
s+Ht/2aSYQ8O8ITFx1e7sLZxd950OltVRX51r9ZEO+rH6vFGSE/eUdf64NlrnVbQXVJjRcLtrwKn
FvLsOS+bSDr2DNBt0gywJAldBsE9OpOFUCkAi3AEfpOMvucu8ctnUwCxgpgyA6oaEyKJ0IoAv51F
6zLsGX0zu5rIrLrdt82Q559UBzXuTbxzy0COiTXXmJv7drLKri4rpueZhgPxzaO49J6JJvxsn/kC
R3VtVHl/XYyjLPixTZ8b0d1dVjy1NmE9y+/xIaV+BabRO3Ry2+b9euvrOcQb2clVEeQPdQKdrlt+
iSzXwilAFDkI+m2KpTRcRRNIlqrhb8yKZOLl45mT5t+viCrBK8Sq4tXXSneJNjPstzglzel00DV8
MKIgvxcvkJrc5vdyBABrsN1RqwKobXLtDaO48cRGq5lT7HBcnhPZEfrx/dMck/PPPrBtmXAaeC3b
5rcTfTwsDWObSOo99Lz7Vrz+yhPXM7r9W7c+iIzyFoz0K33DQOMtCMGGHPzHPoAMvwhXzQWAVY/j
KQ3yjHysJ7VEZs1uMj41e/DJVXDGbCJhBT0SKSB85LQWCsw5sgv7SzesqleKTIaeGn4vkOFizBiy
FWeQH/sejJf4YZ8C5JOh9Ps6mkdwLrNmcSfwTWZziGxuDiqtdQtZTUyDSOBrg8MQh/6qfhOWUNb3
+mp7PcbKjKIPZ+fLK+96fDzRDHxZXIqS94bedlDRGpyWfvOwqYziGlxB9P7wEGLvc6ipsTS+3ND/
5iqOPvgiPbxkWqhFH2OyxjVZSvz0JuJTmhYYLLm8G9tNGqJGTa3en+YD+EL527LlwrpHwGazW3Vs
Z8u/G9fgsf0+s8H1yZT3OmHHBTddTHgv9GPydH2Tm8b0dMMY0W+yXN8ZNWoUgQi9i8Ze04opQBbv
dOrhDVPdeaDyOkNS3hp0NRZi4vHk0qQJAEiZ6cujhpNRsFAIqB81SKLK0xqMWHdUTUK8dVUk8WwC
X6VAav1GdU3YopDw4o0nRinoq48Kw51/4P4a8qXPyQvfYCWagm3e+lmOPaqrBWYkZXdRVibVkOGd
zlD51nTPdacGPsTH514GYSudqn8ARL/lQVXMC0sgeZUkrm4Q8wmxhFt55Kh8HwZoRwqjON755rUJ
esrCUff5j6npKnzD8/gI3aM7Gr59f2fzTgAS3joTPZcUmDgNS3LDROmzv2Lf23kbenoXjmbuUL8V
51UIlnjZP52RjjS1feds1yZsrjPo2M0wHoLiooFWplzS4pu56sbE0yrJ/k2XiStKny8nDC8B2DH4
a4yU0/v1Lyu6OrVh+flX3oRQFtkRDM4F7KuoL3PZJBYA/Gu5P1F4dQVXirqbYmipO6f6qBXOIvUQ
FcpEsQ+WBiLCGmWM6rcCNuhH9LsbOjritnSmy9D5obLCOgctUpXOtGPV5TWlcEeK2ojZukHGt8XP
VykxpcMdIaN3NgVA78vocs/IH/qInfB2AJmbeqBvx021yYE5fKoIeAX2kqutVDBnG3V4KHXplXLB
c3iTrjVk1OgzncSQZ0zjYP9d9xbL7XDtqeaEfbKWxF10pUYnD9EcVWvDfziuI1bsf/KC9sdj8q2I
prKq8hBSR+rh5g+3PTZbpcsczErwMmKLsG4dcskLBaKIVz19n4eW/Bafah0ybk+uk2yTVHJtntZu
NYzrdlLbKr2HcmEfs5vLHoyacittXYYespO6y1Vn9RBhwHPsf1oTfkSlOfaJQviXw8Kw65/Na7P6
J7NrTfU63kKGTqAL8QHiblv0rwZ2NvILhWe+GAY5aVzWqjjilDPnZouJy1ZAWchfxl+LFTXJ1UDt
AbThPSewkD9cRP43Yo1FcPLcdp5k7SydGHneHS84iDQYIF+KbmvFCNcWbH8b4YlAclsIKNMauxbh
dHr32H2Y/rD9LLjFTs/heZx+VWwBrPsv+qeqMXozPl8ZIMiBhfeeb33QG3oMFQB24pwiIkcwsSFn
YxnuXA+BV8jJPcoK8WJr22S7EI5Z6KT5nAcTcvtaNga5UC/CY8G5ntCpoLGd6klzF2RGqZtAIkeU
LWnbCbDjwS0+83cXmxFJ142MGMS6ycYTJtM54odWxOVBo8CdV/FjW6XaIveVipxcQEBn8CQWS8F/
WKCdB+kR+8+SE+isJ3wOJGOH7qf0lQhYi2z4CZQ41xy7vvxohmcYOpLJqX70OJusePtgckGmgAvF
rSPY1OVTyX2ybP6TGP+uMTLh2aBD/D8tguMpkmdb8ayux38E3mC4kWhdS6fehWVFVXKOJYcD923h
7evnA5aDERX+wQcl/sxdbXehWZt9QTeuGBH7f+KRtZiInpv6T+EKTeuAqg2abDBRDyMIOXQT7jlF
c/sdJ+L5MSaZ9QNB97hn514LHoTSjjwNr3yTBg1zwigFk/CxHxc/tMrPF0bIQBMF3RQCW+MeGiiP
XLK1mmNF9XSaQ4LQDzPilBJAgbPUkqnkgxk6dVgPQI+Rs234Qct3sF+p2ASb3aTLjnyp2ayxI094
iXaJwTHeCAkOs26x4WmBOjjEh2S+PRPci3smoGd3mGHuxxfhoEgWcRFzqtQ6cQeB+BdhwqH85vSQ
uKOusR1nmb16xWEvynHp6thYH5C/5X3EchuPnV58t9FfD8moGEzRSK2oRzjIBGIC/vvyIxz51Z1Q
fBmCyNejjsh2HQCqcY342tUqWHS37QTdet7xzt/sI7xJEkjIG9FloBn71GAqNyzY6gWrjGg+nqXM
4cq9kEhDvHlVAwhedq+VUAmkPDIEl31GItGcFE9wB5NjZM5DLmmci39qq1q8eQN2KsCMKIyxK23+
3XQGkt0ojRJXwnX76+/6lxvaLlsYpiiVyrJxpL+f3zwoK3HKeb/So/HCsPY4X3YBPhfGNs2EMPi4
3FJDbKmXMYxR7AVLhfwCmkaPdjmA9pWyRvoX2DQalJ1e5nLhQA2LsQy/Hadd0qO+iBafU32azLwE
04Jl//A/LNmiDtw2gcH/amJcHl2d4N90FjQvaP2iQJu2MxRoRzW0CaeTDX5IApqm1aqSPWIB/piC
U9ZH17Ut4JlB9xlD/Nb9ZILBo2LOeAAQvs69IJyDRkG0QVMd4H6JOaEArAp/o0lgUHjpx4GxEgR0
fP2szr34PBqrFhyrbMc/UFDJRBzzP+2g6agoHZkh9Nhwmmn22AloS7Xpfzn2O15kUD17vbRsNQ5e
iqaGp51vIqniOQ5xlFAS/X3L7X2C15nC2bkzCCpYF38Lwd5kpAQdyj60UzzbKKbo7NuJEQznAHiO
WlySigXcaNrig4u3E1dAkrv07XyY6X1Y4bMnYIxc4/qwi1Qqrr7iVjnRHZ4V19JneeCFtrW2tbS9
vyF1oMvyY3jpbSSXzae0fA2H5lXAiUTmo+731UascaKLn0/a5FVo1Vwx4VvuDcY6Fb8uQOMxQd/1
M+CL7m6tAHxjdntHbX7Oejhr+a402RQUtL7nCGfrheDFQrctnMHTaoBEHZivw2P3rzS0RRzBU+51
8eRc8zsut4QTmy6VRy+o5npQHieQtTEuczW5tlCu3D/8HPmlZ5FNH42XPMfrcG9mbMlqh75QgBaX
lLavVDVTKvuPC5CB2xfqcf6u0YJBd+G1wRPjj14Zk7maRxEMpLavuPEec+1K7EjDpTdwtTKjXJjd
enYK+02hoIe6za5+yHSj9ec8XGkQmj8joUCKoR4c0l4paBpN4oVIIRFZMTEsQvCsMYjvqgsz09cA
tKMeNiERxhJqRvGuvl5+IzEOcoVqNxITaDtaa2PURhGAwRRB6wwAkTc7lk4Di4WauyyU4b21+AIs
92RYkjnKyksK2m1CnkSD/Ak7QI4asztdpVJa6F48sllbJbCVb+UzZNZ7rVfrNQp9i4ZMIrhNUMiO
p23ysrCYj6Qfpc0WFyhgF8VAd//aavvQaw3a0Xbtc5N5TGvHgF1OZSv1KUagv3U56AxqX11U1WNx
Kht5JkX+yUBcBiSWB641leSocTgW407Ct5mReAvp4KuAOCOKdK5GWNg4GLabLdohkOWNtHlpyi1/
+JTGbDKFFBEEOYIDQw0pFxFr1y5v6glGoD6uCLWeHChLTusTNQjPCfEC4ZVsDuNg5p4N/2U/08O3
pD3WEd9FLylwK0HB+EmrPUNIqLTLkK9N5U51bsBQfa7ip5SSxjxpuaulUXhF3oYj7stfBq8qdqeA
2vNWtO7X3gaEkpvgeyXJiRjXkwdtxsQ7rGt0Qle6m/IYt5P0SBzfQDtjAOkBjiNuJM1ByBI/oRuV
TFud5o2sLIYvVs5/j6zwP/vIaYuQo3BTHe0SoDAqv3dqxJx0GA4fOgRBCiQhMZENhrSLk404pj1A
4031t03U/+KW3pTH4qtO/4pq+jhRiq2xeCpajTN7mAbZAltsyCzeubiJJ7dhehmHvnDIbtLYWlmY
V03/qY0sSLye0B1QObdkLe2MYtzkuIYppDhkwLOYKUY222gn8FRxqL8vTocq8A8map/nfICywAMY
URWdlg1J/j1MYj4CI0SB8mOAU68Gfc7Y0uCdkroF34El6mgWt4FPT+DX7B5BkIZHwu0BGwm8hc74
qLS8n82UVnMQh31yagO5eqeIA1VSmNkSMzA0awRHwzCs964bNwzioJzYI9sECf4rhsBCcJR0rC0i
ktvVnxSYEYTKNsDCyaqVe2EPQnvo6POrc8/ZiGGwiD/t2yQ5UJcGI3/zKPHOL63ygy0tsxhNNAbG
L2T/dvSwk/lsuurF42bCzk6BS30ClQ1jLtw3J8E0Mv9sH/IfWyi4v/aqUTZ4zo3gDoYYtUvKzGcb
ueZegeK0O4R7I66+R6HWeS9a0v2ZkRM6Kg2ncY1YgpSkREHHPvrrVcRpkXob1SXG6BfAC0vakEEf
OXv5hgo/0HEtnOb0bV3tLHQvWmlnFmaqRapCk24Fqm1ruvB5y4WagR/tQOHQv06/NPXmKuHvoY5N
ecc9dZYwx/hMHJdV5R+gfO7Eapaxf6XMrTxf2BNCF4td2LltgDCWUT0GCj3CT3ZwF084y0biVF/+
w2GewcZt3XDxFfRV4JmEuO6eWQdgdGJMcfWT7G1bUcBXrKdFG3dzrwtIVr7D/kPHb/QDT6tdsYNW
59fpoPyrVvFRxGEO6gfw2MenA4L8zph5GlI8aXFRfnj/sgj7ec2rJ4Tw5A57GXeE62dDtxCyFX1j
2/okPnUWH8rGtcMddfKqMbD9KnzEoqLZrSm6Nfmq4h4VkXERF+2y8NYK1uSozMLnyizkavpBViRO
HBO9QSSUf6hVvQyVecavmPMy8tzNPeYDQK3T0AOQIGJwjYS09shJNrPI5UpD3+NlkzDgTURgb8oV
xupHAAAGhavQCm2bwV/+lYDy4gw2FEQGFqqXSemoqaD7xrLUZC4RTzAr+9/N/5Q11jN/ZpAQqqFN
LgfCEDm//OZBmRHCpeeGkjOoBIL4pNXhbTzDVvAeUNgEf5Z5N6OTujOKxxPDRCZMd5tBARrOf1YD
DlyqZ7EuZfys1Ej/TLWUlThamuErBhZszX6VbQkhP4FByyHiHtsplXpI63HY+ENOUkyhQ0Z6ceO8
YlX9tqL0HrFqafQ/JoXblqXmS/KYTeOttJh8C/zNpsAX8bkmiy0Bt6k/LFiGmYZJis1UJxrZ5bdQ
fBimh8nxeQlUWBjqBQ0zCmQIF49R27cTpbx8Pdo4k6FAC3PuZXvUjiqtVioTifRFb4NWnlq6mwqm
WKKOnqkENZlPiCLTg/8Ou6dUn0qA0oNX0SGaMrPAgNaTq0yK+eeAIjk+b0qqhAnQvdIRXfUJ95B3
jRt4SmITnGe9FXNLfAqoZF7xAPXKFMk9rr9Iar4xyz+0l391tVJMYHshOudjiWw20LM0X2SnK5qs
5gr9VRd3DXuJc0tdxwXzJvhY3v2tw8rTHah+xvs0Dsg2zY4MAau4PI43c1bMN8GfrPuafczQQ9ab
57LbARhr2rbr4mh9xsVRzk6spHzo/nCMAVtvK+skLXQvkuKa3DwW78xAfgI+odEa+W7K3Ijk/g2T
G9jpJlUuI72UpDa/PeA2OFsar3nfYhp5Y6tqrU/RjYxB5MZzCbJBJCJKiLWcLTLaIzf1px9guEms
JryfPpKEAoJIEPDDlrSNqO9ZTUwsSAG8B/u5L9Jc+411eNfO+qIgJXgWwkozmMgruGce9Xoqdid1
v0a8ahEVG5KINkq+jZ/3pPvdDResVMOxWPs9kygOVS6eCDpWu+t8lrpXK4H2L7O3h/x9EtC3ujyM
WK28uqicOAPqLJLCgfMKNh0gMgr1teZBMEr48j/L0gXGxd1M98NzH1D0/OSpQ3eVCzRgom8twSZu
09/DVmS/rd7bX6BBZWPhrsvfyiPz89q5pkossUl9JOGoMqs7fD3uY2ujQ21PYON+vfp+yqoy5kme
rDo9EfXkB8CXf4oYm5vaa56Ugt0xVQZD670bMIG6ftrx9KWSaa1J4nC/W9djAYAUeG+wi9KtoSJD
RV5J9erc0/FtUxn3Cg7+7QmZZ6nIqPZgQY9ViJIancU58Qj0mvg8ryA6zCPgqkmFE8SZbJVMcBcj
/d+nT9F+vTi42W1yr3b+GkgZaVZ5MGMGMlTOtKiDo1dOdzsIcTKIE47M7IhJnH7eufCvYY38gOko
oqis4M3fqGh0ccCbFg3b3IIvtYxCkS5S30d/kW4Mpv/A5kc+uv4ywZ3TPSNnQ4xS30I8bMDTDP3q
/WED1zzXdRmsisY/aNe3Myl7/5Acr2MMk5JHKoWYLclsLPa5T4aeoP6pRWKcTfcQrk1u4dXMDQfO
+vEH6swoDqceX/isZmIn0II58ebPQPCH+IYcn1xScB9fNqVW6Y1wgJi581E+dBpncMqhFz1ykzlz
HmKzfXWa/8igW0PXgnCZ3ryRUBdEgCKvEyoUgSPy2NMSuBIpUx1rUgT2yN/gZfnx3PMMJSUhIUa/
3WCCRDqiPqyxFUhe0yhokqJ3hRqS2Dgvv4QvNF4k1Fx9jVn52kLLhSq9QOgne6sRe4UQVmXDKjLp
MsIzhwqwq2LoOcrz9mHtGcFo6KatWJNsTkIj+CRoXnibmAAxjMj0Sxeyr0h/NoP1hYqnMfU/nCEd
J4guxlbidiUF0h+vS9Nsi5ClJvvJMXHTtk0VkQ1IJXgM56bIemwHXW0Sv3el1iBdSjW243DMA+Af
a6VlM9w9x5vZK84lDz4j2ZIrbV9LjmHqnUR8CAMR+rODT7lQIZ3tLUTZujqXDh2/M+oKeUlzW0f9
LUyM4Ynp4ZvdYUnil0Pa2t3+QGd4c4V6/2t1upQGNqk68J+D/tPb+eGYEJ0/UJFHt1Awbl7GqGU9
RIE1rhqSD5oenaGLwqcYuqL3E0VgwYhB2UAwpp5QF4A2lQ5BhVNyqQH06JIGC0lXMKNov4HtlYeE
R6+vRJmNz1Swpwr8+IlGJ57AwmXfc1/Xlyzu6cfp/UHz3zKWWiaPtZmwsaZks3rndvtOLXyqTqfb
ajs9EizvvvsBfe3hrvnISnlV1aUbx2nakRAI3aiirI0PJUsYnGlV4vy8TH/Dy9KMvdvNUNHPDZ/D
pHQTAe9/ib5JXHF3yjWGxGK7y6LL73YFUAefl6V1DaMQL8VGd2hdmSc0cK30u53XE0/enY3u22Ij
uKk1Cw11AgFF9muoZuTgvVb2V1SyLwmPnUvgYwgaiIP/iUSWKVfipJ2l3UEk1Ak0oC5nXYqHJUEQ
k1RJ4h4WSauqL9IDPCzp0Z5KaEFL4QtWXr2UpQmz8IxkF0EF0IozsNHOGdSPOQAbwC+rhvgL376X
AuAcOPtCjtM0AhL60ThDJZpYQvJH43AvDSlKFWEH4ffdR+rO3XXt/2Stde8jlcz4XYE6KpLNnV2M
yIOPOmsxVPgPu1Ib5pGW2/qs0T4TPbD4UqSbYeyo4cNZqoEVXAgRE2smOpbUVP68q/iT0yff2MZ4
DZ/V91DsOwCHMyXGFTY4Ab/EhWKSr51wiokP48KIjC5lk7+lO9Cl+TkDYJ5WGGZFYrF06eiOxLF5
BS1tntpriJ31BYsovuQ+7wpvFgM4+h9FZX1LoAGjiiqLejqcKCvYnqAQLxhIEB1nu9yTLAw51ddz
yFob8Ll1/vj47FtHcrHYigaeGZjy9yAObGdTmS+2SMQ1xhkRxvibyirXA+Cj4doGvjR/ccxqHbNC
ulEruCnYj0v9mfax0FZjAeoNaEv2I2WieRjyrSn2dk0y4MPTYVBkMUcTzo0S7/SI5iVezgcYd4kq
YqAP0B2SlNQpIiem6nw4IBJzKURHqtSACmsLqrHEQXGxF2Yk9xlr0aQO6FmPciG+2kjjH3QGl4ff
xCtvEP/Uw3XQl0/lnQbVvIsaMggF+OD/G3DiqngsdcBolBSqt0sBeaXafZxOQ0ZdKZpmkRuzWzzg
elLy+gVMM1wgtiP6WYNjhwfwdXzXLWO3FVYSSJEjITUKmMdEeTBwMLrPYK0LWDE6xYxn+kMhOdT2
GTylPyZToVq7JGuolTAkX1A3Cwzd+61kylhnIKKec+BXCIwppppy7uTFsd4Uw9BrcIxAjRmwpLGO
Yx6ePMwLMs/2L/N4c73euI2DLC7P33FHDiqV/G2cKuvTiTpsfGWuLBpbYlYxH7Z9He87RVKPm3kJ
0ZuSi+djfqFnpVoZoRBZZWblJTD5BmuQAQpxy2fT5a6hNx72RBSbhULzTwkfskD5H0FYX78/4ROp
scIvundXgBS8AU0sgv/xBMs4rW2kRH02m0l2ps7Tbezoz91S0OHLt2JJ7EezR4M/08Qb0oZiMJ14
kUCxD080yb4QrdUx8nK3LY/7BtVufoAtbIu78Pk33rKDW2fbDnQQb7yp0VhI/per+ZpISE9CSh19
MlTBYUXr/iPpQz86yNdCHLw/euM21oQCMJnFw4r3mXpuBwyWcotnoCXO7XYXco9XUwkBA687GsYv
Z+R2or7wZTIeqB3fYe3kUX9SBO5wWdnVWNI2Kd+CoCDCKwAC2NIGHLINtGUf4Qeper8jpZ/uJwKB
JDV3zJ36pENfqZZryFkUsThipROkr97IUdKr7BCYwAq8EeAO6DYBjgeV+maFler/nT2LnHr227tc
Ec9dyh7LRllTIT8OntGFcD4ynHKcBtD0piv0mILCnOufbqMZYrZBlamtvBVvhC0qvytPUBrhqUc0
Vfn6vr0TCU/OrCUaUh3JUO3qbwV4tnu4p+96zm8e9nN1QXWWwlKHUQW+7V8OBe0DCk+X6egMtcb/
lmjVVFq0OsCQyUMJdeJY/6zR9fObmoyHKHHjZ+4YvndzIgGyoUIaKVeJ+VZumKlnJH08NCj+oqTe
7VwBCpJovni5rZoGP+46R7awHa1mYoe9GTvhWyfqBCk9B3QzMR+mRu2Emaq3ddE7HS31F3os6qrl
hhcC0T0ybJLz8MiOKGHkWfxMbWHD2LGXAdGYTZ6CKTOCbNciomhSn249lW9M1bwbY2nseLDwkIdk
DyVSaC1jK952t5rNpdpSb1+hQ5HBPjw4itwguzOHWeVzEQg17+8FJVgrMrnhuUPwwwypDAAVWeWx
Rr/a+sRi32nLvsOqhzu3i7Z6zcFQTUFPzaUw3diOfX5T9VZOD4GkiJlBj27umEHsi6O/CSDG4vya
z1zx4lis2+ZUzOsM3OUU8s3nW1zVSyqdzoSeo3GRe/0pclbg+hBXiNcwgWS3O8GbC31bYzLKN+jn
pol3oai7hVXSRzjfFgAQU0HFkYaTnVCN1wT37fQxKKJPPz/RAywJPzB2i10/ml0pLJr2mSktvGUw
jcS11zwD+kHgjIYW7VhjdGjXLV7aZ4eu4sh1PZqM0RyXDg39foJ3iDjgiKuEZn+D/tKYe7TquJF2
T0YBcc4W+ZNlWkyT+fJrIUFwj3IY45r31jKBCv35tLtzKhB8h51u+NQgba4qu6XEMOeECKgrqgxG
L57/G4su9Bia8Rz1TKWrLcan4vt7UeTq3kdEBX5uIB0doz8sFi6uTawoEHCR98BboP1+I3/AEEdh
5mTFu7EGX//tBiIaFoKnuVQBrMdJ/KcXQYv9cqR4d60Iy6HV3EOCnEOispWcT0ixX1rJC2FVdqGe
xZWVWwoUgygkku210mvwHjtb3HKNT1vVmWptfvd/OQ7QMd6JrFFMKUQNTnNEWQj6+GXRPMyo11TR
uXuQ8ARJD/e5Yld8tLdV7l4G8r+VCGsHTShUeKCm+HwN4GeCOHZsyYAJpkDwOMO7MHTzWTldUJmd
ln4y+yghnYY7vMZCflR4etdNfzyZeD10tNv1UKaSrFH5hGosoY58sEQ6/6MUBOjH5RrUkk84rC0b
vMdCczsfLAk6KWkF26luYGLc7I4d+FXzhxRx8fpkJk1GBCq3GGIuo38nGq4OcubJO3mERaZaB7RN
PNMkRTXO/WaOoi9tMD3RZ+H+ktkMJjeKPPr9FpBPJc2nIXufra5a5M9jgoPh/ESPUsstJEThpp8H
sLjr7j4CGOHNvGH+ZOGMbQutRk9EtYtwiwY6bT5Di9/BEbPZj6QO/+htJPjmU0qW8RfsT2z5LIE+
jJH/gv2lEtMlTi6ryFQbpcO8t+ihwVtXsK+sBnV6/ynvUBYJw/rfDIJGTRw9lA3QivV++O1FAEYw
XylchtY9PjvnOjDWUzYv0QQlnPvUiy9X3qzACYYEzcz3QU4pi3AdLn3zp/ga7G3+xvO5s/RSOHhX
cnQ1FQglovTDsZdkC3Dv+8zQSuULdhUE0z0JL5dYVg0f8GE7AONHYLypkwTEOxlfpC22X4i3/UuS
O38lyVy0wwCEiRsKXvkKkJXbNqoebojMIQltC8h8W+dUlSouoyFWdLGg/eETdHZR01uCC+yT+TTc
klCfPGd5L2i0pBwxPiRZ5mU92N7XyqBrCX8jJl2/5Q3VOwbbZHLWyXLXwCieq2nl57bQfKgqjA11
XXfT2tpfqcTxKJnUMlBlj5VEA9xsNaWpLi/nbgO2ITar1tYI7vGGxneu9TAvTUZ13VWiOaf0wuB4
0tX1ClDow++LMsVu1l/oZI5AWcrN/0ueznmgtWqpR5N/3csELbLalSVcBrPCouJQt2AqD5gAzjSB
JsWUSRFYCzKCV431Ycc837SUfq/CC7IXSya/78DDo+nVxu6QyZe84Ak5hFVtlZnVwxtwotnLtPmf
WMDzhfZtN274PbTwZUijfTqoDYE+56+IIbV6dkc5gwHTIBCcfjh7563+A3R3RrOsOr8qaxVVKhtj
7ts/GiVnCg2XJ5H2k2buSysA5QCYfz5c7HBPt4RCtnPxsIufpOy/y6WfHvJzTGOExzDZYW9cpdrJ
rksLBRMOJBAmnMiMYtTqspO83i/FNdzNng3phcjdgc8LSa+JZkxUv7V0cSykYbUTIiaRTRSW/HhF
ZUIoVGfGgZCitIH6yMqeYKK2X6EZw4nR27MjprW8bYYbKLkrPJ3yEbqBa7/9kbtWnQedBmv/MjZh
9M42aCX9tmz+xvlgMCzNLoPonXET8eRIvQz1UADtr6MMieNW+yy9Rj0ARWaPux51SADdUYIaOOrn
PsHusUJ7hIMNNRr8ewh9FvMXL1rZsi9et0EWUI+GzDspr26MC6ffHBYmAaDugfX16juTMO7ZnxaY
DEMhd5wMpq87ZAVRaw81FHfhbln/BqU3hHUDnRUDsEQkL07flvqCFg7mjLmUMivsTowzfy94dl5e
M0AClKzk86It8rHSB0K5mXnUp8jSWp7/OZYnmJT9EuUAlnFNmMrbaTHJr87N8d1qY6BrjK3dEgwr
TNaWoMv6QmIXCltX75z4MVrswNl9guLpFB/8KjA2AYsHHjXLYOmUedWfxlT8tgV4qGn8KGnsIY4t
SPWzVlzaCSCkIvG7xNcQo9Tdx7cPmR6aJO3waGQZ0f7a22qwNjfc3TiMUqAnM2NnU8ytJFp63Yy5
iHOBK1WQKdi+yuCx2mqbUKcoVcPya1j0e4fTtnZR64glJ+WdXpW8UTvmSQrYfwsFuA7CY4PPZuja
Hc10Mv2Cy/ziBBiOAfzhAhTB5GwzfyTDpmo2L/ZaUtNzK039i4Jw5vZzC9LmyswAx848Ep0C6JdE
/j4K7kTna+QFjY/J++w0g/+Yi3+Wd0DYzgy1d7lcp/WiSzfKVZUsjlzCjQ87glYOtZI1f8UyH9Qq
PvlvJejWjL9cd8AYgdbs6TXKt18sCGnbhhkVy1mMg1UDmfWvtF/xazQFgAobRzTyfPJIa3deSy/o
FESUa9H1adIF2eGK+r82hkpj3l1m8qcKcvdwRgbywjLCz6s7JGC0Dq3sfjSwik52tp1u1ThevJEj
Or0k3mAlYBos1K5ZkGqU9pQ3MD2/eCK16egbW2nuTdjhX14zwG4yfQ9V96EsP5NVVmgHCUX99iAk
tACfTvh+NdO9I511hyvc++RtuGwnD8nwUILSZudVIq8iIQ/iFcZ3Ul7jhxHunjeFaD7gVjt+nNF2
EAYV2InCJ3/KU9eDZIlWMXeMGGzxQRqp6LlCdXs1MGe32tjqnjGrf//Vmnq0U4EpmG4LX8l496eT
F+BA83ONlsK3KZumZTPYMhR3E4JIt8CGKToWZJntiphuIUeL72o6nc89WmKN7RvPMuyRE5Qauzur
v0J2FVQ6K0JNLfrq2O2NxFS34e67mPKXDrL94pryMGYepj6xD7WrV/LW/1+OxeFL5zuMn4n6FWSj
ryVbcNFqjTgdAk2B3r6ecXwsTBs3q/T2rWmkb/7akC2An5dF4dDEo5MtEJ+1qlVLivxqEYpnHGaW
fyqU6/C3JDfRoHWEEoLRjcV9MV4xucysEc4kwuS8c+wroDGCPt/matqd8cvyfdMxodzKFNkIzFUD
Q+DAuQYPC71PoCinIgMWhO7k3s1/s/SMiB7zmHLJjiIOBnRdq5aBdE5xF8kpiZJVx0Xq/hpgc4lY
m3MWu5zrdiKrH41GxttBWebVDVKRY/jaZEa6LrAs6kBYCegYNbDs/wSXHWFMv5h1zQwTtgmDKfIZ
MqKc1zy4UGGPMp15ecz5U2CQ5ZuK3ezoqDnbvPcrm3MMJ+nMXml6qLFGZ1/6Td0FHU5N6FO8/Pzd
mzi7ldRAJupbz6dM3q3LNOChTRY/mH0XX1pt1X083SrKRekhvNlkgcGzeTbduszX+9uV94PcLVpS
ObUNNRx4ucj7LKmLiasKxPLQk5p/fX/PiVbyCeUbbxnl0jSulVXW8w1u9Cc1JOtmSWlmdGeALX8g
mA6y3mq6a8lu91QOR1yPy33zSnqaXqc/PEyUm4kdPPTEA3C63gRY60ar4YbdgAEdGAja4Hyq61gp
fAUrXDWYoccxN8lGt+EmHo556weZ4vePu9LJjA0+fitnzuGNhD1TxNqVzyASzoUJycncF/KpVK3I
h5THObTASSM0CuRS3j9VBRHWNDJqJ/YT23UZj6w0OXnfgjKGU0frBwjgjW9Z6+wdwGBo/FSn/RjX
qkrxFbfOrmw/zqEeoQ54huCsaQElZBgGtf7/M8R40uuY5wMMRvEaoui+nXtVBtzelZf0u6P9aTzZ
BWZ6zJg1w/ICFbRcSsuRB6/wchdmf7ZudkqvM1K7Y6skoPoCSJlBT0UD+OfohvEEmx0++1dl1DaP
U0FDwk6kl9Fndxndf60EKemav4AYpDYctiG6I/Z4ZSdHC8vMI2EhokuJKiIV41U+/WlVJyY+SFVI
/Yx2w05T7FWlprFTFb/E20/PFDEWI0eNoNoeHivfQn7YUH08rNWeRRFZJSM9pETcamVYEFlrJ7Q8
jye+zDd53Fxv8FBI1w9SHAU8wAHl1SQcuI7nHSzqmgvQYc1pM3/buR78dHCJOiY0c+roZ+m4J4P/
TpsB4Yb4PxQidL8DYbXOtWnhpvZE71xnpCeLIXeL9NE0Lku8Rd2uU+/KaNb8OArrN40qkNPuVhdu
u4iNDQ5aviNcPJhHdjQ3hK0rXF4gn94KIt4SEtqiB3KJSClvbuU0TQlRBLQM9902YPtPb+MfCrsU
E5/+pL0Z50hjDIZ827NsduzoyyhZFbhBnyiRabYizKz8z1YhsN3tIW2tzBR4Ce15fPlJVDt9OFqi
BbksHk/pVyQWUv91VhWwgouSmw2NCLWwWZHfuLGhLhfVemuFL5gQ0poP+giZHyFVzVoTjCHDFtEy
kDzKFg8vN3PgNAXuOT60SWwQjlAZ8uAIXyCAgQh9n52rFSrQQZJ4JcRtFEGUE2qRyUY2B3IzPJP2
Irnp7sXbikLK+ARBtCIKWAUYno+MYN/pib5/KFCRqOma5tBr3tQ2+2TSxQndv3yUK3guV/yMAG7a
ZYyvNmueAYjCNQVUy/RTpGRYfAxA+1TzigkRUpaNKQMov/keNYYncxwsELHviGf0D33VFQ68MnVp
T2E+l3HpMSfnc5Ft4pHbzepvRFpORpADceQQN+0gbFmcKWCILUirlF3lYFcoUHyFD/SCm51E6O1X
fxf41U3oaB3ZbIRY+0POns/eW62yZqEm+Y2pdnjHT/usOWlA/V0rjfSeWy0AfeKqUeJ9tnVwDekx
AYtkQXsbkhPz2ODHphAtWhz2ltFEKzjQ6/2nCvVPjmYozrnWgQ2cuwC6hvci16QGARCDxAW7I7/i
+eBLDqwcBsD/H9lzbsmIazu8kR/XgobN8d4SujMFJBRM9H24cZXdWJuii152HSCT7PFaEWdsS0Iu
DgzYiq8zZkG6jn+Z3yCwa8nqjIoDrmJFKpwLFAU5jUhbxx6E8/YXqGODyAo5WbIaQbi72zzBLmw5
ZP12iimAMirv88w5QjjHOqFN93mVEDteqe1Cr85oYUFqFme2T4lySsCmZeLQz7D9QJ5qu/9Vw+NZ
lalT3VsqxffYlEExtsNb+saC3WlVFe9Fjq0uNpFjPyPN8uv7rw8krAWPfPMUZR7ztA/TfHqt3cHa
nzWKTUZAEygTPNxDfr0QIqyP/+WWEK3uQupA3mo2agN+W7Ae2/VNba/XZj/QsFORAdzKC6tqKsTO
jlw6ryqVowD0uWWxSLaChQtYiqtZYHMcF4Vrgfzwl90FKz2mmKYExJpRhEq2iBqnFtbNTQVwcYUb
dLgZYKThIECC+OykHyZ1MCUAH7UXdFr6whmjzG96qcoTwStaTGiCcyKTJx3hdDO65Xf/BgePdLQU
kWjDuYOB7qfe5nPtAttT0mpYOzyC7e9GjW2SlV8WBrYMqtNIuSq+F7uLur6E6WKzDJrQiPbnAfFV
BONYZGnfJV162rHwArzrdeozzdZDRQb6tPbqrycFIm0YeizwyDbIUbee+QLe84/YXgmi/NL2jpBk
VyLcoXzhaqHabqIZjEQfkcHL5yBvKDUZbuRQG1VzZuxt2jn8kOWl+J5CAj7Ihzr/FMTbzujyMhnA
T0KrY/c25EG/NQAvqjITRqabAA6j0W6LZF4pvI4ASXRbQcYmrpZHBZS5/5XG+jR+c09lLKkCzot8
XpKYdjNOSw7rNJpKhHo/OTatjEqSGDrCB7VHXC/FXoNd/W+kQrVA40v5D6yR3VwAa7l8peEX+98p
70eFeCnO1FdRf22abpE79UsZFZbzkVzgQkAnxFzfndvvAx8Yi13jaB8UahfQ0cnfHMXl3GYHuZY+
SSnuwETW5VJChCvt3wQrW5wNVUCWVl6lBIn1Das/+s4hofA+JXQXMIHIMUUAcktvLn5SKUHkM1lL
JXCpkJMTFaTIsFFUzUs1Aj7HJ4eXcS1E0Vr4WiS7TW3bOobD1qLfRvyTV7PNg3ySbJ0pCqCp65f8
A0Sl4qoI5ivz9IAA3PiUSkCaoQT7enB0ObpFAOyOjE532hx11+3UjKmOQsY/iKh1nZNYJtSZIzWc
mSHKD18XbRC7GheI66S4zqedfc3T6iza9cWfl45lqcdKBrWo4+914BQYJiWsVsowVvitJVNacRy9
Hr4OxQHgVw6QpJtbZHk6+tbpYHRbJhzjuaNZUns4jSH4Rz4I8JjBqwTvReEO+BgZg2p3hylep//T
PGvIBjN/75aIbncak/+G+FiLcdSPzPihCrMFtMSzbQBqbJclxGqSCkhIXo8PaERFlhcghvDYZpOz
Yqmwf0k7DT+dWIXx3bx2fG0w45LJbIMXd7OKc+GSWSL//Vm/F/RYUeDqiO6BzJrQbQXzoDVxTpk7
FeDuP75lrZvemEfMhDnQ5JTml/RhsX4TTZ9tCot2Gbw2/XLugonnS3LyMs3gZFlxzzrG8+6ipmrI
L/d/GEDQ33YgxihGGV7a4l08w3MCjadMpzjDiQqGI2hPbaGCEmqXFBVsrg8FmRW0IvbwHxR6ivzM
gBM93zz2Uc58Y9CEVe9B2SxRELdG4bWfKgY9p5MxySCvEo5RCkOf8IVcMHD2dSDcJLo8pTakhAQW
ESi0VrwY33YyLfp8BJvLBXboxVY6QdjbakzC9hCMbrZGp3OhpT9hr3aq2pR8o1XOdLGUOrLK0Qk0
sn5jpaVxZtsaFqPSX8pyd2qYpTKRdTw1L8TfEWs3vJ7uiSxId91rH5gWytUkQzPu3qpmIdFjOuTU
hsNHWZQ2mMoe9fSpwWA2VqFJ4TYNmiPP4DsuThO+XsGKSUKvdtSxK22XooA1OIMRcXXE3UKbc5i2
rDVzJOWSqgxu65whugX0wo2IqpBVgVvAOBTc9BQFJnCGaXqIw8ljTzGcJZ93w/OmJ2rWsh+Dd2f0
i3PycT36xCTt6JgmIk05UhsEtFfQ+xVlCklvxEZRnn8c3EjqJ9iO0EvIS90m4oIRnhZ5m5v3SxhP
FKoNiHk5stcWVE+N9QDDjWG9k3R4hgrfgKvnPzrncXbixQ1NM+n1km8lJR9D/gpmMyy9X7LeKC9K
kbUuTu2nK6cLpvNpFTN/ZE8khKWzcGei+cmUw4lq3gFRYY7N/lUCu1XG0XEOl3d5781SJd3mQyvB
plwSUinjCBkgZdQ1aTHyFbpaKk3bJ+v+59HoE+nUg/rA0r3MyhHb2O/aLdpZDbfwB3mLq8BhJN/s
c6WiQ6IcbhahkR21UIfDKsDc7kP4bqf0LjvzDaGZK8kGmok+Tk0LZfUGme+gqgyW1xf2y3iBkGxs
JrcnhVqIIDOYzqKpWBSN0X+LYtlGm+hasLKmgswfpT6pDNRXPdx6CIOO7s4ZkvA81eU5IfJZ+5kd
RJaj2bJEy/qaNVJJdZTXdrlXR7U2y17Wk/j322tj6iSC1tJe3KfWnAkZEad4zZLD5X049pztVoXC
poh3yV4DaDOkq2LxxvQSSfNEuKuewydw1DhO2JVlzghp25vWwdLDfjYFeGXNjtlZYp1KQMWKyPTW
+DtcDbGO3si+fhbKYTlZwMgxTvEdYjEB2avcjhzIHvJRjxVyQpp+tH8dJTZVOzrstLSlk0esNaBB
JFM6b2q5mzXdMY2jtaw8ctOlTf6vB6ZQZCfHbWQ2BtAiRJiRcmDrzDsxeV8yfpzQeU8sqQJiWpt1
a2V8jta8qatVSUPliuGfVh1zs2Xqnqrdw/1aH0XM8la8Uio11bKvVdLNBEn3k0GNjGFgm4gGiDqY
2yyij/ouO9gh/GqJscOIajxutQ7ig4Dw4zaZRORim5qNbpIgHMX45ZBj2wXJcHQM5tiLrPd8Biip
Lx4QHQDcswqSYnrl/MElrDMBsyg5U9Xiql9JwBlD5lPCk3uCJlE+vKGmLuLvCWo+/QYHipkgbY7h
PrTJH2mIiBCaZdJSQ34VgKizo+BpNrjYgpyfrcdGDmSqSI8XpHJPjV4t2gYj2qbPJ24lB6M2kHt2
3Qz8fuIoJx/RHkJWLv3gaGINjhZrYRkHtmDhFd5GUea5dBjQNqHHbQnY9kNea9cH2EJQ8swH8zG0
u+hzoMFTgJjBW5ic3hoM9hgfN06SGU0yreFDY3KzaJVvezEJzHLfW1g1mvjCYrCb5x1LDqyvgTGx
+UqObs5XsnHgi1i2kUmWJKNjlrWpgs4rlsUxq2J9Epazj02traf1q7NpdlxbO/FRuWByd3i3G3Ah
72cOihPmgYG8tbxtGcrNUDExaHTCcwlmIK0wEcgDRYL/fLmlvjA/n0c5LuT1yldMWqyzT/gIXdM1
/DEP1ciQaUA/iyALQHssJi8FnbbctyQWswnA9d3h6AVm5B5Ah4/Q5+Wno03xqolPmxcbxrocU5WK
9BQsbZ7fWYab86iu/YGr1dqICIAoli914gmWdg70p7R7KMSgt8IbzXx3647E629btW2WI/vWvlfz
Xk1VLxPQgobLp18VqY2lwVE0r2mCFLGuMlfI8IPKts5NkrWje/JrT6wB6NDmpPMCj9ht3eYkLVVF
GGsxOyLy/FfEdC1fiqHkIeFN0U1MhwY1bjwzAJo2zwz7rzb2ZBq9t5VSgCA0wghYojoh6u8aRxfG
N01sGWwjH231/cug4N1dOBZyHvavuSBRW+Yd20lgsOZSTr6ONSsSXKVt/RFlJcCobX4KkEx9nJ7n
xUFT8K9Mxhwn3iyBl+Tpc7oTFS/BJsVhncLicCm1g3h/x526yOuX/lTK9ReCNqsjiHtxbqNa/vwJ
AUtEKU/EwOiuiwe8YrTNiobsALhcpb99gJIqKQvDcEcbYLpqMQ1QZMpNQi60RSG1ouiOX+ovFXYH
Mpo0zyUc23du6WLCKJ3E6bOwTxERrHR068K9UM0SCbm1S1DiewCgSbqnYmz2JJ7q5sw7JmpIHnGZ
IIBhRO2Zi+QSZve6OqvcARwtUnWa3845yzE9ntqVmwTHhGojjOBco+QGORHyR6qlsC6zM8PIEHqe
shvfh/naz7/KnvXXzDXZPPCfT/507FYq1SDzgxFqqbVA2xEJOgvcijusJhZS9F5hPlJC27JVvjXF
4rDVPAYiQS7sNFGMidtpKqlaiBOuIhGwIJrhnbPLJ25zyDD4yShVi5kimn5liRqKroWs2Faz0R/h
LTZoCTLrEZBtEqExZ8whtIU4HetaULJUBFF35sQkkVL0zZ2SOO+ulJf5h7fdliuSZddUmXoGNhrt
qV+UWAULzBd3Zk/OxZufWcwvMYoF5n3o/Pl0lrPlLk6NtgByQgC0wUIe0GdsdipucR/eiwJg28nK
6r4r1DXmsHhd8xUHB0sWk17bJbj3jVGpeOi191gTznhrfPubgIOVeVTdOTdDmFmi2UPvcOaoXTco
kn0BoTemdCTcd1o9pb1Ow/LO1tA7Hh2KfOX0JgrrXA7wX3MVFBsd/fw5PckXi9PSxwsFab918qaN
Ko69MtHsx9Ds9K++SQoTXgC6ThprvM8/WuWXAOaniWHSkZPywP3xvhZFej80CPCru+rSRTKGl1PK
moZNU6B3+TeKT/rfvfnosD+ld8JQckdq6YzI8z+fyHSN131aDn6jhA5FXi2RbHodGXH4K6GfyrMH
/x+mb/1LidROTKMAZi1vpzbiYEjZFO5E7R4DbePNQ27F5XSOQq7fRmKTbKaZrdJ2R9lbZdC59LHG
knisgbsnau82bmMzsbB4c8aIBcdKfVcIIYd0W4Edt4DBqE4/qVcPxapp1zhmSwFozPwcbNWjHKXe
mZBHChGt3/w8BMgIR3sxUnrvJVaYsf7u/jPkafP+JUazs3uF5GX0/Tbk4cdFgjtsRkPiTuaoYpJL
SQFsDxXcEhIiLqRfD83cbBGKKKyrfMEtctaaMooTpaSbDW3cv/04vH7A6AjrifjuLMC87tFUs7OF
N7ZWeEFhM1U2f5EdtfDJIB4QrJ8Ic4U8afu0Q+KgmtCRu2Ctc/HeoTCkR3ZHFmLJO6Z5DO/TQglc
+wrqP384wvWkJBEA5dus/v6yVBbKUZwrW0uDyecrDTMyD08GDPGish2RCYBzV5XEf+6Y2vD8m+vq
ErtfCw7S2qxFTIyxivtUHoSmJCMgKxs1NcMTSwXVHlsN3mqSmqrPiz8W4a+ZAaLOjiEPeFsYPysW
q1pJFTKyU82oXPveTYUq/qsGP3MrlRoK4gfSjwowAMZy1AbTtc+Hk7rmdVUd2BMcDYBGrspeioW8
zpFn2TaoU58RuuuJwhbCQKts4IUq0Ps0iYCaPPLnl71m/W9QZfU+lGMP78a0dG66dQbKs8wYMKKB
c6MXKIDkHCEhj3X/1ihS+1qnhvLeq/1BoFGGtRhQRuYVU9k+RbvGiLcgNyQH8iESiPoa2Ue/LWYD
UucGmFKE/ofixbeFZE+RlYt1GKfBn2mrCug9ZrSI+vQJeRk+Eg4yc4I7+FxFeZ+r+L9N29BCk3PV
1Azg8lmKZnOJck5wWmACwaqOV/7oKVYbGp7kMaVNJ0hix2VaWJYcrZmr463/Jlr/qVkXckp9vnbt
oIfCo/RKnCscUCInjsduwLCEyXIhrVLwqO8pWMbb48HyGZD9ydeY85Yvhq46v0WIwUEoCCHMavI4
AxCP9x1oRFDIAJ/BkHetTSVu85Fpxu+98oQX5csQ7+fCIegSV0RhP8RpIT3sSEFOuwmbvzQK6f28
3LcaWmb4uFdpHP+n7DbHEaSsFGEDLd4lhRuyD2FfeqlWGWP1Ele6RzlaFhcvs3lbtC2alvgV1JCz
BUinQ7ihSGZNcR3X5KhksEFs3odLcejJgflKlz73AF1moXAs+p39Zsc7MlM6Ofd1+rZBKOOTdyF4
D2me6lZsDr3ZLlxGE21R1C4P/dgRxJADU8aBqHg7t69itiUv5YX+3Fa/mQOCKLvUG1I7MKObaRtF
hIb08ki1Zyw9zH0HgW3RREwShMsdIR6u549bbVNOGYx+kOuBfQK7NuJE5lLbj+Lr2Y6CClb17URu
vhJpQKQiTn1mY5tcwWpfeAzWaYqkaqsvaXtTRD4NMSQsrLQvFJxLYP+zebo2FTzunklmP33gXDH5
rn/ExGHaaGi+YDrU8Z7eYwBkkQOQJWpQg+NpdF3+jnxW8idcyw6GOKBW1ExHHeH/yLMArtXwX5zQ
30nrhtmYjAdPy8tGzub/xxVNQJX9TE3E3MUjxG2R+3EHBTdtOwqqLsYMj54v1RMWt7K3LdR5sTlf
gkMf4zqzovLimU9z7JkSTMEpQ37hHRdyX2Jbug2HqU08KZOvCd4W7RG5b+sdpkfAneGfJTSCtcaT
iYqiiM0kRENV2Cd69BfZChl4oAD3fBfQnGelfKFOpco7B9AxpJxl+k666t1it58mD1Q/Cf5aMGLZ
tpOg6NWx92Zt6BqcC7LWG3zsQQSVFw1dXvE1fH1b4eeuXNVATv7dRxTkfmoDsK+NOBHuc8DXJaid
7K1uDIMDfnVlk0LNk8/StQRi2JN3id4mIFZtDp7gUIX2CQo8HreDqHYNInNOzVS5uqoPxvH0R9Lz
kWE0DWTUrdMSgiqWcLYh3pYTmfOTeyjF6y+A/nGI8tOgmC259GwTa8kuRyeS9FLjpC9/wg/LIFt2
egQymdzYqH/Q6A17qjaVHhDjc8kyiFrqNKaRYshXCb+8+N3EM+DAB6R7VUsH09VjDAotQfSAvHGH
76q/tHibGBn2FmDl8Vazz0mV4eM8a6xKSsU/X/u+rKjabKMv+1gG65wd6+EB4tckucggHDQNsvCd
rlWnljS+tjUh599yUz97o3mqPaQGyzIAz6jZ/jMHS+IWHErqpc2bLemFemCy3mSdTBN3Vo3HzQuV
uQnnR6oxAlCbs1tNOOn1mUUD0JBMicXEmuZ7+F4Oo1/mYyqeU12kYEZcOxD4rDExjLbYUXqpjZv+
MNPT8sb2MsXmKXZMCPS6Cu0nJ7ZmC1X2f9sG3Vd0MRSjNxj4I2iNfkK1DchrM0uGdc4/gmB6BWtt
pLtx/eBUz+tKZ0fLKYX7xmDfHnf+VdrZzl1ZAqicu5ODO5l1EtW0U4tIJJYAnO5PQ499gjnOiJoz
YCcQ59cssUWfxqAGF7FBulv0UJuQI46AjOwVOAEJpKkzJm4mCwODbnHTNAoNypP4VcsclKl5b46Z
sto5TJEAzlsIZtPVUAGJDSfDLppvKr+c18RoTlo/1JKSyTNkwPF7t9aLWrIeTkyo2KYGH7fBV0Uu
qJNAQ081rWGUUoSFITaWL7RPOsCS4rgHf75LrGdLRs5AliUBw4jih3Vm15bHD2pjPHZXa9H9X2KG
juhWBRl0FUB7Qdv2Kh4Lwl+RzQIdpBQPIcM19FN5gyjyqAskM26vCLoce7lkdBqh0qXttU4Nm0Dj
CGxv5KRqF1mfTPvkRlkP0/Xu/k4LVobLD9Drp0cFRpPqyMvdPV5iEvalsanarWFBc7VybFN+1fHJ
rY3jrsk7pNm2MPQmanvHjg11/1d4iKjRR8yFBhXzCdy44eGylG4xKC2/xk1stxwCGMmNQxIzXz9U
PYFwEsPDXl43UDC/GBStGyPlKXASe5tLSnU0H+xzKfI2UUtMA19H2n5D7IgFlsr6LRiGZNqx196S
4ZRcLYiPnZ41qbnJKWkzkNg6wEfThQlaVAyiDJqvGoDeZG9l7ZPNMg05nuh0Llh4fRwq6Z4mDddb
srZscYAAS34HSAG9S9bkQorznaM3Ba51NQKIFM42KTcwH2EdYUKylVGKszfGJwAmKG2g9E1RcoVE
Adn+YbsHPl5V91RuOiTGS5flxhH8fs1mVJDCB56/O14ubUgsYCN42AVGOFXignYoW3cVXQQ+zBSK
y49Q/fpA9x1lnyakFKwswsR1GUlH6arsKY8JIpU0m2KnEXJJglFztcDUI7WSqcoWAe/2lBvhFQve
kVrsrE+llMezQT9gxx0mmKItcoj6RSxHFuXrgsNoX2LtzcYV/RjivClZrF1Eo6wdzWjjg2/i+5pi
8SHtsNMYgWoRu+wkaPMexa7JCco8mEdAF16Sp/YyafW/PDRqbRQAii0CiUfF+hEdtQ+mT8+f8yaA
q6j8NugB4/RyeUPL/jCatSFdB3GGSjDsB2oOW9OGAWsZKti+5cpT0IzWczJ6b/TNc4Q3cefsEMv3
ZNbLsgxtvvPI0NBC8LLKP9Fp8AM3jK1aihLAmhp84MrhNTMlDosrOihKxd4qKV0MMrZw0raXKfD2
5w1zQ9IfgiVoaDY6nc6zlRQQYV8bq8IKIx/xYCrUg5yNIEMOzzAMN1FAF7dZ4E4H96yR7x1yCAcO
spONqVQsvHz4ZnHKgZEJX852QcUrdFng9RyEClOZf90OwVDMjudqn39oRVXVrPtTI6sWS15amU3r
ekc9cymJB7/7N45+z/x2zwRbByf3ZtWr6xO3qPd+LehnlMvyPbeCzYqR7U3gEGAOlyGmEAJjUKCS
XhnsrIKDjAtAmEw6mVU3FS4AHjvZukdoNr73rQCbHJ6CquHjBaPZ6RURumDf87bk94pMxgBiOCX7
iMXwPdCdPGhbI1/l4gtwixH/yjIaeZYnQ6BJs52hCT+osA7ZZGdSgvqx0GLdrDTTCYZRH5bQWelH
35ZCT+zlIu1iJZYSbyjt3ISfOsuE2F1ChL0kAM2vCqUfrc4vJZnCZMkFR3wBvOMWi/vxUTtWuvx2
UUya0XNukQyaoU5Z3fs4axKFBROEz2ZWnUugclcxiI0klHqzn05LyC6jTZVKhgEwmDIBC3IX6gaX
rG3H5OE2Pu/IdVnI5130TF9nmu8Zftck/86GPQiP4pX00Ki9VojwVcU+obeBegqUVknMR1ptlR6U
MBoE/0FLoO5GZGujfk7yadD00b1Wx1ZTROV5+x4KIV4r2cJAvxTsb242VXvbH/VMo88H/w7lEUiD
/795IgyB0u+ENX0G7VIhM3tU4aPPhtkXwqly/Xv/4SXX/M9ZLVHkDUpLYg9O8CLZWGog4F2nf8zI
Rv9rOYwgqDatVZusiWkLonBPG/AAhB/Hi88OaipVec6zWaex1F8ELp0fmCDnD1Lb0RPqr0ww8fxT
OsYYnRQFxccvAU/GFwFL6QfH+OCS5cQH4S/4UGFvHxZuoP2K/qao/Dhu6ACgBQntvcL/GuTFxKv8
M+8dL2URAVt9wC00ywifmBvLA3QnZ5xsHCT+m4LdIyJVaT6agzBSz2DKDT+O4YdBHqQ3FB4D8UO8
Sn/gkYtSUhBfaOwMOD1/UgUOwkOBI2xVK/3a3tV4Yyrg3HBzGpFIc667pQ7qwNoCTFRgUV281jaZ
tPqbfm+DEB2GfA26SzlivTYMPvVwEBTL8h6z1vTJMVzEQ8RvMpayCWp/vnIgeD53jdy3tWu/T/sl
KeUo5mhhaK88xQ/hdf/4gbRZ+aWcwXNDFEB+thNWU1o0ULux8clmWg4jj4jhAeDc0evnqTiuy7dn
s4UAtGCQbnebUujIQvu/0ZcTj/zRIQeQE3wevydHF+akGegdXUGCnmcmi9ZXzSH4s6TaiMfKjF3P
nmMq/FbI905WQWr+B1CxCgRQ5jM1qqcL4OmbTjLSoqOzhwnT9zsPDHLYXP+uyQZbcFFpWZKnxdOB
/1EwyWoGXF5H5XfBnJaxOLYBnTTptMddsAHDIpPBt/Vkq8H/AOfQwd339bHawFM3YtUQiKUzvYR2
5Jc4IPanfdahYss1McVBKenFlNkHUZa2gPdFBFu6tBuo5eFr4vFYBFC6lLLUhgKu5BBDFj5C/Ual
oPNJCFQebALVD1EhJ4o+Shj2qvIidl54JJdC/qe/KojlZbzVi9E21YooHhv0hln9oSFQkV1Gc8fi
iCzRgvraWZn0doujUSxBTuBkBrTBQkZOtHF4Oy8sHlSmwZKa3+RasnmkOvzMJ48jcv0Dlb+8ZesM
sz87sq9ABJUeMMS70MSRiuCjmdgyshoFNVUXRc2JU10xFaO8AVZH7QlFZ52Wp9oyjNn0clWBlfSu
QtfexMkdIzyMrz3H5ZOC5qlVJ+cOHZEuU4X2dYhG+ZKrGF9yMq3hyQcexIuyPYPqx/pxBgJ53xch
y4dOSq7Z02yNGCrJ5kgKAM+PtuhRlsMmmfxP4L+vmF1jzPcb5bHfQ4S+2hA0KEKGd8vaEmYJgmzX
FW8YCzgOaEAGI0PYQxXB6/Fx1Lgc9ljeEgqfSGyYIpB984Xw1mOMSvRtLt/soWJ8U+1ClXhp6ZDY
dUltXakjuG8upVhumeUDXt5/B+Vpf1j1KsM3oA0/q/GKR0i9eSYvAtXcqkUlQd2IEOQdpuarGiGk
IlwRIybo5j+WNCQ8tRzDsifAcb1wz0yEz28GBls0LnFlm/gPfiz7FIIznQfUgdAfxn68gHhHlpSG
slD+nQSiw9YalGt+47kBw29z8tWmqzrgcJxgd2fjVDxwlf89PEMBl+hGyhK02Fw+HnfjjSVD8Viw
DYqaMRGpmkh7T7Y4sguI9SkZlru7x4nv5AlIKac5mqAIlAR4WSvaUtjTSGhfMph6E3sYdmJws7WP
ORUwbViwS5d+26xXnC7cD6N4SXVbweH+ENDfIHStozjpAZ1LGAGzDPFJq8yvUE6mTUOcOzstyBPJ
nnlMSIR9KBLZw7EDo+owuafdmBDUfS/Z8Ni+bHXsZVSmh/R1DgLVj11fOSojX+2ffp6L5xurg0lb
+9rDv313NWf5DnZvkO2kZss/yAgBU374xjHkQ7s7ZW3xqe0GdI8HwQNQL5OheVXgu8auaGVu7wVE
esZetjCP7PXDTNvwMxP5bEIFx1S3VhQHMDrTYhI1iU442ZMDflLcELzF1pF3RyytFtxI+HUZK+0a
RrBO6+ovEI/1cPl2chLVC9GTdzySCoMzR0ELSH5+OwWZq5Sn/JpHJS3ClWlOb6Tl9vX87C1GxMcM
OPlTij9rmTMBoXrD5eod2pRdyBd5ic3mAyH8vDuHSTt38FC+gt9mtIr85kt1gC7ikVwBII8MMNm+
i03LDvyGO5RXJZQ/JAzwOumIE+ZTbINFMeiznF9sHqTuNdZDWt1gMyW7YZJBw9GFoKVgpXNJiMAq
Uwl10usRqKkCI8FESfw0UJ8/U5gVLepZ5MdSk6/OngGyl6BdH4PvJ3Rnp0z1J7OumASzZkEvBIzM
lqKjtJ3aQezIyFoby2WyDezsQLq+ObirLgbffRa/MXzxXPM55Zaoqg8KI6JB67D77gxRZWYYgR5P
jtoZRxauUO2x8Vosv19SxBryEt+X0mgcZm4J4fTpV3VcGVEgdc7XeVxlR4BkLcxlr8Fnt6VHYU+u
j5f3MpaD/uaXQyjLOU7yaJEzP2ku9kZSw3bFGjHBr0nH9OqVJXqdTze9dNqf8sZfMiYht+UXLcX1
z0TI8UffyWmJLrbbLGlAtZINomQO878i2Hviqx3GUPwlB+mSzN2V62ghajFFARGxZMUYNqzE/BHp
EOMMchavSQ9kWYmGklZxX11RYXlqpLhNgHOX0OFZo7/UQRHRGHi1aW8zXC5UHpPUrlVZ4xGjh+Jk
mlkf4lGKN3Vrxzoe1Jr5i7qGXT4Xv1w225bZ48WIVIK9wh5WTWbbGlHKXLM8HInYLBxBcfd6I4LH
WqK4aXG9TlQwZAzcI2+z+MZzU/h0pZsGaC/SxkyLQ2Newa5wwrUYlQpAhwgNwLevVtxLmGqDOzgg
Cz9YqhlzL3bmHNwagf+PCy5P52k9dHkywFlUW67EEIgPMPHGgw/aqUYpSrkDyWBLORTaS9c1m2Da
0yLsLYWBmt0t1aT+1CuMHE2EdX3/9SOlKnAHOfHS3934suUpAuWDWnTYhL+IPdPu4nHB8WSVNjLO
jfJw718tFTcP94lYhrqxsIEVSzsImNktPRNFLkjsXDC8cu1kesfeaOXjvfyA9IbaXdL5B8PJGwKZ
ilYFwws9ViesR3xfKA5B3mVaClX5fT6YPMpqACNXooTcwfpsoK5T0ySzEZ2iZaa6PTI8ExSiwPkT
++0S+fQPx0DedsEVMd0otmVex24knRMKrbSgJwQmgH55kseFkdq843wHdG06VJdwbmpca/iN5UBe
whPhhfa7P1PM+Ogylf1yTRtB1UCSU2W0qUnm+eWk1pL38EscnRUkmqy6u320NcX8sOEgB5V95EsZ
CXvhpGGNYjIMsUQiuV3MHNkzZbebJ/ktNhgFNPQerATjsVVQ3/Ly3CYah8kWvriqBYc1uJOpVQtq
DvK5ow0DFNm4yQcUvWFkRRsgPJXiX7egMNm88A25lNe2f5zDO9fwzm1qaDsSR0Hnh13Uhg7N4N9V
pzUHozmWT3nLnXu9YqHcVzyTrHPDxL8OF3NM7e0rG3VPCU69gwaFF9eiJf0GL4TK4TsP275N8gij
9LgVToIwbNFhJFvRs9+UmzSg783jeuXFSLSUj9dcmG5/Q1WHcxbdeeteFtGnpQ5do2kEBo0oqBJ2
tWmr2CC3ixuyAnIKNaDK4xI+kESUlDY3Gr5g1YufG4k3dsHPSPjvyV5R6sg1Vzc65g8uP47OIti5
BCU6trrLcMz9wppDJUAVlpoMRwZvLfWcftxIu05lBdxLK0SanGwj+IZeaxZClj1cuu89Dzh3hpyE
jZs4CtWsRFN+gjb/c6mmOCXy28ZEhFsctAFl0Tyav2+DVMyBZjFBo9EM5cGCIqIjZbjX4Eh6VOuB
GZLw7ciU6Q7JUc4LBBESje6R6aaJCagC/XYhC+B88EB/tUpvAjFJKb69WTKMexsQjA+NiOlQO2BP
ZiESPbCw9YMMSYLk4vLxbjoXkNUQn9FuVi2qPNm3D/OIh4CUnEjl6s+sYJFu6myZ6WszGY0qnmVI
FpXfyDv+DdnPPuNAqMhcs3KRA7+JsYBwJiWlzSM8xzEhyduUFCDZCHj+bCAp/jSJcWUsp8hr9sMo
1T/66sH/YDA4MejpQ6foyO55MET+JOPPe3LdB1xdDWrKoFbzE6sU2VVm29cYgNat1cO3/KVhwyAF
iFwdhd7a0iYQpFqL8DgjOMPBjHjEyXrPfrD20c40nKYrob9i3ymP1GUEueoNAZ7f+2gHFE8CzfTr
mfNqy7XCGylPrN6BIDsZ3N6FE+jMukk7qmi4WTOfHIQWjm3WgIypwNEWh+4SNp1H1eekcG5y4FQ7
8aNzmGRPxqsk2UPrwK2fNmm8QNJchs9Ygi3VLQnsyEX/+U3HwRQMmQz0WxJrX7Uw6LmqQR2gFSqW
7Ka8gIKKcDp3Di9v9M8KY5bBuQ7+vvBum6Wk9MbpX8AnGawcDJnsjwpNNIQOlokiYOALx3Zy7ajf
A/5f2F7ER076RwxSqVqSDFxJ3tC5Ih3iEWz83YRFFYdb+Tk7M5BdmJjnia0qXMe9oQbhPrR+pld9
ZOK5/2LlqkADkjMDcUPkNsmrjW3WkNYG/72iT4M2FfDah+NfbMtxRnc7GmXqgoO7Mk3LlAhnqb18
ZCmQYZ0hjEkE4CVao5OBQBC2JL2A0E/p4LgyX4hgFUBQcid7Jndrj8psWZYRRh0bHUhuNpL1gjtU
k10SQEz/ZBY1NSZZMzlv4HH0cYI8L2t9AmDp7nX+Nqt7gCKas9TQt5MaLUiqPRCPpBAKYZSsXGKc
//eGG+3192IvD8xvoatr48eJl6n8W1JokJKPWZOBJWP2iiNB5IqGmX3h7fNaWbmdN/N2hEddcs5c
GmrsPw21rcUhW47Z+KUj11vpZafw+wF1P2zZLbuLGRxImuBqKgpOuquEz4UG3PvHiIo5VX5eNcer
n535ofZoAv7Sa6B3MEmvfKCt95Cea4AzuUqZp0SE3SMhwWDv/X33KxbE3kc9vNEFTZwUiG0BnKiB
4+LFJ5anUif38Hi/yf8y7F4Ljn26Ky85T11lZ00DDOh96yt9P8FjkknTIIfFBZJcySNRe8cg11aH
EGq1NodnAPd7vCfW0VTdC/j0/T45D1qVb3DkNM+bNiXNSMTLeZLKBXugjYfFVp7xmTKjyqeyiLDl
dd5gC222ZnHcJm78jIAGdoOzUl5TVIOSSGJcvzh076A0BqbRjHbNV44fg4nxnuQcy+Fya5fvhxie
yVhOqE9MP6baoKQ4FxQe7C9TciT2pJGZWTbPWbZUvMk+ul9R2FmOEhmebxOlUfyfNrjPJLm0btiM
JXYmhubzcI6KGhgZMnEd6txNn+M7I5LhcRqpo4vFQAtUr2WlTNi3z/6U+NrxgnQ/062PaMacG2Pb
i/qPFtVUy7PtG/JsYEfEamvOLMeCk5B/3nGhddfW0wNWQGtbajQPdguH8QsPbE4IqS/r9QfR9jPg
uUZPJAU2Pz4HI1/CCQG37vBzqxU+ZQI7BLpBwtF90oEJCYT40NEBn2D8C1PnFU7YdVK0NEK52/Rv
xh7SIo6NsrhZzdKtKTZgYvqp5xZ4Z9RSLo5RasaA1vJsgxKGuLupEwZyMDMTKCd4mpTW48UKTFjf
XRSvHFYJzZZDq4VFbQ/HwutnoxwDjfAAVXiIFA95uzzuLgqIa531FtAQ7/8+JPKQP0RInz8T//+u
1VlZPvlCZILO9p+cmcbphAyD3CNjh4C8m/2MvbZNf3prdD6d/CYnsSIWrrpCoUx+ucBYG5XW830N
hK14MSsQiTfSweDXXMSgRmBUgy62u40XlzsFj3XAjD4kgqGjA+OTqlSTUyLrr7u70W/YXNFixV+s
0q99l/dsWc/4DNyiUiL9poAYHY7udEckKJ4Oxq6+ll2bZGhys+NdZxSCfZTdJ2qhkPM1LWH8dh2m
S5VYyFveNl6sKHqAbKfYci8MnlJcZGg7Xiz27MnL82DlUDFz5dl3PaK6/38Nx42o8nBlh19q3iu5
q14c6w+eDKGwG1cdzKrPQMOK3atnJ4d8zZIZb8GCs64MrbXfDVqLisQKOIvT/8qnG+RPPxPyWIqS
CIVm9R80lYrkV+eawswrkbKHevL7zsqzK0xzj1OH7v3/i6rAOkOa28MRnCtjEaSc+fnTnTlhr74F
Je6+zqSk++fgTfHZJwqv0elC2+HKS7UjgOYTD0Nve+tbeQxDRbtdDb+xo3kjve07Z9DxbSSb614y
0cbnRYdig2grLGgExFuLmWG7MsBXPLl3aQAs8GKZhdRSwV+vp1BRPr//2hIY5abY+ox0X5efzRb5
JGYWK2Vk4hBQ+lCYHsycffIWlIdJPYj/CCdruuEHXL1MJFdPrxMMb9VFHEKIeHDI+VSPlgt2Kajm
e6xQE4fkFl26NtYNNJ/fw2kIiAiqMmAX4br+Kq1OuMFiS0buvdpHUibXYGK52CWnS+18yNPAfr+3
AiCcn/E2pTx2+EyfMERVL4EltGgA8d80O6sefTbmS29etWFnxk/jxGGTEe/dTQzA7u2AQ+9eRFTp
aMnpzga9unm9y2xBn2n5a0dlFUIMtr5Ck/PkU65YIlBPla/WaF9hc7mOYVPu+S4NMVNJhOpYWa2s
M+BwWCj5X8wUDoNkrTn6UWHKWxioi6Rpd1DqmM8Z2qN4zT+tdc4XGtvFLfMSdUDH6YCpBKZXhuuX
BbSU94+Rd+YsDmcn0dNR13xF4bLaSp4t8bIo82LEXS0MghuO82pm8RUtcu9N5cRuJZbXrz/ZaD4e
smjP4mp83xLel5wyaCKDrhBxI56Y5Juq8w40HC2be5C6uIysd56G4ALsGjnqcJIhVGjM9kroEhUR
SaEyYaB1gugo7jIM4eULMmBWe61rNjTP1oILvFuvQaZK4uHkwMCKGsfd1zh+9KLPmmGC9bAWlA82
URcs4wnrGeb9tLeTrNP5QKrxTTPvIzh5B2icw6YpaHM51eLGY/lVR5g6pHFzSdarQeIMWzGqme+W
Yrp0uKUZflB11L/DykyjiIGI+yQos9UQ5AkUW64yh3Y9DnZYgvv0geCXFVDOmiW3Ux3ZQZbPgS0V
iBK3471KGEj1gnkpu6vkY6I6XKXYtX0tSOFwb+2A+SQW1V3nnmJBC4D+BfasbqScDuobufrdUDrw
Btn5JFaL0jFjSGrouFz632BP/ZWO+gx9CY2iesufEtHoT93vQCP8h11qR9phpeQEthkeJtWsdJ9g
TAygMy7+b1nuoaL61vPswBeWEdp84ud2vwW3UCFZ1IDlq8M+BaOKjZicp3bAtiZdyCvYQZb7A2v2
QPfIAFR0TPXlaOxnfN9bummzIxqWnONsbf0GfFkJ+a2GoZ2CkInsf64OJV1AzHh3Sn0+T0V2tvdN
4TGnVjY66yWfAeEsvTBjIiod6gkk3E95ajxsrVzD2BAoRF3Vt1knIFqjdLgpdlFWor9O3bS/E71m
wCOvDwe8M8Ac8lO46F+5Tpv+RbUeN8xHnP7/8whhVLjbu5ZVkqmexK/BfPABFJjyfq3svb62azC4
b+d9y8fs6vQihNF03hb9h2/9WkCFcgPfBRBF1Jx9vhCcn9eHlzE+YqAKGpoUs8RNHXW3usAl61XN
55bF2nBBWYlhvSGEFv4t46kon7abpztjyAgHq+iCXpAOi84NzI2MtLE28u/NPM2TV5OUxKsGg6sZ
dHra6iGlyxbwxKlBx71+clTexA9rok8UIDsg7WGBKPtxYIWbrfFN6HCAqGJ/xCLhdaEhmEn21hae
YdBJejMH8pSCeN0y6fdfbncXJ8W6Utwxy5RfSgJHjFNqpr5GMhOKANuKayMcVn0c789zBSbz0JsT
U7Iu7LFm+f2KT1dmsrZxrtkb1e2wMjzS3TJNu0y6pbMP5xbpJqKVFcCXQJwYO3HpkrFraznMaPhc
A5AXTJCytu3hvnL0588ZfnJmSL9/XZ9ku4iViaWdl4pQYrfY43IeMVIwgDPe6g4FchfLK/Kd6PzX
thdoAhYX+LGBLFPL4H1Y0+1j3hjG8deYDbWou8xNBfk8p1GWjCEFDSVvA7Yt83VR/djBXcUXMUex
Hf6677QNLl8sFGT5rA5tK8gmyUrX1X1gkvHoL1LQyhjfjeblPmYa5dLldIpFq0iR7p8A0d9nvZ4L
NyAkx/c6p2IoHrhwxpCIRJttGXWHLmIa72My+6SGY4nRjWfWuXXQQGsXIc65ZP7CuWpD4LfGZDB1
BXg29na4ZGCk6Orm8WnQmVwPBS5KzUuu2lM/s7r5Bxvc1A8ZBFwOszJLuNEeZjx75Hg5NENOGUVo
CWpUix2rksx9k/RLtISuEsgZN5lcFOUzm5mxWiev8bDJP8cTgEaMO4d1UsPKn5tsgTRqdSJK9/0X
0Kw1IQu7WNNk5NQUqUMLF6a4F5g60wWJyL75VrHEDFfzj5QCSogBqeD6BH12teZve2+6SIifZT37
53yoOhaagwDVmE1+pwAAYBm4ioqZjC9mgoRuGjQQlytXXbSFBQ6TPSjfYgRNvKZDRguxUThMOBpK
zcQDS7d7Bf0cfzb16mm1Ol2/wnsUJNTAHw+knUUaIVkWP/g/8RpAoSFD/+NCmQJSdKN2TWUfUz9f
rsfHyRp4+cS9iiDGsXamEoy+Vss1sZkKt7szMw111OA1hYtnmrA35wCKyW3WBHN53014HU8saj/j
QkwTsP3NeLK/hYr4WjM/I3ANDBCYjdWhI+x0bRlIRmC6d7LnZ9nNJV48R8S8UYA/xYmO0Mm6TXGM
0jQSqLVUtHpI7L6BxsW2JGEMgJiorMcc6U/V7UBjE35Mk3c/TWLbfHmZhxQBLCLU0mdCd09NnSES
eobleviZlOPGjacWWM5EBkqZzIxgenkWDiZV71unh5z+JumHl95rqaZoBH5QG5yvosDaQI0XPaT9
+n2AGaom4Bluio3acBTuM4fCfLzjA+hE8GGsFLHg7UNSaaVlCRuABES70/nFIBuRuI30UA9xtZuQ
gCzuToaxlWZr0ks7WfXM7jII7HOfdqV0CAUDcGrnh+T8BVb/G6or0kwTgDT19zcB7TocOIupkqku
9Pau4ZrXtse4aINcJF8T0EpjhHx/U4DwVCJJjpXqavDvtbT1VxqmtQyDdd+aYymvVsbMkhgBA1jr
/CmvMvN9neMFqGMzZ0P9/pOJG5tl6rElecFhswxf6LJqe/ERqBrKau3/VOmcsEnbKRf3ZSmtveYv
V763PGeGuwiYXdce9kwvZpq3r4Co+1srvcyWeVds1DJom6gEmJ/HX238hmftUKdhk9StBJUdEWXO
k9GVLlcQGHpf2fcyoutYpXWJcSpPPW3sDWD67RfhkEGiRJ/ekdK0m+bwTAhXrdodx7/ZpWQ7bmH9
cdXHH4A/23z+j20zoqM6HH2EjpJjn1UuSQjO16QHIctnO/O/QBJVIiIhIYZehJLQpyXFHAa/NAPv
gyH7NinNgOFYrzlQ3x647JuvFy3ALOr/JeOJtBfn4z+8apvFXSOv0XVa8lERBa7ylANovLovVCQI
mxjhyPzcG8t6iGmXbprBHEeEQpsRydYvx2+whyVQDVhYgVuKWdHJOf2qTs3g80zNC+yjn/qb5N7u
OSlPsPWGD8lm/BOx2zSnAvEU33Q5Y8XgXp7GcHZCE78Bj8AuAudSlUgdbUk350RQ1Ru+DJPECZg2
/xYYD4xsM21EH0raUc+gAKxluIDv7M0Q4GEGvsbszyeEZ/NLzklxjzUMvo6cEAX53cfSRFAQUjht
Vaqm+cySSwyoW9sNzx26ojHfJAjplR6k2hLSvG2MpiH4d5xiHeAeLk1HB9X/phhHaOoYhkiVhldz
obHcg1VdNYCv1eXiLLACauVoGJEO5NALJBqEaLKTKtoGZtBhwLA5KYNESk/ojocu0IZSQ9ifqkd6
cjsTkcqp++4KYgEl5w03XB5whnRD25ycg3px+t+9WONGGB5Gbzd3ggMdN4NsQlp4nbouKht3Kosu
zltcYh7mJWsh8PxIet1X61zrZn2zwW7g0FAWnRnLgYpx7fp55TgYtNeqinaNSb0Q2d0A7A/A4h3u
Ts8q1sGqEICHdArCn1iWua0NCksJuiVG6GloOMwlu/pkgZhhBEFN/Op2C7N4i9W0m7jBoIKKpyxR
q1DHtOgjDFiOcptKIUyyZlFQeSeNlAlqxiRjRqjHTzYDUPs9Jqs0MZeBBAKRRRQR92D50MkJgLPp
XMy1bEK4cbSz2+jlLaxaAJfVFpjI971lWNeI7IpSR2Z9D68AmZzFBWOyzIl1Fzqm+7B18/hQ+kz5
F3uQVox30An/J2EFAblKMLFmmqnOZNWlfbAd6/XqjlWMxf7xKsiIaGyIBe/BdmF6dYy79zkDmJHI
7lXzmI5ZxiZhMMmqXiQqRqcOH3YodNMzvQd8k0zm1ny6832lNI6wRSTlP52lKwyLRxB8R0r8UT/N
U989R2dyso/WxdLlcJ6lZs+bYXIMcVvD8wd0zXyBl8wygpjgjkSlnoQxdgcgdr03asZ2/6wIZaH3
Ek31SCXZbZOoRJ4BVcbW9/jSKroxl6RHVu8EEaeXO606w364XGUakWGuKkfxXPdh82znryW57SCE
MkValzhn6WHENpjvJNY/ewyUr26CZkEyrKNokJ59aO2+nKSf/2wEsZCdQ02fr1WNGmhmIJ/pcjYm
Mh0vuil2iMUSlRnLjT2dVzRaomNd1l67/NzSlwnPJ4DTGf+XwV+xtQgYzdvcctrHSSk78v3o1N6j
1rKL0WjnExLoD7u4jyUdH9bmSKTnMmelk/LMS14Jv0OCeMgeX8w3kt6+OAhY7AW4qhK7pmE3hfYx
wqEip9lDHKRLLJgXZdzqjOCDWeCLyQQqEBlXcdwHCpK0gK/1H1FmsSjn7I8snBdwBIDSGxRedwEe
cPqBDf/scRdXD4/vWO81UjgUOe5vwehn5haF6+0LqU9DKJc1x5HZVeSYSpxAG9dlufURCD6m1AYC
LaKB5vsFnwF6j2i7eHmNnGjGU+CN+KM3xPOFjRVn1djM81dUrrQONVyQA0U2a6lv98ob+hlvMU5r
pMvDOLLH52MTBsttaonKG4y7b1aAbIZAhtGy6VRjUcmGpKJSgh44+rnTr6ln0q3EFcOaamMFBRsx
F9ENaWtDAQBiSQr3P7RPff9yZ+VOcTborLA8SpYzGrDc+7vTOWEGI0jggAdkzWYmCiRFVVQh02es
e/zL+1NNXTjADCbK1CDqT4ZPL+ClVw3iubKtgqmuSUjV3k93Yx4+q0BTJwXA3QTIc7K0t1X7arX6
RiQEeV2FQul25bJQPqBk1WsZpJn3FBZsmys5wHLpPCRNX+lsz0GdCxs30r7RwF/Q5d0vARBdUY4V
/uIw9vimEjEdsRh6YURcchKVFcdifGXtr6Ew/q30qck1g+2epnwsp5ykjORGsV48IA1HGtpcAbJ6
77yzO3rWqfGjfqGxzEl43v+dOlnj0XkJYep4NS8I0rf4YTBHZ9/Dhl3b9ku6bZY1ZiqVAjPF2BEz
TGbrWYNfZTAKjgVcVk2x7g3Usyp+uDj0T8hN1FH8UabbNF2J6vau5S7TDN5FSuDhm7b8c1f5b3rN
a/o1ajjl/+JCn0WeX+yhlSjVQZvTLt4BXZykLJzYSwALMDHRaulg3BJ3xYXFDFOzkSiOrDM2QFHk
bOHhONq0+RKHO/dIy2hIdPCw+fJTM1qPYe8Z4ft2vnjN8LBGo8NUEdoGaco6pAz50VK8589X7lYp
MGLCCiL0H6CjbgHria3VGE+3oSjl5M5V6DU+THBJafsUSlEah5w9tQWVZFGmXu2Dy2q8jglf1sDP
seglwz00Bu/NVD6UGD1MBHNRDkkviRlwR/LW0sTWBdrdl2BarbB/D1PGJycIbiOu3ZuLvet4R5Ea
KjV5xsVAS9BjP4Hx8xYVI07h/xg5bE89KkmylrnA3fgKIQ6m4Hva5iApRjglFUkwlh8RYtPpMs/G
uVukSjzZhfihDQwYi7nlF9ziXFi1Tj4MgiEkBMjUdzx6M0ZFDSUoMlkbd3oYAUxAHaxJPtLejnjv
NQ6e64fR6LQHo6IyyFKL/p1l8qTQhvUAPbg1I2AKA/rkgMjRvhqh9F/u96Oyb6Ox3s9rjewwD4hK
6oo1EZ7pb8EUFhHbRLErX1jhbkU+BN67SvKLuQtwuF+2VIqLd71dENuJ3YZkohLO8gzaBpAb4bWZ
dwkckzHI5aCKYu3TjdjTV6X1ecfjdCa0mgoeW0LuTtVh2sNktC0GVOLwUIHYcWRiJ/584nyvUiCH
pYYeftJEaqn0n7gikB0/YM3rTcgKMDSWkYlOctU9qj3OAl1cNrSyItnMZ/TWZwxKwcqw2vbaUIwS
dRWvzQbOZ2Nf8yo1lTqhJoUtZcha4nvZAp/9a22Me0wet5F1HcSOLvAdx06wddAPAV+5Z7ad0Bvv
Ii1xkH5y6g3zOnDz7PM3jgtFqbAueDIDp/mr09HPfibaYm7qb1aq/c5izYYBgl+jNkOYmJnMQKBt
ZBgRj/4D2mGcV+jHjrRl2JfmqQviap/Lx7xYVGmzPKv6kjoalXyA1+OrdzbbAKncU0zgKlkFTa0q
DZsI+/dF0Igdy4jZ6MXEFZwfP1zODmgjYL5NrTQx/8dwEQtvKOePLJCGoamRY22ySXvt6ClQMS8I
fbnbT0QC9wyew+VdyvCBMlGEvpSWYta1rE8/YryUzXfPUeWaufDG5sJ0cZi0/hsWPn9RdgN9XRjK
ecBMFxwXEi6fDZeif8SxoRQuLtpyzhgB4WbwjkjXKP4zPPjk3IraKSRhcaSrTeZJDVQrzpzWwzV+
D1hoXwEous3nNiq+Ahmh1CtdGSYP++t5z+Bws2p3YmnkKdTOflGhwrfZpcT4h9nzvlNmHmljTR0a
D7jCxCf+4e98IhGDxigJOi7Dqyk+fH+mhcoxJ1Euiy8r9F8meFNe0T+DX1Qi+PG2/IMCB4ojYjM+
kNZPIA3giOwp8LjH8vNwXem5jon1VyxvYpH5qhqFmDvnDNXHMcy+1pnYb7qZtpYaKP+AIV70v4QA
b408RmdhJQKfJdyjUEZgdqoXTlbkfJr+rNcdhI9h4VFa+vSRWXYEk0/gFtlFpxoClwXqxq+vElij
uC+gDLtLBWIN/8FCT2aVEs368KdW0buzlZOIawNTaMMGtH4fEa7RuVdcBmuv/8lVBUZfq6IlG+KE
Wsui9UPFyeRr69897gljb39HX146/ZPnFgRLg0ky+H24KWzfA493XujNv5BXjrrcnL+c2q7o3H2g
zYF3SLwSu2wIfcgOgL/hAOr187Jg50mE2v+LEixdvikXhNd/pZxKs1XA8DJJEQ3OtO6G6UJBnfhG
ze4iQcVtA8PlQ95AOok05mNQ0Ca8LeYFZZIoIC3a+zuqQn9f7v0SdmAMhNnMQNCqX1BVsZzK51WQ
aZn13VyZYdTSBZdCBqArAxgEGTFjmNbMRITx1So07cCYcAdK7e8mjLhcBCgoALF0KZ10pI3FHHi0
tyS6RErA9FLGuY/fcVu5IDIUVBR8yAnZYimXwVc4T1RGqQZEBvtCKZc2mF7Yq1QtEIEYpf9F67n6
5jRaljE7qlCPqNjqieFkCdrN1Vam8DHWi5CzMA5nJxaG1vA+KP35fGWGPrqixTJT9MYKDD7nD0uh
rE2GxUYlf9yXrFSMyVtMrVkqqux9jNfj90OltmiYODd8cHApblg/EiHLEx/wC9Di6oWeNZfSqiGx
Rc28JPANf/oJK0X9g/WvFosOYHzegpUqjMvsga8WiZQG/UA8pVrgs8szjtZSusIrLWQbXs/PD7+e
84T/QDKBryihT8EL+GkPXYDArJLrg5HXV/5OvYYQMgu3SdhDRayW2pA5Zq3O0zQBZap+UbafIpOA
HRys86MdSEtT354SrsRsRwJoA4YIVI5uR1ugZUdLoHZmScKmPF6G8zQh0oWA587ej/JayeNg/MX/
vRM0BcjdngoksxrSTaoTG0PKKjK2iXRdbxDttiD9QrQjz26rwFhVbdAw7gu7VbJsojP0mZoPg4HG
ghpPW7aZ9vJxXC5gyKPIzwdjnVakUdBCZOc4C6gokyTTc4oVRAOiceY+cf13pYpk8o3Br9IYgcOz
IlyWn/fTu2sHg3Qy+vU9nHBrbJe1waUlANMbp62epjPIsb1860AFFx/8hosZx8MX/wL1XJzFbD05
uhr/LN5oruQGSF7BDnxUTkrGKHvKY0qQYYtoBktZR/ehlNbCOCz3yMtekiCUNdnk+tgKPBG6ZQ+j
fcn4enqvNQkJJpusJwiW7/HXnZWLQaAtLxOus916zFso6tV3Cjs7A2v2Bdue9+jxXKo643++r/hm
XrQMz8ITk5/bA5Pg8H8haPHV4cuzzsNZIe+0GwV0aoJyfsxe4Qvi7ocKUFoCmCqktXNrEh6ghXXW
GIoI5+00z5L9Ok2T3EWvR9+eOtbEYzELkmFclOb+1qY85ErcJuW+qpakAVBALaCdFBhLVieD3qrY
sjr/FDCaikxwKCCqFPY4RxViTOIKaE6GfD4Yvo+4XM2pGeSRJQCgxcQ0WEdDSrZnHqR6ScFHHGmB
smGFG14Kc6Z4PIlsD9KTieNGcNmrpbNxOSh/s/uEyrHy4rh0OZUfJ71Zv3/QW9Pg21uCBX5l/Pwj
IA6AvnzYknY2GDfAeZg1OmHydsTwU9Dkqhmks+EAmFoIxNknZXsM2l+EvaiVkbEs5f8cVM8hJhNu
ee0UFjJxAZH2u8OSSVJpKg0K4eWoOTew3u54rWM3CWBunOLpqthVJ8Ar1ZgR4rtpYE1mzILauDPY
a7lPKOXU60i1uaFqNYA5s3TKaCMR+KStpZguzjrh5gpO/8kYMhZMeFqtzqtawZ021DpeOFxuEBm9
2KsDDFIoNVuJmWFP1CyjJuQUlzJHBZbQ94/J5xqiLjmHcMRruhp8LXtbLrFJAY5qL/d0OTxuSCTt
D5R/sDpOXx8yMuWbiM9k18ch/jnw3ldKATR7fAhuKJdUvbCC0xiNcKkO6ROeFslSNE0aFBnt6Ikz
1qza5uq0q4rguCQNfB2mfvMgLTOs/FKc0Yl6ygub2TDf1SzGm+v6zFl2qjgA4k96n7RBP0ReeFd/
ZPneo2G4PofbFY/PAa+VJAyPSgTap/xlOyR/u58PfyUlhBZ5jHboLdNFr1yjopwI0WYck/pQHP/e
xfmabxlIhInUkLkfmH1IsmOLqHm+iuKK/Q8g5JfZE/g1XMrdrihWKrQTDpz6zHmin3JbjzXCPJDh
Q+YptuwyydVDmYYZ3lJjjmv/yP0G1kzXYZ6woMb3H2fO/0MM2vKZZuPqh/7NPcDavyIulPxTUi2k
IytZOoQvGpzym1JjBWuZqGpNHK6xVOcYO+BDMcRmGC7viZ9lxM7QlP5GRXSQCcw22pmGpL2YuHK4
Fz68G1xzo+8Sk4Hl3HZIm2pwiODPm6D3XvECejCW0OpZZsiox5HKFkYcbfI162pPhF66d6sT8HR5
OBTh1D/gAUrdUmQZzlReqpPKsNJLoH4zjft/Jyq22YFK8g+bC/B6GHuK3VxQWbkRQY2PWbgaoLbB
wmANKRKWF/cpdg5NKkLhYdJLRQJAH3B3IEzrETnGfJjvVaGrcsXGK3JFt7+mhrfmNVgKQza4J6AT
+9YM4WFOC211A+OSpLD8i0szxiOLGfQi26QyRORhhOY7Ce1D2xdLsCjNIeAO3KqMP1HvkJ8TuzVM
mwqeV095CDWAHMvV5Um2hqZGJzvkR/z3JrZOPi7SPVevbG3vQaMjx4afs40Ka23D9j4BJMGx9IBe
7QoyZ300GdCc0YtGP9wCLOh4HXarjpLkZ2dUH4AG737rs9S1mti/lJHw1KOk6aSlXedBjHwSGNVo
MmiZEeLrVt2wsEMJSamMwR270Cd/PpibnAP4y5QWMKCj8CpZlIrM76l3m3IfEaGl0qO4OYXO8Djk
lj4iQlf/BjrQxZ3p3l82CUsFvqmfUWGRhMfVNOtyM1WiAbH0HO+V8gGXi/fDk5SElwuLpaREgoL7
AznuHksotFuFdd+gwgW0Cb9v7kHU52no56TCEWphhF8/Ey3dPFwSr+xDCjdBI6Daf0uRzWMNK7AH
aWg+WRjIFhuh6y2g3W2MA3mNg6wn33c/9ortGJEO8A4UdUHgsBET1fenW6EDxojJLpr4sYboVYDd
/oaCPYnUEEVS+/rXgK/oxigzksz/4tTavbWr2mptEINSrIa8+tLIkTceH/bmYXXe826dLI6dj8a9
WsAtGBHOil3O815zjE6XKpeJooSsZTfcEOQKv5Oi/YCfCVo4IGgPwbYOB5OwUpuLa79yMNr9vRXx
zTIWAneR2iJCSjtdRbVs8Wsx1TPt3Oo6DA/uADmO7QZXzUZ5Jff0BQ1++ZHJO9jKSOVak093xdvE
ekeyL8L2kHOPY+W4PTjklaxR2yX7z/AGqDzkPdVJnvMgg1e8L2aWJ/r/TdlPUI78t4g7BYivAUi9
wBGGZQrViy2DlERZoMLaZdFGu2bh+ekwngozbDZT3SiJXgE3kmOcEkf01p1lSfEEq2cblVc1bEro
moGPqqtr2FvC7ihLIDLQHDzGtI96X0q7TVDfFaHudWjDFRPZPTXM+A/YR7TMlxpiVBe4em0o3Kdm
UTyQvmucStf14Pz8xQd9QvtRL45EB33eEmWey4EUpKX02XmSQ9vhiwqD3o7p7jz/lT5yK+xyZBV6
Uq0JE2IyJ1Hgi+krDZHYICFi/1gEJ8WJjAdP221MJB/iJqLx2spIoR2tT6ZMuaG598JVnT1niqsd
tVIWRYi8q6NyfaA/NjT1DskZjSetKJavjbKkkv07Ndzrt+AKQXQgQT6atxto755ceVEdsMPbqGpR
SR6et+OnK0duzSbPxhBVUE5RMvycx698IWYlRtO5DZ8vP1tCBXILS2nCasIjyCKG7Psr/6P12dsI
t1RnlreJqB8Po4m/yWLlHTWdWkR3mvdgdwVqEBXU1DOZRAdoFixyG7x1AUrxfKAoU/PjO5iHuYhh
PC9lQBoc17m1LxbHT4kJWccU63WwDUZe1O/L+5uu/y/ZhXjN/OQlZe1UuCD1jrgaXPNt25ZPbfM6
PHiSH633BrGsDxdo8TzHwHCmQHM5mbPW68V8T/T0H9IoguAWoGkxhFJSFVCQheZY/hsWSubqZR26
SH5tarfytvzlY3gYPuW8cJu9LK6yrHtFZaQlaKETjI7nmvkzo20cnTbzwosreTeEDAnJr/G7ipeC
oiM/bQzcvLXimvTHjU+nNucjJavBOZ+qRJGh8igRgk/FTDWI/5VGdCIwkZfvrwLd02NBTDRRZX+U
XEvsvfqWa/aU4CPErPskeZJxXOA0wrt6WlHpa83Ji9n1fuGHisrlbp6i69wtnzfQyui6ng/kAe54
Zi7YbKpFNw3qaRCxqwWOGeNukAJ4fVrsvyNa6aqtDp4DN8yECoxogjv7plPMLSHt+1TgvQA7X66g
9rhbDYLcVCCWQANtyqz3wB45y/hVflcxTqhQ9zn8Bl76vfuJBGMOTiS2KGAamWejSg0JwR37FKvB
Ige9Izeu7UMdmFL7xRBrcg1aaPWKnjPqK+AsChFr45lbmD/xYxsVMTWIUQSBTpLXkfPfo+QG0i6o
FuiLfIVi6Wy54bSHMP0IdAilZroXWfDDwt9RJdRWWYtqXSdffQTCQA2KpTaVkd5KyLPqwuCEFwBx
FIo4d624K/Xml7cmzbMxPfYr8fOFOQ1hYfmEirdTOD/xfVDVXJOB/aRNe8/uZA7kY4WvL6HWyKA1
UvyC4PFslYE/o3kqEzofqFwMtn/+MwL+QlktMKxzLLKBuuQA5qhtEHEStIFGVBK+LCcnOVabwbc2
w/H+IEpdf+LEkmE+/xnFnXeOPAWNNPF9BYeaAe+Jld5/5QNba5GDDcwEyuWriODpZunoLqO/DFWz
8HVUE500uTGplUiK8t0lgv037P0dtyATX80NUu0o/IZ+o2fkXkfUAmjgAPUH402QjtXh5g7+zA5P
7E0vy/JLU/J6chMkakCSDNASPp8zYEtx8f2lPPA7mvxxoGPfWs0xEfxtINLSXiPm2TxRk0aKqPAz
E2u3wmv8bqPC82haoPFNBKA6EMMLVFGg5FJxx+nWRIt8h9qUXvI+9xkQNHgq7Yqs6AYi8OUdDlNq
YZdWxAl+sx3tsAmciWwUbIDzhZRysjk3Zi2bkOos07kwpGHIs71szgXl8EePRdE8CvynvDOBTuY7
6TXP98+8NKRJPwSAzdA/Xb4hpMb8SC6x5TVcELQ1bjwnUfcUoYYj3uQk7OXbDIg1X+OHX79aRjM3
HbXL+2Xkn6+ZcA1kQ/hwOd5csIH+A5+GInU73e05KtdS5GvCXSJdvFnnqRyIEexxwUyjbp9N3h7s
07QUO+ipaTnly7Hb2fdMzoTB5v1VuBXER+veqYyH23XHNEYBgwSk9xYR060Kl6pYCxDcaBBjaK6x
uulQKzliK7yj1OHaEd47rOcL4McsfzgDYFU29jPVwOBmbSZOMR9UdqJMtofKNjAHfz/STJWJgIDF
JB3s43lf6OHWjMSP5LkU0XTLlg9OrDpIUPT4RijFYI3JCJZJ/06rK34gd66OzzstYRv1Z9G1u5q8
nSlYPp/+NRWXxPEaRHQsh4kLgsAb53CykJQeZ8KQAgTr+TmPLAjWqXhCJl5gEcCQrgWZ0D02O67Q
g8nK0nFrgOnMwoMcUtfv82xfBQiD00D05BZHSuJ9+8J+YEwRkt1KD0R7eAqEWGFwOxwiuz4AGECh
sMUHbtF7LYqVb2nDupy2nqCUBdYEawy5LbkWnIXCTFeHGojVHT90RPTmXoKsqFKJGhW+OW8fFG//
EZP6va79r3nwYIh0Jjukdjbe06IPt+A976sfurhLpCBfCFX3ud1XPk2syv+KmRJbokx3n3mKKiaR
zjRHLCNZmRrpDjaGJrtkS0f6MapUS2212odNQPD/Y7fCiTEe4dUEhz7/0e7o2CN7NOR1Y2XiD0z6
PRTxv4ncgTI1XPozOcdIcn0vdSzVXUPGsHy/Icdeem/nxio6MZTEiS5IEETrKeosO3vaofPrqU35
4rjW08BlPM52mqtN3E2qV/VGlIDR3CbKtYG4m7/MAsx1AJp2r65mYbkMBTd5/fvrA16ElTVOieX6
5NhMI1BqqvPwyoN5Om/i/E4S5irv9bkgEUhPZCN9KjnEk6s+HcpBzQZXT9cZbTjtaeqfsZHmTTIm
AiWNeKeqVu1jUrrk3lHvDa8coewiHxug7Jg1U1BYA4/gocvuB7JZByiIU9N4DEETcUXCn4fyYv9u
ivo+2E2cHEvF20naeVslved8vKTv0+ozj72xSrdSAcSwkXVRAmIfnmHtRBeNtjUwH+qTD1ffcWC3
/uQACjXGhdO28pDjteCpfcei6MKfwphvJ5SFXvpyDOIyo5TugtF/YnR9WcqEGLixYl6oYDIFv+qY
SzyKc2f4ku5CT1VClCjmNkwq8DNwyvmhcARKzV3CrJ5OR9gKnoua++ZiynHXOHB2MrhxbS1m/fde
1HHY7UfC1qu7btTreZVw5ALYJKi/GhP/I3s5wMWsxlIJBOgUaEh8NBYAKumVCzQIM8eATlhnfxpS
P70gv6DfowuK/fBw1RQTRFuJNKTGM/5lhOHGgR1wLdr5xeSWNsdObSPjdvd2ED+EUvY7QusmFbF6
EDhYO23HOTuqTXmRNAklJrlhinwcxqSds6OPZTgnXHMnv1b57+1cZol0Md1HyFzxpV6ZWxhA1mOq
lcNIt3BNbv72HQk9C8zvD56nFPvieJMihxkww0f+cLD2PvyCAFXjimof5faUb7dscdct8qDia8t2
P+pLPo/brBrn5nevKn3nA+RHrgzvdeWvaKC/M7IAGIhrAmxXcNLn/PaAy/RvKgs/6jVwprwsiR/7
0v1cD68i5YYb0MiFoqPDMXQEAl5jKAV5HtuVx7b4aZBKYlC/wdGXCXMcJngZFz2fx1eWPJfLJ+un
Fhv0mvWskYOLQj/59rUPtruHPlojiuEJp23BCcTfpn9a1S3eAjrSHcfwsauOVAmDYDvtUIrXgdA4
Rjr4+wRm9UQlzGBproo3OpGmYLKfPlRr11KLJt7n++FwhZShEmZfnNKsN74pzHubFQCjoqFYEMfW
m1IqCpUIoBS3Dt2c7i11rxJefv3OGHVEdDv9u8Fx/qPUPNpQHTMFgOXDqu9RMyGicKLFwzR3FeAj
QppQgJ4jXzC7uYYzj6eDKVDsjGylBuXEZ+1xj4M32Z8nhMjFIgGzkR/4gEJLk+8eJ0h2RiAqxod+
LolI3moRQbRavkdrf8d10mb/SXh0GZg4luWzU92y4cdHzMGGkMZvT6zi1EUZQb5ewZmCKSKay1S0
e3ySKkTMqHxxROow4g5Xw9PB18ns0c6UeNPdASEgus9H7hBspgRMEx1XL/ejVxRBTd3WSX+54i61
ZTQ3m/eutaHydHqjG0Zysa33ktFyugRncPfWwItvrwbhQl4LXxURoaQwEBso3n3770/a/cXm1EF4
X6KE034AK6twhCNcYjl9zQpXPfEuu0lwUD0yFEFKcHbrij0hK1ZRmoTfnHsU9fhGoJuHU9R/ij6m
4HlKTlDHW3BZc2tyQMPCrdu/I5RRj6YhRG2h4OmTFo3jjlk6ZIHYM808z53Jx26pTKAE0EnlA12j
jSNbV5XZ/W5NV+1Cjlec+tWp04pmXuNzxtDzgcCsMZNR1brzXtliueSoWU+t57t3nBxs2c4WoFnp
BUSaDDcf0oAnhKIcn6t9QKGIAZI0F5RiXU+n/abcprHETJ+wHrnBC9DqOiHLfC7mgStnOpesy9kV
OWGRRnVBqPwtkby0eOlzkDDoAsiEkoFD3VqAiXmvE7IZBpFUgbqKWjtB2OWXmDQ6GOwhUDvmbMH0
KSNASFZJ4Rou76eC7be+gIAPeLbMI2efznT8b2P8gaYGoMFGtmGAQm2XAYxPKjHOFn25xQMhkk04
DdKct7Dpys/xi4tVIQXFWilpNHqmk/YlS2CzO0aKE2lwY9fq6vemJTDafkYGDl/Gv4EhawRWQzl1
eo/0h8M3tbeY8LlA+AdW1pZSyFEB6G7/tuvaw2zAUpWFLaBk6CJxzKx0n9zC/rMaTDZm9xTz7FPn
r8DETF5sYzTpVxE6390Hvd6MKx6gsj5opxx/SckspRtbTHinXs8OuusVXwVJ94ApFA9kAlMiqMDm
90xkvGJNHUsbSjvwIl2c9U4RnP8AKIhho6ayqnawW5+IiNFPLI2dz9GUvqmr9zK93T19L1DT+EmS
z5M5wfrJAAxXu/1Cg6ZWckZtV8UyAXbKfgdrUtouZGkIYC8SD040XEbZdkAhPlWYTB4YinZuxQX+
hIjJAVNUevl0oni7DbZ3Oh452Et3BH48RK9PrIiA6X2TO192h3a/RtqMnwWyfWWLNEZf835ZbvA1
Cl+03m9cZ3jTyWQtrQlwcgze6CxnYO5H/CpZdKFS684RdWiIOKf/+eE/JSrnKXY5je3nnBCsN9/V
9SRyDX/mLaTI9i83pOyRB73bH89yD7cuKDFtohyFYI2CNQjcAQI4Nm0fBhGXRDSB88kowV//0r9j
3TBFZpiCrncJyn7OL9Lf4M45DCBfziZCZq3ts8HbIqc8TDEM5II+F8cILLkOabdR64b1O2quw2nz
PjA2iJsA8OAVCVan+u/+5ZWsE4t7wclCwd99whW219VftxqHiZ5xRalCId3l8WRK2JRVxZbWUdPv
JNidXQaZFTDoOPhRwZcWfIAAMqe/Nq+01/ljtQe/hL+QLGpFyoKpp9jYVFr8FT4A9u1euMg3Fkuh
FaaCBGpQd2t6Q06cC8rf3fcxzZVyxk3d5BBPwg7ffcuaFS8KZFIftWg1LRwGNaQHOVb2TWEUWAox
9/YNtf9W6pLdeomPKdsPo9+1e/IwDMnN232BRBCfvRcg4G6jNjUuwL9TY2WhEIIIeCMmuhfFAdsN
6PmpIyziCSJB5TYek7W4Z+RdLowqmYA0QwbmWlNEIyIWlgQX0YWJF9Ve4q1B+iLM3fTG+VNq2347
RAkH8itBzTyN/N8ikDHc7LG460R2SZVnv6cw5MYCTQltW1WsLBykidzrt+hd1qNQ0voPPECTtIeL
mAmsUKWtszdTJ1ZIvWMYn2IavlEop2Ig4uNIM6y5WD6mCbw5xgjD3GlEm1RjK4q2tXICnfihjBV/
QXirVf4P9ausFoEkLD9uec5NzlBkIYE7ZrUO4NqMnVUxhvFAmABzXX1h2g/naLc8PXYAEq1enRa9
Ap7FDe/QxEe4CKcG1NsUTvIoxBbz4L3Y3iee72abhYRh5rUC34iuL0R/wmz7zxtcacVmu5YWmAw1
NNWt8yuibk9EyPDBvwYOJSE7oOKUBVyDqZG6gc/Mw36A/g5eoE0P+MwjHEguXy7GnpmBjj6SVJYI
vchSMQqUKms2CZAgDflaKjIlP7WVjS/RJjm8lR8WkhZcHCWkWynD2xdLHIPwm0lVIMUO/7xPwFde
IETg77uWvzjk3UqVnpqVUjdsegYjEl46greMD9fsc2hNgjhHID6XXGIlBcczrlnZosodwlEwgWfb
n5ImnDcxXj1vXe+vs1g6u3UGGRgSmqpafgFtOmzJBKacmg++3YyOPml1G2EGhEMFMfyJRSDvfAtR
H/8IfVetVWUu+gsLKOSFq/SVm4ehK2e4XBVYJ8FrWVEpzAkqBSXAy8LgWfzICoKGs03e/1j5AxGb
y+BMNmdRlc843XxjL74i/cvqVL4cNXzt+LXP59PvS3iEy4zssUw0qvSA6lCljXwASnxqA1lC/2/W
2TCG4P9gF/HGmI2PHLystO6Mm6yz2gpwIQ/7+6qKcT3GsaFqyFwKzfNY5aKTg50qHTksKT1ArJpz
7duhZLXawcB8hRQmoArEODiXFqfWwk/R1Ef/9N/vmR6SCkeTlAIVG6SC8j1NT3YIYywfnY9KHyKU
0QDi0962pSweiWgWq3hh5QyYHGQQNx7Ty3Vkkkzv7G6Lkx6LA2/kQom+JOobxGCANumIl2Zfr2sY
HbZX96RuvewSn76qmtt9Vy09bFrd4N/6C188Prv4uBKQT7e4xI3WrYz4R84T+Ox8ESb6xykRcEm5
ZeSRlAucP+kVzdcbOzFDx5HXY60BvEa27nRQXVKJBf2Glelcj9zucnygPGnv2FA8PV4vaYvkbK/V
oEnPrJ5+TkWeDw/+f0dLCPxpOABbe81Xp3B4BAfbtaZ/T3kgCcZYy5sZBap/E8En7Gm4igwMcWHe
dKaGPuPcf5/D1i6geby8AjmQtONryHSMuDtxl3xwL7Sw01iHpNmYT9ZVtSE2OXndQ2/SZkYQUX0Y
cOGUMbiSoYZempLaaUrWut18T3X5gikAhrhZj1kPkwo/0aimk/dE8SYdQYjEue7bs4l6UdbnWWul
bVHrPyeMOjx2JDuIz+9wKcHlm2HoTF64/tLyJW1BNJh9p/H7c+1POxg2pdrTFagJ4I2LxEVfmOmd
IkRUSONWXr4IuTkN1AbvLZJ+dsu6s7eFC8f8P0BAtookbCD6NW4Ltl5x/sFso/CjFBH9FYgqOi3O
ig/OkX4uJbwYRW3/7we05wR7rKO1NK2j9UHaalAh7y6WZ8hgsM2Le/FBvacr44rfDpfsASoEulgl
ZpvbA14Yg8lmkGHF7nkZN1bQAhg4GlZ+BQSzGT2YhMdKCH1QllQrMw5YnRZl0wAdH0fIbbU5rURY
+T9P6SJzfWwMjFrvHrCOs6xSKf/gTwuhKpMhDApC2pn/ZB8AJwWoT3687qzpMpNEg1Q6rE7SI72B
x83AsDoY6vhRLyvofoTIcpbUXZsQoFdWvoFhxCY3rkNHRBuYN8D/grmra18eqcz+JHhkDslfvkjz
yZrptV7101UlnhEcXDlef0aXVm31zKIv4QDZBkxJHX5VJMi/Uaqv7cBbHhd3/NG6Cs988qDTFuQU
x08Iyrvr+FbC+Bjd6T7skKxSIye0gk7Me+UiTOxRGbX9uH9/lQCAaUQhSMAN5AuBHdgI2IrdXC9l
3FNlUhtiby3sVXkmHDzDnrzT7GaYb1LDMAfvmUaYwzNSs0iru+gNLwJzSk+AYRzSDA99wGzpXt6m
L63gLW+rqPagNabzlVhMFMWetUM8IBmBEZ1x/bdugTD7pKLZO+LtL9v1cV0Ar80PEFTKeIRHPbtA
ZfpXBpGc01zpWcbouZRqa8uYcbyLuJLQ8hOPAmG1DG1Zpiqaf7NT6RnDBZ9it4bQc6g/pwbxy2XF
3EN/0igdEkTqY0B2gGi0LCzkMHh9pGpB3kjq/Lm6wLC93/ldzGiyFsFzb85SF+9bUblySBvvEe9S
PEySKgr4W5d+CcVuHpdGKRVU+DOTOny4ZA2LLr4sgMlEE9VGsFmOnjL8EStbbcM6Oo41NUIobMiK
faCfSj9auZv/k57P9nypqE0sxbXkUP/43z1AcTYLd3t8mPG2lAxYvHC/uEJhyi2vyLH9CryjYk53
QGStiRH4NQKZVzke4R6A2fLANjdT4sZroK7pT1PtQOYfpnLXr/E/0kko7IXztgdshFjOwCNOb/6d
nGG/VbJ9q/UPVkINLeTP8HOcaHV5hBX84kIlvW0MgFKKDUFvO/GL+pSVaNW04+VyK5Ec/n6OSiPc
EcFovX1HNn1EiFseb3Q+Y9RlZ1xxzTQFdLiEmwMeouDlG1NVJKNZOXpf/Oml8P0tz3KWUoum12ci
Lm4UVVHeoj+2KIJ/MFh8k+NZay3cRw39/S52JXIgSlWFmEYdjM0zbpEkkvHyeEzdimWlNmaV7Idh
X+2yWmA4FzelZWTwm/nz5toCwTsVAgc49e1MuTEXYqZLAf8q1iXI9IeRsFxza7ApPQa+sgVDT8P/
B96nfRaC1r9LrfYHjCPQNvOMufPDsHEL2igXoBt5TA1NfcZBgpXCPuIR8H3fpft90s7QBt2t+5ZQ
2cayYNRktdw79W7jssiremeFHz7Ufpw+TIbNvwfndoi6KMNzoZQ1Ji3BvbQm1rftSrXl7GqYtnL9
wQSp77RQ8oAoXG5PTzNEPNOV0FMPBqNNigXkwuECtIhlOsYuG0MkvK/lCjXrcfnF+MwjiorOIxxY
PHtUDk+xIay++fyrHfsdK/54nKDaoXcvkGJkOx31ZndtvBWQFVKlnntjegDfgTaNK9uxvAR5I0Av
9FyPyHTa82KsHtquapPgrVKWBHqveQj/yWA5J4+8snSFZK5uxvlDwA78NWupsqOw4Z/kr4RKHRqO
gpmk6kTARoGPwuKgVONUr1U61FmdJsR4dNcWyGGkSQX7SqKHGFPzStHzJYwqpAWl36hMTAy/XAwa
jWKM1ubc8e4gBuSOk8PKQXDc6Mc2yy2ys0ksj42H4P2QHDyZe/OUnhQKCSFZaPbOTGDNEWjHlFzT
plRmKl6ZVmqwC6AezFJFFukjp0LXy/DS6hGk1C6hZUXm1pJPn972UwA9w2Cc6lyAU6P6+R+D03LD
HTJT7cufRgcES9ePvqpBvchrEXqq3NlEh1lyO6j5d1Yf2gv4F+HY3f3ZyzjChTmZ0uK/2LobpVM8
tOwq5NtFUcZk97jRo70rZUxeAcMz2RYBS2pt37XAjnLex/k5wQUP+2soOZ6QPvmLmXtwWIGEaov8
pfXgZnS752gn2dpzPN1uFFILHFlxjnPDWAS87ah2yEu3brfMG/2v8OYT0kx5GECgHpjrsqXu6bzp
kW+OPyr8ugBy74/FQpyJj13gZSyG2sNp7QbNHG1SI/ILgZjpYJ561qTWz/NTMVyW4h5xxycDx/uh
g6qVR2GlQW+bDrFZ79DMlbv95bpNvBvTFBcW3p9RXK6gx0yAVm6dvNvaPtA/Y1wuyQBqj4teh9Rs
gqmbNCli/yFcm6oFxJS9DNmPKn89vgAcDLDpfmoQLM1FUfUhqRTuQtINr7IcMVSNnf/RZFG9g7wq
EB5eKOU/ZxL8+A3yYM99R7+2OuJ3edqw//XmqUODn4aayZDiWKjRVH65bgVLUuJSZWVRDDrYRlhD
kRNxEajZxFZ8nvdGwohlgZCNjHQW6O3s3CYLk8WvXDX3fGKRDDFOXSa3QV+Ww6Ub7flK5TS23UFk
/FYpZvZHCy08Y3t78PxRz6mDpwpcnj2qGYD3nUL4NqnfFYF3Q+3OFJ1R9X2tBTMUOqXoCqF04lnE
qTBQbQGuIVphY718hh3yH/8tn4mzbcO3mi5x7380y6leT9AZq+zjrqUsoc6ze3UX9xdptp1F5xT3
UgO+slziYEJax9Opn6ttapLaafkkGXHhT9h0/JfPbySEWJQZO/gWINTGGzgzVNWZbQdfJtFjUEbz
gaza6i/y+HCVOqSyHMyY2lSQF7Bol/irEKTsSkA30+dvcyWpm3o2xqvNvLX79SlC8csqpEMpGGoj
seEuIUDSsUYexfh4FTeJELESuUXCMLC4lUkjL0zCnWh9z2cLdeuEryEHJx9I+f3JQb8VPN5wiPEb
5vWnbFXB9Bb51W6V5DbgF15rU+wzoX/Wrv7YQ+UMTId262wevUKoOspBxR8A5llvDt82PK64ox6H
11mlc3ptd4mwJAEbkCkAV2rDhGkec/1gdD6wdEgBtUkBYPuHCVtPuVwgYL+3dHITlzg42NG4Xio0
+ZYLzZGysWqr0N6lUpvyttBCu6jhdlI9wcoTH9QZ9gOXXT+eRnx5EqCnASt7DwrXadLKA0QAg+yL
X4Ec7J64o6PqyvjgT7OCa1GdTRTBnINw05kI8u0gj6v4pvw0AGy390ObrA8A+UNV6Ck5nf4HJpZf
yyaqcfnPYo9cUpIhnu0u3H6C1ahfpVWcL1W9GyRWnGplTTFmcmakIpDeKt6fx6GpGbeiAJ839JAe
T358Zs3NNvP0GcvfxSqoKJBsQ78n9Rre3xFcbmiqUetaO2Bxs3gu6zzI1TTqJzn2+o6g6qekoooR
uYTEqam+WGHjozMMGJ2/G3X6GcedSqRocXRtWq9/P0thJwnqXGn2c9mpcMtEqzWJCyiNZR13Hw9o
5alXqD21D1lZePwUDqEJmbO0upSqBnsIGGL9RvkQ2tJ9QY9Cqbi2/aOUXBEhm8SSFcNj16tdOcL+
djzoYyMQbeiXAmcPoWg0LQLyRFA7B2suGoXYK0SXgWSyXIYmhi0aOIv153h4PnBs9Yor1V6y5XKi
g7WFumLhCBis658LgRlZhIiKbWzZFyYVMV9tfZ/h6+dRsDd9vfsqgLeE4AV7YFKPf3WkWc1TZL+M
kov9/ffxwtohGcMEzrYLzFDHgPKKsmUKFAGNktD3q9MbaMw5UuffVfEz1AJEQVeYHKmkwcIkuk6G
0640qr2YEP0PZBk3jCbCwooo9eHFuI6+SbdGIkNU5OkykOnRfXK4/5+bjBPfsmdyZTUykHFBLhne
WCPRYQT3PRQibOxrY54JhQuqHoEOUrVpe3vCuhz0O02u7AW/+Zf/q5TpR2xPG7RwWGcaa4xzWHjY
Dm6ye0gIRYw4mbTuhhq4HNCediQ/7CYtrMIjjRioSvjUO0JPfXwUP0e52830eeQYptoVVKyXn8GX
0pxfxt6BlVIaPNw2L08icbO6AWX9E2IKBDE8lkkt+rDhLxa6T3ZXa8xT+LKjaroCH9pR94ceeN4L
2le7jwL/K8TMrSsFHLd2ap6YGqccK5x4F6CLHq3EP7Oh2F/9aWYrIK8YnsFosXaspgelHxqZpbzc
LNL0Bp2WjhsSI6ozFAB/XvtOeZM7YpWmh/dDXAfnfk6tXNNYNPHm6e3Y/AnuSYTMQL+hOkU4k1nS
Qr9j61mWQFftnMd/+puo0JUL6LMjJ5RW9HOk54ItM4RJMKhYYvxgptHaHuqgvM0UqdxwiXwPfrpF
dNopQyBdkbFn2rvqWi4ZVtXzJ/smB99McON5kwbCztKwPZKK7goqmPLOE9TbFW5NQ8+lrNNHxNbb
/NXYwid9A7fEmNOEMMg3qHu+Qz1HrAx5l9XrR8bDRd66SlJ9Ha2uHqrsq1AQM+MJTCoNxP0SoH3o
a47/okEejKlEgqmUHM9jHMOSV02XbkfVPublozYEi2HkkTm3LJ9zDNYCYDQovG6Myrp0bydo6jUR
lwT75okK6QO1M0920ItINvCcZ+4/4oqtOCYOKnGbEHcKzZBKraNOH4XyFhW+hWo9+quESddY6USp
Lsl8heoF4k9VPCd/pjuE5b3arj88yFT29Nq//Jlp8TXhhTu1rzttqWudSegY8vpbXRWM80Dtm3J3
uKtRq+Xc08Tm33JLBibARqzhc0hlkVrLoIzL4JcyA+S/1cFmEpw6s6KZEckKXGO/0vumYEmER/62
3zBDB5D+2lwdNHt97Kg9ulYpi7QhXSX01ExhgwC5Clrh5gd1APcTqxp3y84XzLyEKymLdyyRR3FI
t9MDpDW+HlurxMbPqt0Bjt2rdBb+uXD+4y6VflHcxlvMMl2cAGHu730Xo9P3BLN/a+OVpr1C4Aoi
YBtZOSjYyKqOCe6uNa6vUiw8d9jmNs8Ab2KSA11kqNc5GGCGWMYwO0oqZyoL9gvq7aBHG/PdvbHc
5CJd6XzNebdLM/dkZtm/UAQRETyMC6gtXjtxLlpRJsCP1y79h+VTzGuNIGJ3exwYnnoui2rHnS7M
T9LPL79TSMM9v9KSKxTruDQvw0E8nivJQ81F6d9vd83OlaAeSa2iZ8Do6Cr1yYIzMLK/5vwDBeuA
zR4lfgbOZdFH1LPPFDxWkRW9f7M9OHG695JDYlixYVpfuNgx8aS/18bUWCgZMIVR/WZK5G6JfU9E
0pA9ycql2ff7hf7l+vjVTF2i40YGmz69fZAzsduPRp8+SGP9cCK8vCzwiTF/SfC2AzBjsiTWxYOP
KqTfCFXi0KDQACB+VtyOour2DwAP6lDCyKPzNWFZz4FDY0F0VkYC1SRP2u2NRk9E1KTiogII/bo3
pze3iCPg4El6psNn+G0gT26uou2Wvhqb4jmyOQANdaYvkSqbXEKsDNnBuaDWUy/fN+YbUW/IOZFZ
HenCz9lYk9AI4YMLe+oldyF0rz4y9sl3XBxecFEMTQHMoLYo506maCIOvfomDS5RvFJEnM/+tzRr
Ik3OhR9OSlk9Enj13j/C1yq8PhInDCWEao9nP2VUFA4NVWuy2BThcclBOl8/pscEnXSZ41ls5yNe
F8g4FrP484ztpWLeRx0enrs1SHtpirIyoBP9OZCqvEz+QnuVzQUIAgyWh7p/P7a1+Xgy9ANLgUHZ
MclZu9sEQD/GK5BFItwuRjbGKwn9l4VCMXgLLn6rbYxsby5THjpQsvavslRCZQJn7CkFDX8neRif
cKyAvE8QgM0W6CutTeh6I4XKsUxw1J7E2jfXTvWkwDGHACJKN8/Iva0Bt4qECwKE+++tm7liLPXt
5nWvfcZW1of22diSPG6H0QwaC55RvLupXUMVIAtrDpVbyeYstH3iDlrLNfdy+dR94Y8wNPphHaQu
nBIPTZhBjOLvkuHyBuejdDHRqmKUtIr3KaZha+Sk5jVwEZlpp10f2HtqYBABf+HazoCVRTxJ18Dv
EgEe29gDx1IRj8loa/MRgqMvZglvuMj8lrmjIqT6H5hMuVmEVq+FY0DzcgS4pGCfuxiOczXJ7luT
shIOGNjrHMbVpqCp9RaXpfKtUyuh6K6sMWaz7Pw7RbNwp8lFVvChGSVtNdoI9FzTtSbrTbbsLw9r
z0LMTfvjfxeisBHZMqnV9DBV+0BANn3fURgLg/qEJocnTPzWN1fXlZF2L6KdhzM0tw7ZgxPr/6OC
yx7BsEXbFNK8noiLezaXWAfAiZwoI/zQnHea2B71ULzlemVx8ilzvUC8JCF3oyT8dfpBLk3k9pk8
inTKxVgr/4sNhoMKtzZgs/6gkz4ZYs5GU/Aza4Hd/ayGtNEconuTGHIrD2IRhg6wySRI7YiNFWLt
vRUyrg6dIZrI799WQxnqKrmCOwFbKeRRqbt7053WzGQjPYNCcZ9VY8JXzpn4hgb8xPxdqV9eAyY9
HWx8Rki6AXIW4lQhnBJqNlLnX9vok15WBHrDg4F0DPm5FwhAwLLI1YFiuLTRJUcasBFY1YBzoovv
hl2pLyH3uhHnsj6qn7jVc5Pu3QjREp5/wCcSuAXOdoyigPBuuzcYeoxY/i18yVEKuM1sRQUqFsWv
TqrIa3s1rQiKvjKV5HTh9K8D1yhwa6Q/L0Bmi6EI+tZuaT3Wiely0RTE5B3jfWZann5OqKRZps+q
g9CtJnD+ucascdEJuS0V65534ZLX4SyB3TZ9ovFu6JedvEolwF8zAdxv7R3I/nhHoMeHJTMYuClq
0A7SxH9Vmx6xDwGXOn8GLe9Ib0DrrpTUteKrtMiyuejXCnE5l6Ne8J1goWVQxN3hLdnaeGNtDxJS
WaG0pXW703orzRry/tAqFpB1ztfVrn3O0Bh/BHrAlOiIQ+rMjjH2kZ32F7cRdaQ5vaLbiZII42lr
jXN8z+cfXAtrrGplTONjD363YCyiMjEO8hKG6tkcpUrdYw+r1gzP8e2SeUmUF8h0IgxPAmqqcSvX
+qie5/sZhxxuOXainBlg7FT6qNAIr7OuFQiQekxbtlMji8Swnfs0ffbgWwcsaR+d5vtzdMzFSoJV
xnc20GP/1N4wwqp3qM+aYYbWjAuM0R9nPTtvk6Pw4qL9STP8TsoqLpwYlwDbncH3iZ1gA0kU5IDH
EWDad5vjwNkudpmhMINjvO1FG1dAjXGpxPBSmeb6C88Z97H2lycEEFw7CKK1xjWCvctzEjQ1dZLA
gj5yzYGvKX/OAw56AMbe4QsklbF0TusrfuIaztx56GLIG7DSebw5uKGwr2rs3q8kD+yZ5XeCuWhC
3HwRi9mG0Xj+p8NGRN+u1kzqqM3t2IHBOdFSFQsprE7QZszFUyXHUSibfk+ARUwrL62kRSy5+JKu
aWkwJp9SwMRsJosvIa0id/gR0YAfmckk1SAn2jC9fjhuaejhaXEITM0dxsX7zL2sHG2NfX8NTDLc
oBx3oZqM6BNK0WHi9Ltw7lzqYxv9SBJ6ie8LUvQm9s+fhyiHouwLYJAXgthrAcQaIR5tBsp5Nd1X
uUjSXuAbWsCHt+Y3TeyPg2yD50NfDaeS1u1Q/ke5Xof3lqX73laB/omzcNQOwuhU6cVy7fRDr6hd
WlbOLDyigtUavUDpxVHwRV0r4CMZMxrWVXG+vVIxMI6n4V11yyu5/c1Gr1+NFoFuaFlyCwOn7g68
IkNmxyg7aHfEskLdhnA+L5W6wCiSl6fV8y1IW0xLY916VTts0fBZzuCuor6TpJbhCU3s9X8+NBXd
5pB5UxQ5v8uZvd76k3tnKEu6hANu68GKU1S64UZ1dukO1vty1+Uc0o7W4bwRw25HTjSZ/w6FaSwF
Ng1cahn1ex0zgtCshZfjwui4jitEcBPMoZ7KZqFXgaoMO72O1+mvTUb59Ok44NWffUTFu61KjvJQ
2ERlMQYLV6n0v4M5YawckznUx223zQCmlMaKgD/qjz/MOoV/yoZHmheurPv+I5zupwCL8om4+jHB
OnMhe38NQw29cyI9yi/4Y4oM5cPzjGzH5w76T1wByOqLVfX52rCEXItEhTykLD8LLlZbj74oEPIW
/k/Q64RSyPCaWI/P1pmfUBCOJAT55baNlqI2R/YEHln/3cPXhuRn37gY0WBRcyLdrGhSTt4sgN4H
1ulSpjha9AA6LmF+sLvnAK75ZmOQPv/PbDx2fPo4X90Ge5XnY9iue02Kf1lT69IbL275/vW62KLQ
YAv2StlP3AHv+BIiTfbNVS/5RGAVa2g3rgTJ+BvJLVuvHn9EYsU8+rGm8VBAYDjBNS0lNaAzC1oi
H6h09NmtviLAeN5Qrioz/nIvUwVSm0fjwHopsWsFIprWF0K7Oho0/tqWenr+jKzxy291vn0PQbd/
qcqGRbVv2PijWNv6ij46VF0wOl272RRvgzHM0dm+scQIpcQ/9yd1/mtknm/tOitI6rFmgnQr3wYH
U/kKe4z+TvxJurdbOyVdV1ArioFp3sB8hLAbim8g50oiLDw4P9Kkgfzp2g1pGpU3opDmPQ41E/x5
de9oqhu0AvCvm85MvyQ893vSP5TCUUeZTXT8XV77MgS+pYFNkeFx/yVtx8zDZ5yuFwCzLk8Ow5LJ
25glyVrfoIet/TYhdls+GTHHgkCqUjyJXfkKRHKOJpTjm3Sk7jbuoUdKhadMuScoTIj+qZhOa2zh
+N2fC/ZNh3luFm9ZMkkGyuQmbJg2jdfgqqiDLVhbictmAWJz5K1g6QqakSzhwwMlKE4J6vA+Map8
Vf9qI56PTH+0ACP267KKwZ4Q5fHKTNbem3MgEDEfQOGP2ogjS7yuuxHL7l/Hos0F3Z2E+5n5oS3B
0/gW5nmi/q9sWiXs5/g+Qi6AMl9NNMrxNkJEK6WLZU5MffIkSuzjPc0lPZNUvMa+fHjthjQG1kkv
m5ujauBvBUf/3tioTcOkvvQhABMXTOfQ3o3GNphqlhwo+NKFUf4q+z7YtkDrrJie1dpEi7547rBf
X6dBRiU86R7e+yedNg0ZtD8liN5HgBYwVpNGIleT/DiD/OOShLLmOCHdkOVuE1/HeuQYs4F7jQMZ
XZiUpH3DWSUVDwh1lb2jP7x36XEKuFm+2kPD3BxPPoIAarQilSoydaxRZYcirKvjH9uC+B+2rslp
dZM+0L6k45CpZy6wxw2vplNCN8Ur1U3V5UrfI6r7LaJ2+D4V4vm54lDqDBhnsEV5G1TanQ8YggJh
x/USIfnCQWBztw4EvdQ7ZME2rNfyUZIvxYcyMEVpDIVXS+KW3LjUvMhHXwFAD1RCXqGP8y5vo2RV
k5PF3kf7FGxOf23GxnftDFlCBKdW/m7+SP+2dnx+qFUruG5loPT4ibdoyzwTIhkTmdOSU7VrDiLB
ypUxzpjr8QjBInKCn4RmExDSZ8WLNJ0lbo/hWcHEQwRGJRAsMWtJ3uRq5HjvG5cLgCYrlzvm5039
OzPEncTD8cRk8E1chJ6HSm7b+yEu3u2iVlXBe9MGkfBRxHlhum+YBfnICVU5PgTBgpG7schpsZhC
zWX750xRcc/+FUSlx7KCuAFyM3fvlkX6Gqa2WS+D5dZ/eTvkytJhIdtbLIu0SSLqO8GcH1HirIjQ
RXGO7Gcr9vyM2G0MDDQaJN8splyfV4tKI5PnSOEBu8CpokA2WMtHBSq0hGiluMno6EcjGbDDEg6d
IGP6YKAVdHHv0Xe/pJ5TaR+r9HgVQ0HbesnG9oJYpKSDIUgPQpAcLA7pf5NLyvPnMp/MQr86Z2xU
EL/YBLCdwR1mOxapp9384GxBe8C7C4rkJ9XPWc6IeUkQUxzinTPrB9zRs0VH1+LHmzAVXbLQNDYx
yPh2YIB1RnZyH78fjJzm1HGLPPGzybkcGuzF4OZBzjfMJzTQI30SQCku7UrTHaygT+v4o8Nlcicg
bCiUkNNFly2PGGGE2y8Fw/LW5sl94ZxJYeCAG7g0ZF4cN6pV6qB/QXJE0RlrQAbx1bLxrs9goPjM
ciKYA7BGEd06gvL3jczp9jcoCoIg5ehAejiB4tdIrWKa/5H3yVrLMTaUztWgA+R9SvduoEdVT4bO
GArUiS9GQuB6gbbNUsuO6w+vlLHBVS7Kn78jwSdI1Nxkfayu7S0hvIrk2OAaTFc133AMUyg3Cjen
3oUbHfbopoXyHiKbYPnbsjH5ijKkKDTV2AP1BxKjJ9aO6hLhMJRiMN8J4CILiYIFxDMZy7NZRQjZ
W+rUo8PeWjpU7meFIwxobdCFqaxMMglXdLUgttBkGbfqZLSyPXTxOizHbWWD+AEm1DRskux8zbaL
tOtO7VEZU44b6IWwDF8jXAlbxXrAU2jPRmZqG/xATICwIvdyTGH9Sc0f9dWPBX4I9ISSEjbD3luY
CysEgh4npHtF/q901cC51voFJUhl53bRou1sh+kSnC3ZRNdovryaWKRXrQusvLlBu5od3/iglAE2
ZFjlVX0NDiDahrp2ycjKNQfNn5PcPC0NUMVpZLBX9ahX7Jky9KHxUvwv/EV6SxUaAIrsFtvCAmUv
EtH7soi9WxJPqh3TEL56WYK0U18U6yCnHcpyXeUgaGBc1Z0pygQvajMb2wsN9sGaED79buAQ85fr
hzf1r93u5cCl57RfvHVaDZN3lQ3eL3pQ15AKKWNMjz+l0wMhW07zjOPTi9kxTbAqC1/bTbyU27e6
5qVh75gMivbe+lKDBTxP8ec5AMKmq1gvYOuOyNWkiVzhw6F508oQrL5msZmilF0w2TGiD0FODTI/
c8mcW9pZjSrSYy+hqZ6X+gdIKoIDeukObPjJIFbG6zplzAQ5H7QmA/vKGHFQGm0RYeDmeHuBsiEp
R+gGgQkr6WNd8w2wOVY7+DIFCCf34OkskpPja2aPc6hZpOe/lLp1Ey/tNvRQShM71bcFgrhAfYrV
hBOLdxtniG0QNwWBjvuoiROlrcdIAIjv7/fhCjWK0HX5xy9d6HULfxt/bKeTesTVcU8uo58jCi+r
yIPW/VXmkrhNMmTA/cjTMUHRWB0ml4WK8VnUw3zmB2NVQF5mrMMdM01BB5H3ruQiQAqyRyEuBs5m
NjQLk1zDKoGHuw16OW6xCtE/gZuOOQCSCHyCprGtqh8RsPKRdY0qd/Cj8RGA4vo47K0rfjmj5mM/
5dn8FmduSOYraakRHYlbzWLZV6bgNgsMZoIuQffKwPKtgGUSB9GoYhyEtQZymFUINY+QSSc11DSv
/uT6pbImyTMtaIHHnj5FPH/BTRjkxzEK1PjRqqCoMe2vQu9FgRjgowENdG9DH42cg7GT3wC611XD
het8WuI1hMHvoNBOXKHyCjukm4swomq61W2E3g900MO49AAGg6coXp4hQfEaOVrKwQGjlmXoJvyB
MSCOwFEzslF0+oOw1kryN7SkQduA0q5ouY4BXtAJtShsNEyXnKLxvcHRqUHxh1uFSHVbWZ/6rkx5
XLi2BiO6zozevEsvdmB0wjUUi/KW8zFVsXSNXRl+tKQveagTEuBpeA7MZ6/wjfW5I6s/YKZ1B7mh
UHSAJ1fvGvcY2RjnP/yQXgMgn9NlaorCSTmn+soiAefKWIirZj/Yk8uflZeMKJH5E41uAyGST8M9
ZlTWxjkAhFpkCbIZ4jXaxyjwaQVrzdFLv98cgc+4jNgZQHArGh1+ySB9VkNswJ2lMtZV+Yjtujjy
hkbM0nbPGuv3dSG9n2emmSEtza38voguRWxOOcJVmWAeLghdaKPGEYeGbdql6UFVQizrqlR04Z7o
xsKwA6RrpkelKymEI8emH4zgKEolgksDbWkpHBecvoBi0mi7qhTpRVbcylaYQyqx2A3xU7wBCyzY
arxFr+sorOfw79zr4ZCLZ6YZkDckV3I0ORubyrL0NLJ0m262tA6M5Z9gJAURuTeNasceVBXah8VG
2hEKyiaHG+ALVZWIEalGTgLgjPoeXRulYFlyhDzCev2IbDg4SrrDwLk5QhXQTBS/CtSzdxRNIGD0
oC+xlEa5JV88F/8/JbfKXTJDvPysogOrlEN17yR5ThI7uMMwvpX9Ay64FSHKXaUSS513XWpga75F
yG+s1vejS//o//7bhqdwAgWU7g8/cWM8TG3i/AL4iWi3hAeapQZ5U/O5L0AMtISi6gmfgYn1vDTd
7C0hWDI9cy1TcUbitBWZ30TM52RvjBsLxPvA1WIE1bAjF9gZlubJZPsa1q/W5ReCjgYDze8x09oS
VQ5YpAkw6WFdyWDtrLdm6sNyjtnzvT8C/W7L3RtGHRgimNEfAz675e/nt2epIHA4XYw93jLjx6xe
RR18wgiyx0gm0KkcSs6i8e/iV/LKlt8RZzacLhNrlfHuUyR0RyJq0/te3hnsCWNbSr8GZPGrzBdS
T1ruOcNyuJsWhshSMsXH7DHQfCdIL5aOpdz+DGQx+tVbXYPaKFq1xlTABh5YGsxhxH+Pa7hjB1bZ
JG2rIb7OX64JRI+3PxhZFP2A9IRUENcZ7gBiwkK9titn+RnE9BcGsWYHc6vuWR6iWzJff2pnCprS
4aGDoaidRf4JE5+9IWYZmG9XRkTT2FDRBTp4NldpUDPVZh544vH6zwaDxb2GqoMk8m/ZI3vZ2rw+
/m9D0rNpX4S8IuzV85EbaRE5gqTGY08v20S/3hF2CAFW8eOz5Qdr8YcI7FzKvpVE1ObpmAyiZEat
znZqh/+QyggtmCVia2CYfvHF7eluydam4Q0SsFMifOdfRSqr14pZRRApZ2oD4lSxf223c+f9pmr/
q2Z7IuBMAwqRPSf154RYNJMuXOi7lh1DSNyQVvcoXB678XnsxPxGzGDuhJqKafeuQbZEZLLmdECB
ULBi50yZGtON6dPo85lAQAyUysz+/bH4Q1KzfwaVJ34QArITjE2c+nx98BQ+AADZUn6jmMdZlz4k
BtHeSykKUOPeMtO5QHiJGHc+3C2VtrANJ53L7/pHMKZt268CxkQECYEgBVW8YTrqSRkFRwImaaEX
gax7oT++KlZtLx6DaBk8/yQPdTTaNWUvE6wNGX7+FZoAfAI3IOZRwLb1jAz/S87CBHTBjVXeFrER
+PFJ5uj0X9xCuSX9UtVH27VKSEvblWqGhItQO4SjYKQNGRbv7adfQrVJuzNwMNTzBJirHiFYR2oY
iDaOeeS+9RRUqDa2krepbVTqli5JhbXZuB1f0bwqDuOpniscfmKqSdY7v0t/WoUbWYJTdBijF0jx
BWuIsbPzD1RGvBin6hHiWgndePbBqnDzf1u50xG28vsp2OCSX3jkQl7hMIEZcRXzNmCQzj/LioN+
UHfHlrABwp75EEJxaMdOIYT9XSsEDFSPndFC8AzUDgusnw1N8VEVAyYy6VFVuy5ZiBkDvyQnWKsx
vY8zQoLI9zrGLGYnjy6WezEIdjX2wxa3f+MP9Z9HIaNu1PM8WIYtBBPi3Yw8n9myi2CmVeBdFzgT
UTWrDPYy55Gv6f84F2ez60viF6gXzqjQfcZ3oG/fTQIq/vvb2MRjIZDlgn66DQ4AT1Dd2WH65F+2
9RCl12rim+IOeJLvzz/ufGnUZq4nLm+UmFWUKslif11MFfOz89CDbo/BU+ypZX67GZ6YZQ3RE2ZF
HZiALV/C2VGR3zhN398wNlBik9G+eQ6adFU4u7u+p8CYqwN199u+G6rb1kASOvgWkFvJtpwUilEO
H/3rvhXb9nNJvkahdKz+z468YuowrCzD7l3NGxyUKee4cmlfMBPPmV3Uwi308HV1DCs7Q79rItCz
hWkY8hV20t4g5EDDecwUTE+UHzp4bdNHKFqJIJLkxo6dCjbiPSwE16/x8FqCFoSqZ5e2q88hp07Y
K+/9pvrbhz/VGJDqcKd27lliShPrqcUAhgzvsqeMP+0dvYrJAawxuoZQwmOX9e88wQkCQbVTt+jv
aoZiONlMj/w0XdqRLxq1zt5bQ5BZWlUlUI2f+MjYv7RxHZ4ZrHQ5L7wAz4PctwlN3NZR4ww6TNJN
aktSf8DWDf5QcgiFSQrUtMcwao07aV8skK0RLWQiP/Bnq0VDjrSeJI/MIxFMhdPTNsZYfpKw7t07
oT95XQmkcHwj1I1Egppcpnrao8CWfwVyhUmNU2lo7Iy310ZHhMPjqV2zWbViBwPLg0YZJMDfRcJT
DVBYPJs2hlxOcboE3Atfihxl/xkhjDad8EWBSKmrolEuyol6sNzcuNljww0Syo2miqSuulb76Ud1
IagX1XzMW/f0dfmXMAc6JdhwaIl7ZR8e8NI3Fd8riG486LZX2s5Yk5ycekkDvyroQ84twuTuSiDc
Js1xfyqj0mg6AJJjcIPYt6c8OFEQflp0+w6V4A9gKbXYL0JV7G984lKKWBmWKq01B8r40kr3oGml
CP9vbqzbrrxYKBfv0Qnqcpo2niFSJplGvc4gv8PD2Q+bs+S0gDNzYuyeh6I/DpGgUR6i7T5/kbXt
EmdMaAVkQDJG5WWwpRxVgJ7/KUf0NFnkBxxwmhlvu9tevtJZVHwvNqLZ+rKZaCRKF8On6xbs2ntf
V/329NOGyTroO1TRY2IIX0eZv1ctxwjsA82VXsP9ViMLG1TwGQ+MLiT8O22QFgbqDKAUqbZ8+Uim
2Icqfvu7tJ7VJCz7FFFMWXYolVC+++u1mehEBSa05oOihLatq1Q3fGmrazhZlyz27CPUo8PbKBt9
XwvbpShcedJtIGW/DHUycI1cpPGvvnRvC0GYh5h2wdTF4m3ZB+KifqfscS0LXwidTAscfvkVvIYf
Q06lD9DP6mDer9sb2KhG0cz/ytfys8VTpHEXYTONXwpgEazztLy+oeneHtvf4qV1wtUxbjbw9vN9
C9GnCrRn4RNcu+mpI0ClXYHKDQWQwUFWIIiFeawhBYq0FmJv5QoA8zdHRxbAzZhn9Ymsy4XyTIXX
YC1yn/DzAQutY+NWAed/4pfy7Z0WM7lvScwy2PekyyVr7FX89XXsm5u4/LaXo6UfL9wXY+TXsDKX
QKGALjosBlzqD3QGV5pNA6XAe/p//3LIc1KiC9pByW3J9GQ4joeR1xG6uTMe0DYC9XPivmUjN/7O
JFpbJpvZTb3sa7tn/zbicwluD6UC5b5memylh0k6gLTNz40TkkKF6PphWbach3YCKkQVoeQshykX
fzB+V8UhdJn8HOun2DUloo0V46LYkvbCSTXgmKke9qEhaeMRcKXBffJOY0rGVLMOr/p0lJKj9DFJ
mf6i5g+YXxSnFVnd0r6264xkfZ7Iy69QCEzellkEe2Yr9+ZCQ/4sDRjnfPGLDaWAeOIq926sU3Jf
cdl7au7X5bcFNrSuSP5XL8+d5iuTOQYcEDcPwR0cZI77kBJRj0DJqlCsOT0k43RGN8fx/UTGftLu
E/wgzjmDybjl9/BTyV8g/EDohv0X/7LlOiqPPofcPAd0dBwzJhCw4zlBmo9i2BjtQXhf5lOjWMZ7
AeWGX/CXFcuKt0Qe/X9/WAAyc1pjFt/tx6qI2+wFIngT2ILpiU+oo4tlTbQuYP06qektqilPAZ5P
VAAUL6q9EmQhJUvrjlidBsFHRXc/ni84naBaknQNvGTqXO+Qu/o1L7tiCaPXyZlxEBCg72D/mZ2U
XCw37eXtL/Nq9BHAoqiXMFz9v1TAriwyrvz2kz1/Wc83wzJQSblc/+hxV5XTS4ykwgU9TxQ3uAo5
0RWtirTJ1TDr96LKpajy5BIs6r3bJoxbaW7Uxuk469eblH495HBjJ+otqH1j3xCho4ZoTPQADT/4
+pETqo8Rm9nmVpwx5rpCby5E+qW4rivfixW7JgTl2eLxpGzZgTk+S9NSFPmaTqIaGf/MOk9j6Ik5
X/bAaEb9IyuwPlPbTBAM9uNz1Ddi4amd+fyXOWz8QwEQoJCZlaqM5T2bPTrh+D1gQnm86/hl+OlQ
OEJRos7Sl+32zrOxEBeYqB4VMJCvhiitnUiouqhSkQNqaL3f5nFO/IpYYIKHO9XOJRc+NV7gtADe
ODQzFhjJoEywGg9nsSwlObelzok/TE03YebeJSBG9/VdkXtc6bNDSe14Pz2yB2tl2LhVy/ngJ/2g
3m6swBMW/GkpmHOmpxI973z4thgad9G6VDcOXYPsp9KoSHaEx34HbR70M9u948cOLx0C/GHnPCI0
Pheg1kXk/M6bqtuJ0bJ6XcEX2kO2vmbtCv5vEPCVpZcy3L7TEfFHDHsxxZ0Wc+mxL6QgRU6j/pbG
6IWvDE8iY66QXyLInihSv5Uc/Gh6DiTPdR+u5tLlmd3vnqM3oA10Zq3Y4JA9OzLL5NhtoE2nid14
XaIJsJYkyGaUtas2oPJABcJewim1fiz4Pxq92pvhanFWTFr6PCUm3LeUFU/lScfUrTuQ1TgOOskU
+iO0E+O1u378YOcLQ/hf3Lvvaek3UUaM5zXRd2rgGjUms+PcB7gZ5kFLd2/Jz4ic437Npe2Yku4d
6dCq4A96BlpixRJ2Qq7ca268RWzv39l7Gefa37hU7h3hLPH6CL7t+JMQBt4/AlR8MoiD+jIQDOPJ
fI6CIb4OvsJGfTwH55iRNeM636xkocX2hGRg4edh27sxb1B0XkxuiQrfRTAN5jt8Nu9pbRDPLqo7
mZTiZPVqMMpPgiLiSdTPQYEVyDAZRj0/UI6gN4xRsU9Rn3YSDkeBW5QbyEQeqPL2aow4Xthd9/4g
wr1wxXVsDKulvPEfkHJw/V86QJvBe/nTlmX/ta0aQmUiPaXPYBXU9v6gUtTu4+NjySDXefoOWMHE
Fmesblu/gQFQNRQBPzEU34HWssSjX75t4ZAWitHyUhIlj7AYLOJoRwM3CxTXkW+1zWloK+RO0kXg
ZZaWGNgOy7BpowIg8efqVrFdbUuRQyuS52xVKyWDxA8cK2MaVtjGoDl6O+/c00NthdX7hyd1MY0X
zk7V2hOBMuWFWHjXc6BiuGjskNnJQwmstqwO2Gj8jojIyiyhs0BES1vEa/rWn4ScUwu3DJ5IJOZx
CwEgP4ELJa/0WLNEwUdgvY3XAMWY0sH3sXX7gE5D4UsGoqOki2/fVPcdETk+XDCuPprPyMRrjJYo
+o3ZcpcLlR+X3x0sY5LTsv3tW6VbeiPUYxmp/zwtrW7TuTol0Kf+g3du4MMQ0NjmnrXwED4CV6Z4
Nxw1GntRpqsQ6+aH5sSosimeos7sgR4GIV6Z4ngJbhjCQVtkb2tqrvZMSow4irrM0rw4HxNnr15K
iKbyXlLus78b1M6axezaxp/WloRWI3t+CnksBmoGwWHdZmaEPyGZP79ZeMxIJ5LuyyPEZbduELdx
n1slfJ0GqxbTKLkluXg2GkDIT19tGYbRs0K6Lh0nVW0y9peAGcolGMemhPrNd5uk88XqDwOg1l6X
riYvE4BfTc/LrB09Unv4OI45Ss3ngg8TO/bq3sMerzFLJ4fKig0I5vBIVTBMeNz3ZCqHdgTufMj/
WbNZz79pttrQSkzRxmnv6hB5+Siruuz4TqvZxmdJwBHq6Tkr5cX0/UvJ1IbPVeBhfs5ZPCM+dXG1
/pzk1svG58xHJcpfPQi6Z9udMeAGDArJUb7Ol/BNxYfD+jivpZ0/ol8BH4oXvFZ6FLhaUvjShdUD
BwxxefVQ4DASWC6eTYbne67iv53pXxFvyQ6COi0807mpa6hsgvKPxGRdCj9WZOUXXkxK1L47ehmg
w4iT7n2pnXYJyFn+Hc0jSnmiaRpJnHjo/pI+7Tyu3UXi7nIGiCrY4fnshAHeeJdmx2aUsaddNmWT
0C9rx+buHCsqje3m11YKe7SM3tjvkQE0rmGzoR6FJQK22ybTPx7nR8ZMaCXohijkFQtOeatrXZXY
n1e72kRgqJT+D8/twxw8N3TBcrZfcYxs1j8embZCV5wJMrXpxj+wjCn5WOzZ5uOoXIoZraggjvOb
9DXKUmyFu4skC7E0BbFyG8+tFgMQNXuF7aFRQ4R1QcJSsrosYfHOoT+2GECox8sUgGdEUZPeGcAq
T7Y4bKwnaVWgCGrtZuJI0sa8ky4ebT/MfCq7aRsVYodqAD68+BJn+4yLF31epaPDv0MBiQbwEzc7
3/Qt8UeVrQweSfrrxjlFsduwgTCiUEyXRong7Mu2Ff3JyS59+NO2hBmSjHDpnfpTsvsTHv/KXOwu
ziJDEoQ577280rysZhVPrinb+hXcGQ/aG/VPhaTbCNJxBjS/rCU0ZUYirE9aGORShdDWc6Nd+XA1
VZVHFSRFe59sVFCv6hw7j1Cn9ABGuRYNJ6fFW8jIa+ZJN5saz8zaEZq6YSGoscwd9yKxMTGYtSPz
JXdAfq+MoXIV1+NioR5Jp4zjpr0iLyrHcfmn8lZEUJWwYrDmUxlSKYD+t7bhhnkiKls9VWpOUUoV
LHoRyvoz+YxTstOW0eD8DqTt057U6XNBqtsHU2KMEntV+bWUAe1aveLqhIgCkxV/YIDPWaYSf/mu
OtJn8EO5G45Df45K252Pb07tt++JM4q+OSW4GtcEGW/mznDSinQe5RiMcOr5jGaehdN6A9pKDVCP
k7WS87vFFMylqR82hcF3OQe2un1VMsKlWLiz5PYaMVipC98HC3M58sXa4EQNbM//3z+qSG9COu7j
6lAIxQrDcUt35oLwNBoWZpkEEuOzWz/l2r6596uzpsJTsTAPpcgUcdix7anMZLKISg8BV+2igrqM
uFGi6QFL7noVunWJVbjGk3GixCIYWt7UMdC5428Zxw+jwZDhKEYwhRQu/VSKNGbFXlsQv5EoKDtU
bMVSywrdZTHtP/azFVEx1nT9hFXLcTBagHiy3VJVvFLO9t58SbDKHoMhE2Q+So2i/mlsYpbcIihd
lgNus0hZ/lZHmdBeUZIxxbkGLGRM3Rxhd7OkVoMBP824duRMcwdX+iOj6hJV6HuvdeGi5c0jZ5eq
e2ZwLl6ZlTYQHewhBTCPgGOG3ZYxCjOGcQ43C42UiNrdeH4d9vQRt1gUKfkUsGoV7Pq+gQJq2kKY
nYTk0Vp+XSa+hnmSyrnUK+S5lGDp34Fx79pnHR6YidOQwytYmbAlzoYe9lj32RkRk/iDPGV4MmNm
Hm0PPpSEdlsz0fDOqoxwRFyW/QDeKDs7ffBRf3MLIH1gl6MNE6cVF23UJv/2O58PTdL7EzcH+Kpf
Bf3qTS+6bE6u3dMCf8FbzNxWNNPLqYmxV6cKZb+//P1iz7HIZwRhgHY9yheWZaVUO/sa753IBHrm
J4ruWIPCYs9X/GRE/XBXDssB9mcKdBwla6Fxnpu54Kfp9gkPJrMYE8kwGdJQYv2RWo+De9GeFalv
EFHMCAeVcZo5vwSNct9JMAsJBJ+eWz3T/u6Ou7RbsGzax4iB8FPS+jWOGZsnqUB8hIFvK+Jusy6G
zV+Wzn2x2X6/H8ktyWzYGIJdMZSDIP3wbi++myGW0jsG3fhYn8+Typawje/lm8xYWEB3slUrNZxk
68VlVtInTVc4gQVe4Qwi2n6nxWIRcQ6ITHae7Etk1zXJHF8Zuj49Qymk6FeL5xAtWGQwhW0F54ls
Y1juxvWXhY7+aN32c1eSONsfS8mcxBVV3bE9Ub5hVR7wsnW3PXUOboXDxII0zB85Ra3TqKGzo/t9
bvn9yPLI50Xf1nNv40Paatyh08OQ1qI5wdvYqGHIvXMx/sXw1xLMAaIwxVcFWG9Ca7AXUsAFDVV/
0m+nAukmy7SbU98pAAvcSdvx8RKnXlTe45KHoFCqnc1gDBLKLVTh+g1HdRghITuFe0oLN284u50u
JyG3Qf+Ztrox4dKsPcEt0AizQvcxk5E6bzutY6zIGz1Y+HW+dEzFcMp7uHQXjbzc5acCael4swsA
z489wHjMjM2KU5jjfPQLrFqCqXIUTRLVy0Nmr5KzCAYr2rMwcERsaZWkSEHqSNkKXv9Rf+89Ozku
y1PIfFIJLYMHYEdCb1kBJb0velWzrSBMbaERym5F9MiYI+CNDwWF33bMp8vboklAbaYk+gDnqrdN
KnS5KiNLWgkQaysipLi9pgS5yPRF5SDsUw8dyHwRl/tjJM1hQn4NiuSft7OnQ31/94P8/8u+awX2
LEWNS64JfsOvpYMwn5w/9U68JOMEfCS3u47vNZLwcsmwPJL8bPg1qthbdml7ocm2N2p5nDqHMjzi
Fm7c4eDQbziSmoSavS07D1fSmYXobNXaQR+FEYqX8HLdR6H7FWWguFtleG5VHCrdUpDd+y/ntoS5
NTgBDwrNNqF4s6x8b3KDPzyTvS4ER/fogYAK38QgLDaDK3xDEwJXV9rvWEzksNFUeIEPKFOjNf9J
uRoLCpH3NYqZ+3CBeSQXHSGHUKeM+EmJHorPzcRF+l+HVbZQhJOyfqw7qZizyFAfS8x8ixty/CGh
sUGDzlOQbWPvxcXqLQkaaJVUUwkRAdbrWksUZ93/9UH1iQHWxi1h7msZz1bzODcLmw+wsXhhwbPZ
CeHCTULayQ8s58nAZCyLRPSVI8ssKtR1x/eNtNVM/KOhpazIat+CA+hNhq8rE8x8rWqtWsbJm8aH
ja+mFHdeUY2ap53ADjULyPSgsPvorAwJLcRIyLgWyk2Tap907yGoWY1nq1ZDkZIQFGXipsYxl78P
NvWm8phhshokZEMylF7Qxoz9VHXaJVyVsNoYFH7RO8Bme0YPLl/RlhVelTpO4hxiYkRYbZiuvgM+
Rpd7buxxBcLXNF5q5ABqOyk6FRMFufGfSAlRyoZdcCYpKOb4hLXvmsue0p7c9AoNQOc2ieFP6yG7
HbP7N2JT6wa2XwU/U23mahMUi8E1CWhGh9QAIgL61VyZcqHqugq9naFJ7QcaaYswRaaq5hGcHzSX
+9nzU+R2dwDinmg1fu43RYyQY3DW5WK4iji8fDreMRJz2nmFk0HzlpVC2ugWibrkhG/aL+IrDhw3
WdsrIBOdzqDM2PdCfvwq2jQFA9er/Oalymt/lX9+AdQ74zSSDj4/IYkwqq/kxUPdUNyUUvAGh4gF
v902EGem27nZd3gLffpgRffTB2Z9aGj3+s3pyIYRL/b8PvRjNP3CQWT8+MzVPH4nT8PeO1urwVOb
RjZfhihy3ragr0YEDdb+A+eC+g6GWGHrwvVYX05yVwv3EybfMRY/L7alyBYDHfKRjbvh7AoHn4Sm
kwknji+X2pFP8wpSxxZboSKrmu/dEkDTqxW0vN2BsNw9JJOeB5A4322I7mH2Bp/VV87S2gEfhxfM
prRd1KkYOffyElV4hTGsYrhIBWVjuktHL2uQs5Ey5CPXeJ+R+T8nOUcyXyHOphNkAS4PEetremyo
GQSIVO9KC97nTBQW7h4dGzD3WGpM7DecGk6B1fOjqRBLH+pPiokKwvHalw5dPV1IHSZ1rUTNh88Q
+9heslL9I0r32Yc51yZrh+lzwZMy4LdQTjZkrGyeQRak1QIoPTtxM+p78ZUu4HiAGXh/ew0GuUbt
sJAgWVCiWlQoHjw1b4030S9mHTyaX0cR97HiPzV3LOUNrf8DAAudqwtWoK6VIjtseDYr1vX0NsQY
UXFphaQK1uVDeW5cr4Ec7ubABe1U7IbN2tbCpP94Q1KRWoNFUu/BfvaoR4osl+IA64x3C2aB/y8F
+3J2Bz1xkxCegCmN3tmgyw6yDIsg0r7UR/6PxGIsKkUaTmM6Km3/SNOW9D+FYafzXpgVxpcwCbIG
9WEiPXuKV4wQOhDV0M0dZ5spWS6n3JCMl7S812zKRT/1JJ4kbATjBB+ZQGNa/OVFlUq8vVrDhqJp
X7NyAFK9UoK+FNG0sUstTf8zr6CfYpWbohI0LGlS4bhmKHi7jcrwILvhDAVLOZeXIg8vJlGmV9Yw
kp5U6OnmYciccN7xEsYL/fojAYajsXzSR1hdThSJfYHjExrxnb/mofWC1wtYAu5DUmBW0GAJM+/9
wQoIWHiEFRmeLbqU+wkh7Y9YQgo4Pqk5qo2vViE12JGw8YPb5kQKYwqC3B3AXS/0nWRquBkKQ/II
ueL5l02i9Hd19OHbGe0VlXLlwYSANctOMWJmSBUO6N1nJyZ4wzO/fuTU8qLESqVx+DMpSzhNY/JH
X+PETAcafvq4UsQaPl/38AuTbjniXV+eG99/2uBnpde0lgV6XVDfyPf24F4OI0Sp7gJBc9bXezKR
ylrDpUskf63EUX6tdMBntg58v74+Npv8NGl0hiQN9y4Whn0LkrgyUhx0eEOC3lWa7FOlXnZ5LpTt
gCUZfXktJXTHHmZpy+1IjJRCzhRj/jrurRpe5GEPRsur9TIJ70jJY+SoJ54Kb2SWYmm7ZrmaCGNv
a4fqz3DehnCf5rK43IppAh5zVIFa6WUCPJ19haav3z3DuU3ehjKJ9gOiN9aGY7ZEmUoFf0LZ9DiC
uZUr9GZfBhSf1MpF0haaN2IcWgA2dcG5edD4ezuFo5JtoFyOuhOUps041A7us4ZQxGaqtoFDdMkj
Sp9niQg94ak9xIBuaFaBY+MV3OsjcgiqGJ01BjoRllltc+1xN11VsCCJph7wVanYGpNpEGy0jRLd
7NT8LrYiqJkvC8AgzczW5FgWxGqwOT6fRD74yx+nFbNzQvLGdRVpzpTcbyQ/XOg3qsb/66O+BWUv
CI7Q4et61E+CbegtkGeRGM3H7weNlY2AvdtRyGAMBGDIo369rm/dThQ5es2SYtXJg/RcZoAyzh3G
a9d32vceBR9rguRGC0auv0pIt/CzNJbosy/A6bJQZ5fzJ79HxdDcnwhF7Y7SIEbXGNe8CWiMU11p
8jp/8Q3OQ2Y6KKSovqDccy41R2GbL2cAFCh1QP1YE1ST8Kd6PN51INufMZ27TkyAN+JjcbsoIy4z
kPQJ1YxMTNplbnlwVNbInzsc2n9nKFFklCa3lj4Ixa8sl12BKKPBNFeqc4bc/PN0mcA/v7G9YYb9
Uim7MEyCH0cW+L5hCnFDH77qhBnICrd7yxlpzxEFLYsqVhKeFX7AdYvRBxP9EY8zFi6PMjBbk/PR
vPkBNP1s6OrnPOx49AA85BhhwQqUtimgLEFlxRkdtnW/NSByxS3KPbb8XUE4yByTOC3QAGEIZoFy
Q+RL4HNq+Zomsr9shS8h8XCS4bOWmtsbsVegf4taeAf4r70kd/VkUj/tRSittzZTzIWvfHUdEIx6
zb1mglVtgxcciavXXl9yDVLgcibRkRX/69Z11cMkmQbT6Et6xIA7gf6fCPdWciZkjI+Foj0af9hG
8hf/twjqI8lXcp1qSpSvWz5yl1VFmQFGU6wya99/h6Aoa609UjyrA4c0NR0CmAzIzcrYiKhtMFF4
EpFRiWt1WvL7lXdXcMy+r9KIAQpjyjXqQ85TwO9cf8jF+6M4AebgcAyiIezdFjkJQ/RPePgMUYMY
GN1Brf6d5ZIRHW8xkN1mXbji0nBkHH5xOPNjLnlBw0WjiUQ7FZoIGwGhGM2FPM0YcftMvrx0zzxe
FZcMxU3RS51gEnm5q2ekX64hy3X5hdtkFh0FxQLstOKP3UMFMvq0CU3MXE1JfPPfCIzKn0et/2Qn
9/kxzLuuRAPZEqCX14wBLPJ1g5e1qJ6s1XtQp3p0oQ+5WzopsE8GkYaaru11lWbB/ITe9gVfLoVW
E0b20Agk78Q37wit5Pa+IDRpOo/huZiq8v46TnGGoBaKeaO0iOoCfk0R6s7GrdJqVmekKu3t3Pia
Mk5tMuUWRrLobCgj2Eow5yoDPRrtp4CT9qEB0YqFzsVD36NrAqMNEb0AFH6WW8p/rqAK2/ZJxHWr
BG5XvwNESmhNWnw5BpmS+xYbEdWKVOETk63L1iQ+qoPrmgI/YoqqSFLFhlyOhmiaISVeMg8cBKdS
rqBgxtS8ShUr6VUh+d+KaNiQqonDG6U5+PizoME7JfgSVXuF+teKqhbrSfp8BrQfRBh7/d0Yo/d3
g/KMCMhabhYL3eNHoRFlI8GT5qdaS+BjlFxnogl0/N4zKNNe6NlhFuQ9/CZk5glfFbwrRYDgQf6W
pf122M/Vr6nxY2+H1b9DoJSFL+cg6rjblYF+KVvyFn38nd3UF86RTwP0kfVN0ZACZ+6g8m8wroxS
i/qlXMP+zn6tNaItwx9Jndl0SaSpNkva5ZFxZGseyiL/j+30OXdFvaCloNFK32xKl3Zbs9i6Gu15
bvjxettli/sXKJqPS8AcypzThVXpvDvoE2SJAEKXG7NkEWzkDA8YVjBGly2eDZedtVLXGAfzcMnc
tShyT6Ey7u5cl4QFhnYWorQRG/vQCGTG5CDJqzP3nqK1sxyNs/qFQ5gS617Sc772w/IGz++7V0Wj
NttBVmUjVUEqTIgKRFCY8RqdZFeFp/6rB84GS+vGJEvM5m8B5/bZPmA4mzDb2Hf7nrLUJOisKhdu
aBx1WCx9jOlwKVrkmXrA4RhlSf918Md/d+HHYxgZvCVoOeJSsNC6VD4AnvX2VkE3A6ThNNij0Fme
yhfysM1FYfEJY+Z2FyXEgnTDrlUq3q21RrlYgz4NMRhHgQJheNTcvL9wiiMBvJIhGUuKp0F1BPZ4
RwhosalfVOGNqmYrOvDPzTIba9WvERM3kmL0sgonn/HcBmTEjPmdDx/Tz+QOjizssMiSl/oKe24O
d7vnq0sWj2a20Hs2tr2X3KdkDemzvdePG+X6jIzK1aM32jbHijdgAtwkzVAt65bnsUpxF/E6VxTr
1IL3cKOvYIV4RHquMgLHxU3W50l1J4FOqc22hCG3CUDVyaXvRM/kyNzkMBvPhrx9jo/5pvrSw6Py
3Us229Fnj36fGnhKQeMpZnDKFlElVbMGAjdQkl7HVUn3RFb4YNCy2HfPUddI4jWa2YkcN2Ol1WeS
wjF0n7BVExKgdiIIdpk2CLDMzzw30RmIc14cuCmXxQH7XyNg56B/lrAWW/6TbWozuDozz4PDVSP8
XrJw92OjJVQEgQUbQ/qywRM89D6BkKpPkmken8AcwSflEszhJAcWXHm+bmFB+hbkMXWdhBytjtB1
VL+erqdwwpeXdwtFl+op3SjAztZ9fkSIvWXZjZaGWjQGCnhL/b9tf3bPXFhgay1WRJpskyLio4Z6
thudwbzvZzizNG1K9nafCgovu3zOsFApQ0edMWR5KrQtDO45tRVzke2jYVEYFZH3j5i1H2J3exLG
vOoA+DqpTsHGJzax3NoxIsr0Cdsk9KVQll+FJv0Kf2NMnQdPBT+gVhD1+kmCQmCZcmV5t5sMuTcw
0HECg01DO763cRU5UkaEMcuzY7k48c2JsDoUp291jSKeKVtqfLadwe+PD0kIaOz+CPRZaCisBdIZ
qmwuRtaqz8kVKP/6kHDOgdBUiH9oUMIQHWyQmqb8BOIJX9JT57jIobpmfBegc4FB78gDWfFPsVh4
7FP8llyOe9X3rIQT5IZdDypMC7n12GnlEOJRgE5a9X3XC9AjduU1eOL1geasF8vJWCuOHYtasC+u
NMqV2kmvI9StR8r6xswsUcEyfVzFv4l9CEsediJ12rNl/x2vIQSm0pc3Vi8YjQZ48hKmJnrC4hGC
Jj7pmJG4QUgtpHn+6y+NDGrYBFWseEBPFC61zbYxw0xYPwNpn6qSGhbXowtraBRnEsCWTti89g/Y
sn+kKXr5lbKt6CrSHqgVC95KJPz2QYfPaVnDhlBJDjEjOmWo1l1M+ubHJG+AhRzH43DVMt8ONmKb
aDir1g6nY5sYbRLbUVs5kcFvi2qog1UTEjAQpXb8tb43jvbIBtUPQ6UyCF9Mrxk5jv/WiDEHqXQZ
ZBxIVvYuu61IB0M+y9ibDSl4Ird1zuoRum57LHQ/xAxKWDZRBz0F4OaJ9YvouTCbJbf7uXHdw3Mn
bo/Hv97cl0swrPBOyw0i6CjkpegFRLlD/nUolDH9idcWl+qIAY+BISmZLLGUeAeTd53erm7eYW+L
O+iYFfilvbHZwRtuGixOBhBemRuuSi9E6UqtQifxvxHUTZz30klvtWsg20X6jCdJFAi4dBTmFb9v
deUcUSXhj6DJ0sniUI3Zlyt5D4ONw2kJSMSrf3wUJ8IsFU//hZqJWbznwLTPUxi9ykDEx08j874e
ozeg4aKrd1P82N/njCMaDuP1TTkFiuLCTpOgTDmzPxwD0130rdHnoqun22WmVNErvW4TqIUEmRzR
/I8r4/WJfFaPrHbNYUST4KppSOAiRVizJUYSubvoJt59d7gUSbqf5aYJOC5Cq9himvAPv9eYEnBA
jfezE9Uc0fbVQ9meZOXw/J5TFrX5E1LIYdaUwcfHmeo75kIbolGn6cLpU7TZuduXEdH9V1LceHnU
eaLoPlagwNSCCsRnKcWZmfDwwfjlvD73oVJe+Lqb35ScY3KNa4A1ivsegB+Q0Vafu/tDKNbAKerm
LAyJ/jEnSYb7ks/w2jzuqX9azLndpAnULQoPyUCLskPrbcXTx/UCKuEOOEJxkcLUpBzhVmexx8sV
VO/DFZCzSRNL8XSRx5t4tBjjYVv4DCdtPGPd07s7MdZWe1zzZHsguMqpXAoDdRYY9yI+Kgc5xerh
cDsqG4UmnevdXnRrOVjVuj18aFm1o8FRnWwdu5pCjU2Ez7ST66wzN36JSVCKA6xIOi0PAXIjtFbg
d1bmAFI40QtrLqE3iNuEShoSQB8ukrFXfKlZKvGtTFq46gzXFUPkAtzZTWSiEju8jReokexP0xlp
ammPPaFNzgAk0+FifYQckPj2dsE8na1dK0P5/3cHAqiv6ckvMP1a7SMUtIzv3lsFM8lgiemeG6wz
gAun7E3JdWV6zIyf50nzbMiabBAUKx/nXQokPpNsDcwlXgl+auXGRqPj3AlGtp3MHzWSeFWbWJou
+0ZGlezSCAgw2KlU8ky1JWcWZKCHB6ERAVIOoqR9UEvMEJXKBjfBmhDYqTo9rSHOuySLGtTyVmrg
mo4mbwcfE33G0gGgcncuGiDiBRlKR62gQilmX9sKqTarB8vm9pQR25GwwFXDDveGmWUm2JXlb3hI
YxtXDuYgOop4wZKFOzVVKTaPqBKdGAJKwR4wQYn0PE1WhdvQbUTuinIgbBUVjUFlBfe6Wp7Qj034
aPwM9gaWzgaZEwadGmiaVt+Q23D8s8r9jhgSbjCrmgdxMVDdqroVE6miHaXNafe+PTJiwdHHHKeS
Pio6+PFmW1bGuZC7V6pHabBbCVSViP/oojzhVAMspPaCG4aytITpk88ic7wvwHR0CD4UTk6IBAjS
rfCkVqr5wNzOVNCdOJEElJWmJO8f2APRTSY4S6WNCjvDDDFnbLvftZPxdA1vLtia/LMPz/waiHbc
Fjp40VBoIagXU1YGBevUEZ1dShLsicV6VboeOKVRNP3dA085mZjsGOTyhEZU42dOrGlKNxyvGnF8
Bwv30nxu2HEaPRQiiskBMOOV87MPSNMKyZVMDwLkMrM+GuQeUqwV8FgoiN33RFpWSv0sMqun8+LN
zXntLvXQz77mQNxLW2K3VBaC+6TUYd4kY7/4qxwUuD9jSMfzpOAQSWs0k+5T87/TRREeNiLU+ZYC
8t9FQ0+t/PjbqKlTJ0Biv6kevpuau9baWn35+E6z4GnVxV31sfDBitRsz6yGr8PpsH+EdUwuFFco
MvjlV+Y+DB3F4NcdByXMaUonj/sVMadEmgIN8elU2yBw6axv8gVlZA+xNYf1nV12SBZ4Dnhu3NuL
eIHZ0Vaasd0iLHEY55iAacICJi24XIKvTmDrb79OQ2xXnN2ErT3HrTkROlktzA8S+ZAfglOIyQ7A
YIXwmecpSXV2dI9EsX5v0Kj70RYiiV2jlyLzUO282Yv80E6JfcnVn1loz00u8EHFtiHZ2Dykb5xu
YS4GamZLUU+Ugc1U9fpXLtopybUUBkVN6FjwNTwRFPvEQo67t+eQrpoJUnXlDQcsw/nbaD0Az5tf
PCAX2eJE8WgIUQZxGMefLaSEaoaJwhe+ymcV8v2QBZ965wBO9VW4rNbppYTxxzCRs5aCnXMZMQZ/
ZbRObEicVkW7EZRR+PRrwOfc5uEfCx3oVEC/1wPCCx8ib6NrzSoxCzODaoG+xhEjdIkDWIyotpaQ
Q9R9v0s1ZflTxK87O+YoJe9lpd/IgXHRIiSq5DaMo9pAGSXNkNAiossfm44p/niSev8Gu6fwJ7uM
m2BIIwa5GKZu6RaYx4Y7LLLU2y3PFNscJ4Ce5i7iIZdPmT0dpFxLWxEfTyQd3WZfUuDUlLosL6NB
dLJTGeMye0no6E+TQ0XmhUH0lR5BjtmbjPOo+ftHyvuI1vYQjWsgz9vcB2qTGB0pwSX0MYTpXt9c
PcJDXNFvRMVE4B0tFIj5+umRFwEQrQCKfe4ZsrGuWi3A33edoS0L7m021Dda9Fl4f781XSS4+52J
Bqb92EvrnPF4xdtdxs3hEzbUKHk69UQ/N4MtqwwpG/u4RnQgFN46ln4vrGlG//2uZ8IyprT60Jii
HTeB6yUyTn++qJBsn8u6zvufjmbzf41TiP9GbgvcmtDoMNKAdd/qUE1VbOMNV4Jvng7zMZKzrYmN
w5fokU3jLH1BDOZJHoWe+lm5bXTaX3pIdOsSuTsJZqgZLwo9Un6VN3P8u/Srw35+YTARJn9Cm+8X
ApnRfcnBI3+kI9qWuDnYu0F43SAL9OlryHE3ZQvWs2JNoV2TYwPqrhEqwtPifgy+YfoUM1mRXktY
TldFQ8EDcnee9bfaiuraXj4swNublRiEiFogxL4sY+lOsUdPlxyGb7btrPKxgFZAtnSUCBKj4uX6
uuA+VgeVroOnD76aSO7Z9ExBXWkcXxF/tQeG9MnSXwUpknEL/n2pL0pUEbM47aVIwBHfUABCRrqw
DEH0U3HPQtbk39676NjrrCcGDTDAJUc7qp+SG8WuL5NzhCZVZo2Enp1HkHj93vX89UN15Q6gjO/f
GB10SnPQhgi9v8EJcFeeby9GdeX8mSkTnYShQgiIE6RH9oAlLlQPuQ0HkVWO6xpScbfOlcZK9EMs
tK2Sg63k+9k8W9G5fj3eDK75zZwv6SbIr8rlQLM1WbiojlpbK9X8b5gk1J2ILqkLehplf/FoWKCJ
JYm+NW9VXczcy/ZzHPiCGMOGlor4l6qwWN8uZ1Y7cnSqQF3ibQFJUOxCPJrX7h1vjK1dCiTWqq8d
+Ebo4OVTgQi1mTq10sN4GIDC6qah2SbxE8NN4D3j1xr+H+cALFkrwm4fZBx6jR/x/pv/a26uMlfi
5HwnBEjDG9agGXwg4fLfXFlWTt1ZGrLo1/wRggLrRQftIVktW1RqiWdwBU/3WIM3NzmUYEJcbmFw
DeiP7mcj+9SypHeLubYnz8XvXfvFegH7kFP/OjiXs9knnwJgL8JiaR/gCmM5PbekbJggSiYD1K6A
DsdOht93khrJZkU4LkekUJpZuchMm/qrnfcWPqSkzi6u/DTldBdv+H2xpnGwH78qcYQ1MrsF7qCm
Lkr4y0jjCsaqyYDKIQ+RmOKdos01QZ2TDuQIgYTIcU3L7DN1yHZluzQxyA97WYBUx1+URt9XGypm
IVT1fnHcBxtJHbd0khX1kVyLCkQJAGziBxT3Udrs/ipXj/kjaL/LPYZJr/iizhDWkNnj1vC4lCQC
SWwNZ7enEDD0QxD8gYIhs9EtvqUK4Fpxy0w0hzT9bFFsNzfLNtSK4nReJdCGaOKFoqw21VTcQEUf
cb4NqD12owc6sh2PRbTYcsYN4vy+MH8XRVpsrLjbouUxmSCbhlt1rIWaKnBIrkSacJ2QQEs9z4+k
II7RXtrr3d2UTV/cEqbkiX3fmBFmCXWUjQNYvEMVcfOd1V87TaYI2GzhFdiHM7sP1qGcu0rcXNPn
yiAfj38OSna471X0+sdcLz6y4gmGcKJFccg0GfhmjLN/iVHFkMmNfHh56HGroVF2dkUA9UpTTyc3
c3rCUkgGLHvJgFWkV7YRZ9dSC9dXEKObFwr8honuz5wAFotlEKAmnFn5H83CajSsiBnY3X5KMN7k
DfHhRBKoZviuOfAHBzXK5lNf6HtUTFskwVtI04XwbTl3JpIhl9RulymDZt3zpddBaHV7J51IgW/Y
wH1aoMAyqco8eP17DQcTmOxHHAxCq1heAPoFk4f4CaA56kZ1J28KEKvCTHVrfoLiz8uX0tpF60pj
S3aDf+A5h0n+sIx4hi0cc4e4Z+Hg39lBk891H0TljsOqSWiWIRzDUQMxkUMWZsOUyNyN9SUNsjDU
p3W+X6wE9yBzt71xiwZNDIB6UBgBq4IOfNCLQF0J+nH3SbdvCjzY/ZwqH/TiES9sFWbi09lfbSu0
cNX1JSgJdkWSH4+DM2z5aqN3WvqTfHzwoSz3j0v95oWQ8Yuwyx5fG4DimnqaJD2sJUmVJqisrX2D
Jg4dYfT9Su9ijdrTBKoeyI+8WeEttie6NXydDwtvw0NdVSS2K52EeOogLdXnUXQ+EBDI/FE2tm7j
ybNW3ejQ9nMzkJjXU9Ec96U976tHOPr/Akol+RJEdrk4K1gzVwiS3kKZajVXO79KZJvhhb68sN4d
Kwh69UVyi0JcV+lPJEAoXriNYLOjGnRNDhOwQAlgbtMTR9w/xuNKJw6pzoehCyXlsx1j3DAMjMQG
+3x1WMYLd0qq7pTLfflfwrim8hWZ04cWvjnw0ktgbCcXBWOMX6GyitufoDcHOvUrzQcwPgwjOfdS
wXK2mlc16tz9NAzzY8QAbyYgsM0zoa+mqbnc6jQKd0LYtob+z8yv4uma3vSbQgiIJ3sHJ+IADsu5
M1UZx+v4pMPUFWmMMukc+e238fFFCHL7++G350Uf1zUaEGdfI1sptoUtj9gWOQZ7XVWKyPe2wrTd
1ESjiTkYv50h8Zn7WPfbJddVlVAKMv47UmZ7moba7s+OJS+1Wa61xr3uC2/T4tw11leeSPcJYNgu
j240ceBwP3k8mqndGCuXWQg1rwySKjZKrL3knwmFwmfWkHJUopr5Z/tXREk+/uJErGVkGVqGbXqr
baMYCtaDkhW/2My4mYJgKfX1fcNFHXXfYwkj9fr47O7jNf7jMBUTJPJxdDNHFw0pthAIctfveJhX
+SWBqLd0swH4gSar/6ocJtPgonNg6MMqS34dQs5zXOmYQr+ABPGmVfGiJOE/TqbbBlKs5uMxTsqP
0l6MmgXWtecc94ThZJBpUKmUW/lF/H33yKX7EzVyuwsqEQUGQXMs8dgoRpyulP95Drafdqoh8jLP
Fi2nN9DmlLyyUvA/LB28ekjBxuZyoZhxzqb2GNRh+vE53AMHC4G2/DS89BxQeN6jlzwztydF8WJx
BgFEfnN7g9Qa7zd1MiXk1PQlj7RQ24yK1TFO0ns0AnA8IMgUrLFHoXQ4aoZKkYKCOSWWXyJ8WZFe
Bd5gP1FojAtQY5B8eUp46ZJZHfHZT+CKZRQmPihxG9Ymqd1jwVEP7QUza/zLKXy/QLtz58fKTVf6
BPnWw64c5cU0B2galRE5IrIooBsR2PUVybK29rNgtY1uJOjwMU1gWot1I0gL9AhJJDlxczgnvyxs
eNMEHMdQ/aNNQzhsfgOtFORml0oLCqXAZTM5JeVzQre0OdPf+u9GKEJ9vK7sNF3GeCq5ZygjBznH
mJyXSvUshvsKy5wOEWOkdq0xB3HDbw3cC3HXEGqleWuuNIzfAJg6tPtQxYQFcybZ1z6so7NIj2q6
ShlB5jtntKwjugdCYKuv8mRAYJWBr+GrXge6VBZPwRvxCXl4O0L+cSTCUAkGxD/nddPAgP+r3RqM
B5ncRoAjYSePh5jLOUl5g97+HTFsKcIBiDuPBjdp4ls1FLazsnlpBKHQcw+3RC3F3em25/Qf1HU3
BPM9U8z+9UTu4J2+a6+yLruS5Acetp+/aVIiP0/UtaopqqhSJdccwog+qNKj8VKS4BXgWKUJ2IPA
NZsN+ge5SXqC0jlto7Qrxyk632xKxd5ujMvGaQGAV2lXY0HyeaUCyajwWIubmmyftKVeIutHMsU+
QmYKSwxBSofeVoijcTSVhFh+JOE3rovXyQ7AQ0J7+BHqNKvYAtbCSKBVZ3L3V5bKkexogtYSrpeC
9QSMU2aBcDK+Cec9vToCgq5iYfE6m+D/Av/55RZZUmla79mZ3+oVHGZBr654c9zu/8rj6B/tHkIa
LmDAfLRrKcnsdfKsQr7CzfWY5FSP/la3lPbPVS7BJPUX42JBonF0VUlcJwQZvpKqZUPnt5o3UBe3
E1jRr5Ltm/MLWAmkKQgVW3P1CM9hL8Rgw7Oc4C6FUANJo4iueeqdotsmdLfGndvwaZkJMJFxUxa9
6WtniAp+aL68eyCaI3YpO4oJ0q8sUshqtDIWzLenxpyRxZCbIveJjEZ+W5J90i6oyxRiekoMedG5
vYY4sa5rjXQ0kQgxzvLgOfjMZYMB79e7IYFn94kMoSSrrq3ps0REZsv9kP+887Yhn8dRjTnA+t6S
LJi2aKBuPAGLO90IWmYBFXgsX7MrWzk7ZqWozxmpUCtQOS+FyS7osT9kWwHVWxqklJiCbuyPMZfy
zql9JmLrzrLD17VoMyB3agAHkJbRRWcdJv++OuhyUnttWnECqf/GSY9CJtXFdi1lQwD400fYiQNH
Mn1mWeROM7tMP86Rk+lgv6EgXDTe3NJAzrvGS6SEVL0Dw3LAIJoV4chBlppk87u36hGZdA7RkAaM
LpYTEBfhszbnOXRy+P0pJOH3FRziBWNwcW0Nkt4DdH6nF5yTnLGYW/FXLOXbtFgbhtiofiufulSe
9vhPQpxry1VyeAiX3yZ1H//hcNaXHSuc2wpESXI0x+JSRRzJ5YPQsRaZYqVUQ8MNBS+poYFZnUdE
gPXG53PUSqDqL9ofs5BUTT3iDgQM/ALGhy3qa2zHs/8gnCisKULRAJ/tEuy3HX4uiOemAIe2KO5T
SAcPlkzi6sswDZiQqpcT586iMtb0z7nT7II8dQMqw27KlLhUBbiXTTczdtcUD0lYs0yOBvmGwYvc
9KplvAiHQv8f2ZQqmOBSppjnKXPdEgobXXMQUOYhLxgkTf5ZFUhOdZwT0ct0h5Cl0IlmrTouMo+W
Srsv8JIyX+26mUIAnC/rxtf+oTyYvf0qkjNDb6wMuLIGRdMVBLh5tI2+V/8FAvNrGIVcOUnONssR
W5kGXFmGwA/PE/gHOUJYdULomgWXDKEinpGzpWuUOKpUZnspCk7gfYA5JFGZ4cFpb1SlwDRPeskf
xPWxFpNn57Q3pBPC2TdihwN8SQiQWn3MymCumAu2LuHG+PeeVg+/ye0t+7Vsi99AUgr3z33++trH
MGI3b6Qfd9lgJ1f16bJTOFBUrcnEz2qJrh/ekXwo5J4lnIuuQlhBU9/kkDVm9CN9OjpsiTXLR+Mk
jjCSKdp5AbeeWjKzygehGcRrGLTgvF2pIe60sqZAb85M/k1Km6mowzATt/hLUbaiUA5keYKvxPNt
/nTSakWrlzbEqYQAhdRwyjnwlgOm65IZ/jNiwrGwGwBCzSFz4vF9Y4ZGMEG4t6iz/mwQ4aH3w1ub
4GFjBqdJ9R05Pfcs/coXKhLUVEBKAfEZYUc3VYHkQ9XrL/JQYT9bEkLvHFsyWZtbeLx31m09UP7J
sZnt99KjEQvTC1c7S/B2nQP1q0F7kP+gR0jhp4sEsxKyhVWv9IYTUmtCVt8uptxKbnxe2YK0ba8i
mC2mYhPoyFeVhgvhEYt0WAFlescitwajiGGDWL8wQTS936BayOcaSo/9H5rW015aSkgSrrcHa3pi
6XrydblGJfDuo8wjbtPQEQJAtcsEbwb8GJ5SrND/O123Z8a00QQDF0O0fuuqi4PWEPnP+JTwFN7l
BWH3yZj2ikYH2Pgc6th9qWotIzwSys3XJQvp2q3DMVaa2ZKxkVvfnqEjgswtG5CrjvX+dPv9rkCu
VgCdLa0WA4hx73oCPPbMbsU+dW18YBrGOChQ3vdtUz5lTGM/0/L7jVJE0nSaMkQ4K3wiL0QS+FBA
YEwtqNZ9Mtqq+RS9cPwx3NEJT0X8XsERPnPH/IJN3gR1Hy8hC1GganXjCe20gAZiIJyBrIT8n5E8
KyowylDznZDRQITwHKI9vw2gy+IoW84A9XiHHhiejjzP/fPLFQwSt+iSfNntHC4OJygUzcYLfxP6
jBUwIEdxXyRXTwCdLHm76L9DGvJ6N0OEexuqjwZS5/GP4zL3EbfWftDJE7rOt7i0PzY3vz4ImcXJ
1Va8FU1d+6bYGDJKSbk1/LLRiIVkIL5NSvltFWa9q4rc5BL44RZatPX9eHENwW2tJiwht1tJwQjr
sCttIBrjfy3h7ViK9Lb86Iks2JkMEdxC41PRHm28+TjU836ABGriPRaPf8r8SWiYZSHpOEN8OGQV
rBArx0XdKTUb8VMtB8jTZWUEk6eqhX1qHseg6RTCf9inhsvj5X7RRJvDo8/qbKBpqnFFSGTdTQis
0qt76g6kUo6VMEUF/g4FIsrTkGveHtHrL/K19o6IkCCWS8dKhVqvxsVsmXb0H4F9Rs6gp764OiAO
NX/r18dHq0ONhZ6AftqpCNkZUOxBPh4eT7/1PP2u642qlMh4lITep8LYSvhBgLK2tMIXtkFXfTyv
tZU3xKhyZ20a+yP0MtMSwot27IhZqZkfchAsXOgIDWhffV6Lonx7NItdv2JJrWlZMyN5Sa4n5ICl
u2nzWfX6f712Luh07TlTCttFay52SKMn0k5n61+mOWNcg8VNy6iVaTqsbuBDmvgEVSK3+asNFVwy
MbFTA4onICU5ukGIhf2hQC14M/yxxQDsw++c2LOkeUiX14Ogl8fXMSWB0B6qoepw1HY5pT7Bq5TC
Jp0tNW/nspFsbdYV28srEpwdCMNo71nHAfgwHuSM3Zfj4l6sWEpm8cY3lgpjQLPrlM2kayWZv18f
rNuDzmAk6ak0LdRzKtIwWbaPoqBg8UqGGEFLPY8xx+vNtZwzx7GQ72hYoEyLMZMj5AXyyXFsmJCD
9RjEpinrkjRn7uYrdwOzGx5dcLLoukJx96vrDRmcrgWzTgserKnmlte/VAgEaR/ipZ/KreQrEiEW
e3NUXC3+XM6sIDuL5q0PPizpFS+EBvRKe1poJFU/EedLEuHLPSsixFqoLHy0Uq3Ck7qzDWmsIjtR
Ivz0DcrtHPpixX9xPV4+bG7BVREEHEAVwmg93nvTiT7eyjL+hddzeym7ds/vNmcI5Vv0ChBBN0CN
0NhvB8uXKHBz/fW8thkI+h1AflwZinhpFhKCHlQhMMwgWMHiedEgzG1lZtHGgSvP3AVHy6ZBigQe
tpEKR96MwhOvq7Uztw7+Wq8NZEn3+UhRXPqs9nmZhPR/xEfQiq8qhNZ9Bp3icRdEnWvK+noT8tT/
8S52QYj5QqQYBV156Wu//8HyAergVoh3Xer6dBLD3NFfDRBTGnjhuA6VuSDsnRdsd15MBfZaOwot
Tt70ylbkEw1R5WxG0iPOzt/OAgH9B3UbolX0azjn45/0Pqe+aMhJqldV580skMfhMD2UfcoyuDTx
pcXsk6eD5BkAnQVlNT/3hgghr9XCpExuVSXAsBGs5VuTUi7gA8sDVkpomSYafoN9TrEXwNiCbSia
si8tJUdOQEiMrmKtuExft1cMepo4mMZufajKY2qIhR/JDrHjMqZNetjE5LKYjb8BvAlzkKETMq2B
KIWNgS9W+ZGLbR9AlSpnuICl0Hm1dmxtBCLcJyZmG2dRzLaX+LPdDdQkel/pvOOHZrP5NGBrQ0Sq
erVrQTzHhNipueRughrlg3ZfXpzze2ObrxYs5B0eYb3EOYzaIeP79nhHXfpcrjVdiUTmVs3sOLPH
z5LDSZ4WADJLUrEfZE/JvqPmSjBDe4SUaejjDoh8G//wjtA5dRQ34WreOgAbQJSSTSWCuau3SbFX
jdkvJY1n9/Y8mHoBSU8FD2mE+QkWmxt2NV0pIz/O9GoMUMCFcmUNC7sUW4Tk2DftRRTAO3gTEpPE
K9/PrHPTm53VELd1TXlo/hO8HdG7F0pRGI3u8JhmmzFbrbzCLXP1X4TZ9aWixSrl5BpoltkBhiwU
8f3vjVyFDt98g2vUAXfPILkEAvXXK0otZKDVnBHFp5WlmSEKFVrp4wvocES2sPdCn7zHy5E0ZvJl
7D4Gd9aLkDr7hmnwAsy9NksE2VD7nDGY/9oCP4u5mZx/nHtdZpZry2N4lGeROS4+NROgaWaDJ6iJ
2brIJRJTpBOktFqU7s2L5TLAZnGqxx/oT0/tlF0lAoeTD9ar2bAXlurTIPBO0JjUHW9yyZRqrkgg
cDOUY2yCMJ+s+2nfR8LIBLKQnUpmNu620ZEJJc/qHAJQaUrVRKCltGYeMf4cNo5d3wpCsN++OTe3
GK/+KDvPyN1CJ7YQdXbJozPXVD3Tqrx5ypJEW42ZTrrcyKGuH2kmxJ3BjauTeVU3CdlXONg/0lYG
WdqWlsRsyHbsI5n+35cH+Ti3umqXyr2p3kJz0mVscK1zAXDh7UHzh4jpRp96BE3ks5Xhh2uQOmPz
+g+Tee30HbykWesPlIy364DR4kzsOAgDXJDyJTJDm1HrQyumicqli/Q9yOdQqGvPhU2OmST0nt68
gdqEpo5GWeMS2T6MWLKzMKdRdamGA0vzcpYHP9MlggMxQyRec/AALKFLJxUT2GZakax/kOAOMLA/
tWzOY32CyhEoE7VZWYYmm/vngEid6DlBJGDaliSjCRCKiEVdbXUrztWYmTCGXEJLwLPFgUsUPHDm
qbHvJefAIUdXX88582r4pgGM0VPu9vluZ/d21NvVsAEu2RBpie6L6mUM+J6EwPql7IzXg27wjBEN
AG4oAIMQ3EYsDBNuwRS4v9pNN9wn4F25EOIA5JJSUxTDMyb/1zEvb930nuDGa0L+sEX2dDGJoeHe
uneUwcym8CjxiC09ZCAUPAxqHZxmSoRNDzznXy0w03wb8PogtsBCVE32NKJk9oYdojispqd2EKsR
bWM+RydWox0kf13vFqzF3vRir6E49lPdl5SiNiKtKzi/ftpsX/AsqLZdJCesuEl+deNcRB1XdMZQ
XbqXaQjDACVm81I6f2aQEozA05A0jVnFGCSkBW2pQdT81Rpim5uY/AIoyWQHD9/Ba3z4K5xJxtPa
B9PWIT8EmewjmX+5/3qJrmo5CdOvc08hRTYr0xjUE0PJcx89dZFIbIemcTbDRMHX9ci5I67ZbR78
UqC7HGMTaoYRthaTLz8ab03e89Iztl9T3QwNvvF4QJe8ocWmFKDtmjCRyLy+7ULlssUEyFzh98OO
Kh212byP/cGGQtnv8BAmSbIevkBkKEzVY+Ii0FahezwCDx5bqSh4eVSyfd84zRnCT2ZqkqbdRPBT
j+dDHksoDYG4xwMVZGFIJ7cthkHNE/ZrNRQawtGNlXqk9xa/MJGPap7MV1aKbmJkK/YiRotM8IPx
abdOO88Yf+1kvkrLxdAcTgS9QCVq784CqardbC1qcfsqmzg9Paf3HCWzKgsizm+a2dcr4rGvkNl8
sC89wL3cP1oCDL3C7pOesQFaejHzGwHpKzvUi+Pqf9eRvViXyQ+9Xk5NZuYvEdUwPVbSWVz7BJoJ
d5/9BLO4SAhDMIwFi5Y47B3uYQJ92OD++VzedPf7tgCr/EhZ0nRpS6qNYFZ81meiJf4CXlbBAKpV
jcxXf9YEvzZO1cA0IIBpmpHlegfHFPDIw3PrnHIiLO05A+7lzQ9QYzrw8ZVdSfLNvrSKRLuZpPzb
B/kfNaWcoHKg2+hDoFYFyKJb3+LzuKs9tmSkXDWWLypDNl0qAk20ooTKMFPPqyPf/9wayk+XPMXK
G4s5IWmfGajayDx1r8rpzGzvVbCxQqyN+hGqYkwp3jQI4Tde3UaNWN6bucmOfC12f8O8CGhnOVcn
jFwbKFrjgDpGqKRAMSxZIcyVoTBT/HtxI3+7NVEA323OK7qgn8CJTZJdc7XMT2rUaPdePE+5HaJJ
dQozo3Eo09xO+07vmXaAfMJ7wmQVZb+6yHeia5/axvjFtHKNGgBr/7j7fec++LYSrkLd8ZJfMaES
hi3D6+Og60ecNL4mbZLJpbgfIMAHZX0cHu2k6AcrbcVn+VuJPOgMbwHaQruSQZyYb6KPMQ6Pbzd2
X24zBfF5A19FWWaF85ZH0u6ylH+045DjlL032iWc6n9dVkl2zuOjuYRg6qlksGlBkSJUa12DVEAz
orr8Fs8GSMcI8Hg81sdlfc4n+tf5YJuRUPHT51KkAIhZJmA7Nc0ja0klBtO6saXTQHcp9clTbtd/
eIk2zkyvsL5KoZgrUEFe//UT+Cn0k6FIj1+DpDfyyBwjBqQls7sjtQQbHiLyF1m4nKibk5LkGsna
8es4fcGAuIphS7UmJ8vMh/jaG4e76CBeST+y+eUTcG0ncWj9CzLwMfpfXCqvm3atze+TOYtTovk9
Ae5L93A8/4JUYkTHx/7HLlkoH0Zcdn9xUcVvBWv0mb5fEUuoxzTUYSERK7RzXedjHeBB/DmcHUNV
K4RhYQB2LT31SUkbME06isiaXU18OMXUi2xWBjFUAYkMeJWxlPUSMKNalsohxZV+D9kmk/tvRIwi
uOkaTH7/CXcmpdgrVrSAkcEl7MlYAxc+Xs56w5ZJqqsbugAMcxD5EhFeaE3p5o8mb31dTEDyB9/p
HGC2XTYJ+dNJblFgM/xPPy8e7qqDzoONwh10GB7/BPqVcl/lATPpN1ZomdIfjhZy108ayiEY80Xo
1xXUD1o3h5za1bGWzu9WOA/KESWXFZckauysmlHugh0vRrsvBLBpCYsqjnekOOxAPBr1NwNySV+O
3ksOiKwJobMY323xWqx5G7LUPeMReyQt5dV8/JK4CW2GBnVs3mHnAhSdyI6Z/aDsWX6tmzMyPIrs
F7xw9n5Hyi6908fYnQq/Pso5HncPTAsc36i6hUiKFstemUFo54H7n8Z9HcnjQ60FIGCO1NM6U+hA
SObuWeWgJ/w9YDt991LpCDIERJ6O67caH1S3Qdijeb1sTjcw75chFWxcfwtM318H3W2SwI0UZHUd
lIFyLf0emJ1+ToeDlHUVxQdaAd6idb8Gkm2F0lH9sZy7PdLnviPNXYZOhDtKsCyJ0yoIjV4brbsr
JCForNNZYg0hH1otC28SZ7IyycwrNf/OviV2Ywn3K4PqB6dYO66CfD0xjeLOCqxG2Zi23Hm8G16j
S+1UA63ft/2bHW1xFIFtQTnqRN3tlUJPNhMaw8ZQTakepim8SQlpY9VHSw/xO5I354VKnEQ2Kmuf
tMR9k1ijvTNfrETEig8F24W76zPY7zX5sdL597ra7TK9/KpaYicEhSNxBzHqtYGrDs7Eolg/21QV
ZnD6cXuvuSOthg6VsYhxnCSuwPWA9ebOX0YmHQCO0xw/PfoBgrpCx7OBiwqfIjgnIBasvz0T9Ycv
Fd2xhI68HfjQ9Wi1kSGV/atd7226ZJKrq9YqLut6iOhpM2S03oPn3wJK5LW2vmXq2HJV0Z4yybWm
POFnRtDnff/qRkdi0SELvT0GQZCqEP1DI6HBT5icTyf49WsMwiuiPHZ1RORUBiCrqbMQGzg5TsDJ
qxTtvxLYfD2Y6i1vsxEzgQrRaqaNkUDHWCQ6iBT75826SykHHYeL3O9deZ8rqe3KcTwjpZKYW8YQ
tCZHPJ45SIoqyZ6WWCPKtQLZgzzALsWhhcXLT4FvjsaI+oiMtsZbVSyIoNN0MUMTGtvgwx0S4rHo
rGBXK37ES4tx/yl6qVdmD+Ec/WCbTI5Q/dM7lBZ+otxjbp2BPaTwYWB3x1v1gehvBraDE5x1FAz6
QA/H6SlxXy0ypwUNuDV51FW7URkz9ndSgGRFwCuTmAmbj4748em60Y5+r3Y2yvvfZdbxRZjywmyK
9VWoED8P3rYnrmPFbJUrLTchB0jakVIs90+TXSzwN4Ijys/wZHSRxk4q/KqdNIPfN5Pjd3B8o89O
wN5TaDkWAKuNMPKGTX41kELkBFgDK4XqGFBYAkJf1BFy/YSvH3vYuX+agbQO6frNa2id5BStz+VC
hkQz04OQ0ku6c101PBCyrmJLAQTuSaLCTIv/RjDlxfooLZwQ6//z3wxoKvlKqtO2Xc+sOmLQooLK
36m1DX2+YB9cgKxTTaqM54YzflE8El3ljV6FUNf4YSomLJHk/tTIWE9Jt2KXTnP94uU4rWdn8SD2
G0b1SXV80Qio2D6Yyi5e9lnx89xiPQ6RsVtrVxkvv083viKZvVulRnEHB9m+2Nvii3NRxWFB4WxG
W+18OJOym9XWSS2vBfwKyx9MRcrCiBwucLdPV+rLX89q1pvCr3OhqLFoGh4SvP1YBDrs27kerL07
3zwnF/il5xXUEePKnF28mXn2FKydjJ2/u+NzTn99JmnaVD27rZrRqJ74uM8ioxCvXnXovzZ4ol7h
j0fbNzu+53WEX8ufiwnTxxKp9g+YVTeDYVmAPW4B2noJm0FSahK1Pw3J1z5vXJhLiM1adDi5S34O
Wog26UM+5rRFNAuoAZQEBnqK63IIkmokYOaVn5/vCMMhEezyLw7AdigsYi0HjdP062qZNXe7f7Sy
1o9/w33TZQP8ydSfNJBjNwPu+BOa7Kda6WhSsbOiya/6yO6iBJy7kO8/Nr5PAZpdWJlk8mcbeqpl
Ln5ttdGFBjcC0o6jMfOctxjjLi8Rm9AjyI7jUGwXTzE7wsKdV0X+TSe9LXgghRSDgBlY61clnVO7
oBUDdT/daV2OEC+iU+VtF4w8Je5LG4OREMOrK0YZrK3RUarn1/Pfsxh8/Rt0gDpdojIxQMk2c/Ub
FEZEbAlrsifkw2CCLGEl37/3pprdn+b0TqCfdbGX7OKMJ0hNe4HMa/rLi0nZ6MaJOjwP/IQGlxI0
rpp21A33ngNydD0eRIIVDtPw8oNm8eKRt8iStjME/4q12P7lbl9IeqTBoIkDyQePMFhfdslLufup
F2NcuJ4a8RUZfiG8t0qO+BeEaUQLttiF4A2g9tgHZaZT9ISLZtIVucH1DUb27oQYMe0yTDZpvKFJ
FlGELiSxBhIY/Hwd101RQWYO7L5wdoQ71lGk/DbvuNzQsq5p+163pNKQiZ8nUXzVgdVQoCj3Cz2X
fMlGoBhStbXNwKk5M+9KYMZLRVC7NDG1KjMUiC1hQs2PvCZArj93zRQrzrR8T4utKNOF01qiVCjH
8yd6OQ2BAhRu6uP9QQSlQ0SKfd1eaQMepJXQaVBWxyS20UrUVvwDytAZT8KKAYhS/hpxru3eZN1B
ktvS3atSygryD1EihRRX2CdnDAkoMX0sMNYlhMYClFfGsUEAVV7Ftjr+lyJDIEwHr878zCLX5AMK
dKNXYnB4f/ySOFrEBNVW5J2n6exa4aZtVZ5HRdrl+jpThiq6dkV0mvvrmlM/BdhnYZNxWJSygSz6
En3B+zp2Z3LXLLl6oxMMqejSF+MXeqXXuzope8VjKk5ga3HtXFXzV9Y4D70/OmkLOPnINu1mfUIy
bF28CHYvm4pZhaZQPT4vCxCMoyde9sxOnpxC2xY1a6j2goysVlmniGhO4f45uvVz9/c1Mww7/fLs
R+WjiRyXXihmRxCaKQr5Wrg3VP4HHtkeVOuBH44h3tOnEgwIjCKUXUjE1PubMXT1y7vM/EsLzdNj
90x8MenyfPMyNfE3ABJl4gVycUgjrm9XWbsr0PsgH8Bwx0kyHGbXQGJEwJBziGhjwMdfKBxxkGcM
5xWqbhaeaqWM8leSRgdNHLZvcxWvJ8sLBUFd7E9NcFIMx38EsS8FV/1mZ8z9EECFrZgM9nYUjG6Q
JvIHo4bHR5QH6kcf7F3dHm4lOHDUgYrVF66BEdyYQrAUob7zsE0pj+W253Fo3WgPnGepibDuWZ2S
VBL63V76LfgkpyX1OITB9VsVtFjFhDl/cLNEGcru02IfFcB/ct9y+K/kDVs8OggT57RQDaR7n84n
LnWXMO2hmlrpEL81uPSacL9xrKLp1wcfVPK4fRDwLicPFTIQD9xbWIc1v53to6etwqe5Wh4QaqMc
9Fg0R2UkpQNKpyiMvlQ72UVtMsRkl5mjSuhAVmuJH4LIOMBYcaAdaeOxEHCn7Ri7RfSOev6TxDkl
+SGXePvOUYSAcSjBskB2dEDwNrvAT3m8kMgxaEUT/iz/5GSqTsYIy5uMW0k/Um91D5DcCC7SQuYD
ptokVo0+Cgx58QxpR43gjrF+Ae1BZR1gCNQDq/mdFmgoP4sUaX0kFZxKste3qgu8y5nveV7EOJUa
JW3qZw3bTZ3uSxWhhV8kQXn6uRp9r4cpqWyD/isRbXe1vovSAQbltmPUgeDcUGkJXkghaO1ELDwc
oFMyHlZS/dzQByCIDf7j+qdWufkvFqbG/5bMvD3k5B6VKOD/Oopw/9B9qS0akFpf+RVPJGsp7Emr
i4sO7jYO6TIg8zMgaLR3iWZSn2z+g7owi23KAeUMdFirqmI4PqlfIzNHMqSJkgkPw797bHTeG9l0
wSl76Iw19KV6RPxh+2oUeMPPQ0fmTTMfYIyyq0CPJjjCBQl0nkv9t7SmLhBRXLK1x5Scuu5p2lKk
wkiReoNg2u8MPr1B03kAbOQ600hcxc2zKS9egxvBCDOnrZwxW/xzbVcUUADdTYK+shHciIzlbMkr
zDRfXP8tT/HS9zos7uqD/ou7jAQHUrOdgpoYmmvGkmtOqQ3hnyyUZzJhRtV1hlovJMM7yYxDCdyT
JWjVPD/Xu4dejWIFA6QQH5i6BGjicr1JrZHB4fXY0UjJvhcAVMSeBIctlR8m0xMcmsfyYJsvSc+5
bPFPh4QxmXIfyrcPmLSly9OCX3AbF3O6M/w2+MjJSxs/ra1kx3Bk7OwEAQuQVoJ1Idcn8h1mUxn7
HdRqSf2snFqGzZAqWUG3WXg9T83gM8wfl6VVoTq9CjnEax4VTSL03r4gIPJJ6nJBDic2kxzPDiTz
/HSX63VgRQRpihp8elx8G/BodrLXtcNE1JB00JarU/TSkB433DimC30z4laN49Jy3U/QHUJEEUSX
LI7U+tBZeFBii+IIMaXzWpgDbVKtaS0dQ5H8W9Qpaf3toKYcm1Bk/kfGvbunHMItjFbT6BZVKht0
NDFodavzQM2x/Ka/NKH+vCyjcsouu57ClIwgQ5jsYekQTRA5uWaEwtA8rNdJQrp6Nn7d66uecSJY
2TrLduP9CN24wMp5aX1uePe6uIFUBQmYRFMCLlFbb53IK2wnxEvhEhR4uB1PgrDK7Of1ybiA8y+t
sQ2AOvcVkvWbTv7rusdeNm+nBUXOaJEl4vtiaIWLIPz8Ix77INq+Tqf1MxqDb7NTKzfDr2IT+s+W
hDuyqVL+PvskNoFkP/NAfNJtFsg66LMBsBBCh6GIvrY9j5NsgHTfdShtz6bkKE48J+qRu3Mq+X3D
Bib96X+bYZ5nljquw16Vy2+lZOPTFB/IqN/vWa9Svom+6Zz6krd6vdZm5KkfJdJ34WFcpxOJabHY
Cn8GQ7w0a+tMseD3Eu+qkhszJbVYBwsnEopxNje0X5CgAUN/XP9EE8oa1Zelkp6X9mXPC08Sfu7/
/IFfnzAZc6xTSer1dupPvuAw9HbTCYaN9oom4LlVDhuj52PVTvV4kcE00TzhPm4CJIxb7UfHZZ1V
aoz89J2yHIM5lajWkXoy0LVpvqemY0qmQyjX2Eyty72GnBf5kMabj0rLxD2EmjhbpNb4TgAv/f7G
k353JkQJO9znCty0gFzR+llUY82X3f5FxLP1Xsc21fPPeJzxpOGAobEdZ2/vHNPavSyQgY8oGsGl
8D2WG1hTkCZYPsSQR8UEVByyueXLY775UPtF8XPojl8Bx21jeGgSe61DfzLBYxxPmJl01AEvExhI
zDmL9DNYgC1wD1UyiuicvIeVZQlLwb9ftAHe7t6cBl8LrxEzsSjZwkdoxbCK35Z5yrr+Zv6oTaNO
uS75ZwJTgEHw9wYkHU2ZuDsJuvdfhr8a3j6z0OBTw3GXBW0mNam3F6IUb2MD9SebDqCamnrzqtt/
kVvYq8EtrkTX8RxpqxX2SXDVPgcZsgkI6mLKsvuM+uVmd0VQ+tCRXs2p9aeYBzVb1LJttR8Hr/zw
Tw+e7wtOmKGCoMBOl/MEmQTD5cntO3o2oMa5irL0Q6UJ/JO5H6rOH78EH74NLXqd72VRnGL1NTsp
gp9mA427Tzy/DFC0z+Uu2LAGgR5F70B7yzfEmHYmB0C92q/s4wG4s7ZuYrBtGWyPBZn7Rt10dSSZ
wrRZlYzWW0QBhFUPkajKB9F4b44Vs3mm7b2Fx/eTWh76J/oPqePiixnGEn3q+hIQ5b9+/5YOHKp3
4A20RbAJUdqXALNe/KDmPQ7EfFRzHd7WersiPQ4pWqAd3R07pCF0xZxLtPHfPkTwPX2JktbAdGk7
1o8YBcVfXKpg1VExY87g5psx96lvTz6nGaPdH0F6b17JSMLO6nyx/MIgGG07ueClYAsrFdEtX1if
UockzroJc/TRXcQrW12cb34THLrYGyQ9dny1bbbjMIE7Nt08Lim+z1l0KUZl1p821vCPaRoZae+a
/kkHGBwO1OVFyR7Soj0HiWHSWuGY4G6e/yzqtb56naUaXVnzKnrPcUnPhupiutvNciv6aOsLdhUC
pe56tP3FQAS4HpkSVCrCkfZQcOPqpMDz+u4Vshm0/i+H/fyvtM31JnbqXEwoZmKiVYpO10K38Zfp
8Jzax2VaIXVVeYwJkK3S+UR+kRmobCRWfCjtEmqbTiaGElW6y+hHOEe4W4Ql9HL8zoZhwCAVnmJJ
T6ugVLnv9vAqV63VIKyE8sxBgehG+1kPNS1tQzcdfCa7UnfO/Ri9oRKVrzB18GT9lZl4F/rqLG6o
vcrCMAdb0h9jB4d5wR9qQKsW4kiyU8v29Y9+HoZejcxSv9alDIBUlG9sgu6jVSRUPt/3kebuZ1Eo
HwGgOgKuc+wTujrWwIHPuFcHfOgI+j8Q1vo+VJVVwa7PjqVYgvuOUZ63Yq0KXG9/V0mr5UZmzD3H
GmESm6BLNaPMXYcHJIP0BdaNRMqcSlQZW8V4J9YE6HYtYNp3GwAveScQBLHypzw8cU2GCTzEUiN2
CobK3HUff1gx+qLhAe+9u+d0HgExKQwYeW+oMdRb0YYU+4vgJNYfkaJjDUMgFq7rOVpPR9wDkiQW
kvmiStgrE6uJv6zvD6Vd9bwpRJHevYUdoaXy1wO9jy4zgv7VtVT7jnbZ/dKQF073q/bYS475JgWv
3cTs7Cpf1sCbcnN7Z2G4Xz0fsxEkRogHeXnTPjqVvZR9Wtxj7BP/OPPsXdlTUwPKkYHF+eMD43qk
/eBn4XyoFQqJ8fs/o3EWsOSN2KqBnUcrA1CFv9zknLl6HiZsOJmkVKidp1spluUkBB8vQxerogb5
dMoH2pX2xPgsveTqgTqnwPnpu1JKdBCL4ASydI2c0oDj4QMzgH2BShTD/DIUOO5M4NSXiCqGElNw
K/WJjOOv9PjgloxmUdZxVVg+aJH7eBF9mzHdRbnqNZ/gHchtrLtPkcH3Oq7/bXL2klv9OAwW5a13
Yfo5mmbDUXRoa9Suz5qJOF5U8FhHNm7JTN2UFvAn7fvATT0+sogp1kzsOP7ge5DJyUqeaiew/NjR
BPqp8jP9u+RTBN0glud67Ax47WBhLJVZs86T9xnoMdIy9hPnsCYrqk5ARHSKQo1EdAlpLY43zMZv
1wm7hh5xToApSvfRSYbQ42ELXW5UPFgjcpaS1ruVwExkOIHIWakqkRwMt2xyntv5aVk7h7w9X8JY
kBiH5wxueNAUHFbXN5BJqTJt4qSGVKmlrbhEkdI5SUtBZqswt1gO1JiiXklZNp0e9J1iNS7aBwdI
g8C1Y5hHIbGJhyxKNGGzn6MsfWb/+2AAr6RylDo00e5R4aHH3X/cngASadYs3S29AkU5LfdeYeUn
1RzOrP93L8+wvoZAGOS3zVGj8nSvLHF35FT0DbfZR1S4uS1q3UXNNJFCrd2auMGRQaennEYy9PaW
Hlj8Wswy2L3pV6svYAwX14tCUA3M5KCGCNvpZWc5wD95m+2kC8x+YCzkItxmoH0O5iLzHGVh+AxS
BaDJI3OydW0VOrTXT+I3Xaetkmon+deAWYFBdCGkFcrW2qomCmxEjE96NW6r5mx/JrRSt78uMB/T
P78s8bk+umzCXBq+hMzQeU2g4LeZHnkxw7olDijQUJYyVirnjM5xwbMY7Lvc5IhY8fQ9Oo0JPKM1
OCXmAUcazQOUuLcOlmOU18DB5hO9PyZ1f2pc6F4nctc0tCZbPTLz6ZI8hkIyXtsUwnmhiUkPV+Vv
VkaqK/IITFswIumMghfWVy5wCwZyaYNWQ/kBWqrOQ9RMTDDj7RzGji0lrhRj9TlHJLgjOWu9dXaI
HTwjI8PP9QIgR+bPFyy7Yg0RbMMtgNKenqEI/+dZX3rHiK/hPwOA89A6xf9rsfQc+E2o5dNKghs5
HlBLML8yNotYazgDty7DdmWV844simPH81khmTl8fbqSeIUUQGCwEGXVODRYqNvDDRPQbAEqiUTS
7UF4cHTP6K02NspDDVTBUvrvtJoEHdZqwVT3jvqIXhqy+IfZdOTUfQFX00opsJFFwof3tSLZWIKM
igfr4T99NEBsrvHnCqPdoPNegbz1q24UWzzs8TESjahvAX8m5Wa1q21oP3tZocfxM/nniMMrYytV
Fb5yWuL52MI6vTQBW9kigQny7UDaBV3Ihq5suFeeDWFkx/o2xw+xQgAGdCUwyVob90+I8oadiZkE
f6Bbxk3W9fu5d0TUsycibnkWiMOsndYbzD8rXJiyifZ86mNzm3LQNsLEWz6uHd924/5uQpNuOoxB
mqxKCrYtTbfaLH1latCF7NmXyzZURTnYrJYtpAkj9WRyWpjmYl/bqfbzzt4AMGc6ypqCz5yiDSPb
mRUOeiQ3AuCr9t5LQV+iDLS9t/j+JBYBVOJoNHEG6lrc5Jg+01tTPY4SBwNgtExxfbYBDY017DoK
S2cTOch3hHqv4ImIFdI1vcxqXnPsYzHzzmbeKocQxVAA4E+wJW8FzTvBJWyPuTDxCPH+PbagjMKI
5AnQlPQTBItC0Ak5CjENKoKDDF/jjW/+b79K1WQopLAFsTYCLIpsZJ4UnQfUyv1o1c4PGkeXYD5r
Z7EPShGgqawGKzaFZikXbntUf7uHGdveXD3cDBBIq8dsj/SKKWDCN0gSx5mRnirAU7vAaPVsdylM
ybPD6bRfZOMAqepKEBdDWvRBC97LyTJy5Nza4ivMunfjUpP2SFnp/mRzm2OP9PGUC+Ww6MN59S0p
aulnpaN02AOUoJ9ffwLYAYFXlTgPlEIrwCuuEWRloNqq390xL+n21wRObZ/zb4bj7vn3h/Y/dz19
iJBCbC0EaaXVRYWG+lM4iGwgKTVu3oRCPWPuauC6z8U886UKWyb7ptOh4FdtdlZ3iV1GGPyvsTtz
O23QyEyZ0LA8nV9+ihzXqR4HHpuxNGi2xbkQYIejeNxYGIhJUuxZUit4IN7O2x+LoZC2Z56xIDcA
D4WxN0f/kVE7p7rN1MEzNm3DavI9TND6zN59nYkSDnDLn3pZroLhIWqLf51Yj/65xVX5DoRy2rhL
j6DbVMwnKo9IMu/OpShszfjyzziVsy4z0V3xYCDaYw1rRzTnrlD79jk5AzE3XW3GTyTmxHXUll2t
FksVqdLOu0H0NNxeQJr3LmfzwI2G5YcVkixcc+wvKEbgYMBl2lt/CleanjLGtPXcDXJppvSgsIVA
GloCctPbFYg4zTcdjAnRmL8TQCk3609csdpeycx+oeYLxvsdCf0goiDvRLO11EnGF5PJdIbNHlkZ
3kxBeNIDZZeY/bqSmxEXInhRdWivbaEQmibIHHYirKkCvO8TptcfYp+7ODHMh+05bgpR5kQiYKFk
0FQcQ4Aez0CoWPVgpHCSuR6QRwS/c2ftUYCN9GN9ro4tCqz6uX+DVykeox92Qyz/H6BlCih/V4nt
QFoez189qG1DifYYvCIzIutLVax05hRJW6nYGP5vY2g/9nWg0urCnhAvVj2fkE7+EAPKQw5+UPzt
K/KNyLbWyFGs+NARCBJQ48iro7ITKbj9NB8k4o17qiD7m8KLzWm7rkM08M6U8aZlh1mK1xo00gqh
NtisLM2voNIuTWuY+qqGvmnTKoKTpDbUS9CA4U9bZPgnPG4+0ZBDeWnHXtOiuVMvSGMRpjUaevQZ
W7jE6biCvyzVUVG2OadIoA38pMrGbfMZP1SG0zvBR7XjewR4ogi8JXOiojuPjROOs0umuRhvyJqt
gi8g/vhphDcrOEuaezqDt+2E0t7MAxdrvI7PFon7FXcanNWUVW5vg/Qed5+G0JuQ9qn2c9P4z28J
NjCkXNIyK0jJNyRe1wP35rfyxKOl4fEkxJPmYNo83xQUS7f4GP13TKAlOX8CV7LhUv5FTw439b29
HlBekeLybfij5dn84EhzsoKLMzPIJKw5OGycTEOn0cgCK4p3z1TjvbWWtDza76D77Mimi+2mU5Yx
ZZvmnAjWMS3/1bAd8tjEcHrT+CCaBg90JGj5gUIffFY9Bhnagti33sAJWwsdIe8YQbXNXoydL/Vo
xyzz2colsIxf+waFGl3xZo5qHGelxBuaJ/NgY9WZp+8luWKiJuJeHOPD7oDx7h4gObQx5uxOt6nF
EgUl3SstCE+9jZ2IKQYekkkQj40U9iYRrL+0mpPsvhbtVCJqMu5ExQGIltfk2qCjrzALso21/6i8
WvWeHUBH0G0U2g+InHnf2fFEg9k85a15AoBurc4IasZ1GtGRV31hS4MKw850g7ZtnsMVh3YFEKSK
Gcbfae4XpTl3q1NXdFZ/KXGXP/GGnYDXPp+RDl/ZCRzchrDtmkCFxiFalz1L/4/AoN5FCSteO8gh
1yL37tW0KIVk9aqfHa7RBghWorXXHM1fbQVOZX2ZwGyy2Wf1+V/CYOMVp6jp6r/Bs3S9mk0Iwmt3
3w822PbNuIYWEK6wk2//qfklpEvRFLlxIebtu0QyfPRLGi5p4N3FXqZ4MaVVrI6tI0tBPOpVxi6C
PQJxJ3ylnxnPnVjPK67XUPDqZafc4ro7kaX0qzvEZ/E6HYtzUrVZaC9+LlGGcdKCasA5DM/ikoKL
QC4Dz880jC75Kdl5M0891yS71/9boj29b14Bdne/VQ4nTOpvavPjAAi3y+w9bzSwdwDNlnhCgySS
lcYBecC3gMJ7doS3XnSANcMDse5Gj2qWLp0qRemC77TKLBUVJZdd+zHkE8/nKRu4e9iU9fcUSrHr
Fduk2glHOI+OyVb//B0ZOQmF41hujW0vYPSgIEz+AS+k9CpR44XlCUz+sQEukZk5kcsVakDMNyJZ
6Qrc6Vp7AUT1o8vwZmFG3QdpZ0RA663rNLSkGLwcspamoBNbWSWwRBPTfjKpadahBRP3MwHkb8fe
v/NBrJ8SDgblcWpXisYbBHYpqjh4B8Rp/eHVun6jwttPwKnngjbUTxBp1Oij4H8HpOPVidGMmHuE
NTphK4DvatuiyIktw3jK1d2+vTEHpCKn2aFGrIrukhUGire5Rnq4V7cFGubytMvKUUnTRcsGfNJe
iGQBaMGo3Y1POeJxoSueJWno1N1VtIQ1HHrgVej+kKzKbEgpc0KSwdbTHbbGYO5ekZ+RdfrxIFI5
wWdTZnRKmdT9r/ifttRCG1Ph7FYPFE7PFE0jPgV9rCR2XtwkqdKE43SY2Q9G7yr4dP5WwI8X5Mle
UaRe9PkB32WnmZYPRFgMhsa7B5xvQJnobcddPTIPdZZJ2/Qn8KLZe47cdMaYd/ZYd32ynaAxb1Oo
zB3aTG1vqWIkaWzT9E0DaNILhD2JSMdWDl4FtweszX9cuzwFB4le4Wrk5UASG37iUvFIwapCoO9a
mh24LRhuQDTnfDhHDT1Q3xvjEsedtkd2g12pxuRFPyyapo17ZUWuecWvQt/oRWLPAxoz9cUFXKMe
++tSrn6WVNsyxk3FFtJ5t9SdCKghlvOdPsVOjTroGBNj5N7LYl3JoEvLkWez0Xx2zDWic1vjEANF
XLzl07OQhRlaK5mypoPkaTi1vQXCImL9vu9GGYCMoxlF+CCIMHZASfAn6NjNl69mqudx0hO01B3O
iRkSixfUz5xrlkGdl9J9DvkIguBtBvGqo9R95trsgyiPai/NPIkRQ7zbfeIp4t314kdEJAjgoGEV
KFYFzzhZXIVCZIO9aZYZJreXF4jKs+r7tGzH5z3f32htOTk3ksLCThOEjLQhalhw4CKQsayuMx8x
3dQqXpR0J7CdHQd3CJfG6hqt/Pr9CLYrgBsbMY2eNz4rf6v47SULayKFWpLmt8Ny0i0UfHqO4iqy
lAg/gxaL7tz0BxocxzRd2FQyY9WvJmTKzp3QFJxBx9o+FZcd6cGwzy9ma2/uhUUrQ4XgtpBf8Oth
Ka1MnvBLToBpPi3fwbR2MGfODK1tSNGuQRWrdSeoO68CBKHUSDKx2IK3DCIOj7mrr+Vh8SofP5+z
sx4i+3WJi/hm9PTsgw4zWP0T785lHno6Nc7+l/f5vNIXjtwBzJ49l2fvme8f2Q+tmhXn0QBhOWVk
hoS4eF8Wnzepr1CmL1HaKAy8yFf+q97VKdIfnIYLGKdrmEO/7+AOallMoLIEwSm77myqbhc1/qAN
dxmCHQ2Mo83PoWf1U5y5AnEL3UFpbvyHPPIvQTPsL5pWWaIL1o7fQBw+COEmcubfxSbLqZa8JXTw
wGpWqikRnlLMf6SHklemAQ4+eTMs3wZ3VB30M8Q6HxcN3dKq3i1tudDYQ5ftHQVSSvez7WzWPo5/
3mlzqxnam/6IM2UD0PzD3mt8qsX9rfLKKi7ICjqLFkbfn7G+AEKbnh8ZMuMXRqRQ3gbAa7vIBuNq
Q3z46slImIL8uHmieas09khts5fw/F45oU5uR/i3LRbr8KJwbUObYIABZTKzwrjLXBcfMBI1WeVQ
3uoull1kY7roqKnnRIP+mzLlIf/z7jtPAuuZEg+qYCttnLvH5t4ISQ8c7MSTHiqWySnwRcKhAuXe
vlbKYbcDMTzC+MSt0No7yhOhLeJykLipRFeZmBwjQRMPhI0ppsAfM+//R/cAtd2BXDU180gOL3J3
257XIP4yruT/oLhcW9c+p96cbxJaGBaA+b2oBBDsuLRazwPni3/ZCAXnzxsxPE3FZuN2mQucOisz
WFOaePVt+uM4X6iec+3PCs80Mh4OvMag7I1s6z6/WEDGD+i3v76Z/J26KDYChyChHjXmGnW3cKpp
Y5NNsfXDb2ixER/NF+PSKOjdRlEoLGZmJ/SF84XQTEM5H1gpO7ksNIkqiCcaGp/JcSw+AlDySNsj
ir+kN6ENu1Rv1r/k/erkMQ8dUb522ZLQ0g0Rm5A83XtrWspp8NW/FOZqXMQG4i71IEaTgBaH3XkP
n0aYH5P1BEXnNEUj3bnk1KbNj5SG/HfvCy4URakxBaUFJLXXRxgWx8HBkc9BZIGFTyN3FGvsopsD
cqeSpNCI10p3l/FK4q7twwMTDxnDFPp5XCTJPwWjZo4sSFhc2POge6a+aNRAkDMJrnzmE6GnlZlW
78anNW/ElaEzP25rKG/EOhuHqsMaOlfVH2Q1mXscvzdxdyl5tmBrnwFBPG15oa0sk2rNYAhHD5AC
cr8f1ecx91WFpUzfwp7S+AtNNYSiqUwbAyHGgd/zQWDltK5s7LF0vNFA2tUK6kEezgTqMJ8hdaQP
U1wXqWVQxiV9Ayw2CWar8m3/y+SyMWTO/QhBk3kngSfNgrhoqQMlM/p7y9+zrv/whJZO13v+Jcp8
aue7Mr78BXGGoMu40Xf+GzKDxWjrx0zUroZwopNdcwPsUM6YGyfnaxy1ikVOeNjoVUpqs9xUEeK3
IBHewtCjATazoqpZ/VYr9jNTiRNUf1dkwJbDsoD9V8RCObXfhqQQ84tD8zBEIEghKLnZsJs14rgu
ThZ7KS5ITIv4mJW94v1OU3yuMic/NYifUyj/awwSnEaFzKmT3MgfW2ddMyrIV3E1hsBY4tyfevqE
toEgHBCgWO88sAGEl5/E3T+dm2XQaxgqef3Tg/uc/dQp5pimesh1jv/T3Gi6QNfxYJqpp082ahxv
HE6VmJ5ZYDOgAELQ8VIIM+ujr6usYtUr7vAV+eBGS1F2dhFKOe4al+trJegbTjFVXIAEXbJlI7ov
GxGzlelpo0/VQuchPcj+s3weXpfJukH4fEzK4tZXooH04YWx/P/0kH0Hd3fnEiC0gTJc9lpF8YbO
SU6ExP/pgTnBQYR87dBekE6Uq04pc7WALeI/xxB5+3s5I4UE/h4DxGTiv54AX9UdVh6stNPUyXnD
lGrBkJyiFM9RZcZipnviU7MGPz46O87ASC8VtVnG2C0RnGn8C+DzyKXaDoBFiDRgT/EMe2mFZvRS
EN/LKvFzqgNF0X97Nu7dqQVCFrpqlUmq+e7TiDdyuPuDckmZ1/XHVc9rzxW7tRdTM2PjFgyzkES8
bEFrz3lx8t8ED+c64BNV4SXxIAhwaoNfD+/r42ge3my+fRHeGbh0uMdm9hiGO1ylC2az06R5t5st
d0zZYPA8X3mB8reIXE0fgG8hTfhoRuTsZPiok+3QHkLYLvOa8zIaBn3DJIHY6/a0gTylEnhhoJds
CkwIEtV3Ta7COY9xfqZWNNVJzSLFDlmTMVUrpxDf6Z+V0+UutDBXQ+CI/rnX4bOeVNmahI5lAs7o
bQs89jcoyJSHO10hHU0f2oTRlEbw0AwRQDiUQPmZYxclgizQ1urXvWdSXAtSWxJlPZoB+UmOZ59N
Vkl37pcmNSAnAysqAvlZoNFSxL1aw0hGHt9KoigAuq7z39GfFnqcGZf9s1qsneiT9+oidz+IEuFO
k7yVrq0YNJQb2nAo0lj+8/JXkvEhvZN0uuzMjELHDPf/KNMnhMD2bbh/qtsbmPHEY702ULgi8FbZ
76LPz4dhDKkLTO3RXC7OicE3HcZagb26/UJWhyIaJA5uQt8grFYfw8IJQljLmt/FXXJs8AqBfAP9
hC8P7JwkE2Tenn1aUCmKEOsu5hcfYs9tFFVMuRjHZKHMSzb8NnGVrmhylGPex+mDuUCMUtPcSoRj
lRudXcLXWQcBxplzpzbDMuWGoGO7m6vdjJC6rIRnGyitM4m4kkXb+UL5VqHDitpRNjzRpK7vYGkx
1xNY+I3ua0qfljEXwaGIW+zZlY8vFiC0sp8YrCScsHFRCVh9a/9izwu1bxroCrfR+t1VBDsa6Amh
6C/VZyEU2svgMzVu/UYJsK2UuDdTmXawWw09Rv0KIwprxvmugbEA2zh4pcGCd8Xbp8mX/LFUZ9A+
eJl2YPdXvsy4qIJqhwGtsgoahZeXPPmwfniFRuoBf8EzbRXKBtEMVF4P7RhepqaCRoJUk9KlM1t9
bDEmyU60exiDs692jeViaI4T792zimPYFSQf53ONo1AcovIG9n04Lp3BtEkjx9TwEfX4AE7Vno5Y
NVSihgkt4cwiudU3kns61KQ0SjqdX76jdwp0KDcub5B3aqRixYhvAHEKTI/Hxke2W99AagHOv7L3
m6bj67BaMwFL5KefBYMYYTEp32mWOyKBs1PJquinujSl3mxJth2zxle9XYKw1CqN8DrfLP+p1L6I
YjKkS7lDlJEnmu0oFi+BpMtjzweozVrW7GVrLrzXtbQ2xzcTHlm5HUZw0G6DMcO1xEAttscol2hX
UwiGPKeqKm5vL39Np/0gA6zDPlgiv/u/ofsmVUI5HNgCtuimvSP4TBjTRrNtjSe6ILHWylsfXP8b
62gCLb9IFNfZozxULlswBz6pi9Ufb+/f5jeI/7AdkfwU4JqnbX7undCH0w3MSpqeo4/lIjpO9qtr
rfUtOx94q/sQYZJ9qUYRZTVzStervKhGxw6HiJ2hot4Sgu1PxlHhu4j90wur7klKX3hVMMv8c+mD
hwgEJ5kqc9gE3ANGzxOPK6oWfntfQod1dtr571BDAdyWHDegXZO1xE8GTlnZBwum5DwPHUhLlWZj
zPsyLjyZ8SZs2JByh9CN16xIxIwpKjA7JOopqQpxVMj99o6KsXBHwCrIXUaZyTRursfpZgjS/rn3
zLDUJsvdKcf/ZAVl5fbhTvMnqTDnVhZfhhDC5wi05j5ex0EufaPFl6viJfEmf72LSSiMpOSrHxf9
EGCQFWLH3QrptjKzA+9G5S0hb4bdBBoTPQTCQztvr5pQhspvl0C9QIpN9MaOydPYs64YNbTW3inh
zC+zNCcMfxC8jhG9edxba2zxiWeiEu+nE613AM2xH1UGUSo/tMmfCSNPjLy465RGI9YHDuhHu4PS
vmN+8l9Bskl49mNVGqD5jSfmSgtNsZES3dPY8N3YbXeSgAzicWxElGF5Jf2c30rqZnTD/5H0bBIo
4N4lFmCGegjaQxROzTZbk3yPQHOSMpQJ3EPsfQtZVepQpUwsDs7e6euAynp8FdpuiY8iPVLzoHm1
sy6xM9KFVzHppzT2gcX7KKBQMpT4VQL1shg4Bjm6QTHD2YMlH5RlIDKMdoEvFwj/IT11DS/ggSqI
/XID/pLmh8wrmUdfS5FDvSayc/QPlhnsugEOn+FQ+cGmH8HxSfCr/Seu5dw0LyWgv6ldlhZ8i1a3
k/MGUozzCw1ZDzu7cNovatXXlCvgWkI4KhOU630mTScYg1O+Dco9fLVi7RyvLm8t+EzalhzHAqV+
gaHqaEEKVQav8XV93lXtsax2/u7zcOaTo0HFyzbNDgy3ZZzGSrROZKXQKOWgyNunwzw4ot1X3SL/
j6znP5GcwpJydJXlRkuFC3S1sXPtAq78y67vErBjc3yJHi90kvuIlqaT++EaDz1NQgC83TKZ0QPd
bjNYMuuyDBLGUSYKV2bIMLHfSK+fkB5jyzjRaiaUTazsJ5ghI/hJF0Og+ZdxpxmNHu8RxQl0Yu1l
e8MJ5u9yn/mSsu3zj6FLrWFJitwzhqbM9KAblbsvJP9Mfdf4/sFZfZRBUl6iocRVIOOaWx2tQbH+
5XTMJgJOnT2l11Pl0pnPIMaW8DizhfwxWzdkwLEbF2mqRhtXj/RBrpmbrqgh7y1t6PHWhztK+qdS
IUpKHkpGXIoIgkb9XS5d887XHEDvQL/0AoHdxDBeY8l2JzHgjJ9QnQR5wa13km4AoKMdBUZAul4R
4Ym1cZCmwtXwUAZE2vHeuYs85fzWqo6a9k5q+PvJ2g==
`protect end_protected
