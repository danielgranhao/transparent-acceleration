-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
SnEH5osWZ75QLB+zWvD6o0eH3g3PAOSfiSmlgs/ylVRp1yJQsXN0Cuiw6EALN81E
ExMpyymDe30iqy1uH+6RmkRvRPZWLmNDRpGyoTkgw+vG9Bh03p+ZT5lcFd8H1y04
pkdNtbjkNw8Let9t2e2eZh3ZzZBe8Afl5Z5uTws+UGs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9479)

`protect DATA_BLOCK
PFpMndsmCzNyurkjCcNio8xhG4LDCW2zcXIGIvHl3SvdB6yfWtBvQ6M7uvY10jHw
vdUkmVif8SQ+tzEyICbpKssMfv0X0KffJ2rO71U6vTOAVnglSyFFnKE0DK/blTaV
CnBv1Mb8LADwBR36E1L8s2UfnMsuuvf6ap5GkYBk09gUeW+MS5M+hMkZbn1b8KKX
V7NogoUrH5nI33YlKfPaNjkBo+geOOLD/ru6LwIBjK7p0aMll3CmVjT0ydu0mPjJ
5EIXptmXDXcbBu6nOO1xZ4JNq7IE39otQlEERAgOBdc/KTEABmMyl0ctg5ewhu6Z
GTfDgS+1NXtxcya8DmwUyGj+ewfceqTkyeUPa3qbOXHcHGY4WHjCGfQXJg9Vw9W8
RugIe9ic/RT3uK5xWqVaY3pYO0/r+kxxl+OlYkytrMTXLkl4NpRuQcbRf0R6sHPb
c6JILTZRfaz+eoJJpNbv8KIQq8K2rCzpevPXfJH8EbfJOnczqWXKlQ+W9a7iHNzQ
8DYA/wvlDHNZkbBZtiDSXVD/B75kgbvbpwZ6sTSBm7t1egRChdIFvRgJJ+EyBXSy
7FGTp9Z290xJB5OrY2FS+nbArhzIhMmwKlmysKrsXm+k3kYKGGeK22JoIcI4gCz1
G7wq2TPsP4I/Ax16tGhw3IXZw33ZA4edCmJszUo32QBNjiD/T1gjA/SM9HNu1VWS
fKhwibDgAVmQ7XUcFwlKKlmHnjp2nt2o21G7Qz/g/ZipSfpT9xJYdscOWbH5ArCE
uJEF5NMZwCOqy5ZjYe8fqbYQ+ogI7J3LiYdrLj1QAbfJqDzTk+Y49ykvSsSEgCap
dSoEEW+FySxL5+3n++6asXP9OzlY6+efug/vWq/MIAnjRYaRAAUUXFINjTBJqUsG
+tyLl0aDeP4C0NqQfiy1AKozRFNGKcz8healufP3JIWcd+1tPw5HSlA9l9qMYzqT
mwQuaSb8qJ8aXkdaVB3ksAUIoVdsDqRL9VvMepTutlmv/NSooOJzrmtcdaV1ifpx
nLYMHDYJm9mgwkn53+TLwy/fPMlBfujlDvNvanCiIYCg7u+jFvo73NfiQ492ZdMi
yMNdqm4Vow6SauF/AwQfZqbEAl9+ZEW1fVAT8ZkaoMwYjBjDk0mW92XeNv89Id1t
iAz9oq+H+3RmpNcKy6apWFiUTqwusZ9ybTMWRvomtQVDy3ql7R/CyQAARlDYad7V
oUwtyCaHigCZQ4qCFCjmqkJD59yIWuIDjh8F2hn+jHI0Sk/3RQA318B/M3V49S7I
8Je3V38Pmzh3d47FpEjN3JJrg3Z0r2/wtDUVxYX0MTeEDvSq12fIUTCqAZ7zTL8Z
PS0t22lBcDcdsyc8ooCDA3/zSvwh/urhD+iA381UVi146w38ynWVC8/VKYQD43yW
mKciX1VaOpFBCFrlCiot8eAu7QT8QTQcHx0K6S3DQoy6Odvk5EuLK6/yhYHJ9XLW
4zNyBXgFviwlcvHAVJpGwL8k5AWLRjvxkZTEKPx3wnBIsVBjOQQFQJbpZz3D0nPt
Z8WBmFcybgfxmbJr29NBMFHHefXq+Nuk9U2vxJPta9SV8HBcY4T+7kEu1SLevXm5
q7xvEjpUdHwbbuaFLc8HkvYivzTWeahj38r5I7cjfIyLxoxIME00v1hbt1imajKP
iswuq1gYZ2HzaNhXF2CAi3DqCmI0l9fKMdMvOdw1Nfz7tBElYMplMsNHELspOEyb
Mm4NXt+w/Y5cVZmRBouIVh+3QjQdt3aJHRTir8gUsADqatT4z9SeaDitQ2UM8YF0
5nidKU9ob2rCPuNIzXXXz3vYKsAgLOKGW3pfW61KV3YJ5jN036ZdAoI/u/l/SNVs
egsTau3PaqJUPzfo68mO+TmHGFy3OdOQV57B30cSHgzOyEkpQLVFBcxDY1B11Ssb
+rn5SgGFzHR7C4QPhS0l7qwZvkO6sI4WbDY/JpM6+mn6lrRKsTnb7NeV7/Yq7Tbx
XhLw2U80zVjjbRjQLDGHIbkJcYk9ymmECKgL9ucFVWwZV+Z0pAp14WLhaE0RWDaV
Ta0VNXZVtj9HridGNEU6p2oHhNUEsbW/uaVbvYt3MsfRO2aBgZWSCOuoUM0Eiwop
4jBvQD2LUGsaCga5aB9RpfngJWhQKniUyHr+CTbILIGlcFAnRUGv4swVnVGFoUln
S8UJtUsmzlBUIqFM04uDfLe7DW362FH9rsW0qinHLw7xuywhdaeohY9b0ah4/W9s
eE/29GNuJyiW8VgzunenXn9qTvjqrc6NrxH16P45/Wkh6iz0EhODjUhXDZKfuq40
mzr9KkC8rZJH4+G9lEu/fSym3qeJVJtJEWrPoXUMHp9cUBGPuoRCmlj6p4NKlR6B
RGkl7pyUP5gYCRIUiHOB0MgRp1Rpc+3Yt8Ga7JJ1heE0QoAT1WKrgHIl5/syKdpG
s0VPfe8q9hx4EKtSja2pEdROWQGCf2gSWnVpGfbx4CzTh38RmDwLEthvcwpkrSAy
SVx/mIw8Pno00xDZjAsJQriYY28LzOc9V4rrYTVBx0OKYWiqyFWFe2ggLj6kFFHP
SB1uUDFrvukNKpxCqRwYTttTGFc2MtopbA607do0hMKXFnU5aCGU/LCIZw30WXCx
AfJVP+ftJkuFCUBq0r/Q+0qidypk2OqwF/6wOtGLJJkgDzQ8cEpWXXvgxBOxnVVL
USaOm5EkWB7UhvIEfeMV2EWdhkZVz1t0NKwBCviNEE0dapWf0D7Ysr2MvZ4lJ2Ke
nmi6S3KfwX5R0MXXqCHyTMjD3kqLxU1tjCx3KwD7GnMWE7ZLImn+VaK1YlfVEyzA
vf21P9L3bYlV9D8cCyc8Xfk8aTbgrwTRAkMrvTFwYInrbLgFLA+0AGO89GPrQEzU
UxYgl12vWJK/yHuVj4nygsT6zWa5swoNrEMwzA0LEKFeIAVcj8bQn78ZcyOE/dMI
el8KXSYCe4bLGfRLnX3fzY4cRugX2R3OCQHGNCJSEN2oQH0mKy1PdDtWnRFbthwp
Qxs3uJRfwuE6xReZ0uLCNPM8fM0UyKVJ1x/4AIyJpSeDLhkLbwSR2UmFH5ewgyM/
6b0tFwpdbOPkJt00bUoAtOIc9oIdYsw/Pw1L/gHMWkOfGU0r9hAgED4f6k0s6CXk
zthUYge1xuRmrvqt5iwEegpv6vwA5516EJZ3zLcLzpX2m3qgicr2H92vncGdloJe
/vTBcB1olyhgG9XTL91Jb99oGVR28GFo7tIyib+uUDj6TQ6zN1ieV1qRny2UE5W/
84iGlqeg5/Ih5Cqe6bJPdxGn9rVODk0eqRT0GFP08NBBjkEOUZxiHCyBfyAX4nzu
ts+hVxVoqIugmObXCObVTwdiDk9OyZsvN7zYoVLwkqkR51F8xXoL2BHPgLs2uKmJ
QTHSapDwPfSjeFb8uhiBpRW3ssbbe8KktcVbgxHPVRgJXUyA+uFV4EAT6qELGf0e
smEN2KSOcYIJvUhKdyDRTgm/Q347jFCELnyG8oGv5GMEkUmdBWneG1OnRHmYnhWz
YLs/OnfyAmZxFRMoDhM5sz4NtL0OAnDiqhXePrMTT9oVS6QXeHEYxUoomGcOcQWf
8XLdmOqYqfQVjDss7n9eFtuJGYobSGonAESs/wet6m5NKDaggmO0TJYGbqt96siz
QLm8BKj+8rM23mIHkLNKz4Vz7307qCxUyAF2u5IecNOvA3itT/iH6rDfYvjUlNY2
F733Fh0pRA+r7ENtSNoICBr8K/e7OWcGCDYljCUF+IAdKp2MgHP+iPwSSTLl1zwk
d3oBUk2zSHedClEjlZexYziH/CLjp+3FbdJuk31U4eh2x+9ZuQn2PMpWr8IfpajT
zJWNfrw0m2T0IfN02qe8EG941mSPo8QVQ0rhEAwRxbGb2PFaUNpPUqSNDrEhN4Qi
uEdDN1EfkaCUWCfHQfAu+3BPrMrG2j+np0CwssDfgUBxiqUsI7g1aVlMAH/dsN3Q
ne4oUzAPDvm8wzDR0TsOxL9k6KVH4SHqkwVLVF1czr2ZEn8SVh68FqBkbg5YPcJN
51A1WCdqo0SuE1O98i4Kb4176i1nWsaa1IK0/ayjve24bXkZdQu37cpaUCuD8qNT
tHRRpuCxl3gTINnkqt9yB3DaPqm+kJ9TcmuZTXdwhj2oJI49Y+d+uaXbKWWmIDMM
sQPIKtSOUX3C1kXXUIr95j6ZwR+en5BiZvu+T4qQJgjJy1G5SLnytXliKubazzC9
eExv0QJXzoSaMh9uPFLrdjIsUe24W/yH/Wym6XTbs9fiMBATKySVWFCKr2r3zxNW
5YQ/vDsyRUfnWInd1A+cNVqH0t+AhXD9La0ZUZMJ0GTPlQcqr2459u3AIAO8RXdm
Gg3AxtKScs15bENc3dnlB+tVZbBAgkICEigDjv8+OpgCUqpMzuEunYqvn+vzSkqC
V3Vqv0woEHM3aTed8iFUEaTTz97XnY3XnYagYbENUaUizpa1bjZf/zb87QKTaCDA
OvAYEFGXqedeJHjzIiMPfx50LdpW/cTRyVmCQ2xd6i1Awz6/1pY3ESrVzpUZ861C
iQDDilJVXk13oDeh9TP1lwu1JmzeL+6ZfFaE2rIxAcgiYmKIVukALy0hIaklso07
dSmP+XN7DtnEczlvJ6LrskL1CD2dUvXHUvqUGmWppNFAGpPc3uD4k2RBMRpRH7EF
LWoWRbrMM4d7xbbrMnXxywy1hY6WjjMRRgbxmRaHdmnC602ZEJqBmwL0OAkH3jZN
8a+TlKz+FF0puZ0+clnZilOTqjct+Jy1NRakQFNxaXn95BTATnT5euTOBGmrFFof
L0g/W2oi3tiSmhyWPJZbUb6FKosFJfHvKFEl/ZbnVJUrNU5l4PK1SEZuh7H8FS1u
vtLuIpT0m7a/VaPgVvG3SR56qgLoAldjDCXPZwRY3Llw2Qh2TORzAaj5So38Kkua
JlUhc/PzJU4uQS5NxScKCWPJKYpiOPgsRxCCeFHBhwMGZXZCWlAEX00tekCQusPG
MieQoH2IQ8dvhiL+j4eDg/c6rpQXjYNH4S2CbZo4/0nT9ZholpibLNAy83YWGrnN
w+2d/dyqq6TXzRFqxK6Ow7aeVOMhHU55Mo8QBjxrcdpvSARrpS+USXbQAhOzO5D8
0bvx5haX8GhIDDZG6jDK5lW+AvbpX4ATmtqfOShIHGPoldsIsUgru9n8Q+I1zONH
p2nu1P47iJUNbTWq9IU1nEkTOrT9dMbM7mjofcCaYNhM+FGLQgaA030kBy4UkiC8
oA/2Wi9VG6JU0QtJzOoO6Xwa2qBuj1BLgkVLxHJldmdI3zAU1iyR6EpP4N75t6d0
zYW9KrLhuoUiX3ylKY+LbvKI3vtZ0074SyNSK3SzzahSeTDENpEv4gIlyF+CZ2rc
0n22YAFjK15rfX+b9vcJPOLCNTYp0+mqh9cHf0dJm5wljOs96qB7EFQ+yuhWgmDb
wiF3StzrmS80VmV99g4NQCWUSZ2WDVgos78pylFCLJlH9WXX7g7HxaosbgxbYz3u
dOy8A0txEnq0hmmtotqrnAGV85NDJtEdQGdIgORbI/n6O0ea0KGmNCtFyxXM4eB2
7XXAvTxLvYa/vwAEdeST60G0LyqKi4qZoLNi6XhjfNDDkhkQEiB80U5ziQsLf/tD
uvsHQ+WLhdIjkX8PRGr1ylsdnb2LBwfhZPnYXoyI9PY4+solgoiUWlOCrocFSPt/
pTA7IKmDeu5mO+YyinwJkTfIHFRIyKjcqG9jhIBMHmnOCOXv2hSCa+SU0W1FC2ur
7jz1ricrU+9woO/LL/oqCujUouFLCdesEl3t7DEpMjI7hr6YBWqfXPV6X9+MnaFg
psA5V0InzQW1FZfDsqFPkQd1WWEjJtu0VMJQpxw18OHqb9nBreMnxxeaNyQRQV3D
y34GDbjI+LBBJq8djlcqXS5yzzqKNo3iZ4FKUyYi7Dz7xzhV26NQ98x5FYA4BrjL
F5cX51/vf74BGRi57eZP2zsYcfoPN07QVs5LqYMJZwiKGar96HYqG0uxA7AFjUVM
C4JQAUxy1isSIbFCiLbmKNodyWdYBP6Rt3XRB9INpTbGAT1LgH0phOUgE58qL6i9
INo8pdedii0zhtg1rTQTHZR4ZU8gTjg/WOZ4y23wpxDh3YGlAAz53V89rfCk1zHo
4OvICBl/bzJJhz1FTP9+QpzvPOjwmascUS005t4b92d6fGahOd7HFCOoCAagRRHy
4yASgmOdxw/iiysCvOFk8mRE0rMVNnSlkYX+OKf89VY5Yv0AqXSVMtk6Wt6Vnh8f
bHRJ0ba5I1ereLbLe/5EuWi23VGy35llPXnjrmeOQ05GeBNwV3D6dtZXX3NuI4sI
ik+ClN1HNDE0aRByaJkmI1o1x97WesWZgveWkbT3SkbfZ5dK52BWv44/cs8++vsF
ecua2HN7BeumfofrvZEqhldD5aplSwowicbmmo96MOSRXfBOQbArEyeC+5K8rCcQ
K6XlkXYxJYuLKizXmulwPWPXF2NsggXwo8pfKJsIs2Va5MDJRf3td6g/YzuybsFq
32v/Giz4UjfEkupoM42E7IScAMnqG1bhRZeFbY/0TCegoC1B9GXpt+5rrXJFeKUP
6BXwmrIdvH4E0nQDq+kgf8co4ssESJUBHKsm2tHYeegSQwuo/iLhyxWJX3CBLfwB
v2heBQY7WDsZze/1f4vrkzDYFZ1MHcyLWIUu9wz/alBRaFZFq+BkEMheiDOfAReU
bDr382Qoaf+cA7ZwGK0pInpJYTAfN5Dd6Mx/1lmVQbh9RolepEOnzrIs5LAWoRwG
ul3Xui98Gs9cVf+OQ6nYFeM2+hhL95edTGRH/Hr2YyqJspuFMF5SnZ4cAPMUxm9o
SGQmGqhUvVl04YMJkeu05YuZ0UCS4Dn/9bZfYI1B4bIr6aGI6DuNPfv6B4JB2qTR
Cu0FMl2rG1w71jHzX1Px+EaVOpFE8w6dO8zaQpRm3dD5xHaWFPTPvlfBWy9Rb6tF
PN3kDfelr8vFEcwJNrGmPFrIbTd4ILdRmiuxFgu04qI1L/YVLhUe8whx+lz4hvOQ
HHvRDHUkSTvVagRITaKavW/kAcedOtxWehviYRic999CjfZCip3f8pt/UHf0KYsS
CNm+q+gWxo1OpY1R5Hko2QCEtxTglKrVH39gy0AW3uO/XRIn78ACkAD+ZAPdTeW1
nAQBh+c+1c1bIt3RLtIYAC0mLRrV6HkOZcPgwFPmqitGuxrU9ymrzgWhQeOQs9Vn
K/du+Hpfc5+IUmWCUmC+zIojehWevgBqowhL9f9HCyelpJx9GU7K1Mw6q1y6lEEq
JfUk1mBtvWfkd6/XlzDi9MV9cSU4+nSJQHdYL1X4jx0rymX3DdF66Tuxhy8HzKvw
oIOXbkSuM4xwm07t5jkG00Y72eFeCIO4S6pqiovS2hYwCjlSpSij4phLWBKp9l9b
VZp5Y8r/b899z3p0TlFsqnOv3jMwdbCMpHvZQ3Dac/HtVlvAlKbmnPIKROQ2XAG+
F06ToaDeB1Jl5PjA4ar341Hw+xmNGqmX/h+J8JmDGBDtSe5UYl2uCSuiM3c4ajV0
HzYKOJcKMtAGTFRAUlPkgfvW8oqnsvV47pvvrHTWIWZwSL0ZcX75UZ+VXN9FUX73
YYajUVuGDUp5CL8qc6N85n0/axkrRoEH8A1COtr/TN7lJdQ/NjOxOvM3eVgt+Z7d
NWSBelYSfHXI1eWnFgI6O16vm4DkQOV2MLUzCLqvG98bqBb7Lcnav63VwNyzoXpa
JrtQKRHfNpqV9PjqQjr0gNqYlMk63ShcTEL75DvSIOjfFZKSrkTt66HHgsZrnmkv
ePI8ixRslIo3TOk4hQXuQxwL6Kh0zdfcZNitDmRbxnldX393sBR59cnQeuYEEIK4
guzYXlMHel1+tnoRo/HVyfHFI6K8naATycmWFEeF1Q7jgpLpGQDxaq+uEYRwDwfT
S3LHei/P59Ya5pjZayGyiHFQCsJu4IfHmx5dtA1+3Vyqez5oIM+VLzMq1oyGSrgc
TXTZ9nlwHxaNS7EvjG4smMNGopmvokdJcPr/bisBtssiOmHpWtFNZO2JQOW6J1CK
8zb6oAUFFCi21GshfEphH4VLiliTJvBPSEG9GmjQGU6h+ZAhH1n8fzWUKPUDPCJC
8lL9uMH5I5qzT/cOHoZYEvcncIO40uHKVjZP3hUmspWZz0ZSQbmatpYI+FjdBkpp
Wa0P1P2YTGMsAKwejUXgkAioswSwwXbEykXHjD0ZJBU6gO+AbfJSx5Np8gTgwHWR
N5atXgV0iwti7NR2Lz6oAA1OnghMQtWsOP8V/6ibdZOiUTIMtgU0dH37/PGuv7Hf
8csAWm0FrNvP2KVHqhuiwBe8y8v23pM1J+VbN5M/+sz6HcscPscQuf4y4URi542n
lUHIynJ+nZbWs5WRmFoyFPRnKa6KfJr4GgUBaMBdeyXwKhwJm8AFvHsq4SkhZJ9W
5msOAlSR157IY/W1r3GsWFocqfCVtf0FoT6abew+IoT8VFgQGXv9+Co7KS4Bg+M5
JQQy3dBsKJyDwjGBXkTWVojm9KbTbbtgExOF8+mmd41lHi95Gk4MUHu9H7CUj3+V
1YkBz2Qay/eNI4FOaMw3OUk7peZIFDIhWiwWM3QBpi/zq/5W31A00eK3nHRH6K7f
boBwBReDWTPlY0fJpw229v9/ZfM9cc14wLQejJ6HfIdbu2so9Ei3tPpfxZWcz78B
+bOXGgM0gI2UYZ/X7TzrFr8PWWa7k/W0nlM+THMVEJ2j4VDl9hfcGbIgqt1ai50d
Jvuw1SGBqU+FhxucRE9J01sDsa1zX8F/7kG7AAcJQAK0fwQ0PFQ7cS8UBFJ4J7V5
W9uQc62y3AEDSphD4TtL4Of1+RhbRYWvVnEYMGoefnXdh+oM2VoQUaWMgYPwbVbn
nXgWDel7fkICUS0PM/EErjraAyAqj4GGu6GMUoVbwoa/hqGOndJxP7swRImC8PwZ
WycVTffo4pqxo6STX16SofVbi/+NpKnU2xjxAoCZRyJC0f92KdGSAwm3arl/hsW1
XOOBt4Nz0JB7e64pdScWp5M+yL3tblSySvpJnoL4/o9Op0ISUcA5ciavtCS2DEa7
cT00PLBxUcWyYYqX5dnHNGPNKvsOQJn8KgreoVy0r9mBSL2rN5jH+ikc4DXIJEu9
ld0ODEbQl+BEvvZ+d89PsBWyEQ/yR0HyE6NNM/V5vCRAQxgmiQ99Cf/6iUI5SeyC
Jz0yf0FQnC1yrS6gYsTwCwgsiIHw/BV/kwWdn1bNRAXwVGN9+o5vJE+tWTu3l12A
+fOj91rNEo6dKSoIhPAzXWLSlJ6wHxeohr586OJar2TVcn/bnuq8l6uGyi03dG0E
rvQg1z68xplMI2rNC965h4GaZCtQTwgwOMNqhfKg85af10GdsqWZa8DndLv5/+TO
bm/7N0reYMSSZz+Nk3/BYLRCMSsZUu8AtDLSBgzLLq95TTBSg0vD8tMEc+GOY07j
ByseDJ1FE9tdhg/Na1/2ED+ol7LVwn5D1Z0T6HNgFHIZqJkJhMaRASZPN0csW7b4
DTnIBGoMU1f/5oNVka6G6hEZVz3taWtCkR3QG6meJWI/beDoLR3dVJk7SkTe/j43
6QtemDvz604YzwjVXuSM1L2xvID+qk1k8o631qcOPndsWLVTtwFvuyReq2P+3sZz
vh9kC16NWCJwzP7b3qxmyNVseLUQfGERxQaNpC7Gy3GlJ2mbl3LurFWm8unK4v11
hSFz/2q1bf/nwNbJ6iqDNp+9YcOWXcm2zK/kIR62Fq5Ud9B4FjcXljqsNB+YNJla
Tdxo9rBpi7naf6C+FLP1dtb+WTCzKUyFUI7gN2nHMaFo/fg6Y99QAdrDi7knRyA+
bI+gQYdU9Mt60aQpn+3v7WE0xopKzcbROZ9izvSFPHg60fkWF12Sgi37f3JMExuB
WEPMi4N7UdYUDz1zsymlMjPju8La1FSSRI6ULDkzqPoSCbaL0AMf0DS15lncuGO+
9czeSBQCWwfOirSXHjY3KiVG4iAfcxjD3nSt10iLs1bbdi51mqeWqUss+xYKBd7/
pT9pFfmHbrRBVKI78RxQ2w6wPVRqlxtEIj7SlAYc8epPW5Mv3H+GlJT6gl5PIaje
NzaG7roffRWFq0g/XWdR/aQiHey4wfQXnIWQi/oDlJHKzreOFjSIhfXAjxMql0GF
LOvE3VdMEdVVjii7FdxPixPallR9NOmTPq7ux+0H0DzsoOrJ0UHW8UG9G92mM6au
mGHUw5TFK4gFXh/0USd5+V+0KVMBSFbC5T8zZgOK7vYWTItWaWjc9ynY13o1fsm4
/aQ54Rm8Gc37nrqTynBN4AOIe+4PjwMMLOuiSSyliCZSoJEa1ju5iqGfFMEf02XY
3WeSVN2RQL6eRyP1yqtzZOVVcsCZupjAbm6vfKWBvvrO12JRj1VaKKBEmcmpJ34B
z9Vjtj9qSaotwwHgB4SLqmex3mGekHkOHMO2RbCSjXWGyye6iwoUlgKEBLvzDoDD
OVs0lQ1agNdJj267JFIcrwduArEknXuI+HqJbzG2KW3IFmOLLmi7zW8DyxV2Q2tK
LqMdlqY03QCLteird4suKfJsJFyg5RVi8MBAEolJmm+yNIbZBXZxxLoqXJAG5h5S
OwlsZ1mGIHfXL19RC//fUJloYxDTpd8QHoau7sJJIUbUr3Vt7a6YuBq70NLNLf15
L/CbIBOal6k8e7TrJ16ghnHxT7OdThwaeEC1re/isx3xri6zR3dLGAq5TryAMYAn
mxkllgbaQ+sb+kBIsQpEYQvjmvnWciFnjnZC76K1lecmxH3STQliN0ZiJ+I26c5k
lCYgGwZox19z0Kjet/LL5DgXkZR+mb5UpkPbyqCRp0vTVDu9VgZTTQnpohdgNdZ1
uSboIrgjrQ1RVQyeKER5yGSzukZvrEEoT4cA3s0bv6SLJgfGSOoH+cYipmARv5YZ
cYChvqi/rejSQxgUZqCcP+hwoZs2XatOLc4E90ayD6xj++vrlIs2jQAWyaGw7nNO
164KNqKMyVH3DwzXL8r6GmA0iNaRHFmBLA1AlOM4dqXNjSQqqHxsQVX8W/lvxr4L
34jgAaOx6XOfpKu2GqvUmc1HC14jlE+SvhOyI5UOf63o8BkBuw1ynahkUAF2pBAC
oD/a2ynFNVemQNsuPTDZD0IGpG4GnAVaRt7W9QspGCsDwHHpcMFxsWkP15mSkyuc
4Iyaofg1hyqlCbb6DkAHU0Lgg4SQb8o6NfamHrDKibR1Btgi/pLHquiojMWrb3ef
U66G7+BDfNynKtl7fL2RkQ0Cg6QwwLPYlqWmmbQuPVPwqXxCDT2rcXxZPhu0Fti+
9zDMx7batLW3PROJM3eDjLF25aW01mDDR+0eY4UWwbnKsBZA1FKlDh0Amur7AxwZ
jk5wTcWxKKOJgVBqhdhYnZU0lX4qfcqHsBehAnEkMeOUptSDo95GiQPbO5OFNsoD
AgXmuF6NXVveZBO5clOVD50DeVH8e+mpVjiMc+HywvTWeUxd5SwvHIicWdSTfbSI
PlBkPhB6otoKck4jSEbeNPUK45ZA2GIxnSJbgWCq6RvwahhW/30DT2fGCprBejw4
6LQrCXrxMnNSpzGFM8XqWaSuKsJ7l70f4RyNJbbU1KoXP+Vm4/M0F5DOz0/tQesm
w0lAkYglwHOM3N1P5n7q3SNqvREDX7p+Uthv3CsO5eDNgG856abj0vUDbgJh/tj6
RTYXi6xYYDYcEjmpEt+GC+eCS3kXyrjg6d/cBskav298R/w/7KTuX45InDmIAtfF
8OU5ZHiEKSl1WsUyofNfEDBwYQadGUNXNQeGVFJLr9U3syGYbRSHVPK6mO5HN0wW
P99K8k329N6zQYhxCDk5tMGJ2gtexq3P0iyOWCBYFwUCfkKJyVhAxh+WE0Wjw8jF
if2A0jsoNGPrXNLOFg5CY3hJ5T8ZQRcjLLpfh79zFIUvOboqlPAHUjvmxaOgEJHx
qBGmXibukuYNtU3x2upTec6gRj0Q0eNcBxr83Ol1n1JMGOLtw/DTqocbuZBPz4ET
0U3j1ir0zjTVa+Ly1dBQuw6roZzrCDRSvQa8mUvMwJoEGWPTOMiiXsTh9mmzSF6l
wwnygbBSFu4Q3R/BPGsJSgvT29BZ3VlVy2+mMbcPFjxwJ1+UHTAnATWoXT6/r4NO
zKFokWdl/5k9mNGo79tKR8GcK66ZePbMuXkwp8W6TTgml7qjCWH5U8/yLpgmaI2N
fwxF9Vb7Ou1KnIqgIQ/fk0NSQrckOCBubF11Gul4idWruBKZp5x/LO5AUoxYoumJ
uXeOxwv7c1qaawH/ygYu1Pubc4FToqcDNS1SIisSDgt3FjQldgOyADg8jaBUjYqW
gnnu28kWg4CftgRYq8hn3SyrrRp9QamNUI0UI1C3dEK8CUl7UvXi28fdM/Mlvk7v
1/0U64Bp0BetJSlcHtYYwu4dNbSM+Q/Y58q4dhakpEed5U2uVW5Kc/drICcNPAXZ
kn7hX1RbZum3oN5BbfOKxIpIHGkK9TCVgFMsQ+X3VkSy1uajykjvH1Zw38SgtHYm
VSgHJtIgtQgRBLX3ta2zQPLRSFeJ3xKLpK+AKPn5zOv9enZA4SiA+Gd7gyX5ieNs
OHEvzuv8gMfFCsEJgWc5w/Br2cCbqkyZGeMwpIMnjKGGLU4+3Ch1r4VhUL+FdCEy
`protect END_PROTECTED