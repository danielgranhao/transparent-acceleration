-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
MRvzMwvyq2FoT6wWaPaJffSBdYkf+Ct31WFXVO+NK9tg1aTAs51JWzMmAirZpUB0g8skw3JX+rKN
tLZaJgvZjaYUGYh0Xnxr4YKzmxzd2jyntJ3rw6b6gX5/FyOGJh6enhw5f3+iWLfDWYN+5Ye/xSdt
42HL4+3jhlI8DalT6I1J8WpfZqrFumcE2TcHn68zlbiDr6IpW0qslq3p81CaGk/r7QEwmyrfCUI8
yLy6D/1VK3G2B0buyr7ReBiPd/s8P2ImKq+7BGssokpI7GmsJdU35rQGNeeGay87xonwc0gTj3Zg
6kJa1gp0Wflbak37ZdqewqWfsPiDNpm+zMUahA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10704)
`protect data_block
WP0FQg/UV1DLCw02U5ZFYAUNOrqsCpNk0aG7UDKk/oXZdA0T1ICsm6vNX3zs0E9zquB16XvPSWLp
2UpWa7lYpObUNvZnd5q3lNUHeD0P0uhSb3uMS4yxqk0iy4P4r1+n9wzT8cAm1NvS2sI2z+NZIH+Q
20ArLaIvJO1F+UjJUzYGbmKIMAKsRM8TOHNAwiQ9O8KD5xSJTm0xO+6C2cfL50Z54AYqXpxkk88M
EmYnRaf5+52gbZFHNwUER2nyfojAvHaVqjbKAI2hxoK2S+DMCo1VVA7I5Rh8gwi2hBlD11hORL/6
y0wSjzdX5pkfLhpt4m8VriCyT8lnvhB8WaGs5VIlbFK1gTEWK9BxJlSwlMkd3M+3mq6lMtbMqLZn
tc1WpUHO+dTy5Zb/yKAPN6T3WcdrIUd0WeKqTQs40XJ4zmh6NmeDWAv7ewKhYBcY7uzq12u8t+SX
iLTfoaS1HGVtfBbTjcz7aFcPAhnKA9rE73OgI98ES7L+crvTspnAcWzrv2iyUWyhb9X5J1yoV+pP
BR0G3i342N5rXizYxK4WHUpJn69DaGLY+7fIasVamfpvMu3aIAboc7ANOj+7D2xEV9Rh0p7zaGWM
JHNBGJzB+t4zAnfhZI06cU0GvP5VKTPXebcPEUMUNFCwdGbHTYmMMMtKz7zH/K0BkBX815uVQFPW
VUbOU8QuPYS05h5W5O2HLhbKckxD/57M9LHn55U38iaerWxgu5bfWlEqe0l7Y5eHLxdg3KWqshzZ
5l2KnptL/NkROJLnGteYDuRq5kOuWWv1BgZ3tAU0mkfGZRS73xwpOnJZXPbMifQjGywIK1i6e0b2
P5J0eBUxwSr6sV7C0F3QvGUf+4tq+AVoCBBTC/BQr9hHL9qE3EwTgJ5O7Wqet+7RqKLEHTmCo7au
oVTLZdrg4v3wNE/M7euphk0srzJJSV3wzSZ9yrWV/L/oBMCGbxIYMaJnXyB0uR/dpXdv+a8V0K/W
aOksEqOWo7OImqajn7ATDRqMO8nkWpA6EgqbW6dL9K1ejwPAHJv1jcuG2e6xvtZA8YzkPOh7Qvmc
eB7sIMTgVrPRcR4nT1d9IySkAVHa/dH6guThrKOO3ddUat8j0XuiJ59mGTG8qkEQUM9ADdNcKpYA
+8oeWf5nQ1AFBvdEwGlOaUuwUJx+Py4LO+/Yao/MO7VYXVo/j8Q1FIYLUnuWCuszfX/QSEL5HlOJ
s5HQ68Wjvyop/PZfbge8kS1iKCvazVn0jckJXAske5SsR3K1OAZfXX4J6lTGKU+9Sfhg1LptJ8FJ
drDguCC/lCx8vWVGiwSxfxSi1USn5xiFEmu8yNYqtUphJqKeioG3UaZzlGXBu5L14aTW6C17+nHh
YP8oKRIipdAYa6Ku9kJ6PY3Ys/R6eWTnUPKSAVRz5fxKZ8oEjyZI4f4F9FjzK7tNMMZMaOh4NkeE
F498ioMKEgbyHaf23wZqZFdhz9UgGJiiSujBNtZc71oWu/1P0luAA8GVlWoJ7oPOeFzz5jthVp/h
cJ+RSraq2gQhXQ7pW04toV98/1CpPEpS4pYEcaOxF5ckEwyy2qnKSlWjvh6tfSg7ufPde1CBLE2F
K0OilKBGCIZkJ9A7gd5eu6SjQNKzNsH2z6+r9VSyfRMJJ2Y/n2kJhvvTUGqtIXPxTD9O0QpJi37H
ar4K8r6MDE7XjyJb2gr4aU0Ka43gd+WcnrWEm5KrrLtq5cK/o7Y8ni4kWQU/PAvluIkGsp0gMeE5
8t4F8w5c+zRLis7oV5UP71HaaSRmWsCd53tJzzHyDKZVJ7BojyC12E62VAVFhaXUbG/uoqx7gpUX
bqi5HuL4DiW9MumhlXufEngtg0lloECmtV8MgF2bMNtdOKS8Kn98Yy6qFAPTF2gsaw5MLkd9BGAb
r/5q6ki1Xj9meLC80fgIcpsPzNSoBQwJvtBCY6bgHHKf8DDGAfyEcKtB6bVsGTzrPUwwcH7DkoUF
x66UBifnob9LkWZJ8EBbq8WOvNePwuNVHYw4SDgjhvylAMZCgRdknwKHazS1auQfuJpmwx2EAidt
O32kqkTPEkHKRJEGthBNueTxxODX+h46fqtqiCrgDqgsSlNAif+a/Q4EfnBBXyN0FOK19JxFQGCh
dEngEjOMGtwje2EGeFaQYMmitsPPf9VEpAm3mr2vPjsFDHgHTgtDJjWnzz5SMuA2ieunF1tCu94a
yd1lXsn/3Q4M6A8IdM5Mo8Vj1NDbxXBs/b7KIv/CPBYLuj2swTwpyX93lKFSViNY20JyBwNR84r/
JOxQvi7GTMoKWhKtcyb0exIX6u+YsQJ3ZE9S94SC460y3spfqQ+e3tgpVS9fk8K9FNFqd+YRAOg3
HXTAoVe40gQEGJcS+1U/8MRxY465Pj13XcXrsGAQr90e2wWgeAVZW5W0F9wDNndohb0AQunmgd8Y
5h319/2xQTQdREW8P6u5g0u26VnTHEFyqcFe1cAQ7MZb2y0JeYb0qKDJkHBt353xRcnl14ax1cuC
DbXiiRTUNRX4A0J3Xoh8tYg4QTEI+fABVeA4nGYBwknLH5OC25nmYapfLPiL8CZQf8D2BOcjiM9v
fwoYhAp8aA8esqhiudg/T79+CCmUU/UbyidIMhwStB6rCrGlbB5fIIoXNlKJhqoKErN++QBqo5Js
4MnmlWZhsjRowx+3G4Ix2b/VbH+249N1JO5+O7zi82fGwvF4+XRtLMz7z7a9I8ocolEz4bXHKLxE
+pQYXTNX9Poks8ulrHTur18rpk1tSB6Zc+UTDofve6L0Y8JwpxSGVVk5SvMG5w+we9jcTz5yLrgQ
rm01I1B78kBfrzkN47mQMdhvAILI2oaAlK1o8rsLTPPwcu4TYwgAPptj/NVitDbonMwOJNXUVjF3
tof1bFnaNOgGhTf91cX9ZFtb1DZ0eQbVbdO466EaU72IOSjf7pLZXcBpQGDhSe3tQRdodHWl1K/T
huCHosPdwXiDSixN0cgleyWvTrZOKjFQjv72rjlcLOpoV3Jlk4GnMiAJCsXVET2SwjvEHo5Eq9MS
dC5ATG6N6rTPPmRyFqu6nsCAAAPgtYxjAAQbk/JnWCBjNUI+r9dkXe0xWhLU/3iffm8C/RjDreQo
nycB8864DQxiJLoaRjd9ahXBCw1d5CFiLUjDVt6NoRzOwbpk7oyQ5NRqa4p1Zbj9wom780dPZb+W
czq2yWIsH5WO3YPs/14KXR6lNaV1KWIfUunGxEicZzIipKUtolqFFYUpVY/Do4OtkcDWP+XYwmok
JUqslUg7oVGBYoaCcgHQIOtIJu7TlL4K0fJZamF2CwMydULKGCzWv/doyiQFJ/uKSOkYPaZi2b5i
mx+SY2yOJduikIdVZcafEhCgfs5e7jmjhURusKdyW5T8kaPr5psyMc0mX7GMBraKcRjgL7U8V0Yw
o7CRphOFGA8zdDIL/C1mrJnIjIxdnn3m5qpTobXs7EfUD13UxdEjHfdB2KpXsaP7tX6bPWuqNGgh
ZYXMTQwy0Jk/zFOLn0ejncAwixCePAILBe4prIXIA+58vszPHsOsUDJk3AxPNZymQtTTOKJQ0Jup
fLn5O+6KOzdWQP1TU8zkpbpqDDvkGCOqE8zJ8akvKomeiOtU9cPtKRjOEzUOUlC9sXVWeh4mbLb4
XqBWhBwELZEQPfiTIp4MRBwRHztsUQvuD6MUgr9AvfjLbXwHBACTAAhao+WmcKwWdMarPclaus4R
1o5gKhjtqXfId5oFWNxV+4+uaaxmUZn+gc1bFq+WUNB+jAQLkUUSoi6xhnK4tWt2lBJPUsAutRtM
g/lHeSt5PjwdANyEj5WWo31NG2yam4bbnALOnB6PoL+WwIIFZbDzOfnKOSNfXcIKdMpcfujQnET5
Ow6tv0Q/6cJf+t5j6xcw9jGoiVvn+ZLWGe2qYcYFaDr1aDTjXCnf9aRxceFPG8INa5fkLIpxft9z
t5e31dlERBwV7E5xUDWESE/Kqg18NszyWLOI04uXXoXDKkuV6lFvjR0x3ROTwlSIYXccIuxEe7L4
zmg43Xgvj+KhsqC1dk1wXc99VTx+Gynn4KkZW/VuUa/xUu/laFDIb5OmjbB0Ng63W9Fh1svzVfV5
9sAc46ugq3YD8+Sxp5GSBLzFbCjwdTVzn+kFTgfXylXggTul2u2fNkwqonJ3RO6/htFzEeiydhH9
yDMAn93RB/zoWefMgmbZdsbSCXr6un5VGu2vmnURo3ynQWRlVSirMIryqTQgWjHN0OjQ4Usy2Dek
oULXr9NFW599KVopt8YNKncEiHs3ps9P+lmDp7J+K1V+WGyGhF8qErayT3e5GUSmUuEkY/049kD4
vgKhUteR5WMGdSxqxDlq+FvKbb0D7OTxyFVSlZolojE5DxDfLsgl64WufJk07wvJvNiZngDclHbz
oZngpfLZiT/0xF8b9vT4bEKBe/7g9VGCUejIWq6hbvprexUvvUSTbgopKtlsz/sQmBf9JLzBA0jt
xAcl0JejdlRQ1L2bwCNp6MQautjnnpD8UVZn6GNGy6KqyqPXrbDgzCHT3qyhHgjBSmeDvqkf9HgD
u9Kt44xB9b/bA4S0hsKcInx8JvpbOa/L4IXnEWj+oyToDSWwl9mST0QSwSa6Yu2bY931fhSgFhTk
tSsMAXFMKoQSCisRpJW9WmpgEW1o8FDGFFrVFZ7i5qEwk2+wy1+Yy/kyL/lY5DgWEBbsNfuzxDzK
5DtpQiC207tgHnUlxTI9heIg7a88vSalNO+zxq8/dYmEQpnBs9qleUytRWTrXFv0oBGxs0zH0nmX
AWVKYd47GqjQGebbBPebdpptfco1K2Ninujkr3hNVsT2K4A3wceWjGXeekH2PpBZMI5GDuPvBs0T
ZNUzo81VgfewAsmFx5ekXdcyJX8DhJ2vAFJVwU7baeWaPo0Sws4TYBvSAVI2jPnSTyw6QJ7/Jle6
QQt+ApVjpY/HsAC9EdXpYE/1/pcDtEUu+Y5RB67fdziP/ApnYNudyJUSrUscBn2l4MvX9aTlQYnL
UWX1TawFE+La/9m5STBiF4sr5SeGLc6q1CrkcD8De1V5vhBV/LvLwMnlnnH84hlS+7D867LUoHi3
P876XLBjMpaIs8Rkoa4tVW7fE71EGTpqjZXYJ/Mi4F0y+sc/J4P00dgRWUyE1PMIOc19JnFbhKcU
HL/tyeT2RYA71ivwr9Li4ETYIwQaBT2fRYLG7+nVI8Ch2Q6mYHqRCyM1/AEU7PLcoAk7d3Olgkvk
H6N54yb9q4BpTw/oReSgeDUpLx1hOeICecfLGmq+JEunqLKS4eGYNGXr3CNoieRADWmzhIr1WKu6
Vlfs88Ujkvh+hbvr4mKQ6FpI42KSi8Ggt8IRFLmJQm4Od+PmzTIaZ5uDMaby3K4JTwjntUzZ6Rtp
LAEMc1Wok0MNVpFBjdtr921DjYqDQPoIxxLVWjCiGUXzuMDMNyMnTorwj5RiKhQ462du7451F/lw
RQiKUxNRkecnY5SGpKGns1SNS3w97jXhF2m7B2+S5ZK+f375k/bWDoZMf8nY3BAa9vbDnylHQiKd
45C5ACbziWTrCliIq/mV4QTIEzdn0e4XXkjbfp9Fxwgf3v3MB057Zk3SrEUoVfyhiBpVsfkSumX5
imB2WA+4kC8PBrfnilK4MzGIYqqfxFeMKEzC4qUsHNAXxteLaD3moDBTO7Lfgm2OhO0yDMbYa/QB
U9iJAnIMGQwFD16DHbHI9kEjZhYpqIONBJehDfhd15zbsprxqVZWC6XELO9lVK041XzFyZmLVwSO
XRuyvMNHlbmELVjb+M3Sa08iiWxQrvDr8po7un2N7e6aCLXuN01GiLagQvQ97vohPH35QWLkCQKF
TNBMLfPUCQE8FOhQ9/LyijF3qVCcxZkFeu63xIy7d76LibLquwYPaM4JZ4wphveiR0jKnpkR89Vq
HiowkIjcKcmqusDe6OPqproD/sLIZIe0XlFYPBD49cioJxzrn60J2jBDElInZIz4VtZsY13HTiHZ
Utm6NB6aOhVJ7CJIZC91W7XuSxEi4hZJa5s4GesJJlc1QNUkVWkbehfbMlg2w5NWts+qiniWK3eh
ed45gH2VxMQgyoJxg0ydPLgbiaPtNMNu4p7r45puLIxnkJMvPr015LHwRgTBVn5F0C4bOoLOrtEf
Q6xmccVzcQnUw45NXSYCDkNhFFvX5mlN58BLKUqQdckWtr17j5OP9+Cbj3f1AV5RD1HKb/+1RWCp
CkzMvB7p5IPy1qoq9+8YMdJyu5suZEPrHmyKcB3RSWsmGw80l9fh5umEVklgK+AqltuFXyLgw0DO
4ab1noffkX2Yz8n32Qvd6PtImbL4nlbe160qXsIa54tumFSDh+seOAsCXEP9ay5WOkah5oAH2Zqq
MNf+/ia68gVUJLTZDAFmJD0Vn5EOM8FyVXKWCYqurL+MNbGVzJ07obzqz54rxRm0F2UyIrr657Qg
R/PBJ367oUI/DZgk5HOhQ5yrO5X4UObmp9WGycQOxR1BCXUIRbNbxYye1t1LLeH0sIyN43mnbg6W
CBajjgVa9BqWKNnb4LYNwHk982y0AVKFEA3nmMlddWhaD+yrMDXpwwgPzuQRlSYd98Ri0DSQc2UF
cyXustEf6dGl9isSw/89prhWYXvyZ+k5LbyXDVLicIc66Cfp5y7lBQcrkRrm7wGpxY48arzz67A+
oBqEfrR7QL5ErTRzO67Jz19/hFYu2LC6wwCb4GCOHb/+2LJYHLQdtYOkYYWoSsYaJacoLv4cKSqc
r1NgYwsMr3V1MJJPed5zi8rSAEUSjpe0Z+GLjA42PTWhZx2YvH9fe3oPYf5RSKkZkjUUUeDae9rS
7TYos8eqlC6fqWwQo5RsSOyUAQbgiHEURCcl5XAystMgup+NkAgMuuEBmXoHxZh44cYa4xrl1AJA
v1sMXRvU6aDltm3PAtJ2BOdPhEjdjsOk6RwQtO7pFMCts1os+3YNvX9bLHXax7GD4uAvYFtSXGex
1sk7AXYc77nc3ntfEoS3WQfYAf6B9c73AYPY/bSxcB4VQz25huRFbMsqHTjvJ/cKxR64DWxoeSG8
m67B08MmoRB/aOf2KGKNKbcf7n2yqf4iChmRgr1gmqDUI18NNUaM2goZxqurxMwZBDnxPxaLF0iE
2EVjcdbGo9iBk6zia6tSTsY5zZHMN8UkaD1yLR7yg1EzjYi5mMucI63o5c/QHbxMSyV4AB93KWVm
zBKY+74ACxKhRnxqqtT+CgvTcbdL9zy2fzLbC7Lszu5K2gGB4WWQFheHJhJxCC5UQDcFms5VKpFE
L2D7LCk/dQ7H0HIJqoUdkuFRzDdhfxM1kUue5eQtBaYOqOyY5u4rwWSm3uSUdhLE8HNJBuApU1cI
yIcfTytoMZdeqRX/1HyIcx4tktyX41VNON3aAXvQBFgVFH+iqagpoH/rsq0qq4pKvfoOTSdpUZ6N
XTOUECSfjvNhqLtqIkCwQk/7hmqD4qF1tg72GKm2tkMrigef27jgvcacdhnQkqy4dE/2tRTj0BfV
+Ri6bbg9rUTXIV6Vq3/mGhguNI7O5menZjEBxWr5/9zeqfVa3sh5T8+wkV/0LKbrHFyIa8h8o+9B
kuvSqyvya6Q/doACJhYtwqP33NumdO4amb0CPkSe2pmlGQP7uSTyfztndiN/yEeEuRX+9Styzer5
Y4fukGRqC9Z7fmFOnUnViSG7L1/TG1XWTXk0h1qblN0+vTCfWjodPeBH8yopB+LT6m4QyT1O5vMj
TyC5RuLwuhO/e1qxzsylTUfXh3HT+tKZrDHI2VmcJgBzzR9jEFcnqTDLqh/RWjL1f2usKg72cQzj
mUxik1PjWnJvcKkIN3+DFffDz8VSuNfdmePpN6cA/UPyzRL6Lb8iOGdRNhrFxb6MQxLamf4MXSQV
NcR1dRIR2EXNZTEiMztO8+aCEBQNkomwmk8hjLAA0w2o+BRshDP1H76NsvWH7g1JitYPHspDmcAi
JD1oO9CS6S2ZORKB/HWgz0c+63teOdGTDWdw+3FZemtz+cOits85qszi0ZB83rGVsI84pGQWWuyu
wJvM0aKPVtrELwLaSWeioI480Wn5VC19M8iRVkPtCi6MMOfEGdrbD11/mbfAdycmfquOcigXWrMG
5B0b0BolYBkQe2TwrZy5i1Bq5zJyHZY/ht6NeGt3sXNm0py7qO4nHaJ+BmCXPV4x3RmsI0v0ueqw
kmG0ytzhVDPrOajPeFQlN6KjqZgSVSOxYcIsxSSzmARKpQmLyXK5Zi12HcUw6nB54lgB3TbvO7+8
GPd8ggG2wk5wKowqEiLc/XjAl0kVIZ0/L8ky0pRIxWCyROwfDe1mQyL7Z+S6NCqDLdinTdbkN8TW
LSMuP9YOOhB3kUdlWwCjA9ewUtYX39BVusYovNSIvmONGMo4ppagBUlWO01HcP9NsWlMoy+Mz8o8
9WCpwzZ3GdLs9BNT77k9ZLroA3zE8g207j+/QydY+URAfgZhrZUhMaAB9GMSAIhqYUPE04G2UhyI
buEDUr8mCOJe9hRH7Mqk6Uyu93zxQwruqDPPBRVtCfj9FpS6vhItoXYSfGIVa6ZcYQxcWVmvghON
4BUh8wIF2Q3kSaKhVrsVCKkIZYa5syYSASQNbwkYsNHO5r2Bp3iwEzlmiZrq0YSum12yR4vcH6ts
t7jgHLBHP450e0GJBOJisoxUfrUnbH7fwHFALdX05/o0W5Rv/+mM121wlx27ZD2B6HxNep8fB/rB
WRDh6XTScaHzfFFqYOklB/363nonDZVczyXpvlr0wHRjoHyLX4n4pIewCRMmJkUHVw4sFCxKxT8k
sAsDwH0LDSooAE2I8gy7lNSbuXyR3ELaKR6jfyKbXchZk54OXFotXJ+8bTgpLs4uQ8fOQsosstwU
41kxHPytDV8XPEZ0kxbxzf10F84OuOPeQx+FoXHBxnyDCU9b9M1t8PGsNcxfxfVvrSrD0HZNbuBm
+rCF8ynFUrfd3JBJMiFJHjn2B9NRzCywds+tKLPDXIJPgSRycfJx3xU1azZQOsdin6SoYnJkd1nT
5t0Jyil54OCaY4+Z2/Rm8quefWznnTRQMGsdGYb6krdV7H4lks2t7QINpQIf6TqywbzGY8RIGlv9
Aq5RgHOMxDCme7ceL18WWaPRiSPgJ0XApptO1sesjfHoVsqibsTtRH+pozykESalqx/Ns5Q6GOCp
6u8e5OmqVyFfOpmKrokcKS7FH8ML6J5E9QT84JBJr6LaWTa1IcJWVQZUVMEFAZCT11eRrwP/NSoy
DNW6n2aLVtlv5nlxLsbuHE2FmEJ6EiBCdSUGWiKh1C/ihsDQzj+Oplz+tXO/kRL3pICC7VWhPOea
6RoOha15lnKXJNjTBbrDVarb9QPmRhwj1rD2ET+Odh1EuImGB/NxdYQOAR8/Cn/O8R1fEdsodvZh
Df7HcHRFXLtyRZwXAVgqxvCcB8mOCTeIy7akYV74PBZ/Q5iyF11k/kJP8vBbATN6PfhtaT31aNht
ZwUQDpgoTTUDQA7nF8JLU9e1dstHPNTjRdV+E7noQYE2BX3eSzVZp8qZXkeBSs/09nplDZmkIhT/
XlWIk4+qcq6ePVgfwVCm+CBGnNmFFlqA0htH5+DeFh406Wra5M7dFgoMRRqmDhFJcotoL5LKw6tz
eRkvRp7cJajmyvrysudXNMabopfzCYRrcN2KDE9qmRfvA6uUhGjMCyKpAexS7pYkcWSEKlp9TVBw
R66uWjGGphZA7k8J4TanOWGZrZU5JYWEjO8HsRpJ3FojntN5L1UG2rGcXSVbPnt0r97VXLV6KIT8
6Rc3cCBUa77pI7UYLBQPB36rXuOG12NYJoMq6DZdOzuynOrJfh+1D7vhDviL09KP4KPeo648Zdl3
qqBn/4DHaOLGEl5oSALclg7zM9iJMg62sEh4wxqlKV79Zv9PugEcTlOT85KNanXuEQPQ1hhPKrxc
zG0GlCTWKJVXoGPpsIhjUETbgyAb/16lTaX6jI7xJP91Bli2Mno2QjBpMOMEdD9szBsNJkhzg9N1
WX+rbqtP06Nv2XfUr74iXen+bl3B7A3f7oW0TgIZpXz8lh+5mW1I0iDYAF6vuVQFHsdplObQ/JW2
H2JujP5O3b5BehTImVAWevSTUtx4A9P/wbouv0uFZHCl6KR0MFRCeqA1YOOjY99fFK41ESbcok16
U3qhQnfVkfM/XmzqPNxCj0+UGsKDmE3Jzvkh+rlHYagz2floyIVv0oOAPYuYfLdKKcibEkkKN/4W
OQpDqhdySybdVxMfsRf/dz8jL4/qOJrfBNTpkkO/k7LFyilCmK0buvlBo16QIzmh9E9hXvknWkLK
JAKoQDwSneNyZBWjzsjn0w3ULUir73DGTAOvNN86vwFRcFvpHQIOlBJxbgJPR53iw+9R+VNQeERK
MNf71z/JaYBTatzGdbq6ROCzlRi+YIDrLW8mx9yEgxwGFy/MffoE2CxdHgxen8USnl101ouENN86
VauPw6ZM5fQs71CeQIrB6CEl+PWFWkWqVOzNKvgtqPv+F0L1HGEwCmGKt+ByqZiGTp2Sr1V2XW58
h2xkaehxArzDvIn+K3/Xq6cJka506qtVL5smqYNR70KkJ+26Cj+yfdavcl9tsP3BohZv+JgYcSdX
lAn6fY/fe11md3cspE1ECDgkm0s7Fo4vvIC91nx6OFWlpEPTmG6DWTo+lH0OrYKJKU1iNygMI1fx
b64H8jXmla6tZ5pii2/LCJYM26nkWjvvh7WJYhOAGtsylFNGYZhaaeB5j5Bg5qor/Ug4rbS+XJtY
+8S8Wan7HtYqKLvFeGocagAIxkq1S4g1qtr8iRm77bF//aJ/T3Jn0JDi2SpffES6+qi8w9Q6UALI
cIyxobnuZZNEfS6jDsbUJ2a/DiXZ+p84pN0esODmIA/UAnVrMU9LEMdYWox00SYQGt1D/QdWAXnM
kptdMHhKxZXIfvAKM6pAODUhrsraAZqSLX9A1h4sOE3r1wWOmHonbgS/3eAf912kfBJ2PBMzsjIt
64kZWT/yjDll3E3CLBCBfbl+w/JDc8V74+2vx+Twp4rBWHi7zPXiaU2FcvNAabuaMLw1sQVdpxSV
0oRRCfUZqLF6PHdKaA0Vuj9Xh0rJEBUs/rqywpghJg49xJrfLBe5v4ufc0wH32VZUHGHiYPhwx3v
U3zifn+IXhqt7iWFQNp7KNNQNFYPC+HWO5RY2opnWBwc1UxwWDtqNqp5+/nBhPScSfKjFaKWmsaY
p2lZB02Gc25vqvszH20PV7NINk3LQxH4kDPuuOVGBYjkrZyoSAyoH0daGPy0HChjyvVoEHZYrX1T
hsluWz7SECaJw/8UyyzJ6br+sUxmk4xLJc8qfsEIikHBLZygOkS+5JraVFtSkWOhoqdZnsvSMP9e
uJNzBm07hvkDVfrZUxgNo3oSbndDIDzZtQDVR35xHr8izngxqHHl2CHin7WzXiTS+qmgSqPb2RBe
bMmYRK03Q8J1Ebv77uiYfZIWokfNT8NlnXE07Q1mLFZtqsfH0UW4+m/n0/Tffiw2SZ8LxTVfY7oJ
6u552Q7L+18V/q2s7Cq0f+iLNdIsUB82o0c+CvoeIcSH0/nNwWFo+aj5yLdq+gJANM4452aj6BH5
okAqnDr4XXCjr49MjdcSaZRKjwXvQBBDfjHcajlAKN1CvrBvIdrX2zf4ogWNMoNjffkv6I/timCV
NWFhwQSnDeIKVjGdgkK+zOWRVRgM14IPvlY0RO3fpONtYLIlI07zuM8S8+jrA99KGz/8PVNJC4zz
fC8+pCgLODOqGUYor/Ii617nv/26E+xep8xZh8+OjpLNTRXgcJecZKzuCzbxmDJZuQu0z4wjOnzk
t9vjLIzyaJlM+y2quNzGSNkWsg7UEGIThD/Yy9Z6nWvBezI/IuVVC/2dvx8yoJr4vdxUHdDv64j9
DXM8V0S9oFDg3+fK8QT3xWBusfJK/qrll7aTU0/vdM3HiuRSq5mar0/xrcQVHcf2X6xgsXlYPY7u
aqMxzrhOjBcZ8S2mTdMrhMutzGE/mb8pHwDWVL6V20J7NDOW+QusaYtytXSh72tM85hJgSnQOeHO
CZgsvmH8QtiOqws0JBAC/w0RLOhxUziYl3g7xGl5pEnAiYrr04bxfU2CQDev63EKGvOF8ppBAH+W
XULJ/qTYTyrKdGRUgSM0PGWFUTu8RKz9qTV1omDQnOb4z8mk2LSWG9Z0A1NBuPbO2zIyHBaHinA5
z0fbimFG0UtQXg7waQSpy6rVF0io/Fj457X9c2w9dFVBOY/1SP5amSfFXo9hA7nzMMy3Ka5g55c8
hC+plO+beuL+fz7Uhpc/j6AshWK3+x61R4nRDZ42By9B/spsrezfTvLaDhoqf5WdOJmNh+j9cqsJ
3W7EDU6X3LSe13p0FH1ABaNqbbPQoBsV2FKI2L/syojLykxSpKCq+QrhHzerpO2SFgGs5URvtG5p
eG0umEDb7CunHrEawt+9y+GQaPkmH9k+IFNqtgQA7X1/O2gaTK6KhdEkUQg/wzBSB6MTG2coMaRN
TgvwcIwfVb5bJvi/OFFC2yPMWK7BlqG34Zdnq0XlvD2CaLNUBYxM+iPtD2nlzfRYuYqRuItIziYf
Snw6TUyJ/LaPoUroJvQ68C/TG5SkBcGzEqkbe9wC7ZbZDVAvqZhxY0T/d0T4CV06AmUF+YDi2sDQ
fYJB86nbdiWZOUVqsOvM5DnxE3qYOZ2UQ0dAAVuiEoz3ZvN48o3cSka6IBZ4t61evyPmE/JNnaMl
k0dtYfXlkTsgSY3SaKEfCI5TL8lATuBENQLbfE8XipLcRac4xpdhFlgZq38hJIaORKnI7OAaApHH
YHS6zdmyTd9jn7zk/iN6/AAxnLz9L//yArCi3ui+RcTtBThIjRFFDOF+4JtXovfrAE4LxtAyg3FR
BRKcqsnpBRZ31S002/5QBv+kC5D4frist7Y/Pcxkd8VJBjHYCUPgDA7a+FTfQzEDt6fC8NIKxqX0
ssg8GBQYgN8Y89w5PskM2Gn4FSzccH6u8Xfj9XeX/R9hKPRQQdngYm5QS8aCIOnVY/Uu4TZKFvbZ
CxZEBkgzUu6YU3PiqzbfT+uvDaFFjxVdpPlfsYo6/l5jZnnSf8IXiTbHkZv+OySnreqReTmzp3Al
t3ktB97+BRD8rot+vxzPKKGuUgccdI9mijv97PkqOKVlt5Xhda5bbgNY1Jue6sutEqybles2vF+T
HdfjH7+z1zpjmgtjh9TkAYKtl/ODy5pUBFvnZWvt5PGoU99apv+r0vu9NZ1nDJDx41UQYbSQMZ0Q
+bte+XpplxThkU9Htl1m5DEIDPHKEK7Z3Wra1g8Lt7zHZb6L20nT5aVPi0LsXa0fjXtb4YKl1vyE
Doq1WqrYQ19dESxu/uTRTY45yaVijhCC2oe8mrItZah2c0Ziyaim4aXi3MvDGK3k7qstXqfHM1uI
VuY+exRKKJ+X8nvcX/buFhRnrIc1fiHGrqOOX6wVhvdo3DTvJwa82BO5taURG4KHxhqS/W68wJ7M
K+MRpNVf4g/xrkGhm374O8552d14ihTp4sua2JcaGzUYgDw+RgEyV2Ae0LIH7SDNDEubN/09whVF
7MYjCRwjCAzQScCm659UN65EQlAl0xapZrPAqTRQXtkbXtnmUZobpjmvz3kcCL/Ghkkk6tyZyMKR
BO0rXrCD4yItIyT/1MtbJ+/Nhpf3JxzFDSwQLazZQaAJKgmvU5xAobROWNzQiBXIGiQNOHPeJPbd
nPVEM3v+HvMi1ffhQ5QJhwavxYPlbKDkuOMQBzOJzgFjpio773OSOxB9ltBi8w81/90wzkWvLN3T
Fyfk86LPocsZoPHWgaySlOsegFvMmuaA+gPFzuqsjZMqG5v7HewFhFZ167Z7vZ3mswcsXAHljiWZ
ZsQJbpYPl/Pv4nYIDKj5lWgVtNREYpoNLFaTa+VWBgOhAKTA6ZPTmuGgZExFa1PQceS/9KSri/Br
dFmNOcf4GQ/EJnkSWdxH0rScNgci79Q94zkpukQhXQuYieVDrKeeAaGl3xvRIyvt3MKRDtChDtFB
uljzZjdMZgd4VuUPkTx2yZJRYncu09ENOd1Nl9h1b73L6sm1vr/ZpHexA3GURnB31SsKk0JMPXRO
A5qGlcYnpqN954Ev21AD6p2RQqJHnqW+b565Uw7cCrxm1vs/E67DibBaSyKQTEc6iPDC0qMuA0jl
1vipDPIbJBGftqs79syJnQJAFvLqF1j3Ce/4NyQPvZnYYjjvg/yCkyhkb1r3
`protect end_protected
