-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
wDT9vrRp4qGBf8ZdTGEPFVT+4JAJLsCvr4IsgsU6gKn6V8RldiYzTTQ8uVuaBGDrYGVAqFFAUfeW
5A3LgtBlcVlBFTlZYwQOhysPW129l1tjGcQWQjAe1K8sRjNDbK6EgYO6wzHhq6sih2oIpYiRxPGz
0J2bVK+Vm7FDhK1To2DBUpeHsTDKG7Qpy1a2Ehiij4wko05RvzBzYeal4MQzYWkNS0UoQGMly+F0
RoqwU92YULAUjHGfhSJchqpmxe3AfPXJgSzA5xvIkEZnjFp+RDo6o03VGUYLT8YsLL39KuEWsb01
F4WEgJareKQ7lQknvueRVFbjmI3jZ+CEI7NQSg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 7584)
`protect data_block
P1/+Lcw5hPNgAJVKX9Nmp5+/Rez3IBPkPpseIOE3jDPxk2BO/rCrIdpz18KwXIlz7m5H9kjWMV3B
1guK6cJLnB5w674wI3IBLy4WUn7YkyySoNF5pcsPPKLb9RlspO1hPBwXMUR+ycqYgVEEHCqjd8b0
iFSoX+DdVY1J2+a/3vH9qwYaxO4UvZDfycJiZc7s5575ymmFGt1lvicVP3ajZ+UV/CfNRrzsyW1f
Az5Jw+c3PV9wyK3lA/UlGfFyU1sCeyMPpPGBCE0d6Rsf2kALy3D9eUOPFeCW6Dx988tiTCKHrGnU
m9DqT/2zollpZ+j/hCnjXQGLVe6fFZYqalWeZ52eThDjXsBxqj9QOEYHq0mFCJaJ+095L53OGTgA
Z40e2Xod4d6eNG0zv56kT46pPTym20YSecRcRhixHBKm5iMTgt/h6kvTDWH538ujSTjjA8QvIREC
nS39LSxGgGzH0UvsQzgHXN2nx2iJ5lqHPX8j5qBKERXDXqM+DrUZKnXxcOIGPdOO8GTn1aB75y6u
9J5BIZO7Bvp8YoSZjWywf9bpd7tPgvWsHg/Q90Vt2QqrJ6SElUXXpEACbKB2VWdN1AHV9x0B62aN
/6AqFEXf6B59NlHbbgXIXmpZ4JH0CAP3SzelVwr2V106Uwp0Pa+GU32m1NVU7NBQ+Ip9/8hfGP4t
OD2WjoEgE5qH7g8AHF7rP7naG441PtA70gFMbrhqNAbBwTsMXSwb0jx+2mfyBw9H0kueQDXCLo9G
tAdikp/AEi+TOWtFZ1InUxB2oeKJ0/KFID+G0hWOoHvNorLvyUe4Pg/RFFpLkV/roYn/CNr4DwM/
Ju4wAnlf0vK36tMO6/KaHPclTk0eOwKBBD239/sX4BBTqvJf//j7/MwgcWdiocOlCORMKMqIiQfY
h8iauIQFF+ZOSl8oIjJjx7RKml9MWk0+JqSA50ekq/W9gnWLBGmVFz4cGi3IufI5i62y4LzjIKHC
ZPJ+EETWjcI6jvIgE/7nl9q1KVbatbC4cQAO9OVwvp1AuZSFJIsPWA+9lJa8QDF4f4z5qiK25xXR
w/qd39Q1FRYtFfTuHslOn0e84lNPmz6KE2ceCjqUskZuGajw/VYs1AabAzPwi0+tr7/BEOp4IlKR
0XPehannJ615oxSpPqC/+IcYHY1DpaLnMC+AI1gFCVwjiGg9+geD/+Ox+l+uIJdC97WT0qpxb1D6
HIjDc7BnE59NSKncL6VWEvc5la0jS5B6+SeslVLWahBw3IzkihvjS7MynB+ON5bXX+EpxIitO+ty
QvElEJNLlyibsRZfCTo1bk/QaVIPAwECBxHTB+LolY2QhLsabm7qV3yE8rM9iQquYpbcgulF61l+
ziNkYbzz+YCk0vdVu1pDDEhRZ9RnlJddPLM79ZKLeoYyuCWfaRMhelY4SSJicXJy/YLyJ8v3ic26
uIIaFFsRFJzEaxjJApGHwGiIG4V/UApF94GBQ2zIiUbtz4OzxkkqGtABATl+D0Aud9hyRxhaSpVo
HBu9WmnOY9ZQvlaWrLzblUdno9uCQyTAGiX926h47kLaL2g2Zq/ZA6JbHIt0q8eKt5ilKmHeRn3L
TXavubDpIETLHWjAx8xzVWp3wy2f4vehUKyEe6+VQmJTuRzwmhCpFPu8Plgwi98X25tjCzvNRa6n
VjAKeDqE+1Y2odvAe5ICj31qpTOwjeFwmUVZT7zoKMN3PStAn8gq56lVdV6Lemjbeudy4EQV+THB
WvdzRn/eiouxyq4j6jGwoVryynPpjB28epRFfmvknwh0VUYXUO3eHsUVQvW5sLShrjJlTJo3l3Kk
PWSSCamJPU+F6ijWHyE/SWiRo+gy1XWSruzZK7lfVqCjZgMc8l4QMEOMlcAhcJlptrwQIbQZxASO
CiVVQWXE/NRTDFWS4KG67AUwcmlMkngzIEFkFInpy4WJ2+tIN1J24gsk/fTM49T//lyG1XjdlLqF
26vuSl5n/jRYbEtYuooEX4/iXqjsJU0eRVnRJwSYT+CJ+QbZDyKdNH/Y0a1FYcZtpIEcnPjw+aWC
QH21gc3FGefkPXEbIZ88ImwryXqp28E05IswEjPA+DB1begFhKecExtGpdbdx3ls/kuD2lRzwIrM
9g9I3jwUJslzd0lWblroUmMaNHFUsvQdc6065Q2QEAycDfzLEctCWcJdq6/IkO7VEillqhclDo5M
wCEasfGkukfVkvy3KcDaSC2N5oRT3fCB1vHvffb2+wr2y2Bf32HZ9zj7507kxQlEgEEZuNZfq0tY
sZxGRQHrmegQAirMwG8X8omEugSH2ppcmrBZ7p0aa6YqHdwXS1seusIh+O2RlrCQ4ejdVdkTZ6LK
dcxIx349oRwZbmD66KRPqx8fZJWc7XjNvlojqaKPB4+Oltf1NVZjnNuJePCgzaNUafFhI/slNaRe
/8b89BSHh22qQIx5SabqG8gvOIr1IDoM12ilvyjVmwwnQXcYHGH/4XJHllAg78JVCLIqsTo+du//
r1wfXoUE4tVmQIkXDYS/5wfcDYBbW8ZUF163aqAm3Ihg4dCGb6QbeWkFqtwo4VaH8gxKP8LPc1zL
E2gza70KhHRI1UxedEGm2demaQQ34KphVJ2TCJfa5AOitqmCSnnS6yNGy4ueTULezv/sDLeKUBpn
nx3C+f+Dpk97sf4G1U5i3rHifc/Q42I9uUGXFXxddB57YW4zcFG8yJZfr76SfWp3svaDWvdhbHz1
voI3yK/mt7FflZs59ziQeuuhi2WlP6My+Usnz1k9rT7cTKhyCiG+qfNpBDW8ftfpavHo1cgJMeIK
ABDCuejvgK5Nhpg5yVMdJ65fwnjZMg4QdfjfIj8loOAWD1fSgBTLIr6FuiAjA/pyRGpLkkorW6vy
qU3Kw19o3MwJlL/XrSbYsTb86OmEebqn9gFZaXNygmdaVnW9EpDnRI2WFPj7qgkraDedHbQvl/e6
d+1yEnDilNw8kf9d15yM0evLSNGBqPTyeFwGKEkcDz6dCfz/ftF/khqv60Y5yKiBLqX1XnmmzM0M
ZfI0c0X0JgFKHcyAfYpLg9TLZuL0Lywbe602ULaay8XqT3nluKzQeMzrMQZNqcL9D3YB3gPaH9xY
NOrT7kIo/9YE9Ur09MTlG/GrGxGxdmxjxbe3H75Q0nyHDRyXLV5DE0+2CP4Mvhvm9mPjU1ylRLEA
md8s4eBv5VZ+6Kbf1lZKJ0HFsphBQKtqpQtX6DWPZlDV1xizD9XgedzjMKFQCprQqR4mTIm4Kjba
BwM8u0ZTlAmzPkLEtVlEfEPJyLHXSn7PuG/DDjCWk/edemWf60UD0EHUbrIyWD+vOx7GgmTAjnZz
HqifdB+jv0Aqf34lyyMC3SpuwVEJcYG01GEHfNQUrH17F8BKN+V2bQUSMwUZO27lA3AC0SumDk5o
fzo4DiDzzala6QhfZVHPYHH9wPvwb6tOxPbSLv89pT/pi7SvvMn5cwOjxlCIQ8AzydCiPc4UslUe
LU2fEhsfdtHoeg9XIg6r89Sh9Z7KBVU0u8NYgHFkT91DqyHxhyVFT7IIezSE2ujGTGIEx7ipIYot
aeC9HwpYvepB7Ld2048wRbKhMsYjtKBYybPPRNtb0nelHFaSpJ8jmDU5BsV/j+FMGgQlJ2MpeeT6
EAMsHMFYNbCkiz/v3kWO00G84/11pfC7BQwMvWgHKa5txvaMMWNorRTCtyExmfoPV0u7A9W/wqEF
MP5+pGd6qwYL2haQOcOOXUuT9cY+0UyRdWfGTCcgRjAGV8j9CSzu5dh6tR28W2bjHkR6zFy1ap9l
y5RimmTmzwHguLGtDzX8obCv28WXSzLVh58EPRahun9Kl6gjHqYvwvSg88KWT03xnNVPppFfnWEE
8ReNI9qLRuGknw10QFjJSB1uG1YL43JjWCi8k8E+MADqckmWBdah+rX+7JNrFrJ8INLeDMTPZvX7
4yTQzdrMfnlZiqzu+A/KaHwf8U6feCcwjN/pzmREKOxLH/7aVMuMcQyxbeaJgoGfY6W7Pxt05YYN
QN9uDJMtlNdDDsnHXC97luLIf2fN6t7x4XxXNuqBYmUqdQZPKumRenEB4U6Tb5pNOTwnTAXvO/+v
FyTUONcsKAHNPHuAIz9N0u+AUTbJiqlbYjBpJzH0vw9wbQSpiVcfPRywq4azXtZNVXzc81yoXqsa
ppS63MSIa/ItI4pKkN5vLeVwQPzcJnzOrxvfciS0CwACksFl6v6L9WQljNwr/Lv1iGBXO9DOsFFK
MxLiU3EOYivuFY/ov6OhJubs7gqud0hmaWiur802zLj49C2ymbCUpbY5t7bBuA+UuRPKwl9V/v2/
e3a/iQr8BIE6MjxGH8WVw4DcHTtlqvRbskRUsFnGUDf3il3EVqNQmj38Wyp9ri/G567ld+dgcqYF
eMgTf6w9KcFOILBbKRJt1bKbkmPBf5b5vrbChiWNyBuJ9kxviGqktqlYO92Br9xH/l7oPfDjhPd5
JaQ8eMVVpt7bOrJT1TkUFahNUNZ6umW5Tnc+O7R4jdN1PtZ18HqnNJca5pGgcmyjU6nKEfK+x3nc
5duYuJjrGxLMzjKw+MkguklBlRRhnuGdNfFQIDyFAiQEIEnO8eZJMRvHYSgbWiU+CM6czy+BdzWh
Nakj0MTkB2A9ueKdJNjCgVTrhJU1c5jm2uNnjqc1SEkneYNE2olknBwd49MdAgumARekFXEJyeix
0OcU0Yh+QRfO/NyrzCGiO/4NflKB7A5QK/QxAUwQzPofZ568lZcg7OLo6NW7BdGG68agrQtkTCW4
Wfy89XBIYyejpKZi68dxio1DMSCnu6YLlmrNeWPBXCeNO58Sv/YGRSwAXSXQJZrPJsYucXW0Nx3c
aTyPuanI/1ZxS9h1RmrScuJ9EoRoy4p4G8Nxew4t9c7OCDiM+3eQLW59+fLk4j7y5FLWhWcERfZn
1b4XuLBM63deUobE7Ygpqs5pzoM/6G5HukF1DG+sacVDGN0A0JjfQQ6EyGfELtolxt4dcYL/ymYl
t3mp4Du5u0jkMNRBbAex5vsRk1YhliQVmzJ/gWC7+5asSvEbaE4WsdlB4gKWvM48482Twzwd8ZSg
Ktxbu7Iw4cSCMkIrGo3Pr7lpfbktL8oB+07FRFKXb8WIIX3/RJtp21evs9cPrGTzz3PZALABBNiQ
c8HuToPeQiXAqawzqE8Ydo381bip1X3KNnfCiu9zR1r+QS0cs0tfqICs4lExbQO5FD0Z7ZXH2ljY
hCXTz4UKZDh3iEvd2pCc79BqxPSi9VmQPxvJCcdq6aWH5X/EvKANABELTMLM0axDuR7ReW+xdl93
Smmwe27Oh5PDhj61WJnCjoGd1hLkP7uq5kFyE7Q4ONRL+pXjVc502Fm3uvu0fiSoI4IpzRX+6hSp
CbedOO5o3RT3cjVKwFCScwpUTEp4GAh67uGlyLjKF16V7LuQo6/GNhaLUDaZqrrEOWGI0Oy7UVGQ
252DGyTHRRyqIy4ywyy6jQ6komLQONIntvugDpJJ1rb7HDcb4R5aWkUO1ViklyhjvhSL25HVAi1R
cOLNTaqOVMXppLJpg2C9qx8ByiUp8ZgSw/AzN2lca6fH8O9tspXEoWrsMyFMf2muMGPdxMrkq9t+
viEKz1bGPSRINpqgmAx1s4sWXVS117yzIHNGdr9+UuEDqp4jgoHqgn+uQy6NpfwTX1WiWolMgVH6
ENebxsgR9xCpqLey5WuxCXd0ntU5aKNEqBXUj4xnZnuGb6l0c8/TDAL8s5LOBwkA+3DYJnwfkMfg
Rr66WX/buVNlTqs4/bBWpZhIUEfrYHMfXDNWQal1zLhvzO91LTlcrvkuBBMU0xzpl/ZX/dV1+N3E
a7Nl6jQ7f6ONUJUTwcx/3Pnpz7KXbCe4T/gQelG0UtnUJwDwzqyzZ1MfrojCMrvwsfV24dJ5Cp7+
jjLtpJ0U67ae4qx28VOtLaAAyArzSr7Yv0wWqI5eQ3ltCWMQOVpsSNWWHUEX8b+204SkKsapDL9E
tBOM1Ol1rJBSevBKBXiebVY5rnJ9bHZ0vWqrTTbRLHU2EadtYh5bDHkCRz+dmw2IWJxjj8pzMa1+
U/DjMeMioybZQd1cvLQ2IDRTPcTdAt+L3qk781pTjZmgDbwSc5gl+F4TqE+u9Ikvc3uspI7ncs29
nEXAEMu+/qpGuZyESc+d6582GbYhrkxtyXeeIMrfMrWnmIZSjuobBPMz3W2RAeyRyBs48q1WCWan
Ptw9wUWVpvAz3Tn4NwycBNYtad+7qbKPytG5y+vXDneJvjJmky0WA0ovNVOtMwh8GJ8NrTOA/q/g
TjdkcCwepJo0eM324UyPl6dCndRKMrt4SEvSnB6gHKLWeLujyNIxo1QcEFf7AiTvOxcM7k+LYclk
Ytoa27Albprl+961Rj0sAx4rSAroFlGnF5BII7CTWZsOSZUc+W1E8j+8aUgE9DaGWcdv5Av2TssQ
U6VNGPjrUJ2fyslsOqgUfsnjZ044Cde2WhZXEXJ8xjYyOieb98uwvT/7iinTqzYTsxpR+9IEXjhR
GgkNKxGEfuyTPlBp5cXA/8VAtONIQbLnfl3OiTEH4Y5knOseFyvGAKGx0cKc4kMvwRcnsAFXIcq3
MbLDDQxDla7zJJp6exlMn9hQFetReafdOrICeuaeXzQcyo4ecWLzf2ofnlCpPq2my5qdNcG/eRBq
KO6tqrg5L3q6TH87mbkdtgFl3Bcp1+t9fFs5Op7TLJq86iUeeJR1tvKcFaxJeZMqr6WZXRH+DvyJ
IsoiBuYUqkM0km+IaVWA9w6ZyOjSCP+eN8JbF6eKbyJdm9NrMeWaOX6fndOjN8GRDo8KI/5kGFwT
fYtbk4+ysDxTXHk2orskjcs9I4TRxLd9tB9skHn8rGQ22qzVu+S2YVQrY/XIxUDIyiAbHhxwVO6z
eDs9dQOVd8Uuxk7jb4MpF0mJtQWZDdwGQMj0m306CKzAlU4Z0v1BcxYS0fu8dtoDdy4PWz9MG1bV
fZYiVUluPAAk09OcYJUfOVai2JQd/omys6HeLn59/6+Jt6ytcDE9zE4HNMQx6T0lW03WJFyLjic2
eTeyRS7Miar+yek2wUMrnF0t3XLPBgJN1qfkcSHOF3EJ4eHTcRCxnWe6gCtRSNT31LsCVelKpaBO
oIbckAsFKXvGYvcF1kI18sX7T8Rr52TRSMcm0QnYuIrN4JMraam5AiXD4YBwZ8h5StOx3dgmsCCz
h79K6VdT7RIxAV/7zde9tmIi6PAbWKtFhgx5O794+Ye+vXSo4LuXiEg5UJzoJPYd/jkAZucv7nC7
HvT7MocDLJfd9EjD0X0l8dB0MQtfS4s1xSYVc4h669AiaIBvh/HMVcyYhJG4zX6u1QjI8xEHZISN
ubSW/wzIztyRsPoIZ2dDHXgqZNZNHKTMIQiI05rr7eMVkdDuk1CMo2aJV45iGuTYSkcrK2P/TQvl
cgKQNsXLHjqopgPQG544D1a+s9FZQo3AlaPa2gdiHFIMOn3yo0gX10QnjyyQkC0bMwlpMY8/tY2S
b5Kw8y/iSRwDQnzAVBAs2HODDTv5Tce0GN9eo00KE34GSQ+aDM1TQ+wSOfzcieNa7b+s9ogghp93
HKK/rrFCV0A3agx5yY+/ovOciLZ06RLejQacbqyunozS0omeYZlxgvLY2/WMwdPsssHkL9zsepTk
duVqq1zHOoGNbMeCYE0rvAHnQ/wBLS84RpXRfVyzWSo8nqq2ozZitbx88WRDnOI8YN1nOquDt1O6
gRfJtw45HHnS/Eoc34/vwF6LmlmdFk8/OvALrJkhAsgcHvE3eNf7rhpjB6iq7Ez8rO4R4hGX1ITv
6VCTKaSV6uszLqUwhdtbd9pEJtVfhFmLtV2kAORfg+sITcMasUgfe+ZZ/F7eRGVh3wYytUnz2NWE
hfMXT6wi9en+dvKXZCBiovSDH1HYh61N/xk1mrjopT4AcJhLJKcCMbaCQIUT0QBVidOygudJuFVG
7ASs9Z3G4qwG7ugcDa9PBxdPycNeSIoyLAyT5FKiyhu2goesSRxOK65EgiA61BA/0FXOGgtHlywH
b8GkOraYS2b4VHZSgGlUjqgKG0FHhxgTn6KRrQAaiyH80YZcY/fFh2PZZChCTothmZmGVYaEFS2B
KiJZYf1ks/sHCLZw27hGd1QazIl4bnZZUWBHFnpghJ/mkPIH3gtviYBWwhxcpxZg2B+LSTuulyqz
O4phCvidowdurrYGOLfAGcF0Olr2mkTQxa+GOwb9Z9RslKt01MoImRtQFNjmNw54hTZcp13MZPZM
bgIPPL7jjqS6iiJAQZKOy1ojZm4eJqYdJ4WbNWIYA6s7qW8EA5Q5gyjfBW+jmTudpxGQx3VbySmG
TXxAzx0mwaTG6YHcJXbVR4z/aAuzXYGYC6TL14x6qHAGlCaubHzQ2QezsE4/EAohtjzk12rAkf16
FRBRuD2p6ax/CR59i5jihZYTtKCrWaQdGVNUJrWYbmt2Lp7fdIUhAQ5x6Vsd2Dz63ZbSsTM6xiSR
mF1XA418eP+33gqV0de27cPL0s0pCAkWJ6q/Ih6nIzfepcQE65Ik61xpq8UmDh4kplkcxKr/2FPz
Q0ibJcM7W2Q7mJP8NVYUhUeStTbvOcNZwjU0LMjGWKwDrQr1mkgfFrli+sF1Wgoi6qo3Lc6U4nN+
zfxA4jNpTTx0UrGs3/LWVhVCYU//fxZ+vGn45DysLKFxIZmKQg3vihjbTTyKhYaZWz9Jo8K3HxYG
Bi1RdVyB+AiKg+q0ksjMS4YaTTYw8JOtnQMcdU1tGBbK0gCSe+bMSORV2gP7To6wrj2Qa7nRVhAC
upDeek2DyvanCfoDP8YDKfVk0sTutfvyQOWoH1OBsA4BWOkK0nzUm9YTG++3CIYc7OyJzWIo91Km
yFRQHPS8RJMujXEy8NHRCES10v0ZG9aJIbrdnymY6aQ2HRaH+lJALad5Wh+uXj0yWfl6+wGhRmQP
lGbQOXLbk3qua0k7KD4YMdXCU//R+HKV4OJNx2uiW8zYAiic+EzbTRlR+UjisgIY9NjrpaNMeDf8
pqq4l4yGC8TwjQaN5Vq5IjLggPnCvPUaxRxAAkP+6NfMbRfOKDeF2Lx0+XLFqvopR0+Xww9GpIRH
/kTgsm7pSkSJP1uEsHuzN2t/u1cP/wuohqkZ7NQQOwe2PTAS2poLZKWPWBRGHFrJFSKVGLHT1erk
nSN53a1tCG5X9eSiJoGhox/PzEcerQuSlCJCRUVDbWOGaLrkrZk/3d333bWVYU4JN6TfKbDW5e5U
2D+Zvxx/RsBi/jyfkrKR6pokYAPYY97/sEocxGFuHaXCNT1WgRHPUtqB3BWCDDgoBCBMaiPEf0CR
r16kDvD4dLhXSAaPWDWbcLjqfyS5i2fnmPuxMeGFIwJVF8KbdvrgcgCBoozxsHFXx1IoQIMjF4pA
8wcO5WMdfSIfSUlQkhz36JZUhZWlQ7Q7gecbRlP2GBvLEzvCs94IxThsLZtGOBo1fYd+a6YQy7Rx
igcP4tP/1VntDdFWNcXK0xexntza6RA/1Xv5TTMA4WDKGKzwJ5MkqbXwNUWJGP2yiGqzeVTyxat7
NEU4u77Nzdu6133Z7P4OrsJ5pEb26HIzbGUx/TFthKwsYubiAJQaeNcNB/+RkXB8ZN+M58iY4KJn
09frMwzglhCLRa2bMtH63tfVzNQh0wYKMTWYAljIGa/rK4705Hd8Z5PpUDkjJ5uBz9wWPBoOEYw+
f7sjBSBuVtya7H4xxl/ZXjmJp3xA7Eh/TVATVkSL1Jo60roQ2lfHY/kU3UM9Ib3QXDoqGotzdhf2
OE8mdFxxVPVuWLd75PtM1D6vUoxNIx0ZTVryLHMoYpvsJA+/u83srdMzH0jwwBYKJkXNsOHuSTjg
UJ+Mw8e0SYsHNl5s9Uo1DTgkoYQV68b1Ru1x6KmRiIJfBscmfyZhv1sdG400FDwjpJELIqCMSQbG
Mj3I44g99HmIs2qLME2zCLbMnI2HeWoIxnNCoNJADDI6JjHy5Fdsi/z9TmpFf6f4+bSAiK2EqAFT
Fzv6LWDfGGzXbHZjMA7DBEV6R1sSXKOau2ingsiNzdwWkpIJFDMgshU3U0tyxz20CqB66K9CxBlu
XBwN
`protect end_protected
