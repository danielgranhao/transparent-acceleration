-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
IFPmznfcBNMHpkQmn7gzHEbetcyK2Inr2vlwbeNCx10IfhMeSp5uzzJIfFzPPqKC
66c9s7qSMKZOT9QZrUr7TcL3JeTPv6nbNCxxJjoeRVQ8QnEqk8aE9WDAcasQ8+nq
k5ueJx0qYJQDP6S0lpvrcvZHb/pwkk2L77l/8GeVpiM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 29975)

`protect DATA_BLOCK
aRWmeTt5iqYH4F6Ei+OYY1pNpUt1wAz+uD8NUlZaETkYLcsaVASf2gdV7wORHSLV
zr+dXMAWpQGfANUw34L5y8NKkJx8znPGolZ1lCju2u2G42NtwDG7dRorN3OF4fGl
QoBDJER4nO3yIfujqFWX+3nWr9howKnOnRmrYropOpO+OO2MmgnOGZ3ff2OJLir1
/oJDqOLMBCVX9ljZ0ujFvqwflfE11FBAYrWabsvbeRZc0LtvsCdwZdd5HIUCitz7
wbsE4jlWVlsmV3bRnLZcPWRh726w8J9qUyBtgtirt8deNoyn5Oh8w8g76y7RDo/3
/mXMH9ibJAdGvU4V00GGfCmqAFE/tBOv8YRraSMATnGvJHnk72J9Ey4s9+UM3w8C
EoFrnfBTGfRM0e7tm4XzrddIkSRbWBFJsrTadZV9xqzwn81jzf2uEMcZiws2qvFJ
GVXSbYAZMi2Hm8Zv+5mAOiliOKGArF/P1ha0ezz/X1/vO03OCSfblzcpjxCZMmcy
nwJoMjLVngOygT6DnrWyPKmWKSKPUYfZYxiD0RtM1QNp+UdyTYGNbFyYB29I+lRW
1bYWgGL9wPBtHsTebVE+Cb2VIoDj8Y9T+pw/EpjLxDhIsmNUcm5fTPLWstdgVIwh
7jd0hxAP8wpc1wtyTcqvfmlqDFvMjK6Tux9QJXz9pK02deax16pici8q1XPM/AqZ
gFd8dR+232xZgNEWrvX+JyLRvkilLnfRuiH8Ii1x/2EkRLEQbneiUqTOa9NOAnM8
r8SWMPxk5qiZfmAp05g5bm9Ny/OFTOoqljGcWSTljWw6IJtZh9TkWL6TBe3zqIhh
uvz+APBd0O4dnLsMqdtvTbKKeKkTZElyabu0gCXI5u0x/UCfvNiU1wTQiW/z4Zce
kamCuoQVSPHoDV42f77AroCZNchkYEFOhVoCVENZesw/Ec1a3lZecEZnAOwNvhfY
/o6Sue9vABAKvnzLdy8xveqhTwa+zx1fd0kC2maOiTd2+eO1Jt0fLhQ5OoIH55lH
KsKQvpQEpO5YTFnqfs41sgLm5hZvu9z/GhHVqeYHALoMpfsp1zksYpXYnhJ8Ka/t
n8Y0Hd8m5iRM2yDFHpU4sXsrd+yLE6Tyaug2PUoTkWeGH3ywIEyMK8bnzzwR+A4x
vocVu5w9RtMbLwSOtCjGtlZ2awlOf3pRH/7PutaUBsTV9ty/WQi4tVZdgNRBeqpt
5SIwGQaInCLqjKwrKmnbmdpZgumBjy4cHk4ucMY9tA+L3BUzqI3zwqgi7tmNHfpu
49bkogfMFseWPHAQ7c87DCBi8XNLnGTS2nyi4I+wan0x6LMHSO6+9pj+aKLGc+LA
POow8H5Q1Lf6Vf8niYmly91bFwk7GRilF+vPKUw83Z04lhuYN5p1fv7c/CP+zNvw
racROx3dxcwjaIarWcReIc1ayUTCO1sKO9xmersNxXlB+pGGa/k4LuflMU7O+z3P
TNTc+K0GhrwXxrMHpszlTJ90BeotDc7f/5VLnGnCsALTe02tG3NBayCwgOcxmqHZ
KfHbmRAdXulXqxMaR5Ejo41mgB02d7BmILm41rwSH2tJtHUkYKtiriWrUcLmVWqu
MfP84MYDw3rKP5xXHSEsi7O5KKCXHQjph8c53Vwyf82d/pJEYfDKaHZy+Q7n7OwP
jZdPbedG9PldpX+0d7+i4QG/pkOZ1BrSgX+7D1MEP9d6OT+8m0jB2TH/mgVFKMw6
976B18JeGPQtZZSH5HdIqJ5HTA1xdgAqtdWtDO8ZUNG7i+ZpJ9Z76V3985yfkB3r
hgCMRPQZASp/ktV6vJE6wpiCoPVujdEUrKOX3DiiLYs4/PehCyL8CFygBQ5ZSXYn
lRJ0vgT2kR7yi66UY6rjOpGz4G6sa8zWYm/gUcih2l6q4c3+CEeSHn1rJvYMTj0I
UiPg9EvyyelTGI22j6lJYz60cB12UyP7fA8kGfwRQ53YqYvSw/EulnB33Y9aJIzt
5ieQc1RJ1lNYiwD/5hodq2k923JlfUd7vPYZhMldcq6JynjpLWcDVpWpR6dAQS0e
uMmBqB/Z3vnIgKezn8XIKKB0Bq0T9ZLAgCITMpbPrkfqk0J1xEKuHsgQqiyjmpwP
Pt7s6EPJq6lWUxzGQyCv/xpcch6n2NkrH4g5lURq5ehfpVqaBis7cmYQXfAA6jwB
3bwhGH6acHsxYQ+KTtGCxvyEZ07mP12gqETI6yYsRl1NJ06k1ZboL6LJ7xWi7ALt
sWJzl5PbOe5c/fbWEVJ7l4c6z3emBTVkxYbmvXqFdr/BNer4rk107h4KP18eF3Oq
GwYOGtiiKLmHfLbrLMPScOQGGmJWTsSfbitZoOLHq+Y1O5hh6YSvF0ehXVH4xiFP
TQ5lEfXQg7H0xTEPgZNVz9fcPMtwnbr1hl+2aeg7y+0b9/jS1iAABNxNc4XN8KDW
0hYZblbeQaKHhpIAw0SbXAMQHtcvnjGXbXzi79K8BcLEJYJ6OgzijEk/deSs8fPk
rFMZSycGnz1SR3zrH71P+8H89/TqI+nS7xILmEPuGgl1qZZF3AiDQUoUeZR2RAwd
k/phtuH7Of9tYR4ubYYzmKxKxkTqePC3w02MiIR8UJPHFuHYiqH+DYy+0KsKgMtu
vZNdbsLXjjp5FEwBiEN6oEbbTKdlimsd7xSR6tj2ryGfA0+iSXxfCWjwYCo7ULCp
nl9CVZM2/bVP3sp/1HRdJb0N6TYLxZAoXnomLdCiWbNlYw72fI7DxluxJ+XpkomZ
Hsgq8rQb5wlw+hZ6+/inc1MUC6m8HhI7qFSZrxzciteQ5P5OVdrsUjOJWfqy/Mim
rrngriyCpE2ggNuIsUVuV/wx8AHSJ1WUb+RfSl1u29GZstOH3bMw/qX9iGjK8BoW
/1JI/qNi57C+6ibyXk5nI6ZyIVMOSmYEzYKwRGWXOGFg9RzQ6c52M9oNyUH8Ga9K
yYFqFo8oc06SB2DXulvUdZtLsFBtTkjA0jgcAXTadiU1bWR8xdNk0ZDVwWze0/LW
WKZ8wXmykLG3fbc0ANoNmOmDBTeWRsRXe1CyIDgaBr7eu/jK4g7fH+5fyTSA3nIM
O4ougVr/FbVjSDjemHt3+CqLb73cUaHbOjhK6fUD9DBkG5xdIZoR8DjMTivyx+hg
adw3vZOdYquitNjgo3JLQhkrpTl0Iy7ULFQ9Wj5UryAjqjMxlSAS6050KiFMf+92
SN3TkrWeaGMjk/DFuIBifzqSVckdOrRZr6jzt40TtI6L0w5Spj8ahqaFpVmaZNZq
AqagJYoLXMPU1csKBvo+OWVPgY9Yp9yBzwJZPZ1v+ZQXH0n1rLMM5oZ0XC57GWD5
DEqjTikp+h3+0+7jKfQSxDXijSfXAIN4dw7xime0Rc5a9pf4j5rlm4t4gI0WfY3X
SoAXl5Kh6d+Jq21zbjklj9oQzcC6qnMxFga11+KDnR0bKMI21c2RgR7/eOCOF3XA
DHMh5dYr3fufWnfebWqb6SFH9LIK1BC4lz25BK/s8PG2eqIFtHS/F9NKWbIDWeyW
0G7sGvmPz1mhzzhomIefMnG8eLj/3MXGOfKQnIR4qzaRjpuZ7ZO73onHhn0FiRBc
eiUuozndWfM+ttgYEDz+plcFzFROI1XLGT+bhzzsNEXkRTmslm4eKmfuwn+u6te/
Xe87lapA6h9nlTpBXakvAr5fwhpTlt/lzTo7F5owWOU8QhLg0/Zy8k2X+BwYqqVS
6tWcnalnvLu6oVZUIgQhYu/dVR+i45Z2g/QosFLgJWkPoZugvMg+5JMeZGc0gRNR
xtXr5LmCWKScJpQI5nrIy+pe+ZkMFs4ngCUzUJnbBVNF3dkC/2TCvgtnfURmsgJg
d9BVK31y5xubLipFudx+sR7Aai/oJMZCacNrXTRMrTLo6SnG14sDGKPjkqKJmR0e
EyEv8BelNkvW67XhiBfrFNm6tGxmkgl4/EUktnpaoYAgRe2conaDZAkjjcn5mfrq
G97Ic6g65vfBDstwHbG/vGsAFKqfPZi2pxWNDgtUkF+Jg+CfNeENxQ0Swzkw/+e8
krploGfXxd8XiE9ULXp8SfRhgFhoPPDzapw3I4Tv9kn95wUTROagUcNL63rg1sUM
zky2P1QW4dluwjs04ry2MxwKtQjUtEqC738tsiMVDls3V27Ps4PA0KwSNziWIL6d
QzutYpe53xwX03pGum9cUqpZsUJipGYCVWHLsFlXbi3uSjL0JgV07O7czB/U3fSh
+BxQXOprzm3mRbVqBhm8QEaK4th93paL4z8Zxt19f6tQFl7MvzyPAVYLqUwoLMCY
Ejzf7NIkV9lEybA6dR0xtW/UtFsKI2Gj+O7TZ/FnYru6VbG/+tbL96BidbBB/vah
+rglGXuwG3aCblVLcWaSH86m2LfR2MGhpsX73KElYMmC+x6n6dfezAPQB74ociRP
vrALpYz2GIlHSFzE96yIT9RKY5LKjmms6h/D31OTWjF2901bhNZtmDXAcwtpCyCS
PZuJ1VNckSVcpE9uos+rVnpY0LicGczbDFb4mzngmRu2xIyRUQbQJBsv/+lhRcyA
/1bHSckzQvT5MJXtaSnDBBqfSIiFT/fQlfge4NDHn0u1EuJ6fZJrq341zLZvtdla
mQvaxdN13GOQBnPPuFoZYxfLDhhdmiPEtx4zdv/L8oVGolyVw+uh3TKyqWe25q/c
ASqk4WX4waY4Id5BipOCYrCpkJlVzShOyb42+VPtU0DdDlFlOLc8b8dvG2Bjg/FQ
phX2SMzDWcTABBr47RkzItg0FFw6jcBkNGAPM5QRxBMe1tnpE4Lw4ML5MsCJtRdC
6xdK8h7M47F1YweIY1GUAcNIgHPE/LtTENHz+2iMC6/DGui7Pkz/a2aSjE3t8nca
NPuNtpjboAdzaOayII9p0qylNdFIDT5AF9L/pto/Gi3EKYlMdQ2Lpzc0E68RDLym
oeQRFFnCb32mHa8YDkOloah9N1Pes0/Fg+V70XoolEbGuIXY+kIbIel4B9EKgs95
Gjx0FI9nLNl8wLaiaFclwlpCPLqnOMq0Fo+/U6lzMaVlGcgfrhA/3ZN5TZkyyCdm
pnApGoM9G/z6VdgGIRKKaj6om7nsyZkh9z3u22j0ATk+CzBmhxW4jos98VuIYOBV
JlnnvE9h7ovrlfeW2EmczoI5EQwt+N60ewwSXB4T1Wb/41fNfztBMZBjM9b13JoS
zYkCgeVKoe3lcaYaMSAUn6f1nJVqTTwn/tuJMMg371C4WGik05Jjn69eqGCAigy3
GABjqvR131+NBQXxmlHnzJO7MfZmkZBH/loqgodEzfpQfyGyNhfNxHnFBEBJu4ZJ
rWXXOFIHqXv41dhSNuCysxixF/YHt7KznvPyFfFG/EcB4nJSLu3YhkQH0fHQasJ4
EkrKr9z9qhY59ACy1mxmfj6h3dCgK8BMA256INs1kILSmtPDcjXW6a2bekSC5SEe
fLhAKPgPSu18i5XtTfp5HoblHq3f78ubR+XKuVqWPNK/GkuLK1fvo9TokrNIABmY
larKLut/wkfdRgfjMtUQ/2bHRY4tVLYLClGnGqLxKPLuMbAI0A+x+4UFWKZiC1ho
N2T4JJhqqXLqorHx4m2DlmuGgtaODiMB/Rb79au6fIVmfheTMH4EWrRKMnvziNHM
5IrtTy6vZXjqazIkVYozAmwUiX3ibmUoV/VbFhqI74Oj6z+o2/0rJykWmd3tDpzX
M8QROYz7IMisVT6g9QBFyMMu+i86b7tsGOU3uEFjcFnKYBHl6R2WUflV8n42sXke
LTJqflJyd1rw4TM/xSwKwwq/xj6PGXivq8ltLesGGs/RFur3ItPwbDEiZKEIx7Zq
PN+aQjU4dSMBpMYkHVzFzf4YG0IztKKDepOy3qO82zn1+CfRXuz+5i5e/jPx9G44
K4WtNcUUwYmHbCTJnNrriaRD986x+FTi44Yw1R9DdKmsBBwPBQ2JcCmWAV+RjkQ2
BgN1zXFjS11NKSpZAzD3pk2Wr6KgIU9prFQ2oI86L4fe5BWBUbHyi7qxvdxHVLc2
aXpMcG8TmeYGqSiYlqCWXAUBzJZ3r4N3DCNMe8OKlFS3/Qw53GnJWcV9AxDd21si
I171sar7vN8cLXu6LdtLLICTPomx/7ZLSBYatxCtp9iCq/4uqR4JfgYZuA1kWO10
XlqD4gbdHZUfcuhkKhua/8zcxG3C12/64ZfcEEvBN2Gsma45cu7S+LDdy1Yp9Ddx
OXR4QI0hQyFCYrkzeufqvDFw+9GgzVIwEFWeJ4UQsY8qqyIFAVFoeTGKj4nCUjSa
m0KmJl7d8C8pY7eiXs1bAkAbXSA6oYBvLsrZOruX5lOFOnlEm8sz4kweugl2M2Bu
8JcugpEEHAUHtS0k+A8Pk1b6NqyiD4SDTdMOD3gj01ngEY+IkGPq6kXe0fc5ggHe
dpN5X8KKMHe/ZRxpzqQBFIcR1X9dH2oimCBxpH/mVIHKnuZG3yBPFIc1+trF7pmO
T5t1MYGaqcGPY0wLrLp4pce55u0k193xtjoMIYxiF/mMMu2ZRYBwG7RJK7PLNOj3
qRmxh/TZTKxhXXZ7lEo4IXkMZDyYtuWRUv6liKxk+rpBXZhFhjPHLfPxNMkFvXxK
K0UYRdXtjmjglJ1dSghuKl+ktb+SMV9Kxr2KQ7FSaVzR1ZZIfYVUG7WE8Zj+uy6u
WfZvtDCVdEsHufkkz5m3z73PPVV+xGbUgDEim1AlTrzBR0sb18HOKPOtDpJruSJR
FSZ4dOJe2vD3TLN7SGQZxRfrC30Dm+JlpV4ejM7sSxZue3gBk8f2ceHgtTJbP6BB
paOLtm9uzAsKpoaUzKTsVlCpA2a5BxWTxd9Q8whN+IGLAjrkBa6a7hRC75434ClT
F7fNNNTF91GyCLr3phy6RzP59ZQLEFRlzTRDYhoBP2iYkZJVrqwMS1eRcPDOFATB
GZxYbFWV4DhdWr7hg8QO62vEkQI/xBuwb+YJL9VllDzS2WHeGHAhy9/VlQS9dp9l
1jR+6jnnZ1VidbvoVsbsyEM9oCJpEKn6RvIJvBg6exvjhH1vUVqLlyfRFrK89aeB
ghNl0+p6JsUNSbdCmUoEqjThiPXK253zk/M5JIxQlUxZtiIaUT5B+I8xmwl3U+rT
Z8S7oUgJ6dfdCZ2Bx6VZKdLX6pJGG8IhmLPVvilhobANBVJlUnSj9ihYpRci4/cm
wrYvLj+2rqeX1cQsLuBl4tnBvXrCSKhNzbmop3oUamLLaOvrqOFg3sIx78onLf9M
fL7EtPFEsrZoThnDiMmsXGOaimI3EYbIUVDvRsDq6JHWT7qtggk/V5Rj+NU8PBwH
5S8ds+O3WF/gsXT78+y06Buqsg9b2SBeUYfjIKNUzNEyKpMjaC+KoExJQYTKpsXP
dupgY3myk/d7/kJzidNbnPeWiaaQyEhrAJaVmHUvWJirogBTV6iXFlsZ5bvp86ZP
bnFQ6HDDNF5hKFILoq4AjNJOj2uTkbBa5+DETb7Y2Wu29WjLai4GHuSWHj8Ap+BV
ZcpBLomADH5qh+mRs6bxFYTqdT+D42gdUSsSCcROo6RappM0GXUldK8SKxjxvaYu
ro1VpJ59dax4CjPRdctnMxNj48SMcCG8Ll9s63pouSn5wDxKg04pA1s35pWAB8Gx
+wKdKh9DkNjeZI3WT8L9NxOhxLIjVFf72c4kWqSQNcrxpFa1tI166ymH+rfLF+s/
Qvtm1v01XEt7BNWJLmNbjq1uv2jYl8o+iygEzUl4BdH3fUk9urPvxVbT6cucS9OY
Wx34sCnLaulziZkq82OxD5jP9NYEi6GCOFL8XvfZbcCYZZ37XO++IvZmXdNXSu9E
Q8rjhjGNWBqGDxli+eeJrO1lJ6o1eJvOVYP4XlImFazzKzUUR/xIOAWvY3FniX49
yECsGGlqE6hvtQuXXmAyt+/zNtJXp7P68gvrezI4lc57m0C4aDcCpAH/TYhhzFoj
hdxcAmem26cHU31We1sf/jwNTtn9mfSZmNyQpi/CA8xqjD1Gd+NpiVG6mnzppAKO
Xfg0G8ibNF5ozSJeK8JbyRy5Oxczl8Wfa0llxtY1cCGLZU4kwQqNqNmJcPCFimni
Bdecz87DYOQ+km86LGnnRfZfnfjOCwsEfL+J6zzN1qzOJCHDtQD11h2s5Qxfplez
wPKimLWsuuA3lsY2XTecxAiEM3/v55k7HcSt+jnXLFXTnI08Q8b2HK++yR1cUnFl
0nOBbawfHObLTDkq7uDnmEq7i+iXGcJQuL2VSebnwMFhHpZ7NQOohbv8d5jsvB3o
g/41MqxIMo1riJQlOYSXmmOSGHnwPF+EniujrP0Suwc6j0uLWK6iV0IWZI5Bh7rJ
y3/C7qxpgsR+4HftjyElo/zqwTbNmFhKv2a3um1ED/aPqB149FOn/XHF1VMbOi7t
dkfCF/WQ/ARJP/KRFPW4CJEj2RKix95f0V2OVp0mFe70BdPLDNkBaexu6sKDaZdM
dYxRQF1jEU197u4oc0jqhII8UfA2m7nFnLxUPIGlfy2630gHfaizEfsGMyfrPBys
9L7FgH/PiepnOfWhnz84tjRb8fBsXiYm0DH+LqgcJEfbGHy6AITBJXhXvsw83Jr9
mBBGQ6xYodqqLibsjLMxqeMf9to6X4qIpQxobtPrlI7OuLxZo15RChRF0EcZyos9
JYDZQnmalFsrT0EJlchNtd5y47RViTpbEvULR3XfUuoLo2UJgAYFKrOGdK3gknUI
NcNt0wvec2QGdk9Gnc1xVV1ot3nCm+toQHmJeiQ/kki0/AEo4ftIKeAkMNkBqN7F
F/JdIM/42fIFG9hDmhRSrwQeUldZTRYnFrNQBG5p115FeVchawMQDZEqcN0na7Qi
QN1Zzu95NHNWPzW80o5gsLuAVsKJ8Lysbx4U3CWgPn0n6VWM4qTmG5C//sg5pkox
vxcgxMFh7xR6o315SYG6XRT0i+FxMAAwVqXDgG+esk4MYHCpikm3DfqEo9ZHsosd
YOJt5DQD6Wy3pu+lVlu9zsMIBOmyWMgA1DzS+N2bu0iRakxCfsmNBS2rWDYPGjuQ
I9lP8mNVsYG1ZBNT1OTdjBQ0TMqkQgINK3NkrJkszEggVzBqFeVDtgI2wxTIS5yM
lFxx9szAaTMPCodlJhyA9Pe6cbn+dZd6zWA0TwWC9bkfoME9KBB3t0O+78hHCRyH
L0DOEa44zcRe+XiAhP5sUHul6OudJQEDD2D8szZL1w7jI+MfzSC5NP/83bJ63Z8j
Bg/LRYTgF2WEjCNmt+/VJ9p0mLHEb5iupipBErYa+a/mDPvYvlzfO3v1flK08elN
RiV0qPdLNWFdkRUjDnjgycrZEatwjiwTnoGeK56pv9iI7BuwnBNwYGhOOr1nBaoq
f7T9HZ5B1tvSZZh/fH4h4Qo2p9b101NmDzV/fMxXFNm76o61A11rU6sj/UdYkphO
xU7/Xrnyt5xwSsty6QrAfnBmxvescHcu/rx2iINnJwzLbEWmLr4T94f7UnNyG0nc
VhQHllKOz2gBQZMm39RCORNYficWKfkiXbWl246EixeRo+t9v6DDMD093T6MH5f1
VfZ7M6zlwAydNdd8jpxa3EhcIt31O0R0bajBn1wpC7nv/nOwIMJ5y+ACqs6jW5bp
U8uojIQhB6iDusslVvinqMObWwuuaRnJ6bK3sAKl/uoYJQVcoYzCVngNreGtum2A
2N5TW/f9p1GxUGqACCGO81rY1uYMSaSdPCN75qt0Y9itfUOCkS7JDN+eVThrRkCG
R2/3CphiiOyeOuoo0s0q7j60/6cO334Ar1cWHUpl92yJhcnVu0cI0l5DN72s9rNn
rG++zJpcvi52gW82iEiyMgNTCxowZTzOB12awgTMGODNKVqWvD9ZqDBETixcdxiv
NqAmGth8TlEY5MSBiTx2UmhyEJZQdK64BXPvxFW90ASAS4Dgpbe0FBLJjZjm6biu
wsFHtew64D+Eh11E/0o+ugZmgTElx8Y2PSmrpDiQ6Bvz4JWFezTFW9IFXUEHviXx
ttUg3Xz0yoHlUey+aeIADb4u+tCrBL81vs01BA09JxK+3wW3twfM/nN6MlqZ4NOd
SouOVuljHJe0gV74J0pwJT4xsxZbbWd9yqWHTV5s7tFHf0Lu57Mt3xHnh7dL4WZm
poONj/84yPgzKYlrOT6skKVjUEC9pBPSc4KN4OifJC0+Bb0W/YkXW7/voymTvA32
1rm2p8S1pvQVdDxumV66Tz54NKJqz30guA7XlXDH1j2tKjlYeuo4Qu/C0yY8IQ+5
sHDZK9DJRdx3INrcCrHCF1rv/2ap1upv0vNQv23TrxhSYL2/Raalz7+lqjbNEuel
BOtlc9s45GYt6V6JM0vCsOxxkejpVMPSx3g2EyPbvoMaGHs/kgWks3zADkjfOYoQ
6enxQ2BdZy67X3nBDnwpqfGjBKjo3xbbSRZocKnM/VKGKfUbkhpthfug0IdxL3DW
Ame3mOAAZOiBh50Ew/Rca6/0Y6X+yN6GWR55aZbBl1WaSXL//XA2CbCQvVnbljQ7
cP8YLGqSiuNfZEx0tWGhZVv9ARLx8Y9DZ7ZcN8tN/libb+YXL9hriT9D6eD9V5vr
AxSiA3Uuo/ApyBuBjI+TeVBf+wje0v3FgbbmCZL+eO78w2L9Vl1TgCX8ATqUwJP7
C81h1K2F4e7rrcIBct+SUeXd4tMSeSq74VUhl8XrJ/KopUOk0kSuXasdOOUF6a3t
ihZ4onc6H1w6/JFRpuG2tuWKuKAW2W9xvdhp6D+ky+sEM8WfOfVmsaI8RH/ko8Mu
EwX24ePkQ1kkiKyZDjLHnN5unDzY34uxKmK4ls/OR/VOjeWOfmM26ilqd/RnwtVH
/jp0Ngde6CuWI0sLqyYXpXPLxnEWobBzr/oqJTg/adxv8Pnd8y+Xv4joP1fb8Sa1
mp3LN9tU1jEmPD042+V3YUeEVP6z8GTJpWANkR5KcMlxsclDIH3PDjR3ThSMoe/V
IuhuL52H3nhHeeuenRySBZB3iw8z33zSS3OefXqDa2Xy2w5KS9I/cUiZg1eWHcLd
UeP6KARYDWVjVPKjgEnN8AGOL0U/FrftZtbuxXeQYSgtA/Hm+iCqO79A8NDq2ztL
vJLbwXuuYVxikCY9ZZOYx2AUOWunThTxH4qQSsbwGrC6IlKh72zURl2PE8W1CXqm
EgmdwUgZx2B1IJz5KtoREpDYtygEDzZyf+QeTzlIYB1kkPhvVIA19yQlAcsVGZUX
KOFMGDeMkkbaYay4JiCI6stJO2eX1tnC9ZpIPIYuOoh24L8XI4+62NGOS/NfmuzH
pVQkTTI9+6YRJVxz2AMbxn3jJ4SNYjm6hYpUwAsn/Qof9z0XlnFExs32Hg79jDeT
sm2tEbvytJBlrHsWCaM2CKV+DqrTtBTAjaLYeq0TYqiZIkyXp2wOcEzwfyvueZmJ
+2BUB3e2S8CO1wVwdHK4ir4v7HoR864xNKTNj+pGUeFyx2o5rV0NKjlOyQbZchI+
KqKdU+0jZzH4X/H5MY4hrEVz0ZHu6E3K+5382v2X7D2FoUKq2bA+3z/VPbAIjEx+
layhJQmZBNenEeTwEYwxSmAIQtso+L+hcyOjdgkwTXJUm8r1w2sYhoQ8nPZh5i3w
nTPIfpQgsncx4WBaZgfeWKK7ctmwsw+LeUEZ/EvMVT5YVHPbgrJHzaFCc3wQZcLJ
wO09Ssl9ujcFkG7mfA/FeSFOLTCHY+EjApGl9RvBrKNa7WD83u1HWbRRba9aKsGn
OEDj4mlsk8DI+f7kjnVSuz5TCDd/vi0gab5qQQsWbBLDXYlwrwGMfADaSphBxE0F
QTOFcV7jWOvES48Rr+mcSfO7Gjq6XJ3WVD1Q5WNfG7aDbUUcqYjQxhHx5Dy5nd/V
wrZnqxe6pRSJiJqMYb2ZxKx4M2jv6pjZUoedT3Yp39j/Pm0ILyU+qgKOKSVg4waR
DHdmVVlGt8p+SsZMzLZkUkHO8z6XLiAjrMr73i9do2mkpoOkJvu3lge15xLqnFkL
t7notR6Kt519I/g2EspOP/kptWEjhfzqz61pLOyN+cXiq/vCUx+O9H+VAD6tTfz/
Uaf5vpZqt1HFFPzY5wZ/hwKHu7xocuI2zHz9T5GcyYjob+NKNC7kbomGRYYsQJgJ
f7USRcah+uytDgZ0Mh961CAEdHPwz5odnVYvqMvlmOZqvXOilpQ/tVMXiqsDM2jf
M6OqdAJPZ1TSRzV0rJoaXfSQEeFCs/V6hgd/X8MbePSG90n6CqhTPQpyWty5m/zI
YU7t+mxFhTs5XRRLaUdz+i3a6W1EMVPDKCUyqIMOp/BwBiJjMbspKHRyHqkEqrlS
mnUtufzLJ+kpvAdv4VVD7VTTYUhDUJZZrS8KfO+bci0LSDTC0Lf7Fr04QlhaIb//
vI4gFn0JmB8GSMRBjFHYnD+WlOOIR3Qpc5HtNv405dDc7PFWuc0Pwzup7DNnpKUD
rvinmyofYccnmfDDT6YCNbQK9vSuvuSAv5WTGgz+vxoHuEyoLIa6uIkw/FlqGPIK
RKIDLBa3+saYKSe6+FQrk+Sy49sEuRURvjrsjWVNvHsgBGt840ejTeqEpXH0iuB2
LnvmMiB/VPfhewq0VfULgRRVkdaQ2BqA/xGxCVsJ/7s1jXFkMZ4SytR0mRBIMa8U
KQT1QS3EEvpF62p6O6eCi3y4CvtXx49svUhkL1ObeYqY9As5dUxHKPWAFPxJ+qVM
xwigTPIWQapFjB3lFtTN9+1C1N6rkMbyzTYaL8q1K+37ASWmgFAhF3/MI266bQnf
8AgyhVAkBE5dknaeJhX5FyCmcjYfAbDaK8vWASucCiE4DGOOzBWmKsS/r2qPsPiY
EjhCUgyL+esLDE2TpM0y3FW7yPJFjVpuCwDJ5PeuVBU8gqpImTSe1akDZqeL2Ydd
KRlIPswQMhWLa/QnUSX2oGguv+LpVFalrZQ4BwObSt2KlT+AQEjaFrvlu9Wen3Ct
bSXxK/pHjO/BPGiy34TqM1b+ncpXuLtG2x5oPyT4LsUEV7wy6DY/5XFbxPlmX7yh
qwUD40iE/9SP7M5Apg8HEoxJJD0b0+bcxHgS3+FcbugiBys7s0SZkRpI5AR3/t2l
n08W4nVmtLbU4iTc05lL4W1OANyO2FpZ3/ifSY7sic6JcyMIDBJfi4QNq3WXs/ie
zsiZVtkLgeJjHFOEEzco4I6UTMXwppim6orLnM8bPFug4HxvN+mk1gewBeaSYM5b
UyDhVB7SJEa6lSF/ikQ/BtRV/8VjCwY+bAMCNYNa0SgRKLI02nQ/tVmTHfQVzN8f
d2qs8tebYe+xxd2vOqk6rq84kcMGW/Cid/fBmgVgY6PDJzd+mhH6j6T1Skk9I2dI
32bPIhbNJdtwCC+GoQxdOGcOjis8dvIjgpvjbwEusTUlkf0vKYHMIxSdmt78HwNm
b/4ShAUHrlNv9jCHjo2eu46F0DZFAuNut4bzombr25uyXU1BC+pvZJw5+5oGjuPO
faqLmLBUAX0UiBsWfNxo3LvABMrNDjxZUlR6kOBrWwUghHpbMDvIExWRxsgwRoZN
A5ksxyTja8B5u9YnrULxQs0uDi47qSrOcSNv8RBfHb4xPURVVFfmqW7R7CZptoZ1
YAxZbU5/5iegu4MjNAfYEu5OUP0aj11b2QLf6gtzZHZT9HyLDqD8YBD1LsoxTlyN
OYva7y0bna/EADNTCOIz/VwvJ2uAWrPMu3npmZQAfxGoKqigfXA/0SkSol9hKDMV
mA82fahwjS4Ve+zGeWUTx+D64/TGACWRT4ivzI/HkPpTk7nFRZrErTOP8oLyUygt
/AS1bAVJaZEzrK1GvMS3+r4uU5sKkYBB/Cc/9N9JlKA6B3Ofpfta6vXK/ISXAeFd
Nugv8qFyVSah/vWo6xJG2LryL4mIM8VLj808j5G7gHK8X5uHaZwwejV2CWc0VK35
SysIbVLm2sKmTs6re4AO1BT9rb6pUHChdVYNjWGomg2SV3HbWcd8OmtKGwUJ4o/o
E63IpAtG3LkbEg60L3CRmfRedai8HxXEQFYf+cpEfxzq4qTmUBFPcpumJdJdCQ80
uwyNODPT59H5mdOI0kv9+MIlfZ2hjPYFMEPfRInddetvDgJss0T13WUqvyJN0uI/
o0u9BL32o/52dYfOiz/fB4uNBnEibDMsnD/3+kFG6M7bhWcpFUkJfizwRC5lEwI8
I38vdZVxuJZmZeHft2LKfDeMFRoL1j+oQGv022Kk/3YywyJ3I0qJnjIJ9z6Majad
xggYnDZiLF9HPmrSIzt+k4b65hh695pF+S+ys4AM7AdWLxTB+zW1CLJ3MFIFdwfu
BZLdr/QaAce2j4DiRZ+iq8gBKKwepQFzfbG00ZblwTFqREkESq+Ge6PfzDTzAtVM
t44bKPCEQyqOrT3xBKOI72fSvXZxqt2LI6HzDXZI5JMbx/WjqXW5e1h6ozL1tnWX
efzEtDK3Qu2q1re3HegMnD4aKCFx6hToyEnjZqZVtJPSj6IqgsZ5k4f+6KdbB7Rt
0/32WtRekwJm3/oQnVArIB2wbVfS1ruqvDPq0DjS5+mNN6Z1jRj2bZ9wSvZVToLV
LzgoBk4p7Vi4kMnV9iy2vJ/iKFrz+Ug3h2uNsLjcqdJkruZPLI2vz5UHuTiHAX1A
jwt4RjSpNErMfWjtu9NvymowMw+rVI7I8aBdMlQqQ2g8IuqNJcsPMq/InpEacT7s
c6iS4Dr32/qSzrRQgprHpf3AEzxTlrDwnigaynVpHxN1pHOKIsJaJL7l0hX5ngOE
CSnG7Y+wVfCUTK8dSjYu1P+gvfTxXzTx4yca1OOgrDBWzpfZJcKoLgxIbzR0rzY9
grJiFbbV2oH7BFyTlTf2V80Xqr7S8ilMKqxIbtQOj2OSHVos0HzVI6u5DbVmdQeQ
GGDebYYKeGsCqzrJUBkYvAJiS64YFW/UgHCJog2M6/F4FJu2Q/3ESzTZr/opDFUm
fL4IDBDQDoE/NIy193fphMn6496razAsiSP4CZegAbGmMrdmS7xBWuKzEPHmAW3P
zOvW/8RQFBAhkkzyUWqvWZe4Bnegf/RRo3/Jf8jxpHodhiezqLB4enQK3Om5Z5+B
qfmx7UgeEzFFlAqbrxx57kY+v2s3w/ZRi4WzlUEnbcMrcat+WDI8nsEX/p8ECvKl
7icZRAKtJLrTznjvpXxwJylaNj+51VAECVy7C9hg8xFeAGQ7k5Wxq33Yrj4DOxJZ
zgYaFw2WcS7sEJDiDhmLoZigL2EUFS4iFI4hSBly93WgCYMwvucgmSwkHrQawstw
zNKZezWPvnKdjDKBt2dNlPcCglrTepIqoeaTjEzsKKkLh1cOqm2EFPomHD75STGG
kUbTx9hBi6ug1Vg8x9PdmzXZIvs9DdEIFUW24FzX+AbUHDmbFG5MftySZVqzK+Bo
M50SpSsd6WEya3z3lzQd+8WngNEeRzgC9hd3dM7YDnE2vKq2RYI6nDpe3bRpL1MY
Gt3EY6gf4+ZKhiQ1dNfwB+sEu1dMHIYrYdYPFN/nbcmKHAO2o38rbyd0/A+Zz3mP
4Ox3Dbi6nBUPI0GnxIjGdS9z+6GLr7cHfC02/PByYIZYS3TU31RAyOe+Z95vFqir
XlzCSDjZmNM4n94FX/28I+toR4BxvK3MvdV3U4b3Ime6+6Xh3FgSZWS1UzXertym
ojFkj9pEZ+z6xnLkXDvvasTMkj5K3GgVRD8hN2HiC9nVFryaI/vpqU+uvhAD/R/r
KUaTagug606Abr19FdTYFD3HuW3QVvoEXTY4+sV2Kzfs5vAyEZx8A2+7iPKI2A3r
QS5nyoP5hHweIDvWrzzdK5tkzzMoC4FQI+U2lrXEquulugrh8kcMHZpXHhz837vn
ctlCxNnwoZeCTn2dfOYguwA+xbu8ncXbkxSp3aljcwK88ZNRemNKG6fyq8mj6zii
rAJVjYDXoanNfijbI8SY4XBX3JTQULZpO9wEYPzdzUe2ruIXzG6VzgbAKzOGdir7
L3C+LYLpH9Stvp6iFHs/R+onYtJfZW8gXFJlpG0s43OkeN/r9tynjHwkqp+jz9QG
HwouvlCOfeTp37gprkjJo9Zsap19worVa+OkQT4sdQH2US3A6b+JsyD7B31HSAqM
tNl0wOvNRflpz7COyPcDPREqYsMdgf1850OU6uHio8UPL7bpFGl2JPj9r+Xw40de
gHQwgzDL9QXBnkZUnbOFyF/KkucTUpbSb2ChuR5hSC6wgZ000J5ECFLw90CK/Cbk
mOBRQGH4fH1cwk3QB1qtiw9xfU9nxBeQwyz96erCXLw4ecohI3LrlS3FDyp9ztyx
/BjwZkqQMO8jm5fx0k+W6s1fiWM9h+p7LVv39PzZZhtv1jbhprDH6BaF57U142GE
96llyLxfzezPULlUD7de790/fHP/QmR470Z50lhenNeYgwTg4fZAsky+fOOZAS1s
jpSAdufPigLGNqesY1S0jpahNmKw1yTAkSwEXO78mnF2Yw032aY38k9voOl0e++c
qyfSBwMaCl5oUw2W2t6UZlKmSBEWypLQN5tytyBZ9psfl72o2/dOOv8zNJ5nGZi6
43uOHCOQ1kGehEmnlZ13/x7v2wvQxjR0ggSaFpEs1PM8OFd7me6h+u4t3HbS76w2
egS7acb5EuSWEuj/s6s3W0yps/xr9DBJ/8aVJyBAfdBe3VnuNG/DGQjP59iQeqci
BIqCruWIifnz9qPT5whNCQxvBcueCZmSWUwWvr+3QYnRxQAKkhWoab5FqbDsiPDm
m1z8t3tU5TPwRvfS2w+xV2vJTt86NhWKB93uX/W0RFnxp6DvRYtCUrCL08grbiEQ
ES9Kqden40xMCSnuKWtENbxFz8hbsZoJ9+/9LQK33oLlBFLzi3EqHEwh/xYMDnBa
Z/KypFHwkv7FlqX+8O8nDFNZApQejUp0F+tsYTqSP4AFdm6gB9h6dOXHf6OCK3Or
yu/xY1d62jMr8iglGEkNbPMt7h8+bT1lSX6DZi8Fh+AGUKodeKOi3/BMAePHDjAy
+Re/RPNCi9F1KSoZoIc+BwjmZEPGllsNcdrYDxf8jxdiSQvujMZlveVt8DZh6f3S
Gh8fAMv++8wAph3ViNI+4viaV8gw1mmrtvonoIPy30J6okYMyf5IJh/ZHzTzLYy6
RPvWIddI/xeVtuMpeCcu8sgJN6o0W33sm8P1/luEJucCRm5Lk0SRYW118z4MoikT
hv2ULR/HyVL8cgKU3qPKDU2TZd6eEJjZF9M03aS9ObZUvbuNvYcd/nz/jErKGRBD
qxTuC2Hht5umTRayVWS2tekSsft2fK0kIhtatvl0y9srCYoDasZTkmsS2r6Ddwq0
pjIi96UnR27dVg3UL1kDN9pAjppyeA8hp86gZ7Mel6ZKs5UV12er5rvByrue50FF
StdVeLR1l7/SA+C5UJ1+ZurIMMSmywKNEw8g4mG5+wjuLiUh91TcTpsXr1JDbdi5
AR8Sx/Pjvxog4XQonroRYF3uxD8WejibXD5viQ472WY8BDqG7gJWu8dZZq7G0tMS
NkC+E43QfU/7Yn7+WYzmHPTUMEerhnKXS67pRIGSNYqQGRTryDhf/AH/O9kQ6bnV
wBM+PL4fZE3knHc8cb48uBem8cwqNt3sw13w+9DWXGFb0Wwyjc47MR0Gd2F32RS/
ikiWJriOxMfzdVnl27n4WW/SFy9xNo1IbLrz7mymrHpfBgXo5isDUV5GK6oMcumv
XeQJkG+5chvaBa7q3VWuBDkf/2pvabM/0xxzOcpwE9Ke3QfLgBJh+BUEFcBuDNjS
WoN+YKygXVniFA/R1L4uIdH+XK8I02NpQ4A1/TuZZf2CT5kKp5B7D5laCHzGPDt+
DJsWoz0ABkA5tRta6HFAWUVMN5/8crLV4oTJ8DKVTCve2EfvhyvS5s1UtZlWQNuJ
NJMJWEmnsCvG8IRuiyC6ep6jLxwMCHWE+LMBZW1ZMB8VluvMo1ALKUV8JPLRP74D
sihOg64IeGgpkTeuT3ynmggvIAoTU29/ptG8mlq1n0STk+l/siC6Omg68uq+Dui1
MilGXYbKGuzM/pahaQJFni7FSUChQbvkxgYhh3wfVny/2cpK4aVcogVkyQCAf7TD
7Nbd2ptmut1WwmX8pWOFFWfv/82vZhhZ9F1aUgH5Lt5sqghInDJBxS0MSQDUt6cQ
ahqvoXSHaXqfow1Q/mDqYEg0n5Rs8mDCbHL/nIuLeKDb3JTKwHB+Zm0fJ83AuLEJ
WA9cBwqExuVwBtIBocr35Bx+OD6ASpFQBT/8Azn8YBHRzh6zRL0YJvbemqn29quS
Gc/WeKR9O1ULyuumy5Qwwz5SdCq0ntSuogvKcxviLdB7FE4qsdPeIts3Ln8NKn/u
1/24BmqUlYc3YdfMBbdQ5sRvCbanXZgB+OrRy1GMw5Ckx/yJKjpyqrv7Vl6dIrVl
gh3S8BqYdfbbCLBnTK8ujUZjsDnidrFLhbBCUegyx7ErYb5ob5GPEzsLq3sIZK1o
ETHQeG5tu97P2bici4mwxHaf5S70GLb5+rsHYld7GSH+aRqiNpYq/D4YuePvCgQ0
vPzvnxw8JCfcLGcSfo4NnpsgaVktxQ4Js+b/CE6tyctyJ0cNanJ0aqrfFOWJwAc/
ts6N8Um1MfqdQDfAKaqKSYLEmRBsDHgyZVlGtZntcXpFueQvCSkuUgEIqGYp5RuZ
5WyrVGxNadIiZ9aqdh8Dk66wcvaAl/JvF+g5elS7tTE0ZIBemnmzJ2Bp0aBOgpLE
l5DCH9iAPCzpAB150b9nKiRhIsU4/V1MZfYkPDdKFcytkri1HMYn/A1eo3Ip+BxG
qU/vISWprrASmhafzNpPHiAILInW6T6jYQo+gsZ8fFBTbdMJhLZK0dKp2afAcqOE
ZVnLKoUehqAlem9fZBGhMvhBFAtkPt1NDbuZlhXH9pJ89Ew33/9HRMiZTr/9DzBJ
WqZ3yQMEOevXx8dVuZ0rRDVtK5wDKg3Qv/cHPIHprwcNy5G1n6rNskxZqJIoJZgA
0SMk9aPTYDuV5xqfwGHTOG4C2MoMywlvVG+7ZoNGO7oSkKHoQWhFlFzH71358vlt
CH/TUSOlXTEcnzENoIAVry6Wq6+WiS7zy10OM7jZG7OAvLGm2lPn78juvnSzDIcM
fq7EB0IvSgXFLsEzH1J4SZhHllECymlPwj86f7v4u7kHRwxs9Pkaq75zma/ArTHA
3cKLfvKfq+/1PMRKiklBGCvBvy4E00psAn1RrlACNFARYZZO7Z3clqzkRKmx8d7v
dyPatRxH8DfKt9Mnm8AvqHoy4C/VYRGTVoTNloudrjXwSqQ+FhmmftVqVCkYrxJf
uo1+1W/pv0E8jA8dHc1U3dKrQ10BzyCz4GlMi9TRwMSrClC4HyWIEbAadZeSlDnM
MazmBh8Q0vM+2qp1u7hrgBZwVStjjJnywQhVKL75ajFX0VKSTbRNH8AhwJh33VVA
RCMa7iixr5mtWx16RKNdK8PA4QO+dfdO8FYp9KuWNALdsUAB6swCLFG7/yQ5pgNC
JjKey/Tpw+hv+QVDRXMIqQlnWBTCTEvcDuam+Jgs7M83LRPn4bfQ+V0XqtNZdnXO
PeWBKGwXyiXDKKgukpEbEzuLrp4qZdEL4s+iMyksZsoccEMGbgKeDc94WUuTkYMK
cHXkaAhxzWYGnSv4ay2iumIzgsVtmDMemPpVk3ecET9D+BMlTBVP+/iWnVmfEwN+
ptbIJF3+CNuWkmIaRs59RUX5UrT/nef8Pe0stiS7f3OJGvRNhD0igiFpl9RCx+s7
pjEcJ2ovEJjktN+YPiYFMwFE33A54/fliMw/hA2fk+3GsSzkgiHu9J47TS//4Ure
+aC4daXJqgP7RzJ2pNGl7KuPQVSh54CD6QOA/+3xWfCzj94thvOJKdm7eab7liYd
/JbqisB9FZi6DMQyC/Ij9G86Z8RFIm2ibFkDaatzv1Ic9jBUCmnMo7urW6w9iPvs
OnnyBHQQEgzTbVAm/zl3KB3pEjVkRAbdBYoh5JVuNZxkmmzwwSSkq7CIYn5oa63m
FYdGeD1JiTq8jHgwPZN4TPA8w23AuJrtVQWsR1FPqBt2f62BhBOjqln2o44+VZCS
EtsYhKAKLx1pCOt5qTen9sedxhhvBSRLM1oxGiBilXvCIZuxwnvGCuvo2iu1A1nh
MCLejE8ujyEktVOEfuWVPNaybt2Qm7d0UjLIsNiN2F23Z7SNHS/CqOTXc0FIPpuo
jAN1hm0GFc4/xnIa0iwpE2T8hAtB2OTJRJ9iIWSAElYXgI8z09RZtiXvDMvH4UiK
C7ieRfYzQvn8pZuj5MIjYY8TwI0CCK8sozMM0qtQjFakJUF4A9aG/WIEEMZRMuC/
nAozwOh8iucp7VJbfD18l4zX+/dDCjdJ0X6XLKvOZoYUQJ/zgPmQzDZPjX9r/yEO
4jVsBK1+1NVyrZHxrpaGcJPx48Rhq2piAmYS5Hd9JqMZJsoo+g+CbLqh59FTL6n4
j1dgEYFXbmX7O0VYeGtoK9/ekKUO0SB2UsAxeM8D95axX4WJudBw21hADhRDXWTe
+hJij5MxJI1Hg/5dwkX08TtTSbb8qHw33hI1pP4f7Qe1CICLuhUy4Xrv9J22jsNJ
9lpijao8BkLEzy+/BdPUO/i1HcEEaHiPjiUAvKswL1QUCGe+PDchMuf7dKe8sgWq
CGD//GWJ7ILxTmk7FaU85M/kCYqw8Hu5zjMZ97qO/mmLdBYM+6czyz2gMy5cU4sB
/TEh7VZlTJABWrWSzgidNT79ZiC5zC7Kp6V2ywR04LsQmKzPNWMspi3AyHZdrxA4
9Lqks/JYqUhYAYeijuoAuK0nDUD52AmkmgQSoQ1FrFSeuOznwuuoiubWeQZY3vOu
nfgmuYEsb9NE60ADoeOulG/ffMnZC9uvD0zhUw28XRgqmVIuD6DfwoUFNcM9KgYv
FLeZxfpSFZ84dJOWAbK5aDLivdlaiQSsdNfcLFqLllEya0XqE0+azDscT3yOFp8R
V17dc7GqMpT7NjeaJt2hGWjn8V5hqcjqSsFzW5OFAt7TS0dmgRh/Ad4zo5Fn7qGN
Sgi2LwPqf8jLW2zYSVvzFAeqjJRZDgSFeC+17iDppA+81Z3+kF0MwqCJDQFX+hQZ
UGtvY9Kx1szlqDgXz7Dwivl0dyxmM1R9NU520l6Pr+XmMIyEBHF0Q6DAWGVVXCC8
lSyGm1JJ/BYd9hhhGDoViASHR+X/cZ3tMj1sQMxLyjk/owE5g6FW1kZZ+FWpOFhL
7oONiEnYisPnZsgg2HvojHF6l3PmgrK0ywSpykbmlaR0NznVt3lWFmrI9G5r2Nwz
RW1kfhQ9x0xVaxfEuOKBYIEiNZju1Z5L2WE1R4Uv5/K3sh8kmTRiWT/5aFnpNiSF
2wtQwIU2DzHkfxXDOtxVh+7ZGehdEidNAIqvB+HEfxSdfsIW3+5KALy7w/9KcoAN
le9DaIdR7tOu9vY8iG+H66VbOuHIrFQIYG8SD40zD92eXiuouj/m3xAug7XmC4LA
mIpd01SL37fdleJcVncKHpNkIfg1E7JbXPjZXeZxBC/5FJSS827Anl5NGS7NGwD6
fQcG1ndy/H3VHUiipU2JmB/Fp+b/YrmEcKq8pjOwu6QxQ20ji3Bn2aWvh5BY06AS
9st5411Y//wVTn6ixImwFXjU2OUIsQhY0Xs851O9bD+AwTU+wynsm+NrfvtdXt4K
4ja7G4oZdoEnUD/gpWSHc6NtlQihRbdjqKwCMY2LOcirzg10HgbAipHsRps29Nyj
/15vMXnei2M9AqElzAv5DuRl+gbnxg9/XTQlkI3M+Llmj8xOG80oGiRvz+L2Ow2u
Cz3atmIp8eLeba+F423pmRdGnlPtoerO6vFbMnUIhoYhh8OesJVt2GnioS0gkoTm
4cXoRKc0hTfBYHjCCYLOnDUQmBYKw7Rs9U5On04zSF1OqQKVK1F+wK+1QmEmrq00
DnSZew4x+hANhI5QzXTboukE+SWB0jYAUzQ4+7o43rxIfZiDLt+65tsVuNop/6wW
/pJkAj5w2BascVE78eEMdg1QiRzfcujpXnZ1I9PTn41faBs/nkcyiTUTnuvxXf+e
Sd+c5OosmM4bEGzy60ghJ3NGGEYgx2bz1EfeZPUqY6uRK1ocAC7iI+p5L/rb/I0C
9Vx46A9P6oiG0N88IY58d7i5751h0FaU3JrtfNgcgYN/DWr2Wznj80RV2fT6FBnv
nt0twDCLWrSgUP8pdtKqBaNj4wLWaaesUA3lgJd6t5+GEnhX8/ugWfHJZTE8ICIC
TS90ZjkvaYspRcyqEBRCOphzkcPeynE0jfZqTv9tYnkbSR9TJKPdnuJqQoAK81Jm
mng/2ugalqNT8WSAMp6qbNCQvm/nBRaoV75pyXNB28NwZTYQzk1eV0DnsU0ndWGt
T6MZB6yYFjqOpMdICWmRBIrbW0iCTSkEJngW5TJB6f3MQnZuFCH4fd/i0iXGJJLs
zFOc2kFkbHpXx/mvNLCONPXhtPtGqzItI24HyLqJ2wbkRpZKqxR2xAAbYJ5GkV1N
SxpOSaTya7VjhKHuZPMEclYNOUCRQnF24PNJHPIO5UZNIzMi5/wIVPP4rTz1jjeB
yTWh+pKiQWtXOdh8/tfZfX/SvVqSiYrxYHWFNIL53I8zpGsd3Oi24yYbIiGcwIdO
dbOZM96d9ih31VJFcNYjFYJUMawcvMD9+SSr5xINpGEHUUKJ0T+HWWqxZhFl6Lje
F7jvRxYt9WhlKPo4XmuEEzmPT1TtEfKL1Z1cIOA1dji0Zh3XOKyGaEj84nTa0OJD
xtqhsSMEvpBzM2IeKv4ManNJlgj5Gl96NcvLbMyW0l3j3cIwYC7CWrSRZM7v0idn
qVzf7mDjLQwTqoGFwyLEAdqrlLAlopROsBpw4HdwMPnRfKpxhWnWg7DWQ4pYl7fb
alhCAKpsNEhR0Nz+8Zmc9FT60rd+MqEhDS4ZbhvTBw/BRjGdMhaPLvnqXMND0pOx
OlkESFO7A9mdFR55bkvUkWT8w4+vCNuibWwWthJ4jtUmghYv2sl94n9khJmqgGa9
wv/Ny/rFZpm2BUdTb2Y8FF4pf9OMzt8BBEgjtGm34r5eSgQmZafk7ywavTXdzW3R
TmIK/qYbIi1D2xoZsHjHV9RuIOCCxaMJctl7BsgQ080axAcZIp7aF1M4ysGSsqp4
dBU07gOYCtSOoAuZod70u5Oxvt5nL5ttvNC1VBKnm8JNSIgDOA/X5rGagWaS4FHn
80HaEE6dF66jEuwgHKCTEqohSVXhN7aEAfAhGjrXQ9XLeE8md9bd3kdKllCFv2rO
vd0Zb4Atg1rzhtKNLIsLFjWlq5cxpUb2n9swY0DguocEXSIx0maf+48IYmyrTGjk
K4y1I7YZhDXI5uabGlPp/7MANnPT47vZY7HV0PiPOKrTgSx7B8O+FHKEUmHhnc+M
Kvx6VVQyIpNPan17gtZ9YTvRGP94YJ/fFxa7Mitxj1Caw6qCX9ckcSL1RoVvp3NU
gkIt8GVOmolvi10xAyvVQFQIjP/MtYU68hUv3TB/X/SKvWihemtupj1qnqh/869u
xBC2xGEvPQHP2w+Gt3kplptdxzErOJ+0u/PwdhlGynah/+HrjuZaLSBGd91ElZZb
y3qzAv/yH7AsiYjA6oQPwS0u7uDkmlZPw9KN+6G7Z8ZjDiuWFyGM8XWO5Ar4GvGK
SmvsoWZ7fO4+9mk7tyGd8zP/jRgg2EcQi65+YDoxTIgYEvlcUuQmzwygi/9ciTrI
l3pn0Mo6Foaw2WpC/gQMbcS/FLH0eqDx2cXBjzs07C3htN9wICyiryCnDXkLvuBR
ep9+ppnE94pcDy/Op693zAXutCdVHf9Cc9fBqmdPmj9wM+jKc5JDB5FL4yu1YEZh
xUMQWg93hLcGp+BoEnrZIfIp+V5dVXK9O9YjhpQ18RWu16Okm72QUwUzJvVqo8OO
BxKANF1zIGypjB18fWdUI4RYDa+KdHcnVuFrsCdYPPqBLCSb8V4t+uEdtcakK6r5
uN0yD4m0bN5K8okrBPEfokJCdlWp/C8FjYCD1BSobhAIIjVsVW9ZDKNq+p39Pd7f
q9at3cO9yLa/QKA+sk3/ExcoBRlcQK/2FsVhrh69sFijXQ4xuRPCJ/IqOWUPHf5y
0TjTgzTTjTkCtlox+lOrSxA8ava7+Zb6rS0J3J7KfHlrpn17aF8Ir5GDTw25VjSW
8gP9+pWjnHn7+HPgwnuljlgKL3nQtqx99Tkf8qDr7C1u3lTPitG3vVDgdYv0MPfo
e/aVNKf389U9pkPY90p1dff5emT9x2FyTWhixKQFeZPNBy/KbN0cTPQCejtVKfoM
tA8rcICcFqrTgShNgWJf/s3/+hFVFjX5jDAC8YHpdSn8MpjvLkqHvKnvBKhrstSS
GarTgHCWQVUVSuISn5PWBi8LUC5rbm3Pc/xb6JWUmGnS799EVNUkMYfqiCCsyiKd
IIFwBDbKGMS/cxtd52UZ3O3lCrPMCO3bIfFdzXWp1wjRQsOJ/bgk/Vv9jbCXAstT
BJtfUwDvsvnv09EOwvXbkWJvpm6aj5kWsKLmRCdK6Dod29sD/KWJmud8jBTygq0N
ybImj2E0mJM7Nz/sTsm1BAXt6qrjvyK/qNCxE89Y+B/IRgJcgg6/COEi4zDbvnV9
aYLs4STJhwlpi1XRV9JvxZJSRuUDo4LC4YoDNwSKcX0nhTso90qfI3jjunsq6GEz
Mdkt9gKMEDbHnBCBj5KY43OEmkTaSTKPmccPBVyd+ACiGjKHEwBtXchZsu8EYrcK
BFS8mQ4hzgXHesTbHpHfu8uagt/H2bFwG4G8p0aZRLbq2kADVGeZrlnUw4AGt4hs
O/T2Hsqyq3qRgTTCZJbuIDqWC2cO1F90u63jIBNI8kWqcgvUV1cGi5SCGO34NAsu
hssQ109c3Qv+LceGR/mPgD8hULayuGCKSe+/cegRadpFqnnbEda4dxUp1MgfKxqj
jatZoi40c7wxsUDWC/hNvVkaN3rMmM7E9ZbxaYZpVj2MqvJVnd0zWpGy+CaNbyWP
HqxnfWClbdc8L5HLWJBPn3ku5C1fbev4ipcWXDpd5g/A980Be1AxaZl9dX3W9n7H
B6bL1P7NdGWVrUXP8LTB8BKKpBUWDwHkSqO8b3y7bq1eo8/dSNsszeQt5iXTkhzx
rOJVVG9loC5mDceQlr14L8BJ9yArnr8JB1nLJUYAHuAFJ7xjAl4K7WzDwwctOKB2
yIZeGOYqjO1j32aGlZrnl/TBlg6rRv3fG8jkgXg1gKsMqfyyc3bcRZBzoUuwn8n1
TOE7aYnbmKQRQzecu+Lwa+EsfGm6AFDkuJyLLKlQv5mQR5N5DMZeAtk4SPXYXhVC
LNYl0CqkPITvPbE+NOmF60h9Tzv9YybVgTU3QCYEO3z0rKJlusW78pqScCTFnz3b
dY8gZAD71dqF4YXeF2mL/Zu2tpajy7foXxV+yoYpKBf8CkTPhkIjwHiHYx68vx40
/vF+5qo9GTADySIDIj1r+Svt4oM7KJWKzLCCf0rr77ZYKanzwr+D/OaLBokYMAaD
eL62dI47MlqzpVP7Sqcu/db1fLiMGM1SaSt9AzMjz9aj7QYxv3oBIplEvKFM3OOe
2COjREl9xGDmLYLmDOrBQ18imhAiEAlzv/ovP+Fg24SxlXasZJh3PdeIZ/5BkMlF
38hAC5J528VwcB++HiTbdUrZ2EjVZDlNhzBt2J4zOGfQv3/nTWk5VEBjrBAH5YSE
fjlq/1ALTaZpuVwVDbi53AO3mbzHltelwk5jQFq1JVS5JKF8xmSthhTUV0ZEUHs7
mQvtMkobYf6zzipMT+kh535pE2wcYzKUBxjThUj0NLf9gRkMZCvl3/87aObc4SLf
qj+1Zc26ZWQ60njYjCcFHSUID4YsJwTYLyyXd21hy33TI+pjGC5gVsWcq6MSu0fs
qqjMoKwLf80VRi0POxTKu6tc/Cnaw6aWUatTGAkh1a0gfl8UBc6SN2hPosdCGcX3
N53+IuYROd6pIxenJskn4uB5dSHBCz8wZEz//MTpJ3v5imsKR0WgxIqgu6Cw+Yps
7FPtKnv0irmyu0cb6CJ01hnEzAoMfwP6H+sHAPwDuC/e7T0+PvxrrvlIypwdNfrW
B1sSQTTH7KQbZTN7hcaFCGjl8STDgkWIXJZB9fAXgu4b51DdItUihVIJWjtpBCXh
HdD0ybVpC+aIR+bD0gs1GR/yO+jsvgGiPEEalM7thvhXhEO78bp/hdJxSg1+JX3a
WK5OuTWto2LrxkJ7OODA915YQH4GkqtCZNU8O2Sr3T397kJR86J4sQJdOg+BEUg8
qMNK/ff1oBkte1bIaQ0DtCDWs40e4JkS1eEGTRRDu3JPRZVXtSnONclO+7aP8+DP
NhU207Ttn31dWMB3CCsRz+OT1zKuaQOmcfpepdYPAcmyon7q0K3Hypx3nw7hvHlZ
N+4NfkdiOTHIoKllmy0hx4LwSLUESSE2wkRgp3Ib8j+borX7EdqPAt+qm2xtRF7X
mV9XM9p/WQXQa/IXlLq6Dr2AxXG7ht4iVx5Q83McQjw/iqzUK48ZMJVV/HGmnxzZ
/Xu3I6H2fk0YJmpiI8NF559dfVgMebOSpAP34m3bGyuYcoQc8CEhP64ziMi0xc+s
6CZx8amRlI0KxS4+BgETGQtpDikUXkkSGQdMC0Th+8uBsAU3nGzp9jRnWr0gN8L/
5WrfHY1r4y/9X9QtlKetJFNoOsnWYmwkkphooy6uXMoRX6tf5KGL9nBd4ihCiydv
e3YYwN/sClW7WXp1Qfozgz4N7UBq1XsHe9cWmU2RzhH5a/6ZAS/GUgpBwdgS/1zo
rmysfFqCmo/STYv9DAU3j1rG8NXj5YBCYFMPslUKLoZnb/ue25M/8MFNYKIVrJ6V
VjmZPR/WM4mvro8nz2a5RlDd7oYAqSnBK3F25WdeB7agNRQm2pQrIuH4yciM4D/D
gp4tWYM+q8JsRLy8DbeJF6DbiVPBIipA5JCZ/v3bj7cAiLY+7ZhnYrIw05sCI0E0
nkXv+005GhH7bcVw2cJpYneMcKIwqXo7Q2+sR0exIycr7lZJVaHc/xoLCFMMS43W
HW/hqsvy5DR2TNR4JUOrTV/ZbOgwaFeo6Oh6HhptZ6G/G643TCyzt5y5SWwxMYK7
dCwftR0afEu0zBqyJO9gqxVIgFv19Zog0uxfPzB+K1MXJtaAGbDi407JWeqQ3y8R
gwE2bzX4C1sWZOu9A1/ZkpQFSsBIizDiDnAkk0GG1rebSFYMMllNasgSrYVglGtl
u+p0Uo4bKKIi0tAO0xKFA4n3kzG4I/0i2KyG1P6yKaMV8DVQRYjobxvx34Q+LhZ+
sU5libbfBaTJDRkY1r0uaTHusjdJbqqu1YmpIfPA0gUTo9EYiiD2vbLf7vlJIwJt
SZhE4/IqgzrSWXGreKqu7UmEsFt3Xr5nIOH3z/ffrfhT4XrNJosfK8wsi7i8eZ55
0oY6XKE/kwxrjuQA1ZaC/+avML3BfU4jbjyP3tSH1+0VePNkkzg1D+bNcNG2jeF8
SIglqVB+8TpaBfMjhDzvjbbi2UIDR/RA8dtqCjVeN0vtJsiBbwAOjWoWfuhfPpcy
4Jzq5Y+TuyxUPQ47dTegfXscWt0TOMptyrbmu12Nvk+vmPazn3XLSzyQyck46lBv
gRnZfQu8MdfFYM39vDkIAUiO3wfVrTYRK/LUYiqP1J8beDCfyKcyckPGaRmVs8Na
KTIykY2+5DtG79CLN9mUs0S/hC/4fuuV2Z4HZk9O8QKJnpH+JcY3mEyzVn50cdnG
LtH3ONB+4aDfLH07ujVRPCl+Bv1DkRu0jOMt02Vny9jQVxCw5z63U7y6R8KSJWIq
zlHJ8343pN3/j3FSp0kMcKBqsngc5ok0uHxRa3l4hleqjle2ncUBasw4B4clxqZX
NI/PA7H527ZXU1z+npcyINVmrPOScNcExAuDFWXmpD5494dZHAp8l4DT7A8pXmqD
wp73Pq26t7DEzuKnlQ3qcO6iixwRF0TNMNPdAn3wyIRsM1ey2bQssKgZ+j5VYUQu
Fyvn7e0TCG2N0Z/VNtyNECCXb3fYmjFUqU57AAKMj4X/C8oE8haS5X6IACunFho6
5am3iE5g7ps4bDKxe0LJrM7FMrah75PMlkVV3GSqWBAMQYvGt8qUvkndADDBVADU
aDCfvMvJ2Hnn/ZXEqYJ7Cu5wlmuQhTsjC2jtgJJXh+cz4W/WZVDWn0DzXwvxE425
JKdzX4x/M1IzSdOPgNrhpoft8lb/3M5kaIEmg0+G5N9qWv7b6HopEWlk/RD23ukl
TbsoLPI6qvnZ4Rj85IkLyQFvP206jTazWmzq0nnmz988y40E2/zAXzPHGgMzqY4e
BY8z5k5VMof1CPSujMftjSdlozTfWfn1Hfsy7I0lB5fcx74yTAjcx9fCfkulGp/y
OmPcXk57aQHtdQQ89sX1UtwsTDSglXGKyRs1Ime5eS1dntLvtGBTNnIhtjxwdUcm
MaH9VVML9hHmaBLDBMXA0uR5U2MwhObZ92Vwmoix8nhsLvwpWFnsK6VBVJ8OvTnV
gswf7i1pOWaUaT6gOIEgam9f+WljANB1RdvPfE8DB1e5F8OhOTExslQ32NnS8PHQ
zU4QxFYUAYGKuE5icu3SCS/huh1VR70qrAZnLFbv2ErLRk+eFQmruRbkjKpbtjDF
ocToMiuodFwMgr2hS3rKo7bUG0CEpibtvlYNjvcoe1hR4buqkCVV+lXPGkYBZMAd
D/oSuv5NlIPc4Kw35lSPqQdyWDmTRDPl79niBmoTVx+bGO9mmPbJZr2iqvs58ycH
rQkjUyDXEL+pHIgAPXp4FZpPQHKPh9BajN22GNRQMLYurqkQ0XTH2pQ4xZCAmaHV
aPG97c/Qzdv/DnTPpLFxELsDXgfz7vp5diN/brTiMNGnFk6QqOgw17/vG+ThKsrG
f+E4OBH7uY5aLniZcoXUbQ9OugpIpBJAu3u3qG8iul9IIlwE9oYNAsG6fmT9rlTw
kF8ghjnqYCZx6PfscDTjHeuHcq+5JNnQpRejkkr9v/TsJoi/PgRKgE7iMCGGZSBi
vhyXL93K2ClztkQqDdme4FsTkN26AITJu1WwzPyudynTxDoauVGzZHMrHXBLJYwx
31tD22PEGXUoKDGWHUvF4nCECwMNkUveoQx2JLyu3a/pdW6mktgEDWIZv/KgUwSk
0Bvhv4Gkk+RzWA+LxsbPt3pGJhKTC+dhpPL1xH+kHXEY5f4QvVgfkdRdAuUi3o6h
aP5onlkvnC9kFx8FtErVltmsbw+jRgxfRGdUvlkyMUZ3s//turUK7y15AY1My2Jb
0bC75xETQxjeR00I6uLbxVVKLNQ6Y3b2cxCOY0vjpqDdyGANKu+ZLNwWlaJ/mpwQ
aPnaPWoEe8rsxG6rwFvMfdyPyP3VfTjgy2GfU2bjcJmND5pNFalGaynTiD6l3Cq8
icUz9CW5AXIHW4oOgh+6EqUxjnDfqQmnskHowsXUiHPEK/r+YLwsDQTHQsAsRZmO
cZlFj9lCdF0/7RIUY/6Tm+Oc6MUKzHIZ5EfsvdPzijcMM0NQer+PFmNFG9vERcDK
63DxCPkwi+X30DMjB7ufCDc3VlYiBI++JgYqkoLYoVzpcJmJu4SeG9VyuujWWy+I
LVwohK/yjYNWiw5ChaCmL4lVL1hiGzjq7FYjhmrEFAcwyfpRyN+NqWlaCTmCxte1
H2Ctu0dp8eq/XFWfzBM8tn+y728RIQZ2rCVInMOiJK+wQtDA3fUzr5zanw5TmFpj
wPN5auAicwkgPZVPR/sdfYihx1c3cnIJEEFWX+j6L+y8TjnP1zbLs6Zi+DPpjVt8
8kPQgEdN1Q2P8Iv8YjbprMFNxIQ0ZNGtJaizhsTlUwAGYftakEiShsGYQKHRkfnK
vBMtNP518OZUkO8PTLyCqovN185CPKlz00UhWbt/ye/YC9Ovn5FMOO0mGwu0ZHqG
fvHMr9860T6hiQVHYP9C81saYQvyTQ0kuRYKNW4SFkxqTwdfTYFAB3Dzifee48ve
EVgjYUiGHeFxiMVFLfDkadxYqg+f4xJkyqcjgBC3UzkyBWW0xi+WqqFVwxeuFvKA
031F3WllxBW6C3Bq7dCELsR13hFPPqL4G4NSsBm3Ys420EQ0Rqdj+F0tvjV/hg9O
s9KXuRuNC0jdqTp+meJiKZFWOGJSCO8SRaEn9B9rlfAYQZvY51zUjjCI2HUkD8Ch
pf3m8dXthVMGe1aQHYnXxasKyPbpFy3r2x65+s2vG+lkNLcIc7fPrBl91HGsVoua
OEjBDoWa7uWbg4Xne8/nusHbvABJpzFNpv4bYhmAk2bybHabYUHpIr/zZic2hZCH
pabo0dc0gdMDCgGeC8xoK625FJyeIZqiNRFUvPBbBQ8aJAdOcjdn8vtv6R8iNN/G
LzhUlloMJTICLGfUfSJ5Mf85kU2ru7m2kozq8YbeMUOcQVvz+56TvoN+8nYUpt5H
U7Da52Xn3VwG1AsEzdJqltLaK6gKoyQ2IGkudiToZPBFUwRAHjWGFPKeEjel+wPO
7Hyh99vZvyMhIi3gfaIg7ww1IK/qTVlSHPlIcl6DE6o/5Xr7GlzWkKTdwFq/plGD
vpmR6IXK22xEJ6NUELTed+tEmiK8Ts0CC4SenQMulLqyXb1AFzGH2UUobie1KhYn
+4DKtGYrPGQBa4ROb9h6/8yRc5Gw8n4/MAbLO0JAdBUswRY1mH60nVH1XWWNU68u
Dxf6lfMHyq4KBYEfvEkWQHA1mZA+1k4esMsjTb16xkriL3eyPbrBvYOa0kiIrBUx
ThDE+k7z1lsSi7C5N8Ztk0gCXXBKs57ANDcFzXtRBBlH+kbtnS0BMxmec2l8n6OZ
uFSxPQSs+Bm2NkFVHv7jyWOP6JfT7Tbpofp1eZQN7mQIEoJyHrWsoRjcQBdr08bZ
tibN2aE9y085r9XBX9JtlGz6Bx7PIIe5wRdXrh2Vi5ZJ2IpywyiztHMNU9jXRMMo
CzPocH28tealCakN+nrTY7PGtTXsqnTkfeA2nhYDv5ek5pzVKvk38R4PCnW1NIyJ
ehbvNUsB3yTMYLtqaQHrppuvdsbptEkpJByOHgTyQ8TPGtBJTmkDizfOLQwPgXJk
fg7thacemoXcackraZGhHbADMXwMYj/QdIKRHaKu/5tGCtFtYgIYGmAQzZUtTk3A
HlYedFTSmx0VoCBRGGBRWAXwjpb6118EOP/Je33NTN1bHNXCdXEdf4RrB9wJH5KT
0M+drzWHbhbiiE5OyQi0zKXTkfspeKAMcX4zGd+94342+zUO/aAaQZ0/G7C0Jh/x
DiNHHHSG01I9VAh8uHG3C3IjuvADFgIxHRyJI08iyxTmfzBKCnvub3w/qmvOC39q
YteDR4SamPQVq8gVY4FhAFPiwlRmSUy8xhb1U6MpzQa5ynQ7h2BwfRe9I3OUFW0/
ULdgkmEphtC2EYFNRTkrvdZhCVsqi4DSTrxP4CJYrqyT6Vzk5lEC2OOF3pD7ct6w
AmZkH+KgKMFSIF+zsIX0rcInUAtNlRQl0OOk9UbJsP9VilG4q6rC/Rm2T7lZnpo5
5/4Xc1OzfP1HqaMjmZfwVHn4zau+FGHkyxgZabWNl5fmcB42gRIimCznbhxOPhDq
cYaJ175hhXJ7PC4Cscc3U3kDZ3ztaRFvGe74rkXMP7vIDaABObPtMr7PPiuAeQMM
EOeOPx/mR03f6izn+PKHaedLlwmAVfXNGZyuD7n0Tku8oeKDNh4TqZ6aaUFnQQwn
Fc1DJATVyHOLsA9ncBl6zkRbhpjHUTP/bAt0EtBtbYpXbzwkw+T6TyNZUW1RWfkF
Q5IWeCLDGoAkV9hRXxo7Oewpx6HMhomxWhWd5Z8ZZOLDelv1LUn6jCj/LjGNCy0z
q3a1W1UoNS1mNhus9vNwcyd5nn3CWvuXRtTNoOp3su8M1d1+cMFvlboP058Eafc1
Tw7nkFT/wmxPyOQ607FnCZYj7BAyWohjb3/gWOLFJzzJzn5gFU0ygSY8EHyU6vCG
RJDkMpfCw8AcbYfFrwCmYDDZeepXEHhlUTYNrrE6LHMzAxpghLoFKMCebWMftb79
xbN6tba9aloX+K/wKX/7pa+F8Gd6zrsjJ69zqzjvICW09Fe4DlfgUKSYyVkcjg04
G+G+VluazDUedGvMBj8XaC7aRG/FfV6zuzRPF+eT5Ng5YQOcAYzVVBvGfsgjvC86
j8GwRFilI0MVuNovu0/ymp5mhrbeTYl5Bih2BLc3Q/AelYkBuORDEKHC6USG9sW9
ZVMbD4zK+3vWIBdno/mqXiKy+wf3hm0bLia5YdkvZJ3IkBBsct/qCK02/dR1VZMm
Sb/JKuZshnlACbfpeKASfsPFwYIPn/3glQHlL1vlU035H3SJyDr5+GxdSMzRDASh
q1pdGdH3hji+jpD1LBoTaFlR6Im63F/uPfPb81II0imloOoFb3bO6VFojeKrMoE+
6BEap08xK/Z1a1BhprcUMvYtk9vzX08LbyL/nqjoIKkiS2j7XKKWLnKTS6wuP2NY
I0x6P8PkyJMxDUgHo8WfHxhQjhNzIzZHe4UEaNqJwo8JhRu/kl05nd7+pYFF3u9f
jOdvaOI8aHrL7gGekh8hpAgtVQ/pUKYjuZ87m9zXgfaDsOxDOhP0tp3U5DvVatq5
CyIlTQ3TnBoQ0VqVHiutCb7Cxprm1rm1wOoDMwUF/3+2z8p+EAxuhwXP+fOmuU0p
myrUMkpakVvqKv4CfIscfrYzxOhgGqhYo9EFbS5MV5frETCxN62w9acRON5i03EW
Yb16YZEVwBLLGGlhMmX3+X5ufgOSdG3sqlPSLE20nyfv4pFBGXc6DVP06F7EB5no
c+DBQQkGKhrHk5/YmtpSHE8w85ln0+1RedmwLRKBLDb9sGLOY1je+DlAq63SEOZZ
m7Z8b/ZCzQMwLoQ+RrEwvKMrYSdkkiPR5JkzOM5rhowdIYGVUDtzmZo8cmPAwuCE
cUTshpTHhrFFSyfBo80EUSM0E85mfwmbTlXKc3ad0ucDxPMvBX8u7tOmqTscZy30
a6LDS8w1TMQddkG7MDdpljTiyB2RihFtc+iQydL+N2wg0JTMiOtxEbCKy/8BLf6w
Ady+ELEaQlnZXtrtI+9BlFzx0k1mcZK+5usnFIzm71SGnKQkJQK69rej8Ur5WRjW
aHKBqLOUKR8JPAgr6lo6zm0ND+aaFfMPqwyKOpItYGJVcfD2liszs0OzG4/+F9El
KlpYE+Rucn6YPlPeZKbiGav9xkbNYn+/POt7iKyml4NKhMCofwGbAMHSRMnVGh2i
+lAfhynprml4BU4C3ISzkMdxPVzC0slF5jNy6yYDShRvP5DzxMvqxlfiiz/NB3Ay
C+TzJQpIuNBkwBdaHbRxm4QPGs/kS5CeoHq/74VeLhTtwMRiBquCtC2YzxRuJ6mQ
uoRACPJ/EFZj/ed04KICWmntuFUSQX0sWO07XYnjUCNo5XEr1MkKz7SajcK1Wz3r
KTtidmiEitOAAQroyxdg3h610uhoMfn1xobfm4YGRZgZxhzJgQIgzWOPVqR+/39i
Ox+gItwsA2bJUigUjJBUA4lG5GLqNkeDPcAhq8cCm1TN7q4zeXlnamgsN7Ki0WHP
ziyvVJFCQyfHdc7JSTCI028LLONMpU/nL+QfVh7aFuHh+IHWYjof3FNC+JaIcWbs
olhDQ9cM+98krt/yMObmWKmGescNLoNAqX5tIW4iPCHIYeuodnDg1D0zLkNXL2pC
FoyTSX0iDlVJzSrDgnXB3NSh3iN537I+oxhWUh0Xet2YXIsB9GV0Wo2jN7bxVTMc
SHGkJKFNM/T+3BYYgUVpffJ8KX7fcUS6gq7ra+wWPItO+XGb0AUUcv3zTiqWtkyM
2wIr8l3hyeXjBdaHqyIvUseEZ7jwH5cFggyZFsALnJ5lSkby1SmD5TfDPYj/XJzX
fQSWWA7sl/vfsXd2hJz7ueDxibaeh3zgG0avicTzMiEnkQTlTM7zxb90M8MwA+Cg
89CmA+YfhCy2utQNkLDXOsLc/x7Oodmcp30rfTW0v6oOWSRqdB5kRehyaEqelzHC
mGghT15vCZeVq1ew1t0tXcuB3k+0wm85eBMOMfiPAG4+9G55qKpHUdIUSuEdzukn
5HRucVIPb2NxYZzXj9ZndY7I276aMPaG5hDE7vRG1Vwd87WL3hqDrS5tTgKjeXsz
TdVsVQkwm4d4k/ERBcwuy/t0pch66Ul3qWBaYfYLem6mvhYtIrGw4akjHHtmN43V
cryTT1LaV8XYDEYUfzEMbWpRGH8sXnnmHZieSy6aGfv+gMEfR/MaPcE2xY82Yj93
H6fnCG+Vs6HeYR1FY8jnt4tlJZcBdbgfupBWQvo1A1F3FBUGBwETZ9aZ9Y9G9TjL
tGpXv3LKGAnoEs0Z96oQVOgYCBkkw59QUQ3RQx/ptbrNmlEKvJj1mLjh1CiaGbbY
xTOdl43sIR8NOxxifByhGpOD28ed2EVYwhBJHRKSckyryW5lq82Et9DQQx7Pmlk5
4yYnJfN5uZmWZcTW0wBrTqq0m2dmNAUtHIAzKDFqGeRadIERAnsQDXSswzhN4bva
P/NfvDKXhQDcBxVdAahH1+ywIOUA3n5n3+GBraoLRaUGLYhlAwZjOWczM6n5jJ1S
iwMRt5X2WtUzinGW/yMgvlwJyMgrnKilhFxVSGFPtBoeLcwQzdOI5fgsZJcN9jad
ux4PwzB8w1zLfNRDdIcosVIT17f2vW6JrzNHp61RGYQ+ZwgM/jK4BhieF8Gy5Thj
WJrvknvIE7rSxmwKvRIhV/+a3KZoDh5DnRH3eGDIkPPxY6krJsPc11T1hnUOq1xs
s6Td/1crNFz/LmMXO1itvnRyT/Gyl8qOP+RUaRk748rSgfiVkFRAsTQl6il60vmi
Qf+iZTV009+FCrSpfuF7f3dRR1v7ig/KtkWlGvEIWbDJghtwXQSTly0D7z0F8r2z
6nVtO9mEuk1LrbdZYaF8BT+E4j20d9JsS2SrzFAj5nmZVDF45R6e1+XpunfkQEez
iOC/HaAbywvBMLyOp7B8vmeDswCMtr7NUzA8W6lGHGo9ZEl+yAb0BIjfcBsxCfYd
e3dW1rqGQbBiqO5LKZjk+gK/t3Xe6Ck/dszHISOV+aoAnQI0nCgPlF/moUWrFk4i
etVlYBdBglXKLLitxhaEyoprOZaQMtalNtF6kzKle09EfUBA2gxgVDgty5N7ZaP2
KgX4ma35/G0gH/v0iCTklOO89jV2mpFXqqRVvVKHUNBaFB33blN5BSnXF3nggdXE
pEMF8AcucSp5L9lLIbwGkD3ZyG6qUpg2On3Y8oThtfsc+nDE8bX/nkCRxFe/whnd
rzQ9w7ys2iA8UnzFMNnLhagUDQjcl8A+UTf/QXNmYXqLXHvK/bxmDEVhHyqRKG6h
d+/48J9MAT/Uex0uQmTZXouNDdggyyjY0ZyvjQOOD3oM/Uptl50+O1hLXUitAqDL
ID3vR3QobTMngWhZVob1cK5IqYJFDJ8dyOMKkDb695W0EYJ164iKG2eYyYXvnyh6
qv4eK5Es8HixiQs8BU5VRrQe2QjRr32cDr+1cQV30fSeJtyfMq/wF9ALPRLCcEOX
xiRPnUjJXh/Lwq1i5QzXIhPtJty4ADtv8PDAIvTrp00KA5eHwj+dh5OMax8bu8eg
4gLWG/iRhFM26L29LWtE45KCH6cy2YjqoNyyaKSQaIJszT+B4ESP+yZ5xymvehfh
wvpGUL5Lr8pyFsV9kBzPtzQdVow/fMbuQwldaPx2t2VnGaYBclb80cMu7sHD0J0z
cRzWl+5eBBj2UCNtVNgekMFfv9nnwf/qGxZIWO3HkEdrYikILquEXA+Q32eNVvBI
y4GLP2vFOi+nQR8IJ2wk/bQb5We20sapiangSWfQMt2gI64MuYh/Me+HA/OPLmDW
cAk9bumVdOgkyBqxGnwcBU/VgzdK6/wCbfbz2fuWiapPN2Jv7jw4EAjfb07A1TR0
3VmpXlH50DrrOHZHD3+lbzhIA1dxc2wOi3JFiEw3XjkO+NFTiaQJbz+BsdWCgAXa
PlDEuv3gizHNStB7E2zEghOM8r1hDvZ+fXg+rYAngRxt7O4+rsX5OYE5lTzMwGxE
T+WgbJJTXUrTONmgJzdogZwjzculhcVmtn8kMIMa2yOKzPZUhwKNqfK6OMHLLNv8
vCMa/Q5YbwHLpn2TJZRprM/kgOvEhKQTZNDBk3dgZQAiYZCq/xT72W2UUQA99tPO
Kik34WE6MPBAXU2rCTkID6VwJ7IUJVmGGLzdohLu53wf0ZsPesZh8pmUvvDQvQLx
rDzXK1/UtgyYdeX+XyXX4JopjMnTukYBkmc6EQrWOoJ+gXel40A/Oe779U9I12ZS
S0dwskTUQEUEqs2D7NxzpOTu/cWHrdeDPV+eMX2cqgTk94aU1F4UpNcIcdPtQVWl
ZD/we8hebqmRzgyKKSdsMYa4nr7kHcN5mzFSX9Mh5RkJ+WtTuKkqDWIoNOhcUiz0
I+9Lp776OyJwWCW0tD1TOBQ0ETDc2DWMPxyZ01lT8or8mrZzS3wxxAdR0xvu85A2
NcW8F+7nt0w7ImQzuTlbkgQmrOgK3NMc0RZeXfmloS0c26BmCWjn9UhcTXscQ8kW
3nAWlGcL8wC4s77LM/xZ9HuQApii10769j3m3QKLAppWjTYB+gXN6IqLiuQcdBs3
nrPY3eDiq8lwaMPMy/3f+nEQmX3pdu7LcFNvkVpc3e1lbqiU9r8QoKqbeSdz1fka
bzNr3c9S1sRkUau0Et+dXmWhWBzmtFjj/PCCZ0OAILXIeHJm9/7r/p2MMz/VLqhG
AamVRNJ8R1nEXpSGk+PhVq+SG/avLLgp5HJEQM/8oJ1eRSoi1v8ypOW2hAeXjhWt
qm8i/idbcZWZjZBh1AObVWWaiyMpFYis6DKodEXejjXWbplPSWSGkfd1G412juB+
0RNDyUFQkB1WUFTiT5L3UEImQag2Kxlw8H7wQXbHIzheac8ezUnDXSiwNX5q1FNk
0YnDuU+T9/OsaN3m/offN1DxDaBxkEEP+GdWBZg74IOq/KMjCa+3FYMq6cYcdY2U
61DxxZP2kYRSy+pN+qY2FYYVazFOVtbB2Ro9/hB81FXQsQNavmyxN9szXISUDMts
/3tNF/zy0iumNFgLyF3gboFTVie0e79DZp7Cm93sTihSh1esMiiYEi/KW8VGH3aL
DrU+BhbLtcQIVhCvVg1mxMONLjExKGoDPW9AxGglQTW2LvmHmujT4ap4v0ghTfs0
Do9mCTFAYiX0+GKvEYphHzPm72nZaRwp+MEbzdcngYsKaCfUHCYzdI6pqcljghnl
Hb9AF5yQE0mM997Io6C1s4nEOOY7qpkFob9rnZ4oXv/mmzz/VZBEshaLo79HOEic
YzuU4HuXfcc3dB587WPrZNHeGrq35AazLoyIUD6y44M0kvwe3ZI0P/y/CBJSXDm3
jzs840YhM5W30ZP3V4bT+0ibGbcwaJlbEZ31rbBtbcUP+JK+CzidjLfPnt35QRJ0
2OIHwPbmFlnmDcm64sNnHi9smC8uVGk42LTMcl3xR/+/3zq6rXb2CNUJvGacHKuX
tsVdt7GQsC2vHOsJ1NxWlqLSC7Fuzc6auMfjJ+r0MiJQFcEpc4NVXhk0W9Nr++Bg
TyGFCM33z+4RnQW3cFelb/UId2ooYRp79cXS2Ko52Q5ZaT4PWYUxyWYrXtR6YYNZ
gNphQvoCitBBTJyaF+NTBAy3NJ5ZDynmRZqsEFAK21PupozLY+T/hDsrSsMKyZ9o
ZMf7T1PhKVI7kKOoXsvSZpDzDHiLypk4dHgRGHNl7tUV8Y3EPAybdIfJl7ihKeG1
+DqcV+Zpl4PUNdnE8y3q4jZKstGlxIbZcLUdgz5o4T7CoV/vvhwSJ0/veRydMxOO
wpcT0AbfSi2x/sCSDrRw7ASybcOWAFsQkQ7DaxSBlK3L132So9W8mbDkGy3AxQzt
bmfXtBK9Tzq3pF+TzYJSlDg9B93c4c8BWAPz0c9ID47/xv5FsQMhlHeRFRoQ6yvt
NzrWfMq2Q+wIsH6NnzhdHF8AWdWIyBomi5Y5iG1XmaDnw1ZbSDi5vKbnYPOEHQZc
hNjZLgpiao7LrojYE5rkz0riIXbtR3OQikhzggrQDw4QbPFzFkra/aTBelvynbLE
xlgyIfSPFW3x27liBDCr/M4ao/M+3waJCO14XGhahW4FajK0ktMoDPmf/NS9JogI
+Vb7YOcAqSxdDhiExFdOFqyPW+ywh8HRH+FNF4Cv56y9jPOb+uOfgvd98fD/iqEv
oi/08a708fUEDIhKJef9R6GtgiG9XspsU+RwnyH4BCajmeyeghNLvupa+mhm8oJf
JbB1npX7R4WlLH9oY7ab4kNj+XUSQXMm4SHJ690XVAcr/QDCftcZy7M9Ot7LJPTj
gXEMoOIjWr/1nW42HQcxtRXtsHJmhG2XKQRZZrQB3CD81r0EoNHH0swu0XTBCkI3
VHQlSRrQ1+VyCVqjyCrr46m19L4jWuFMBV3ZnXNxfU9CSgZPcVKqGfUvOHn2pTR3
EOcs4X32FDbHTlCWpasmeRMOFGtjoU0k27huE1i0zst7NDJ8byRfj14Q7h/cyCt/
CmlOHdvQuqyOo0MTMgkNYathaIlYBKBn6OtgrQbQxUpVtFF1NsQjsFqs1YQCoMST
A6R2vVqkukLEN0dv6pK3bB5n7RFutq1WYQTiT0tUqSOtDw3ZBSLeYLSF7KlbX8E5
boS33cQBwVDq3kgsaa9yHHopzDA8r12T+AqXI5rOQ3H81fqmxtpUkHqUrEFEvb3m
thYIH/2WdncNtL/uNbCITc/8xPfnADJMYd3xDFid1U2Nt7StjhtdF9hG0oGwKTxC
3QfXPe/3q17K10lrpgMLMdb0ilUI/Uc2CqIQ6rI1O1QQmYp1MD9iUPgd1a7NztEM
ZNYdhqyR46zuvEeyTTyoWNmdBw/S86d0bLJJ0WA/LFyQLKH16FUX8T34dlw81C0g
BGnQu0SMF6+zZbqq0kdCF1MJRCPgKR0goqcdTFoX4+sygKZ+lCTcCpbYgis44sDM
t2d44T1AENtgh0dLFXGSblvs8lh4SCS/TCh5AbpRNCe1o2nx+BHFwsyf7W2PlXdl
/xAYjMusW4UlHIvDK7sPUXbPlct/9okkOpt/smZYgyqtXKXMRz6GQakQuGtNfYwV
vh6zOTwgpMIdSxrdPPJjX/KZ48q2kRYxQfQezuk+L9n+fotlxjOptULXS6imOXB3
CogHhT5nkV4Qhzb+8g6FbVeDkJK3bUrl5uOYNozBczoALC/971NxrfyM/xCuZceE
DKh5y6yAxbqW3rEkPMLr9SzDKGhDY8m/4RQMmv7F577rPyQq/041zUCeD+X35ugU
g1AZQdwnPNwqzAl/Aq2416MnOhmjD1pIngxbjT+aAybf17C6c/etipgA8FvwPC8j
C91Jc9A26MpDWJ8OdyUqtcFVCXzqKIc8pWW2JLOkv9IDCHm3tKHSiQCH32rbjH5B
Wz/wavz/+LpVscb3a9dwt5zRc07ZNcXhnL+bPVdivg0ZxYFOt0dZXC+pisNHW4VT
badQROpChkvwvNxdRIlnpkQCqMY2plLtBo3Oy5e68OIlEIlgORrT6UzarXysep3i
KzHm/7Ad9uPlfdTIC2jJht/9nndk4a08Zr/YllZ9YxSIGzlvES9TgFEMZpdpL52Z
PiGHxNQKUZ4fXfz8uXYerIJnj/zroypQHL7LJP+LUuQbDYf4+K7G4vPi0snU7Jel
F2uVtu00AJLuCV22oTfXywJrh+3ve8Vm7cEqE2duUbL2t1+9cB9mJUYFrmarLjDY
1l/1jLKFQ8aweZSnGvqkfdNxnX0PkSNWmFC976X2SDzExqbAil/iR9T0ZT0xmJ4p
d/5z+rjfKp9gfRqJA+iPWIW7yBPRCSW15DQe+F+JyivhZTmVzmuHhXiHbJfTgA5F
zkP10lrS+bIKE8diAatvTElnOFtBSKjjE9SlpR1pn8i3A9BGlt+zeWlNGTr3pGB9
tC3EAoTCjDQk9H1WAm7/dG+f3HK+cy6cZJxn2myNY0nrt1tWl+81a89KMba64CxN
`protect END_PROTECTED