-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
pDxiIyB8Ku5R/oPr3yOYq4y3k8tMWLnqmvhQF/sdxS32q6PS5G0nY/TjlBuPVztN
sW+haoP16IIMD1fmwBiTueolB6G9bthFMru4Ga2ecpRGPpaXTxcNvjqxQW7msEqg
z4BMF/A5i0uKOkVUF2Qp+UsqZ3Oho5C676MLltkV/6I=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5072)
`protect data_block
tabUU+tHik7wPPpOaWSdfBHLfVSTb+nMm+CRxHUXH3RgVTqcOUgD3axWO/PmykHR
K64ia3Zjfh/Nfy4kscJIbU++GA9ozBQceuamHrzEWhNM/uCn/1pWu3FXwQJs0ZNc
wTqR+EzBL7a0Idi8zu5WR/4A3vF1NbohS31hBIRlmJYUJ+fILPlCntLo7iFo/ykI
5C7TnvjD3/QZLmcizQeoBtuna4x38BcucjkVsOt1xJW0RxKq5raRTti5qpZ5OvJb
KKFyIlv9BmceAnrXrbxI13anc52wbfdQdWsOtWMoaUBosY+6P70u1qatIufwmSA0
dpCwvRhMTsYeVuQpmS2PBOgBlJCXd2Vf43aFqyDYfHvjcZAYj7kv6eLGkvxMwsr7
dMcOaBZBv7jw0GSPdrRpmVO6ukI/9P3PfvJsx+pAf6fLLVTcVzXlZMyxnDLNvoKy
fABvuV/R7mQPmjppxbOzSVAYu3/SrGaLsM2CS0lH9V/MZiq8uH3jEQK96LNPiIM+
f8yN6cAVUw4/pd1CITlmF1FJAKrc7QsjVAZGyPT5epuq6LRqsP5w6+kbXbPtZb1m
jywg6l5AioJgJUggK4p1FbFhaueggTNCHoVg6s/wWXND2tuJiEXoD428NcxxafxF
F+8P21mubDOg9Zm3cw+qL0M0nT/5frskKPhkPS0yAzQv8VWRwUGWS40t2cUX5gr2
Hln4z+dG8tCraPh4oHiTccorEtJw3RHHFInZL64SSH+1BdIUA+rU1Mx1LmwJpG6l
pWwVSuxDRPpd/UY15F6hMHWAMehQ7dWZ720P1Bzf3eE40oTyFgaAdP2t1LRBx9eN
oT+j3bOj2EWhXxnXELQhObRiBQ2MoNHFHqCR3bXJ05NOBRAsFoLo7VJn/+PhDrkJ
Qh096EH52ABTUaaptJlY3Eb4fsrqonYMwyG5biPVYtAYKbKUttTmTRgqsqYAtPP2
ehHEkQ8aQPH4MxNPQ/VDMv0tuH7r0wpqrIf4ApssnMfzbe3VdmmBpGGaTqG7MCnJ
nnskP/qYptXG8pytD2tpRUu4nr5vyu0CFW/4MP1YqIP+iOxv50EWh5N/tRSuIe8y
YQ29dqyXc16NUVuaxknsLwN2Xfzjr5LoydeEeUxCEPxsqP4ynpGqVnXB+P1XCSod
RdiacQ+FBoi6bPTQwjnqlzycm01LTnW0rfenp89uqvMkwcRXFWNqyTJ3amZfq7lQ
B9NRFq7uoI655sFvaY3ClHK3nyabvmmkafiDwLp82iqRAg/kLIr5b1yDsLdYeyL0
RyhihZozENQn+bwEglfQ/q/LJIO0wrE9snb2PgoN5JtkylSQhCiIKBY6bBdkLprq
D5lqpfeZC5b7274G8Uxjxlj+idyk/JUJobLXORjL0oD9HjyCmq6jI0Fo0vFbJhA0
sIWAn7VGHduVZtwSfkZvuIlIbx9cLI4037KMYrvAibQoVu+iW1AOTWm/dKssxCPQ
+6aZeTGX5nEx+H3KfEW+9CC0XC7TdOnoVkgWd+5Mxk1VTgxwe3+pCFopWq9roRv6
2fYxLWFl5vm4OgdWus72TRieCRVOU8q44afgEKQU7EWkmT/4s9NePmD4iOb5BYIQ
rGXyImHG6ytgyaF1d15+Z8tWCki1kxMGce3pa6JVoy5Nx7vTyh91O8agYZNxRUsF
TLGIpqQ5wHcCHHLPdy0N0PW+dJ44nxgJdltb4cOYT26UUjxUh0N6iD7ndji2MPFl
LYAzCr31vITDw3v0ybVBB0xEudKbDuWXnNPcgPOZRwUPthDnjC92Q5QvSITOysTC
b7aHCpdJaUPbfUUX56ekLXG37GKdWmBHt7S+tYTFAcHnpFTy02z1DDIMBbS8G71U
jmmTVARz/UL3Z3whoQISO8K62JtGtHS/3MvtjpMiLL0S8RJA3O8vOtKSUmgeTMu9
67omHHOe8jksMB596lghqzhypL3FGTyvZAwk0+Y4GUOp0hp9nSBw4nWEUUGvV7Ga
icmPyLHRmngqzrpCOpA9XwCIGnk7wge7j+GwMTNkKaGw2HSvRpy86Uy7at7P1rLg
4j/OqtctO+nKcBZp59Gqyd7k4TwDcIyhYYcPA+lq2hZqbv5ZLkWJo1XhnJwMEdKz
6nFH+m5rskNrfL9kGO9kb0bPB4kstem9z23mVfTIDwIHBV1jAG3BPABrsOZ2zF6T
mjBMlrhJW9pxeo2rMXJY1HAOaaMfPEiLgUB+kpM+4oZg9wz9dhWGbwv1sXDpDgL8
xW/hk9CIH4gN9wRm6svmX4LtuxxMnFDYYcC1gC7UJj4OKq5JNEvVVXm/hXutYJvZ
0Fx8bkRSgb/Y85zqLXgAFhs2BgfTX/yat8P7+tGKqVmN2FPnVXomT8pGiOY85a3P
kLLHWm6qr2mqO+FxxBnD8EG0l/I2kl9wINsNwCYnro7fuPzdwTCIvAakCNjLSkaE
JXmr8bGqcLyIGkbgVThuOG4K4aku6gbmZZ2BHZKetJLZkHw+MuzTFyIW62n+li6Q
Ugoe5PxLIEfiwPpfpc0pRPNoyUUVskX+cFz+2Ko6Qo8bNS0Nu8GpCs8Y5kc/jVKJ
o0H0LVjdvdXNVKC4csojive3+o+6rBsw+7LveffD2RGXxR0ArT6i8I//Nzjz+utN
NUPaJttHe5dA71BpoMRG/Eja9Ri6D9sfNyphoXIwMGIojmW5nUy8Kc05JRFtkeiv
6guanRWLaqSGV8T+m+fFCCStGdiAt6HAZUDgkcqeNG5/ZpmAYfVDmfRNrZoabl6r
/wEWrTJ/ZOaa0B7XHuSqmnXild9Z0LjqU81wF15YAT03RpY8iSTWy06g6DKAQlTV
S3LqOCwZNxeVDMkzVBLaNMaHck2CWdMPw8N7U+PbeOxlaaGFXermKSATcG5eGxTY
5H7cVzMmVP/rm06XbbdDsv7n+M3qnydX/s/pxwUJOY5kuPyGS8EcpzBoJoa/Ei95
el/HKOoTTiAW7atvsP6JoslJ0arpUrafZ3WThmn/GWtLIojGdBhwbD1BkeI2psRD
XrM29HxDTrJMyFX0f6fSc+bDKPVD2tdRDC+nhIBhnDWPPWXJTARHspRk/5vZIqCT
yafB/vi1Y93W0vDAMPRCjjtJC561gll8FYQ8tM4z9pb0on9HdEgBu3PyvGjkbgug
dCpZgidcbvW4i3rH41SR6uR4ze4kJ/LVuv9/fa1/A7JgQXp08FpWRQBmFkf5ooG6
waQLEyxujEkGTEMgl4/5mdnJvKaW4z8DDe0AhVeUAc8AJJwAzLPRmbO+GUqAdJLL
RN9FFcgzyc9E+TG9+LQODLgPE8Fvm1dv7OipY80tbGMeOkkhMLP7E4Vp8p6lcW+0
5vIUswwpxoQFFmB3bR/EINJS3SlPxnH7f/AGsEL2QgALvuLBINm5lnYZE0M5gJRE
4Yw+5xXEzhlScLM4ICB4vlmyFoWjVr/dp/QIZFy4f+5Z/fAeeImF0P7fT8OTa3Us
9rtHp9LYtVbDPOKXBORIv6z8UA9mQuntNOjztpIAirWnsLNJqd+SgRH8QlaDU768
AJR+CmylxffynrtjElBEAhbqWKmtFZRV+8AqEvqc9jBaJuc9xU7kmoKsNJ27SBz9
fICh6xjOZrOQUmKEmaLWfcuLsp36+YyVNRCXKCdD51YnMTCwBcLStJb1lw0+JX1+
jyy6K+U4UtQf97jNa7MxafVmTjlrtf2d1XheqTUDUljF/wYVnSvYr9TIB5BjFJNs
+I+NGSM4ZhNPWalS8tn1wBkHs+6JQG0VR39TLCSSQU20mn/H/7DxaXIL+rv3qWSN
FGWrbCp05zqVVIbQ6mVoAGpdWANG85UMrbVGw50TvFlyWm4fnwe1tigR4f3sVMxI
8MTrfCNMa7PziN++v8/VXG5/QxYYtXeq3lXsiGA5s1TEow6ACp+f2xyMCInMSrEh
YLmxlNX6jU85U5BDuWeqIZGBv3T+oVoGe4eTT6BqTguGkUzIhqfgtIeBlcqZlay5
vIGXHnvbzka0GbqqDBSfHpNw6jJTw0shbFzHigBtILKB4fZ1xS4Qxn3LGLzPVns0
lOe1+bH8Q5YDHaSxxdtmEtw+HJbShFAUW8U8u7qR6f1BEqDPjS9fEulI3gJdenMk
7bKGLtTJbRdGy9UKsbII+3f5TaHCEjdKn4yYeyqG4XyGpoVNQNo+2D8EcLKVbZyP
b/ZR4Q2e4Zc+e8QCxnTFOlCmyCgwMFZC4My4i6Man8Bumj/4cEOuboHLEqjzZrP/
O6fIxFhY+2cSdLOE6vom7LyzpLJp2ZyJ7hR/J9Pb/mIRRdfI6FL/2k5ait4FsUgQ
0swqm0LGCycWlZUTo9OSqtoT1kA4Imzlj//h8zu+8xXAK4cN5vUhtXyUwcJtXRi6
94p7OjlS5q9CPsPeFoFCzKmSo58cXt7kdvq1NtB9TpEcFnnLl1qN7ybyD2s/Mu40
jtU+KvtQnGMJJaIjZCW5XFowVH8KOSwEIL/8jQ2R6uB+w4jofkm4eKcCz6SGjo1z
G0ljok1HdfjJ+VblSOre05v61pxiE72iEL2zTkFN7wwbK3U2VhpNRQ/takh5BpOX
v/tMo+jPxVv/fNQrNlo+FY7Pgvc3cBN+TnjQlPmkginqL8QsHy4mDxh4xQ43I/wr
jh97WDe67eKR/MJqegmNXlse52N2g08cpE5yu/PYEtYICc/kzO9jcidrayOfNU7H
FC0UCLWhM4n5AwY78kqnasDzQVNqUfpn+eatwOyfiCefjB2kacRgGY3bysg3C3N1
I4GfnEG6pAm1nFyrY4jlsFcu6KVErWDcEJC12cnawQmDlxujGlTfhnnAdM1vIHe5
dF/hbvrhEy9gQB57eKYfRMNliNevEJDYh9qRYBSS+RlsoVb60jE/ZfIql/hR4RYe
5p7E/NbjJ6Tx8hs0tCgX5o2Od+9/t80f5p3oglzGtPkVF11eHl1X875TGh6PRwK+
xMhYwgp/DUeh8S0lGYtNIGtjOIEjIJNpDQiigrBYV6eltzL/5tyUM6dhXwrAeI+e
CD+MgGRXpwAuCEGlao1jN3ttSSpNBQVI9iWI77CZgHjilG4BzPkISdfFOjuxbocN
nOmAO3nw5vbNiC3OdKly5sIznU3+tIuIyER0iraBc+9i7MwwiGTY2a700o3c0cTh
5idBCI/qQe8eEeNBYqiwSEwlCVW5v5llBSbFQ/H2scUyiqtFCv5SMwfPzC8Zgxeg
s0evrnEdT2jZEaR7PsBKlu4EZhiibZ/RYJCtkxD0Vs7PfF2tSE11ParzNWLyPKga
i73fkQnB0nAKITvDizqkFh9MNu89J7gJDiOzn0p1TbgOXDU2QFnKyks1lhWda//L
iA8nRWou0YGrZXdJ9pt2mXz9f6ELnvF23AnCKdX/w/DFgmDs2VOwBtHA5mHatyKc
U2sNcric29mEUhf8vSoiAE4RyQz2akXXt2/4Tz8LuigFh1mEFtK0cgBBEKYWqK2F
2INw800MSx/3wtIJBn10J15LwJPDsIRL+12A8D4BfZWrFv2UU/WjGJS42Lvnal0y
Sl95T3k4LdoZfm+Vr4QJ8Lh/tcQUTKGgZoom39Wi5KXaqEyAWIOc3tEYQ1vxoIa6
EDLhDLwTdShSfaE6KwJGpKPEjCRxA1JdY9gp2rhNYNoYVZSZUzcJVfTSkP6Qr1bL
RD8GPqOQ4Y5qWNSKRNFKkirFcuKAEFF3TG3FyllgPLYUd+XQzwZt9uHMw8xUMKXh
P4yWCkPwSFCMC5VOGpCiY7v5unMq6AQ29obzM6irHkHFr/IOYYPP2eY5+v6m7kjV
YZFappJxjGaSxIOblLbxp2AiSv1YmmuQQ5+WwXAjBNqoUY5oqWZnFyVL9kh26/AF
DSCAUsYBxlUKs/e9B7uraZS4Hc2hO/lWJr/EFoCdB78ctr+gdJZLHQq4xiUxelVC
iXZXMYRxaiiVVp1Hf0PHiFbTXmes0UAjnVpFnQpJoA7H6kQAGb7b8LZrWWySvnoe
57u78IPkpRVRChvPuiK1Wx4mZffVDP4gcV91S91cCrv7Lz4ceeTv2LfXUF8PC5LW
UR9y/wQjILCcZJknSKVN04XTdXyUZ2kYoNfricDVwMzLKnrejpktVKvb+I4rv6Us
0n1g/Jf1ERjQqCtyMZeLXVqUC2TnaF9SEEHx9VRqlRtLxR4PRzInsN0yfMnBFiCJ
gfSLcC4/RctuuHDjTDzx3wm+NrjSNQ0gtqGqyEr3DD/2LHj0jE/YXysmsbPZA1Vt
O8LeMtybCpGWZBl0dANKhBvYIXM/BUkiKxPrXEvbHaAYaEhDHrRxWiJbNTMRxHiO
chSoolbOkkFFffJy03WpVrz6k0+Ljq4jJgGkP38G2tU7p6MEkAup4Hkx05eQpMMr
q6Znol+iJPr8q51XFeTxc/I/kAZsXxtGZWigzuxE9nHVNUnaOgsOEXJP3pEYwx6E
pH782J4CH1wO3I9tp5MwFNmZsTu9VDTUJQGN1vx14xPdgwOaaUpJvxBRaQ9n6DVv
37YKxdFfJWrQRuxoVanC3HITEPbVosyjwvWjnMDt9NbFHJ53NcJjYAK5nueirc2N
3Bbx55h31QOd0jxBDD7IloB9bI5Ad6NnwARJCdnWPLJ6Kp8wB88QVw8GxcyxGgMD
MBsJ7vep6lvUBuFMy2F0j20Cc+59wy95zdh7yOB2sRw1zuzEq6TGuln4rVQ0Ck+e
sOghWPFHaYpXH2282NiW4mfTZRR/v/3SB7FWqy6rBo7trqFD6/UvFEdYHEIoNSGO
OtXaBZ3SHVXHGrC3LLckL9VlUnzF/sRxMtfOlrRLj4M=
`protect end_protected
