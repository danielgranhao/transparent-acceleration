-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Q57JKZcQp3gWHeQYcSsCYfyTMKj5CtC64SVLJPVsTOBLTx3o+nly9ogD30zqVfBf
/nmRYsTON9ObiRdSR/FDUqz9cfaj1LPmicdgxlq6Xo2EoTmdE33rg0B2HT708w+V
BWQOWdvMqaYGRRnqwU5Yqgpar4KCkOx09JV7zT+CsrA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 1680)
`protect data_block
09QI4z5khNMVNqRTbIMKD0rofWA461OAMQsmDAJvEJQgENHriSp/pOB9TJrxXuY7
iDtibOQku1s3NGCeaFxmcf1hidId4D2m6/AEnWmu8GOJTau1xsZy0N3UU5MDgXaw
Im5e1c2TcsSVcTW4vcVUSwWN20rjpZrTW3NGgaFvDgzyjLDfGH6udEGsA8MvqLPQ
v5nqs7ZO1ZJpw4ygjG77F8+LSZcsxQyAh6k77q79gke+jEvZbVp0vqbZbh8JIAs6
Mj9PBa/lnf3dwKqS4oMaHq78xpLAtCJ67rzErjmMFM62/4K2RHWoY/fyjHZJXh7b
4z+FcdaWc28+Ebf9gMUaTslLVq0qfqvO2zvXLaMGLZsot3009Zn6woHH4zl0X0rh
mXqYXWFtPsAGpS5qX2134MiXNmopT5FYCBulxMX6taoQfeMH6PZU248nw6PU4F77
w4EoJGqGYxuySnk8RiqgKlNWm/YJ4+fnEqBI37Wf7QrCEaAdegkii41WpmZindO2
H3Z57l2xUpg+mDqYtn6hSsHlZ4Zsmw906F9hK7w8oYe3Jm0q3+w+ej845ZV2nYcO
ZqsSgiudh1qQnv7Lz0R5pnZauYhPCooPiDCjw70Q6fUBeIpKQkqJNxd2q2PZub1z
RzyRwi0We8/QuPmAFauqLbNwW8dvV619mz8d7Of2Qu51IrxPaCkYPngcBvJQMyWN
wGaGmA8QGkrU14DNCMfcwwpAfqEkAVmj8wYkSwGZv53j5SHIYDi8ZCLrbTfM9RQl
IZ3b/X9dEGrCDeKYfrN7ySy9Z1gxVVkUDfIhno5AuFExgaUVW4z47O84gmb0Oefr
FfdpwG6K5LC0KaPmSEwXxPFhHlSuzboIhfyniE6V+9i23wLvMHtMXLUZvfpXFriK
JBq+50aMPcJTvpifbJ64NfSXtwCVBog6+gr883mQ35B77jpBzGtFN8aXyabbOL8n
Q2CVqJ/djStSxzGcsYhR3LLeMTmRfE9FOEGEId0ZCnXPcKHRlGcJUqfrp3JvN5WT
IaW4DpHUNTk1tCB5JQwVx9OAQ2arpViLsNC5DFjF0s6S/X0Irh8zp7VmnF05G2a/
UQ4ONn19tfU40/Qit03aF26p5dKcDz02XUoKEoPYHvN9EIqipu6rjekY0NKaaLqk
Zu8w5MARuEg54PUwE7QGyHxhab09jSAA/gDFYCTo6leZohJkxsZd2iSSalgtMs8D
5G71SSxmBBYUoPRW8foImKHAYld3wlxhPJI/pRPqn67jUh8Zo4+I6qfJ07hLGuxw
LQprgcW4gTIyoebWDx+0qjalWQ3OQu1w9SQ7WXX9LEjs56vhF6IMHcduT0a7/BCZ
iJI7ym4MNBNyjWslkO+nekfRnufS0SHN3xgKIyQnw6f30JH82wUkuBFUh8XSA289
sFS0l89P5g+uu0q/yDf4YwnEZb5jTud5o/ie06xAgelUetOLjSFbBTSWJd1pzCOr
PZNZEtVV8n9yvIhg8YUBB71zyZwKZ19TEdVRwmHEDn3ZjqdgFif9nbk/w5mHlyfW
6SOx+TDXfod12l9xk44QD33EdRMDYV7n4j9UjIDeleVrBf5y7iz811luokoosf1K
Mh0xkhBiFWUfJ6cV6mwzeDTrpv8GEoajdlazmFJLvRqeg9gjGWp5oUK5EMX5xT0P
f61i12SK7rUy2hSI/NSc52PD0QiUh/zWyR35HoHXuvyesWCCbxWiFMa3GiluE2HV
jWbWZyHEXJd2z37c4C5PHv+/Xt9ZrHxruvFijP1U7RRixIiaEd8PCmGJcxfBJ0dH
ymMC9rLeHY5jZudBdy5ttmUM84aqGSTyMn4uQHd1gOSTF20GhAfUY81K9RxN5X4q
e8XhuN1jwXd3dyQvDgNqsRYpbFDwdRcMVDbvcUTRDt/Zb+wVvo9rIj1Cj1EoMeM6
Stxo/VpLmQq0O96CsbiaS0oHnAVZuKT1D1DUd1c5C5rr9rlx87nDopcGUBpntzvY
/uuoG+IGYA617k4Gvm2tPxhj5uCmceI3f+/iWnybsFFGWmCE/80NZV3clkHIHd58
+HmZYmSw3+EqHhXBI4T0jR8w+frKTo/0aw0XZhtHoCYOLcnZqqoRfILrHBMpBSrm
DfaJ9SBLOqG5XznC1HbsD2qb6SFKlndY5PcSlwpvbUEZ8P/E6jBWj7wBFFfao8rR
ySatQAmlQ+nugMPKOZXn9XA+N++gdrmJPBZ38Ds++XS9uExGK7LiAXhZfVmvLi5L
`protect end_protected
