-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
VSqCWAdPWzTrZl7TSdwN0SGkuBIrXy592qlgPMsXYhEvVo/2PVuIDGKrUxQXboyu
Hx09VjWgxLdKAT4mfkfIWqnRjCFkD2vhdRh/IFaTfldVRb8tiQ5nVGGZWV57S1w4
8sGHzJTK/KZ8BhCG8hjr4C3Ci05G0rD89VaZQa7f6w4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 36301)

`protect DATA_BLOCK
HR8lEi/9ioXPPMbn/bszsk9fcTgqi+2SeVaw9SCwHF/khFe2gTrcCZ8oTo9HGyCD
D2L1DkN1nxL9J47POfsn3Hj6xviBS1RjQN47JB0OT4Zh78AJvHWGOsVRE4zRerEw
2m0TXv7UX0Zuj3dUazyeQRaNGNwx52sV9OC11HEjrfL8KV+Y74c65iQJ3XN6k48H
ZMJZw2W0OlXm43w0YdbPpCRT26jLTXA2PubJYUqZHX+73uMqHInfLjUbR+0DMMaT
1a60h4pE8vcB9Gzwn+2SVHFHZPf7YWb5vY2sh59xO6866PkQ8HCpnwHipH4pxrQN
cDR4WYlDHuJhvxiaS8O1mQBzMgHZyQD0dJ0bQrpT4RjPIVdyWoBEG/yv0dDKQlfI
EO5WFwX/E9wd43D3/7A99ZZ6PnJxZ9nCkS1QW23WV5hrBliHB/I0fQazphOl70ts
1SBd4UYLbVPDVYTqD3E5Zb1rgDzANI1iwbKKRFru5WCyZkJyt0rtsnHZwR0pMG0S
K4LTfs8Cf9I3NhbHxbck65JF7ZjYFk60+a24M+eWpxKvHkqHcx04fK9wvgzTxT1x
cgvo+0KGWkIlBhfw6TtZz2e/NH+gQ+BKnJ1YofoxGSD8HJgEMj52u/FvM2B+iL32
EvZj8+5GlzclqV8I+e0+daw38WSJh20EwYnqnTC9fC8X6r49TLagYKbFzfBuCp5q
XycG1c9GIxeF/ncH5BlMbpYjQcd3mtqf9HtXhRrXD+bw9lc4Vk4co11ZkmmwjK+0
fP+xrw0XQOk1u3EyIxjd0mQdaFhE4hZCd0FvlLTgblq20/u0DJCZTMQRbDRaoA9m
U2IxDZjVGoSHrE4+LJjiUT367QJH0oeXxoDZjdUuxag1asViSm3P6Q/VnqBk2IR0
KqS702GGLAgN+QNO2HCf46+VzwvLe8e0ub5ijJ/IBI9pWiqXawtmis03woMxJUFV
W/vrrRLXc8enIVA8uzPH1uEuY793ompkTdc7LTl5XMGqEgndOrO2SOBR0lxmEnnC
TqRmoy0lPuOb5daqedqCxrEzgveXl4kU98KVX+/yf9m8gdrbHhNIQOUlQT39L0SF
ro/LQc7kafYfJIQY3mj5eFY9eSJv2dGfvOijWCAwUxYeP8C0K9XSCrVUPLhQS1nY
2Fu811RJbnEttjjKqMvWelJIsVsHuI++nZyH/KY+VW4Qetj6c2+NQLIvyngyxbBI
X0hxdGTMaC721mbeurTclveUqswRdJeEqwGwS0CEMoD7FxcykfLj3/pHO8b8WRk1
7wtF24YuUDL5mUf3hDJ8THkicK8eqMSd9eOnCcfuuk5PbqZ+76airuq954/sJ4IM
iYRSul/D64BVZ2G7C4lw5rbWxJfyt9BTau6k5s2e3gCFNxGYoYRb0IBQZr1eWBEq
E3k/4x/ipKM3qY+MOqKJIh6MVMvxfjCXZzCs+NgnKotYNOc9ydzsPMJC4+QaD2iB
mGXR4SFoz3aKqC8GuHDt9iKAZnyD4rvBD2ZOEcoTy1wI5j9pVmaMnmRwtn3oMnf5
hw16DB2XSuzgJDTJzgpkSCd/Vpi82rGtYYS7BWYOWFhfzvrvBJ5onZxXdy2bSksJ
ljReJ9si1Rc6DdCIRcqJ/HxDvLxX4L0b09GVfFvrqYD0MVqr1IK3i1dqgd08vPn5
I6/eXvQvh8Ic6RuLdMF3c4A8dbnBkpUpMTDCyfKSrFhG6S5wDZax8weHguCYFmh+
14tm9C1DYvJoECh9kCTVHtvbYGPJfN2u36y7GlxLSsjXtJ+xNXnXeYg4n7RZjWIe
6CaczOdcIRcqxeikKRLOFwuJcc2kcyCLlImoDN0EzwkOmx+pyoJzgc4b0wBs/czM
wDDjUP6xyiyz+/dyfLanliAclYNzAuCVj/JTgWlHb9WH74yfaZjmxgWaUijYMDLf
3eNOqdQOr5nGXSfn4xpOurn2KR8/O0szWMW45JUp8I76DhzXAohVXBQSOuDFO39K
fsNrL89TTz5M4leaQ7v391OOcJaQZskwHLuWnAFB6kS94qE6Yo+XrsiGTgVdBeFn
smfaZhY4fDImsmrzY5I0mDD+1/yhnuYO8SLOb0dU85kSI1jWhfTiPw3/c872zR8R
JzwLQPaiPO6nXouARMnNWD0Nov2Xs0svoy0YK+akgr01JPyFkNTkxMa7SY/6+61C
A0efY60KmM3PrpVAte8uLApHT+buMkjKg2+ftfIILvIS1qMWnY+vTkTtMhjsF746
V3hIBB+VllW+35nVTrWEkE/9n2pc+mZONgYf/7CVpE2Az//MoRYQKzn6TgEIftsn
pHkqy2fnQCht95m4iENwuF1flykr4NG9Ye+hKEBImMrrPk8jOSPTKA4EediCmGXD
6XUO4NzBMW8PfV4RQsbTl36w24xGtpokqqJLSpYaVEVhNCKYOv93xNJuydCtEZVv
hM2hntisuhoQD5ejM3pqqiJTpTK+0Bi4R94P6HfbpUaGlsLA9RX99PSjGYfzWcQK
6evzlLe33tPFVPfwR8BX9V5LAavJj1Tj+zB1TulNTTuPoGHZz6WDPiv36rSNSTrt
isLApU2AzzWwj63n/OFkv6GIwL0cihEIQKtoYswU0nGcgEN8OpewQT5x5QQ574UG
sTDbzKOFg2A+5cEtlQT+Vx1guRoQR22BlQPyA8YHmfJ92/qgf2VqSpYZK1s9ZimB
X6u4EhY+qIJXPYLv8k/XAUlP9B5tQXEJK6eZN8u+VXbN6Qn0UJbx4OPtkfOs32UZ
HqVH21Ietq5sH8zvNXLNi6yRJVwKCxlkxYwXXE6QbmTqOxM8zcJ8mJMa9Hv2vg2Y
TxVw3jhtG979DlkR/eqCR7B9HiWcc2aVPMO4/07jW78J1LrNBw/sBdGCKDmi6yhj
w8h6xWYBO8SUaaG6MUucfkHtJbcExv3l8EuiOofi3R6e02YlsZTttEFaO+IKWy12
nqPG1a+dfRmMInWRNRyR/b8hltAnrFsqCk6DjMc+qZnmrQnGADywazbQ4O6zt8UA
fVPA0BbQHpKqXTN3PzO9K69pLB1YcxZocUHR/3wMdvP0GmkM0EyVMj81KGyAJBt0
3c7+U/+tDX1eFjEGDHS94mtI81BQxbsnEwMe87qRV5NKPJ+wZqMubHvHRP9/JbCi
LqCTMuvZW5haof8f0cfOWmOLtO0B2hZxEsEdjPJreLU9dNTNMwkpygy8641+333M
rlSQM/AqTHmXJvwXmypdN2ptgXoNe1O9g3ObqCKXo28kVqAtFVqKL7ZP8xGppIWb
rWKQNdJuS769ZsYsXkdbjnzvnKfGZx1DbqftrgsecNgMSO6mZi0+I6XUXki9RafX
q6jU7XhfZvTha7v6XCfuxt4jk8vfxEzOE/eP74k+hzrjQW6N+mBM18jEep/eqFnf
ehzq5wVQq4/dC4WErkZ4W+rqN2MXvM9Ew9Nvsqns4gf/IylrVNztK0P6mByt7s7Z
MLKKx7lDZ2BP4UIX87CBeh4cWH4dNsiVNsk/dV3rmcQSzr9RqhbfJuoyLiv9fuBj
jJX9XTj7uz1oI4X0/Z7t/IKW99HzYrt53EBNxCM5HX2QD+j+yvKwQdYMapURJgGM
O9s63LBF/qjD3fiX2kklQnpmXgt/yzwutpRL9oTvMFnGvKrml8MZN+QkL8FngYZC
WbZV33G/aCEgOJRCmtz9+lgWgaP1h8FgEhuOlTQuowYQeFjtbgRMl+vYNDH/3IAH
la/7YQ2ln85OSjeEEQgO/OGf/8QLk1fD8mObSEcO+8YE9wIyr9f6Ckk7f5z3QN3W
VUypkLcdjlxtnjPpQsrixntI56FwjjMehzPKXc+s188msmj6dRl/Tkx7s6jOvuMA
82HZJmt53i6kycIQU8QfZCLRRHYESStFyqWMuqzOL5i+Gt8DIa7W2JnPFrOXEroA
5HYQY6KftsVYio/+i/ZjKCPR2GM0NuNnftkwgQrFOnalEqku/EGVoFL8ISzdimQv
ebMdDs94uIqmJK2D8TNrPa5ng7VFLTrvUjpDuB+268XbajKvTFfP7gZLJMMpLuX+
S5GO2Vd6EzBio3Hbb4s3RpOnMY73E8LxSqZcuhUemIMcZBGdMS7+umn9RNdn0Giw
W3pw8ww+vhVfV1s0q0QW7yh56NEjJKBHW25QjFb4irTEuKvbUJOZ0oQqxVhoCAkf
XipbZKeL9QDc2kcCQJhvpk0M8gO+wHzNT8un0fQEaAP4KWqYLzO0ClBC6SeVxfOB
J/bABGeic6yPldQVfGUtrvtUb8FnWLX7/VO+yLWEd4Qh+DkGKohR/b7Xg+8Zot2V
Cle1zloDmZSdGHpIQ2bU2RGeplLn1UmzLVtp8uH7tUAxx9uXcqVYmzvZBzFyghw1
t00c5G1D2d06Y6ZdLZrhxdavj0LS5BumYX2z886lXsPrkYSdq5f8Fs2Ak/CALOb/
HmM9gr9vC8+C9mkd3nzf7EBbei1OFLmKKmcX2KOewaJODPJiO0GFFyvqwUuq32wQ
6gGjecZ33tAjjk2WhblKKVqZ7/rwob2eS5KxxWsQq5Nj/+n4ZK8KkqdSWLEBTePG
xZVv4FLeayw2ZkQsDGVmj8v3REKIZ0SHOFG0FjDhXtoIIKjo6CmWl1M6pVyZ8gHP
kJG7UykQ4OLo+yUU7wgsNe9eHAYesIlMal75/BLABigjyJmsUKPZsTh7bwT+EmFc
1vAWzsY0qi8jvuRwL1yCX21QCNC1FEOgUgsmlabFPP28wiJfYii3W0db9q/baIlK
AZKFDDeMcyhIPgtWX0pAt+lst42wskIAIGwHqWIvmUsOsvt35F/vWMl9ziPsc/Au
4Mf3j+DKul+oCR7Mx0dQWb8Po3ZvGxxMAJqetDgqV8LKtxF1389GySpY5Isloj1j
BrSUokUAQ5cZ64yO+CAgBY461rXa/336ZOFMG/UZOqfV8KqsZ+WSZ1pIShgo6Zc/
QKWjMtTES08PUCI8xl/oD/ZP9+o8N9pcX21nV2QOJR8PjfZdMM+gkBf1JAheElTe
tfMUFSSpb7ASZzovHSIZhFUcgjKYM1pFOvN7CoNLbOUoGCuViBqb0fGo4TNrIlbK
JQjAgxqsBt6D2W23H2p0Sp2fBFJGvjRPYMzgu5ysiwLib7kJcYv3Yzptq1rPQI9z
HcBpvM1vo/diZix6G5UWZGf/Sgph6s3FJXL2h/SYMn5jqlmHWjZB01QWA1Q2/T51
i3GKslmIccurd8wIWBU9/+kewTlUFWuR4H8Oy8nX8lv4BtIjlsGZcag8Ek9YSefL
Br/BvsS11YdbW5i2C6XXLBc2kAqdFjafs2ET7n3lxAG7jupeU2/3TiI5UWY0Pzk6
uMoFjM2L8193rvIxay3cb+fmPzHEnUoz7G9jsfxvvS3IljR5csi8Or5xKtBMAY9p
Kfm8iWnTlec6P0H4Xzpzl1Y/gheIQWkyk5vtGBefmnZzKAV0u3ApqfZDyQZ76fsU
/gWhLUdRilidmzLaWZp33Bcjk0mPjUz47mUMs6NdveFKDV00EdjmvpYyHwFy7InE
zwZwsYbsxH5qrao9E7viAlRZ0eA1Tg23/vn95ORMRVrkUuUIV32QpvIEPumHjVqN
C/YWYbmnuJYhfpJvyz+d8+n4okU3L7OOKTctD2x6bimmp6jit6mUtUcnCZyE6Jfu
4yoJ6EW/ablO6fagY25MONWwy5oiPgyLrFeEReyGykNsVivopBiN/gEjfwz3iXzD
Strz7CKG8da74z7p1osXeBruBQZ4/ynjn7M+4bxtBMyt5oy8+yf02PvJKV5wwMND
zdP76jnBCXE9WZk9lCSbQ8qtcCVC/OX5tanJcoVb4E4GIS3uEeut3UwzsA/2wMcQ
3ZBOyE1OQ0COKumuCfEq8vsq+kBEm6Q4oH6AjdJSLrXMi0oUrPGE8MDazHTMch2i
5svwJeLQLZOaPK6dwLjHdDxV64URNEK3oF98njWqm1oQDXAzgpZQ/J+a53g8n4F+
fexCwTQM9Tyt2NytIqZZZoycnFhLPUFgK+EHoB9qht+sebmuagntiVmP4SkmbbY/
Nu/1SjpUty+r80Boa2h8Jn4EdFkudkL7SZ38ZQHOCXLqvl3PiScFVxALTQw4Y4z7
k8uF1/xMtYpLkQRup1Y6xNcGk70D/bM9/3r2du2um1yBepa79Ot90xB11wrqGAK0
iJUB25g9iyrpqGdDJM+2bYvASa2MvPWuZUHXxDbJmh0NHQr+GRDshAggKYMOdD9y
tMcd3dJh+0QQLnHTdOFlclaau3AI+Vw1EJzGN4Z9le5tjFCwzOxVmmsYz1LvoCxm
L5ufYU5MIIC5niNJjjwtRqvLYn3oIIieS4hJNqwgoLYZYIuyI+KzbHzPgGNaW+oq
LYgvNNbydsyaFZEXRemNxR8cBwui0fkbiiBP67RBPWtbdkk4W3raSkkSpMSerhiA
q4dYzqcPoSuf+9UktHG0cXVwjQHMDNcBcFCSmenEOIEgDa3voPdPWwnvb/0M+z/a
2mZ3Nr0N0/QYDtaIqe0/kGgyX4x9GTTUceR1OAHbxlJYTTW8nANUW27XVnx20Glk
5KLEkrngUiTWdOW4Eg2LA4sUCpsRiXxQPhUsF+PVDS3diN7QyS9Wq5KHhB1/wma0
oDLcyV1htsj3gyJrnsNq5C4fQ3p2OFfO43+3d6AU2Fk8puwZ/TErcRS4r9jmbxzr
3u+GrNQ99RQ6P0vYrHGROeWjEfOgYYc9uA3ge5/Q9Eh9CBKax9zWNflR5M1zikQx
neoQjKx7ITsoWlthRCoIg+syXMH+r7FuJONmUCoN3mfvwtEbtDnAOg0Vy3s79wc+
nGizo9oDDdPIp8kSdML2HwaXgNAf4LFzhPDUeJFsHOusoWE3s2h9rGLyKwKCPoNk
JnYfOWORcyCFXlwacyZlzN7/VWmbMhLggcW4roM7ythDs1pUhJp8yH8TT46XDQox
82d68PFvbUYr87vDqA0Me3clG4ZDkEmjP7kU2s1JCsv5r1Jvc4dSMfwAkNunLt96
rmOUdDWGk6XPX5LKp3gTERmP4c4xjz0+JWz2CpTwCMKjWpjurKtxWHEBEgCvAkfA
B/KRPAAWLM2S0b13KwsFERr9jcFRHw1mMNjqdrsVOUrQOQYsNp4fucG/IM92DlXl
9J+f6F9eM9RpJz5uoK3Jp/PEmen2UZ8IgEeVkbqg86M5XrMtTIJ5meqmWx68OVNI
p5LATJa6cHTv32uar2J6rEpfocvTrdea7IZzfT9bJMAXE1q13pE7wFPwTcwOBdDy
6Y/5AveyEZq1qx5KanLn+Y9CRNGGW6Gr7MUsLWVA/Fk55JJjpgnSgGHwWOZ8GFH0
ZfPhvyujtSx5LhKHkRN6Tmhw3HqrvZRpFY+V77wT0K4KSjq+6CZPPkpg+VghN3F9
rka0e+8vSeRPJtmg6E337YtxV0ezk+2+nb6V+KGYMbWPSSosViBmPYhoAnF93OPM
YrlXHBhrZGvU/88AK+kAb4u60AWdRQ+0ewGMnpkh4j+hVBSQpzdiKFJ38CUX70Tm
XAuo/8bRGZruVDDlmcm4beH0ZvQ0z7b3DOOsJsbmycMNdq7gjVu/h5gkUTdV/tT4
FEY0SCW3QWUYvALLVUGlvemQKgDshgj5hcgFgTrbYU+14BdR55Yc6ZNLZvd/+krj
M752y33p/4x21wwotcdGTjK7owfFNow0naiJD/SgnRYX9cI9N0RwQlHU1jMflhmN
meK9vFNYawnPyU6JJxyozwUcXpk9vw1PLqINJjAKsattS6HXKspKxYtliN6ITF3+
3UWB83CFzzRH0U+0hYkilxLIKeIufMUn0fgTC7my05MxuxXC7mWrkqNf4zGgPud6
6ctcleiyX1Iiz2EwsZ6yVNf1ol24TZgvrAK2HX2pWF412VdIr6avVnLPH+RsT02+
JTkm6+3HqUC8e70dL8OREPLDnirQgJRpdb106OtbSTx4bChx48kivdhEfvYYGyPm
rBWE/2ia82dakmeY7noYgTbI4SMBjiZhCM7mHJOqr3/cTTwtjI1958obPmg4xkOG
+vTgtcDIQk6tFkr6UJ7XHv7PwLcr1gD7996HPFl/RaFzWvKXmX12I9rCn7AWcEyL
2mQ6aB6CPdlrnanPyPeTQ0xOlG2xD9skiOPspgxssi8lQLiilu6i3uo8bEJeFWML
RwR5VNUsEEluFkQLoQxKo4JsIeHpYqKU6qf3rIs8g5jEsQhHX2AcPmD7y2RgIHGo
aALLg0n51EZF9BCmiEzVQYRYleO9cO6XZMoyuapoilH0c2A0En8vI1swREbdeiI5
YhUgaCLkx1ZkGQ7VxoA32IJDYduvksh1g1zRSVHPLDNMO9eJmurJYFUQNdsOfuHr
MompRpRbIyX4INxF3sEQKyLVZbOHr4ILvpYFoJK66d8h66k6Ps6ancktMrXHQ6Cw
LQQgnt8Y8t6YJ3S4KXKFMqtZais3Ng7LO7iWCLq4lKmIFNy9VMJPh+sHsAvHngYc
0jKd3iAPaULB6aIp5F9Q2bO9EaBTBJ/8buDtiD6o+/hl/RGzBE+GLzaqtdy9nYWU
GuY8G1qgio8Y4/anhK8bMmnE+U1ZxSGOS92qKAztrBUkYonvd0m62/jL2fBwEKmK
b46EVIhuL74ImVDMfaBtuDRvXRE3NFn9tVUaPmlb//eaxLPRb2b0xDCuMZmHNDYx
vLOWoYQPALzFPW5hN3KNjHzIPeh61Kxy9MeeN2o+LlS4rM/uKIXZRukwxs6zyLSK
YlxeOADSIr6JtpKyNL/2vkzpH+OFoVXB7ZtA0b10h7RI5YbTU4NyaEGMSxKbDhz4
+whS1f1i7BqwhQk2oymkBnwzzYJ4gXpx1KwM/C0er6+rxda7uCWfPy04a4Uav0Qe
qeW4Sn/RB7NYps5fl0mWFKAVrmDprImcVV+mqGXpGQi7nOS2ZaaomwKH0O+QV5GI
SvdtG7AfueNggBgATVOhc1YgWctrAlywyefZtZ0QqlmGo35gszfzAGLeT5TZp2y7
sFXlSmOSeq64FSTlcVH8bOmeLPYWfKLL8sEb9a7XuSZks0cUoy2y56NC8zTF0lvv
GzZjy65h9WyV9KX4D2ixnVCRjxgnmTBQzpIaU4lSyK//E2boJ4uMYy2o04pHltBN
laJKia8seMWpBnx3GEeXwH9qdG7j+jQxKY0lcFSeVQtMIk5wQWQm3IbRAGyQiuB/
HEU1rj93tPCA8W7yLWB24Mseg7r0q/rCXrtBTNqZlhOo9vol6BUj1xZrsZL0aZru
GcQeruxdEW0C/Ki+E3EMP7wIKbL4pk7Ywob7U38E7VAZ7/OP4tHl+Hlo+QS8v4Et
wJJa1ESf+0siQnx1XGnHbTZ5CBaIkeAkK5WjoYN0VYLFSUXDoul/X2Bp81P2CGNy
EPlSnixhKgIcimS2OjRhineTctmznLJXlH1vIjVn3UGyCx5wCbe46Svb9W4respE
df029X6VbkBHspxCfWDkURh9xLanOMUWaYsui+6bf6r47iHqQgLydj+0b6ax+1Kg
PVNuoLks+ZbpzZ2hxqtIywiZre1XV1bkEAF0K86ufl3SzTULVrjykRPvxwJ7cs4i
xFynoQOkk0C8VJDyDk8GGW9FX7hRB6weCO9LcA9flKYJhb0ePgX5EZwEFHu55CUC
8M+OTzYrskqWxy74wKcov29RXXpsZNAVL8/P8GCpPSsJgjFdkafyWZsTNgHvRzux
Du8FvV4T7ZSjtAut8EAQVNFbBd+t8o0XOXBjuVkuO3Vd8SrWX5vDid66dg4ZP6Xh
6RljMQdahWY3EiBTzu228SdQ/hqr0QvXFrFvkvw7qVaIb3rm+Pe6ZcwxJG9L7V4l
OrBvN0vtw4tQC2PRtmuerhcSU7f9oKu0dkV1A/MdxjNzWsOOz+3X0SbVvUqfsdlc
aKUX41B/Eipq48Mv8VIsbPK9dueAYcyyhxpsYzSgPthinI1DocI2d6Zw0jIzGtsH
rOYL2XZtYsqJuoOV9ddSQ1jJydo9JC6f7YEdRyjsaMtX1wUK7gG1x9TrdvRE9mjc
6KocJsu9WF2xzdBc3kZbxHb/KyT2ABa7U/RNixhBM3thIJfyM0vwRtrafP9KY+hV
9M+FxpjSmhV+wodU1wAwF9V/gNH96fm76VrG8rrdZcoUp2kBJrQvVtgUsxg6tZA8
D2Zq3xGZiukzuDW/M9fGRkEvl52x4RrYT8Jxpy6IKE4SCJG5CS5MXtka2KF5wzpW
/CaQq5yDD4f+419nurKkW0zkUSAkE4RPQQgJdS3hUFYcS3IzApXoLuAznFAQfT2T
P1Dc+bw2dedeuqupKZ5/ls+MDMg+npYCCdBGP/L9kZurI85iz5rrDei6DJlMTKMI
xanOPz0daB/11/r+EZ5TotMffF2w/ALl8meSodwBv9E0xp49KGlj/dZybnpB9ybS
K5AXUdUQf27matXLV/c368G/vswiHrdNoymBiGhkELEO31iD6lAexV65OdIKQVnh
6yHkMXkCV9O94OIBS++ZETeYfkV8SYDLa/etWYUwC8IvuibbkwT4OByK0at7u+5v
nzdUWjMCKE4xxjMIEz9x9XwBEQekJaNPZSA7dm4TB9RwiqSFU1fcWH+D2yS5SWvV
I4kugBAYkcviMufFg4UAkiiqs1tjioUTC9BSK5TMJEsgcaLf7lOMfZl8QrupnjJV
y5jQuvAUVGyshlQhXHmQorEuG5vS0SLt7Lbx7Q43bt1W9RikcXWaZKo6L9w3aN9u
UeZgIn+8leQG/fVREoEmwUVa8mzpI48ie6ANyNtY0QPh89p17EddfCNFo3nTuT1O
zK3Bm6Si9Pj9Pbg+e80pMdctRGFWEys/q2YUz2xi7X6ccxqc1rBg58O7TVBHPs69
CkT15d13aUTO5YuxDBrNHt7wPyVw/O9nIMiIVVGMcln+o+jZcMCcDX1qnnnXDClQ
B74BlAOg5CdNpQUBZ/DUJ4aeKKV3sC7SpkDZchN7RVw6d3y8MA2+ZSGdabS3XsfY
D1rUsUmmWym5bxYcW4YusubG7fFQY9TGN+csZUXJtQp6Tb9fwui+o38zGLp4/opN
BSZpKoAk1+GvoZeTtwzx4SH2UOrkXcauGFaFbmijpk0LOe1J4tmcCz1F9MX852Jx
J1bPZsF7ZmJA1RgfWCCQc8GrEgYFxNn3/JmkCdLSJRUGjKtsK2jCJLaChjcaMn+M
KUXjzL68Fis2CR7VUdKy3A6GwOMVoKI/eVS56PSYUJYQeNd7dlZG07FCc1rMQOq9
M5XR83hNCwWVHFz8BY0dIZOoydGYrXdaqydfz60dVnPxqeIFynTDvuu6NHmNUWEF
T46JxlnzU/K4NKe1L+5J+d+h7DRyQFqZe0VvlSzuvVBR4tSz1sOAJxhb9O/YVSmy
FRGYH735LI+VjKa87iU+AJvqMUHCRxItOlX19umVct/0CP3pZylznbpDHHJAO7+d
TjTlaw1VbKfMgc8VzTV5vLk08coRdmr7kf8WCgUNnekWiez8RbESK4EnRAmOtAe1
kyrIYXdViUq3vAMmZWrIjsskx/ZXhL48c7jHAeGJxp21Dj0VtbESi2qArZXNm+qj
IYvMcRti8Ej4avPOrz/OgJZ/cI3BErnEzTeZDuo04Tz7722WXOipCjm4IUqu/UTO
naXgn+C/gz9eXoW6BZtEXQIk5HwcMgaBvV9kPjNzNlDMw/Zb6NnBH2TwrIRoZsto
GewJ8yxbW6nDVrzFdATa9Audu5AuJC9WBCkOPLNGzSNZCEKXUJr9vTFUnD6zyh0d
7praLN1pgWhf9+MGday/Rr19HU+nRGrwye9reMkeDQ/5QG5J2VM3vFpGi7pMFDJN
drsajDeMg5mbTnQfAt3Ad/1QkPYUSB8NYE8ZnOgXHYKzKMhXtfWWF2qbVs9HanId
J4qlao5o6hWMThFxH/QZRT7xgFUr80MT1/dptwppk+yayJT1ep2VESnlHaJLNuqR
1em7g3qIgKTk1qiSn0KLIBlzBmFglmHcYYglj2UC2hp3NHXCvc24xNlJJ3dDXiLc
OrbjM45U6ClKa6H3DXtGfOel1U4RLtyBHssiZh22KxXjXmnEBh6INwnxDvZijTd0
rX802r4BbX3j8lhetbh/rcsS71CHUKEjaCnmC4iFzoVKuAluPf6vhRsAsS95IO/w
3p2fkK/cG8/WAIncSfZeEXiSd09HiJ/a4qOjLogr6yAdBYsac0pSWvZA2cHCY6Er
hMCyVx+G42dLEfGpvnOxrVZxARldBcXrW5yoSjNx0t/NIl2BR7aad2zvYX3pNnUY
tcGSGKXQUqUeJZRZM25OC/ToHe3PGv/5sxZZV8OoZBeIxeEJTu0uIEFO9WhuYuO4
I+PIUysoLJ0sz/joKYdWL8nkF5EfI2H76u9TspvNB6RpxogyYqDeWwXKcQMAnSSY
Mz2vG/g+dclVycB8w7q449o+3c3wvSdS1nnwAEXTPG4EG6WXt5VQ4HsaBNICOkr8
E4msY4CReVs2pibTTZoiPXlAbibS9lmp/eO6Yjw0qZt0FgCdK8/I1fjlFkbYV4A+
pb+0GADlAyIBsNDdupW7dK0B4R7Hnoe7DcilbZZarMlh27fOLdiKVDJ4diXW9CvN
D9kooe2TZhI/LqjWhxBQUe1CLoY2ldPfHzHTUHHnTmmYzxcy7som9CmYVa7rMaCo
FNVZuE8MxhnyRbRyL+Xsop0jkp73m0Bxl3rdu0+JsAiPhcgOkItgNxqUQT3pMV2B
XTmBleI0AYlUYLvrIpg3/2AOmH8+cB08lrVKQX3uAAF8fjzEE5xT98aYjV2y5nrX
W9zg5myZfNf/INaQLAo+fkhAHdn60UZfosPgrB1NWZlB7G1xCM51LNH2BzR5fdKz
lhfUsYWRebAOL1twuMfOBOzhj8p63AvcrlH05AVqHDVhV05ntZRoL+s/QZkGqW5B
x9V7TgN6NzYV4XI8w+zD7+vWS5diZUDb+f/n6c81NH0rnfNwQjI17yCs0MWCRZCz
kEJ9FPyuDjAGXwUxF38CdrQWi2PJp5xD+V/YQ2aVInnZpQLTYJi5aXJZ3TiNCdXq
FZ6SHg4Yd5mZfnnarvs30oYZ8H00Ip1DYnUISNAkavutTAgImnKpXepZxz0+MtqL
kZ3f66Zg6K4NgSMzO+LfUHZeWfOC8k68EOehHf8H9GhC0M+TEW87ZdFRibrWCcJD
aySvfyBlIhRqyLVBdsnEPQW2afD8xBYqFhUyQrxzAuyy1/yNmNzWm1vPxgrPJKSz
MP4G77NpwHwYhi+6vetjczqHpxSIPdta5NSsH6qKYKk6z4HVPfjAA+Bu3I609jua
Zc3bLsnDVjb9BKscKJsAaJYMJfqzewfxCZz4tXvzS+97NdrwpJsmxmxRkzHEvXTA
kwYEscp+nkLdXtcx19bGiUmm2sbou1YwWbo0iUXKudx6S22eXOilsfWt6OhBtTkh
p8dFi3jBStqO5UczUwGBfCk+U5HmKKIVFbwlEoXKA1FH5dWk494knIMwBocDJElC
lu+81m9gT8TA0ecEMYX3UUnUtLtes1cZ2j5+uu9h1/0Xf1Ys42x43YOAA7atj0WF
54Gahj0F/NeGx2PCkg3qxdAITFfAtxx74wnyhoHd7PT9DmTeUdxcd/J6wkiF237H
KptJktAjIdRk3pCsPwk+cveeLgTXALC1ub1JUJt2g1vanfPretxfORy/3O4z5FTC
IoDqalJv3wRrCjrE6hA4vA5ONismz+4ajB6hbjby70+VbWTtqSvDDBG8tPjL8EV2
qLyqeLLf38gmTsesWycLcCTeGPxKs95H/Ovkd/9S3hoEVdeVBD4aS0g17LU9Jsgq
q1vW4+czXuDE0O9gKYzspmjw3atKUPWwzeka2k0iWw1uwRc5//O5n6FbQmozeYcq
KPQAMeas3+PgWlEbA1YJmj2V8MgYahYAIsPZY+iBN0KAhtU9IbpQEVBYQbZjsOfF
f4pN2S9NWAXeAknzh9aiOzW7r2MCGkIrCVzskBo1OW8peZePBgEJbkQ2WeSRUZUa
8nKy+7BWZiCD7Odw3bZq09Xg9mbzlXOyWeyvQ8sS5Qy06WlFI+aZY4kpQsZlpQdH
FcKsRSK0FYWtJZtzQ936rVM7+1EPYj0mIZw1mXdqcwmezoWn8Pc/JpPT87ekm1y8
YxTcvYwnX0RH/h3dJ8LVRSztGetND557iffqtPtTQm/VHOsKHLtuQmfiWuR/3dFI
/olPBcAW4ZsSoGAAyicto9puERwXyRfhHTd37v2qeWt3SkOLUBCBfY5XEO3u9kEU
sv/K6H1yatCbcojtrheEJDs7BUczG+/o/DcvAhl93WbYvLOVCcz0fmLgGet9pVz0
ALYB8xKYCGqGZsUwd+ND7oKq2SqmtyITrGtEeDOqC1Jb/pv5qMJHOiPLC0TcHvND
xuo0rhF1amxWEPEuQSQmvBpsxIN77VdsgyiYHwDv40vI4dcRiJrtUGmGfeNjqUpj
VmdgL6LC/YCi4nRuFlWQFlh5iOm248DBYsHfkwyC/foqKEPe+fSlrjtK6oB4uDRV
Wsm8TaiaSVlQwCRxsmsq7DN7YRd6kfCaSEjWhk2cphVnq8+g7iI1KPDr/6ySvMoy
DrteKKhvUIcU8jQ1B+KL1cxiRGSSP0+MBnACyWMvpJIGg/sdzaZYwCJ7vCHS0QK0
X+jkChC+P+u1SwWpT8sP4ERsQAfzsFxXSwQCv1oVwiLrUxLT4yfRAvpJQIHMNT3J
9V5OEYe7o3ImvmHZaCAhJ5EbC0jc8sPPoHisVS3TH7I5cjuRbhrDlGxpFrMib/w1
HEc9n3Lk8vaLZyBlsDK6BMdhoDNBc5tZfYsWA2QCSyDiuT1N1eb6aBnp5AB6u9Ry
cVdzRLM3DOe0rhw6xeVaa17RcMRHmu3AaSx6sD2uNCADHcczCuzWP0iWbcgjefJv
kAv1tz2gEqNiiGVPvjgnqLiNGGQl60jmp449VbT/fq5J98FZuEAxuaAo5sIwRcXp
ApH7Le4J7ZGYqkDYB2OdyOZp2JtkcnUYlYZIagykVSLvyf9DqG9mowHIHeLZoenn
kvDh7Ss0hAUD3SV3V46AKM1AuOT5emRfubblmfDcLji5TWqrwBscM2gkcCj9Ms/s
34Z6sps5d/V4UM1PzQVLRzTkkYMPXw5JH8LIaVNrBpxn/iKCCiaJIat/hQ53N4HG
xpwNU7+eBTmr847wb2n9U/P1p/BIEVnNIgGbkFGf6pkoBZrM/aOVQjw/orAHO5kd
GOsW6/HSa/Qx/MVw1bGg8OlqSZexnmoiih6uRWY8AexSkySHygd217MtDrE6rI9A
XhrGNOyH8OQT+bagZXnqupuqee148IXO1C6g+Avl78L+RoujJTWzZSe1r1Jd71+J
hiuzejgXdBP5TMAF79HD/NDf9iUxGQI8rnFP11nT6jM+jlxt3OLYMcoM6jTa61sg
EpPs5nuL1ykZpCg+0WqrEbkPnSlKPr6wOj60iKuyR/DYR3ZL54H0ZLb0XVd/krgM
qtKeNSNBjsgMZ0KTbkNklS3SF8TZ4MbVf4cTtmjIJ0r3/BZI67DJ4bSg6eL3V5Vt
8iR8Ww19lCdccedmfVuL8YpkP8Hij5pwBfgCX4/P7f2Xo9bAX5nd81EKhAXCdiEl
q2imjpBxkLmcebqTdXrDCJUxtIHTepN3zC6+15fhMbVeIMBfOvyN87m04BeQKy42
VvPcm76QhY+HxXtG47dmg9mLtxmUuFM9oolGD3TaRD2+5nH6lxOqR7mKi+N4l10I
T1l2xk1ayGc7Ib7ChvNGtl3tG6mTM1yode4GodGNP/GjupTLjC9sC56xO6VdIUpq
3MfxttksHwJZ6tNxerDLD3TdyyKtx1osvHu4H+Wz1ZHKY/1+VUmsAfJU3faW+PU0
ZOGc8qd4VhFMaHC5iR9qQu4TSukHU1ow/VcB3Oi8foADGxybnqqAu7SwhFpJwFHf
bjrTI0z6tCXRjk6bX6sMjCgN0l6YBm32sYPnRNJYlr5BZuxBZkc2aF2inI/lcy69
xN3OWhVZchfIPKUWvvXF4fmGyGppqsSZWQOwrQJ/XdmL4vgQgPZ0dJXpL2QrOVRz
nqMKxmpQ4olMUqzVzydFjPfE31bzQBwTbDqzzrkGk835YgR19SxOdqMzgVTWoves
uiT6nEEDsccW47hifypBlqPyaH0NtuYmIdEiv/hgWZ+C//jmW6sp2y1KSVxjZ5ip
/I9TXGsWxRV6QlKbTinloy4EOL+Aa/RPjy3jVlDcwpHvlUII3UIG4TmTnlk6e+BQ
cDbL5jnczy/zPd7Xr0AeeRec4Iz/rB+wWZWjNJDAQ0CTA58ZEHBlptNdbIYMpgGI
b46ncYT+YFp2LsY7HlJAyp1SxQoBMI22ewd9b0Aiogc2gojy01m9JCCivGYyP7Ae
1A/dy9i26YdQf+TYm5NZF7k3jQNEqI1h0HDwHES+11uMP3c6xtQ+lB9/W1QZmPne
9AY1f/n8qZsT1zE54ryCK0zj0UMUX6ov/gWBWLTKdZT7Ia5bQimmQVtQ41wy+u22
eG7R53CjTyGp4+XtIVO2vNL4qXFNKVI2abXwZJcjuq/2v625NUR+zkvmYVNBr/xY
A7XQKl8i/Fi/2tjPop8IChljhPcs07Oj8iqmth8oPrTUxfU2L7u5Jtwn1SbfWokR
yAvEOryBpC4cTy2kcww5HUC11bNCfmclFLIQG62MiuO+eqYySjndyYcH0CrB+pdM
Y58vKnKRHAI9FK0LJtMvIeAmgpEaXh864qX77V+D9MpZmEUELizS+SBn2nDP9NFz
SIVnnfC+zMlCU82VkrtVG1Na0JP6suS0TXXim57dfhYl7veD//TPAssU9AFRZhPz
WmK0FAbNOGDwxtjnMKgH22ikKMiM2KMxQUBbgqM4kOp5JU3vzPmIIE1Ab7Vkw4ar
dvaL/rL7fG2Ap7qXYn+8k5R6SDbhVM4SxQUFzwaWjN3iFL2jQro3dc/9v1mOsYKk
o3DFDgZuPMOYEf4ttd2Wye931lCFdenFo7S18nKUHomEj6s/b6lzIxTMB4nd/7kw
y5YmDZpoDJnn7H9T/FPmauM0SNHhVOeUOqsZntSDXAUTxr87oIsNx/SmLr+aNAvo
Rl0xgvsPz7SzhxbCtvZh9yHhfmZMF0Gr0zKtkFnGkKW9IN+KdtcQrofs/CUxthFY
/aFOeUFB+X/wVYpSVy18x+lkZPKXtMedrslmbnT8mMDwpXkXVj5HPXS9hCIPh/Bu
hDSQ6sHrG6hTWqJv7lXkevbn1rJ9JPtTU/bVkl5tNIJPZup80UNjqlP3UtR4ixeZ
Orjin2+mweDXS4EbUnqQ/mopk7wOw7cGpu06tHrkhNdixBodnoJ+kOUDBshlH4Jh
nYYKXelUvHOyWkdanJsR21RsOfVxMiKMmeNdGJKswuX5Eoi/oVPPA3EdC5/YB6P5
IHhnNQGtrxCgByOdij9ynti3uF8pB/84gVfYsj6GHaMIj4juXMeI2shUxV7EzCvV
7OTHrzhGgftl88KJYF2fE41oG4F16Uad11JtzU1Wdg/zJVIBgbLO1tG3E5IWcaa4
NQMFl7kr5WThCyiGFExBo9xFYtln5aUxYeUpkNZ6ft6/rmZIIlXYBGKg45l4ajy+
N8Vy+EgIaCi5LRu6QcY6zI0zvZaB/1r2yu9mCpA7CimbxA0eHOpInwg4RjFtVPmF
6No0XF/IblVg7LSgkmOTJBKQm6uAoskO7PqnYj+siGEju8gqb++uo1EuN0cBGtPk
yyZ1T/K9FDf8PsBB5ZUpVgeO/ofxzjwxFSDFdbmxis4rzbc3na9/MZ6iy1gJ6S6i
h+L+MqN+CFA1ploPJ8jhv3zs+ROtIW4MJdBxj60H2+7ObuSMALSfhs06K4UqObFw
3Fgv/ifsmpEflK4gcrXuiOJVEfujP/jui1ltbC0uTCN05sWdkOFrB5yWS0vPzPnr
znhfhBgGwTkKIi3U+YsZpjII6hT7C5GERyXfJUQDVNp7+1jKMsZIbd7q+WtI1Ucm
VmLCbmFSwsoZ+9n9lkLRjJD8ysjzFaowOVUYC4Mao2f5fIV+Go1onrTocyfallV8
WoRAJidk5Myt32kfMAtnsie9yS5bFyATGep1Ctj3Y8C6RvUuPrGKNAxFLkoeR4Mz
IyVg3ADd1ssaFwhdtXOlQBU/mCsAHravaERMZB772yfVHSsEI1iprp/6q1A+DC1Y
lyYvtKiMBalXTfGFkmLtiYcAiyZYzUHDo96SHQVOFzBOYQ1v+9niZqAZru9a15mP
2YD5kE7B92PAJT+tXbAXACCGJlOUHA83O/Yo/eLDFmyzk+7R7inLRw5I4+1RqaLE
evXYauu9yvw1YWFoQQQr+r/Md9KzJ8dM61d7CitmDKx0W++E5y4Mp4Zmz2fGHPeA
UgnbB1l74NyiBRoPwauGEr4fozWWPwtf6uxTy05YJadixB0txCjpzGnEQlzh8DFB
wD5GPosSbmMno6FNtuqNqD6Xb/CLxfu45ntf5x/q7qi6XC0/wHR9WsGNmKprMEQR
BKRNRJYP4oXHMpEexGBrHlt392E3bWYR5kmh2y82AYhJS8cudlYaotDo9ov2tCgp
XmnMH007yVAHkiOhc5YVv0brkZQXk9jFryb9Zg3TbxdL+YhWMwAN51jpVQsA1WnG
jSD2qj2n1NuduL373jQCiZIB8rS5m1bOw0RKUCDfbpdJz2ogFyzqrfYwtw85Nxso
GKQjWqyXaU0amQ9baKgM9sJv51GtKf0czFfvI3bsDFZUNxCKZP/E9O01Pyu4/AYK
wrnY3SJgrG5hYIoC4QlWk5E9l9t0vLexIe7GerroomTXWvPHNAysFx/tzaFvSapt
7B6j4BlzmnX93tvAJuVbv6RoeogxIEQBAbJcqH6RvWzO5Wx3ibqSev2rxMUOubGG
LGY0+Cbmu59bYS6lQWT6flldZI+4Syw6Kao2rh1fRzFH+/igXwQR5m8mHTFAr+nX
LB/yHtutpMuB3HDrth4bnctbXC502EhjY434bgP4L+U4iHROALGHeBqO//1+xDis
q1RSnJo/8xzakkLNt/PPI1AfCdVFuXKv5/nvQ/u8lBfERY+vSQJ3r7eI1VGxgsUH
JspA9c4rRtMrIu408XwDo+6liDOKwrt1QBWEsXAMNnF5h79k8BOk1Zd7UjPkG2zw
/PYbEE82IjJjHFEeTht4rV5X1FCNUl2mVB2OGOjQDw9N9Z4QHsHEENibS0qA3mSX
dnFfeXIo/TiWvF38LsGjhNLXRRc03mCgBYekxjrk9aYxdOVPiUj9bmuIB0cGfTj1
oOazBxU1L7wPU4leIb0QwijJveRFnysJ4We3pMn/HpO7dQXDqPe5gmMehRcErTTI
O21tlNdxKdXy+PteNg9Ze8OVGHeJoQ4CDYEQLCJvuCdWv9nBXbFiDLUERMrgppoE
WTLTNpvAEXjSp5f6B11NNtMXB1YXnvrIovCITCKImwrFL2nxHzVJQ5bUxqfdcXK+
JR19JQyL8wZ5HjeNfpMN7FBacnrUgaza+rqgHP25t+ncXeVaPQxpL0Aioi/AjEhZ
dflrRaLIPSN+rfhpnbJ+ojTimDWeIhljHzrPLCzjZldOagb9ZMlEKvbVnbfZOPWH
chToI7XDnF86H+oJ75ZpvS6hq7DoPrOrDHUodvEnkHQpDK3fFQQpOQGj3leK3PSz
hRkPNASTnJXEe6lYA2VqX+ashvO1ko/T/S18AW7nKg5UAsntkXs6HxaXkBtNcgMY
BKRCEIdFQ5jFVuElKmdYF1hrlF5NFj+hLO4RzgegPgBZ//rJ+91EtG/OHZvST2we
N8qJPs2gfF8uToW2wdmvpSFMsZigLBKBFXQSMrUEhN9Dnqz9IrwkB3qd58QS8Jar
5hQls/rsJ6COXvM1sk8HzTG/w6uWud4jfOfO2AXPVAmbtY1s3Fnu1qzxNQL4Z/Ar
/acg3gAVTAozRuX0PD9RHdaJZox9rdeM55sUsO+TC8xdPC3nG2JusKrmNAiTM5Ju
A+QlbESALtNW5HO8golpV0Kzb5M3H6ASkNEjRxBLHxmDjkHZwqA9RSFm8EAbbRGM
YFYDUOnbVH9QGiy+iCPf9VU/J6oPRixksFui7Yr6XzD/rVmmMsAfECt6vO5O1GaR
hyeG1iNyQ8f1mSVvqi5EYS9Fngq41y6a86x5/nNyFqI84XgAPgYZ8nJTwkmnDr7S
dZANe91Qaa37/5qmL/230FrMzbH/yh+OONijQMaF0QjxoRLz5FUrLJiaARZntRmX
MU9UopFLVgVjA+Bs11+ErJzHr2/wGUir/IY/zdns2u+XoGMqJAJ9x0wxO5/2GL1f
+6MG3PNBZFR+LkZGuHqWRD8Vu0ntfGTkW/giw3A1JafI6SVZvCIuJGjc+gvkB3RL
RN3+/ZzUdmiBEBgH2Snjv7j4BN16LeQN/nuU5j3I3o6ExmZpkHT217K0efZMHbje
oopf0FTkyIDmCF4TYmIUyep2S30EIHCvinZKc8WI1+cAsTDeYpY1GcScqnKNlgwU
csZhoEr9Jk3OuE0hSqM83THfr3n/9qUrg9y1Eo9Z+Fn+xLyDdxAqyc7qOtisEDeM
sB7mJOo1MPg4sSX81lMj06FNRawGrIRwkKIgK/vIThP/OFxHfbyUgAuae/RN6UGd
NM88u8RT7hpMWuSCHGjeCBR9oH0Db4hqLWaWAbpBZUfo7uO2aKylUw7e50rFWzNe
xImwzJHVALAVdoVYqosLq/32A1Z/3ZhoPVQj63G36zK2Hws7EviLM/go1xZAAhC3
TK2dhGsNfJ2eCddvijfqHsxk25dQvjn5d1AyAFy4mAiq8RAfcHCXVvHVvm+w+0hf
OFxQ9mTGainzvU6fm2/oCSWKJ5yiENW5+DJSbk1dviBIbMuTcsDOC4JLHrOE03Jq
EFZ7qQsOXK5YgAGf7LeKPnL3BTNzYDEuca5dfllGGTlUXAvR+vhpnpxM9B0WYm9F
3irbxJxPbmylbJjp60wNLSAUo2WMmBNUuGD6bMdbwu100/LMjlQ70KCUuBpwm0Hq
grGSDQ7WLf0BvJHo24FHfTXJa9nxf4F0SVWwzEYprK7eHKDjlClx8N2n1bkOlgL5
plci0H4MKKx6WdqMAlxYfTnjmAF1ersETOaDdurY0UJu5srEk8silVlCPpv4Qep/
9I6gu1Hetzz/bE9Nx4wVXfl4HPI8gRDByMhiTole9q2ek1DUyhyOL0/Z0QXqHqIJ
fLpUu6qbt60MKgI17+ebhgB/BWcbtsL0R1RZhcWn+6x0iSLQnFEFif+t39t5JUN0
9+PHJw4yoTV5umWBi+i9FPcd2H39IntHO/f4PWzj0VsQCBTZiOxk0A7IBbT7THmn
sqeWe7t5elvqpPy5ny1NZmPgTc6JThiR+rreEOuPdleZAJC6/Vv04qFV3homy/Yy
dQIAoyFdNdfo7wiHyF6Y5NHjiFWHC7jFzz1Bx/sEJtJagW2dmDUv344ZmdMSPeQZ
KACei7xb2hozcWazaoOXhROl9vmqk6IeWSMWD0zHS8PLxYs91cl3AzZl7jmkVBxT
OrlV2CtcGD/xtXjCo+maiH2uWTniAp1EZ27mNYUkoSsgbVUnj2lgih4ZqrNHyBpf
1R8esKL0OXTGraPpokeMf5Sa2YfISGjoBF5sOO+Q5xYa6phAcm7GXA1mZDjuH8t8
TqMOmfZZimHSbUAa2sZ1WCwK1+qCntjl8gtruZcnIkfAlH+ALM6uSiyEIP5zdD9l
QQE94ukr1n+hlzm0KMc4YJL7AAF6JrWR2BSnRh1+PzrBdzFlE6DW08y1tY1/4m8T
taVMs0Brzoom9HMyzYKiJb13/0OGxC06hOyY8CpTewdPVdR9uOnoYiIJcfWS2hiv
WZaqQdUl33oCtZAh5t/aOXa53Vlta/3/HJ1659EXqntFGNnMAC8ku+eQI1Dn43BZ
BcI861Dq3t0daeoC/2cejAOJzRuQoPXijFHiYqE5GRXZt+OROvxDSxo+MFp30dCv
8ICUYYwIaI5MrDT7vICmcNf64aghROkH2LuZX//uIaloaQYEh7bywoTteRHpjXGc
w4IhQ4nfeMkx2k+7uO8JBon8cIX1b0Jjp/JTdSstxCRIyOHGFtSjc9/XLt+7YO5I
orcNiyCDKXQA/43PQbEYfW6b73mi1RbxY7741oGClZF9JPvza8z5dZocNdp99yKG
FjJDUIQf77Xo2LT21RdkzlNQWDwIr/U4JAJS2uG1GoY3cBuljC25pkeDHwGaF53c
J9qh7O326HXPNlz9dgERrS5tbWFLrednk4eeLoThL+WI8CX0E/2KXIXfECOnxKe1
gpPqrpVR6CN61oFVV8dIJDzp44bV/wrkI5AJ5tPLdxPHmcd1/kF6LiTmH/Tfysnd
3vvcxY4OnvODzyKWAgEgd309Zv22h25DC/E3mdbZ10Z+wPg8bfMB77hDnfUDilne
qe26MOZaSDvpt/ZcFHhQJ/W12/8G9MZ8mIbhaGwj5VlkQIfd22Ekdgj7YYqxvRbp
Zo0Cb8LHnCZpGMJfC+veiCwzkqVO6orf8E1aCvVILUKuFfCCwwp4GWhYiksQV/mU
GPOm6wLVB1oRHU1M+7G0nq2Cz0DLUKl89RKNQ13IAPy4Lg+KcIs1CBFkBFKjTwwK
cmVjfZG2Bc65vGVUkw5IDZ7E9YyoMTi9jRhuo7Gz61mpHBLRfe9N3x7hg0em/uJt
uqzKGjsjf3cStMNLOizWrwKdwxr465EcgxJDVc66h8IcJT/1Garuzto4UfmHWrBq
A3J60ZI4VmzYEvzK8nZM2J7gpVmxSTquUT8ciKwxRSO1cc6Zz1s4xiBhfBYEovUX
XYVi5Hrbx7j4KUQ6HrnkNz/TQAR/vgB/QOd+IgtMJbUtljiAKj0An2FCUnkDWRjY
HkyJcTxBeMQiQ/iz4GEQFj0oVMqvo8769Q3vKReLLPs9NNjYXox1b6pJThuUGdM4
dR+KlfJy66BLbKowKRClb4k68ADkAWCGfZQHbMCnbZpx2WC0gqRv96Wj0bTAPWoF
ctOOY3AZ/4IIzsw/UgLZcgs9Nk7/kBUGBsP1gxkhjBUibWgPNWKR7qR2aNJEVo/9
ZQliJk8zJ8akghKXIa6Xt0aNOVC7JEwsjgTdKkEh2Jn+s8H31VDRZuHdxI5zI1px
HEOcsH1EG3qdZ7RC1+IGzObJkRe9SKkkDzSuSCUOIphAcKO4W4K6e4iDlgVZ0fwy
bJDhBE2VtbuJIqrmI2QsJE0MVODBks0FDZFGtBQe/P/ml/JNnzzgkqzOD8Glk2wq
DYK7Jfy3XLFOWhQon0qzs3gDnNlNeOpSUEt0oS7iBb+orSEHN1b7vZXvy3L1Uc3g
e+7EnGRWQZ/lxBWsVya+Stpsxx3+Xls+0i/7hwYLViCyiwoMkb92qEhoOTzQDa6Z
It6g+5ZDWNF1F6nMXnO07SzoSaKv8o8ygHClhQ0W2PekaoZUJBl+SfnqsOISsFtS
22beIK+qtLFURZTCuZ/474T6mbgz1ZMLZsuBfvy3yyOQFHJ6gpyq/e5SdbeGj6L2
eaeK9ZgI9IYKnRKRWgxyeuUVYX1M4tuMMbGZoLvg2MI5pZFCQnpBis8XLEI9Zby5
AOgjMXhgoqKsha2GMg3CSg6wIPrM3nFS65gZXpCBWsf9qno8mC2pqejSf56Mdl/I
l4HDsRXB+5cI2qtaKseDdCwF68b2QyjC6hMFPdyxa0QFeaOR9ZwJCo4sUwf8q3F2
t/IEdKfSZVnfpaJpfekgVHc0/4y9qxtlmYuA4lkpf/fUvQmv1fkO5A8MxsYki2hq
vcw7TfKNYYkBbbVF0sOwsaYgD7f8p9NryybdnvTBq6aVGozmevBQdpIaKQctx4Rp
ElofCkgwEkwJYIIPJOlO2+w5+kWStR8ylMkoLUVLQKRRczqg7PsMBdMiYxdZN7rf
QZGUs21ouC3LFu8mbwrY/VLYZ9qePIkGoEUyKoOuX9fZ8VwJJ3JKRliNwLEg6Nwn
FREzRNiQzav2jlamMomT5XNPg3mMnV2ykwbl12LXAFtNE4/yvhWItLpqPcwypHfO
8KGbeH5YFugWjLo1Ppz6IYHiMc4At6OBRloPKJkTOoNoSHdBonQttfv5Sag2/9+L
CnPRyOs5K40HBjKlEqTVW9531OJXWBTgTkFN/asHzMUJL+wk0CwzD1carxL4DAPA
k7UG8tcqu1/EwjKsqZIEA2C188kIh66fxjKbPHyL/dF+bD7IRP/JAiTO613QeUIn
gzKU7uOJRHQPHIKj/0CeVLimUTeo+nkzGWwd20Q0wOH31gaWl/R3XRbBJYlnkHU/
wvkK+RcDMGtYCW1Fbb2YKHUmaBARvffQ6zdcyGtQpcbIc4bGHgbMbh0/2P3PGsOR
FOWD1IXTPdPNx5pE6QYnCZQgjuDmNSqLh0p1mlj6pdzAg+h4IJlt5XW+AaFHFRaB
MshBCNz5e0QjuF5CoORYz7F9DDOokULdvLCdTtBLXhgllcPcZHATUxh/46wlX48t
Tj3beJAMMbKgMWVe99UFmKT4WedGWjQ6BjuspGF2qlWaHHfeaDXRvrL1VBDz8Lr1
tSpBpWMHOtE6yr/1NfoUpab6NPEuilNSL4+TzrccmstC6P9Cr+2pLAQFx6Yv1usz
X7cKfSBn64vnqrCVk//PDPqtGjTiM3IlbizWF/bQ4rnwvSDW8/NtQBOvNoQYZGtl
jmUykyufiPQtttvvjfuI6ezGoLLqrE3XS888ZLGV0U0VkdU7Y72AGfQFFY9Te9ed
hwylYThrCQ4Y58DeWhY3/ONTZE+jToaW7eCQ6IxONgFbPBxcu9JZfyeSNhGW5vPL
i1emmNJNS34DcOOg/99ovqx1E8VI4pak0jMsB+GbTkZ3HaDTFgo8kuOtUy1gTwTl
kmor5K+kKfjsVQtDKQcKT4QxR6REzTOxnQDh0gdwgPdzijGvAGJBTC21xDmiqgcR
4ocWN0/0nMQaoc2M5OzGvlXpEmvRuTGsu3JjRBd+EXaylMlF/uDQcgGtkHodXQPN
oqckAiGutqxD4DvB8xtWrcHcnUh25rGn/9UlHrVp8yVpuKDDrm4UZyNois/Hq1DO
OwBK43kDV7j3+jPzBSYNKTMeqMKWgvi1pEhK59yO2gTBnjQpftBGSyL0mpcyRdIX
hrhfyPzIRW+2cIOUfE6xVT6ZOBpe4igeSWGrTJ+7WwJgs3EtWHOdzNSCNFkov7pv
38YmaXqggsG4hUPrkDZ80ilN81e1rkiklQD84K+m6UGBDIEk9nuNZfexcF97jnGD
QvWtoYtLP9LFAue95wu1X3dlSPuetr+1qajNgT+QfSJzkYcAFAhI4Uardla6tdsm
PpwrXgY1KsjsfBsBlLYcCbsjl/Ioicoe5tM/n5weKDgtvuE4NMCvhVY2C4/tGvFj
aYUpEO3Rcs2SvvbNcDbTXzMzeDxKcFxD82mh6nwT4KdZE831a7SvGhPbvMbsRLLn
T5BC4WwPufhqvWWszQdTFSb9cGEpg463D5Y4L8mqLO3RVBmrSejZflciQRFvs9uv
Pb87pMqkP0snU9VVF4R4nblXsOusUibFNwIQ4nWANDn5tyD7N02f3GDJAbS/0GED
PdyRKfrjmep5JbzRh/PlMiI6tY+RwSOv70cvvOR4GdfeaxjHTWNtoPROp+sSwhTp
NuK2qC1oDpFUmaFEsRfJYUfWImEvUdp7Suc3LZEbAGtcVAVivAxNKb1ZTyfeM+Ge
RX/rgRa7eGCiCHZaM4hwkA3cjg5VlxUA8WJwhOM4qbv0V7tNYKOFFIDHqynBUict
ae+Daz2KwYGo1CMn0KcTaNUM3L7TQgMID0QY9QZouxks5veBS2IJ9zVVbjWOuaZc
s/oDSnpKT7pTvlE/PCq6CEREt4VJfu1Hj0f6dt0YhS1Bn/Hrrd9zoVOGdC7gqZeH
jmZ1LTyci1ZHz5/vBvcngMM12VSLaqfro0z68d5BvhUvwBQwfs7jgefIea2iP97e
xFtCPQQu3AIC4cDdn39WLByHhTWvkGdCnt7xjQlBBqQ//p+7oaKsB95RWQUjg3rz
KWPjlhJd/qt98MGDUshBrkL5VnqG8VqR0/g2Ou4CACdlM2M3Wh0dp+CDY0w62qfG
dsIAgGdOt//htKXiMi1fw3fVFTCbfgL+RubjHzbhrMn0FxJdrr9oRwtd+Kd9jdsL
udu+E0LBHUNbqqhJTawY+MqndJvKlRIqcOsebcnqsuprodLcaKg8equp2FQo/p9Z
CznkIA2GQGcGqkjheRAU9fVNprNOS5uX4H+H92IFUy9ZbjvXqJv7GvFR6Kyvn2r7
nESn2l/+vCVv3VKZYgMOhSGkXdWN6XWfmTgLZFMhwGsCP2Usd4ByXA5Zz8BIQBB4
h2dXn31t/nEQoGtKBa4+ez58t27uvlcWl9Svo0ATkARRnsJA8BpDHxI+y2lB1dCc
bKeI/clGwqDsscNzrvgXFEvPOSjDbGw4DlYeqXURV3tJXYstFQuTqcw9c0HLwOEu
YBWmVp6HKfVUQoHsPYu/+Nj4sx3mkld+QYSEEsL+CGR9yD+qZJWtRo5n94eSQgHC
B27rV0+1gK8R8+MA9fv95l5yZOqgnbpClHNmlnXq6J4cIsNmvbaV6rrL90Z+gvQE
KNA+67UJI0qfWi9Q0xQ+TMw6qQwJlY0K3Z8v4Xec0mU2uFhudc9KMXyfzlzcmBUg
h8AX96aD84D/NPloBuvc8EDNBVeKKQ4Tqe6zdT4wsbSMmYGTRwa5MF9WxIe2pJ8N
jsRH9qtXwRKfCIL30Tnn2hDjBzK1hz0F/ZJFekELk4rcpSYas/0CJ7yLUAfytHYW
HBIk+Q9h8qIuAtBFErUsfb5wuUJ5NlqTyQ6BAedXtflCMFg+FnE6scDoJGNcCqdH
RJO5fif6sk2XQGoinoOQPACajvBrPjyHGR/hgvYjJHi6zvz0DB+G9mIr4PPUekKf
eaLUohHNxRyJvueEewY7IPD3l1Uwdu9XSQ0kecyA9txQ8SNWm/H0ipFjMtSbRPsW
WIpNG+4Etwpy2mU4b3X4Zvb1EGX9yNRZCEOsz42UQMgs83pA7lJ80KfjwNDLJliF
BeNXSVdn5S+lRB38Wzysgi2uMcj3ahv8CLn/FA6IKmt/fygohEG2TM2zlitYhSrS
Ibe8tb53SCUIBlucU1XTtGU209GdFR5OovR422h0OOy4tfsoabbHOpvty3TKzCl4
z+h9L+v9UMbYCOILTtdr1WEeyCD4r8WVIJ4l2Aayrf/LyrR696x+0zNbffS28//U
KJjpxsJ23iiV+wBmi8XUcAOmYRAKuL4jITRlfVU8UZyLiUmnvU9xc71OJOfFeKjj
CKTY/l1OkvxS3XpAJ8y/tbma1O3wScK4YuODFl1J0K5vO+/Zzbgitc917OIfoU1r
C3ZvTWu9dne2UqvuyTh4uKG/wwIaC+IyHmz5qjXfdZsFAMbC4/dnuP/+y8G7QFY6
50mXylzAAs0yPQqbto9tSL/E4xV+mICY1of8xGsR+cmD3biDzUSqXOLO5OyZDn3a
BPiJFuKKZcm1kSW4TS9u+aYSw8sKol/4Lw/2cUWSoOLDtBPaKvF0HWYFClTbebMn
ZCG7eTuZT2h6n7BJivSxRzKrKuqWiYk42s/owretvS+RaQmS9ahqDUrWFyJlYI0j
GGUOgpqGFPiFgztBx5hgrSXtkMhI29uzA5FJUS2zMWE14ratciW+BL2jM+tbVPN9
VEeNH28pzirdvYmP+7VkpuB8jzgNGCWcMGyWqDynxZV3U/C8o26/eQymztZmgPd6
QE/LlFtbZAZdoutRabzJ3JQ8iZ5wJf81QiKBuSMCPybv4mEPLiaGj/s1FtLPRtI8
5Zna7swxoXxGnKMxoSHuiB6PPgW7yayiICqNU1aOPmdzLLW09IehrucEWKP+IAnf
O1ea7Zyvc6amboUAEAuLgZaiIY7hbQm06EhBlmEKtZ6VPk0a/2QvpE6tSCdcQYIN
UxyIMVMUuyXZTzVoxx/rsdrxeXj86z0ETVHlmpCjok70h3PBtgIEqeqAkhgOJJNB
k3mK32xenTrCyjlhwFXV+ieGE+EdbnIfkP3gzdMVGtpdwXKTma1cdnRp/RaxiIU6
BMOozcN6EVtH0sJPnCQE7ktYcNM3zhzZMAHHdhHmjztzhulTJDZBnjhxfcVa7x3t
clk6cuML2fnMBdqmOfbAN0Wyi9Y13TAYHmKGLhQghOKq06h4K480DxC6MPQG/BAt
Mi6lrO361atucvWlgQVQ7lZ3OWEvdUgdd5ictC/ZZOrOPGmCoNsjqD2o1G2tVWMS
utZfh8Mu5s3uz3XjSbW6oiGi00QeOannpOfb2rbQXwhGQpGXtrJaETPGiB2VG7Jm
LDAOudJelR58xu/gmV7d/Vq/4pvzcqycqYQiswDSVBnMJriAHyNS0rkiLeBnmohg
Fgg/n4jmL+W5zvh76F4RqmyfA1Z0zr/HAFAbuyTcwA/K7PhP+xAO2XrSVU2OfB3h
JaoI3oNa0qoXlmWU6Qle8yD5TzpmzJboczyu3jo9EMUcZwtlPtDIY/KGcM3BmgLB
YLGqkbXWtGK4LXZmCtTWFcVmrD1/tvB9nQzvF4J4EJusve7BiU0bY/rmBIHTwrel
xyI0H1ajz08CbJUA1rXd3IMkrpSsAAf/z5a3MCGfB7cXDwrMvk5oVtd/ek7fEZtV
7TJ2TFZOHu/K3kH7pyExy2qy2U0VnYwzCm1u0HVWJ04EdGoF3t+1lAszDYW4/w8W
ogRa5OwFhJ7HPjiynen1+NvRNdEYP1LIQyw4yYhE0v6HAPr6AkHeHVnPLCreqwZl
iBIKh5gUlPhKLWicS9EP3TdAySaGwwmv1Hvdc9NKPGptiZB1kfejBODTL2doZKxz
wSHuOVNL8gXJJ1nu2Uz/fwowev5VZAgcf328tPg6BnTTy1u/PgAfB3iyXRvZ956U
a2EYqLfI04K/Whq9c/NPDG/9/LSKhXXufN1qWEkyU8WxtfZb0t8nlHy6G5JkX1uU
ufvQSPlG8YcD+RuqXymia6jeQcgUJowX92Oh4kAnPKjeQXuE98vLRpGsC2X5N6vy
6cpzLYM3Dtk+73EufHW+6dinFk+8in+3McKB8uhS1Zdhf0ZaV5QHZVEp7bBRwLAs
K7Tk1lalGdW2EdyKp8PeluKnjohmxmWiotvV5aocrlEYBaOancdu8+u+tLj3bwGZ
L0SMRCCPKDvmCED7Txl1Sdr012g4W/o/b9IjbrI6Lnd9huvQbMkA1aLS53FkE7n1
DRnbnUi/7JAC6g7+GGYuzhegP2BcWTGZGBOeSKFh7TE7zU2/DoYilMfleHKeAjLT
qgp2V7KSHR3FScUZIOk3pDEBFQkt7lnz1NnYgirB++IpySZNxtq/pGsZxm8OuX+D
Avzf0WsKs46RqgItWT0HVqkPGxBKPhdyWq5Z7AwnEQfK6p3yUIk83r9RKHuEM5jr
/3l0LB/RwJrXKwQEf+N+4aZUnxXy1eMqkRVqnxJ32/MiU+uvNkXjOy5gtwA0IZXk
9eYokFNB7FHPCvHCvA6tePy30CpWaKwxUsUBzZT/UMIAAcr8poiH+sgNR8DgQFqx
8ix/TzNofQZ3S8Y6izmCmfA1YNyF8kAguqqhhrnb5PwV9eMHUmaEZCShUAezrli1
3WICcSjZW7HpallSvyqEk1ImISrJFxnOoQWPr0unHZM+AAmPjegvHn/HUuJjyVmU
xFEGYibyG5EIB67gAnI01N24aMV68oyqwKOblm4V0SemkeVge/+mLt9z9eOaGqML
mPIuM3KgWK7k/mfFjux05WOOxYZ2ADFZLcdcB58uj8aPZyfuq9pwhK/yHjH32Ggg
arjIieSLrFQGjyhrDF+1l0BSIikS0bO/iK8q25U/OC5HlvSnks79mxVdW8GMRGwE
CPSfG/vJB6R9BJx70VD6GnJk/UruYmdnjPlDiogAQgOasvGeWe2rUUd9T8rjw24N
v9Zry5cBG/ly0M0pjZ9UNLlCoV31Zj7AGnQGqA8Fm1/ap+87FCYeweLwy0bpgH9Q
rq36Jps3bWzGSyMQ/Q3yJdIRkG11RRbCjI2qG/mn7MIpSTBGvp0QqSyGb1jwhoM8
4RE8nafuj7Y63pPWzxHnC9pJizBp9DSWcnYkxxdhcxIQqWsfbYb7hWJnUdeWHXGo
hdfI1M6NKc/KjnO7c70dkIsp3G6AQIjq6eGXDNQ+4MTbZZO2fK83F0Ps52GARUCn
6uLQGQvpBGLiIWVq9yEY3+0w/5vkcxtGTJTVKNiWMEdNQ5UkWPoUf+upZsRtDwGd
36h4MM73ykENvNSKoxAPq4e6lpo2nhW8KYofW5t2ulcbYXasrzXvYHSaFhYfrlkX
+HdVQ3+ZlQQxTC63YZFFidbza4Sr7Y+H2sTys7A25SUFINN3uUNGgtFHL6rLRL6f
RJuzWHI8+1GjYQQCXyumjpx+GDQXvtu6NMQi3OLpWztu7HKeA09aOd+Spg/s2CFX
+Fn87hadSZ+fSfg2F70FAu++Cjyu2M09ASMTyz3LJQF/c7ZI7DdZtqd07X9+Pnfx
d4r4IObfGYzHVWvY+B4ahtgyS8KTmUJnvq1swxYotyn7c+NXkrKCOoMbNMt17AC9
TtP0QAq8njHjy5xLHwiraVA/qLjaDlW9bXOM6VkHWC++Qr7OiGgd1pF5vr73GcoT
Mprmk4dt9Vd/ejeIvIro4WS6MfTgFXIKBuHCfMkIXzJQbm1ckWy+yX9Wyh8Zr2g7
nCJt7jFePeTUeSgMShVgqQNxsIfXmhfN9rVB1YH7wwNe6tqZ7a8fU4jFQMbEGICs
BasN2Q2Y1kJyvHZBZEAv9RNVpZae9drif+ok6iAmewN5GSy36cni0ak+LZZ9f0LP
au79NP75XdpJfvphTgRyEV5EvqXR9glygE1pwvnAemioExcKm5cdv+o+b/HKGC04
Elzbk3AfNOthvNTV+IGQD6E8U7yP1+Tzc8ADJvVridMsIbhLEx8znqtyQ3JtpuBZ
Dz3lFqeRoPBuJXp4GHpUH9N5K08BKHW1ekc8tSgXqMMqHY+rcaUzZioU4NZTC7gv
cEE80pGjKgnrrIRdE0WY/YwTrTIL/J6vu2ZgX0G2g2qDlgd2ycJ0VhIgeGihHGEy
YIbQMeXeuz/26A0ahBsQQbYHuFo1HhQgmPRUehyQSjUvfA85FG31Kw4qxmt7VG85
nHOI58seVyc2dVzvktoNkTRuS5w7NpOE3F6CFP9GXID9zXg5Kanch5IpOEyGZPIz
3AqbO9g3UhC4b9OK5RggIHfdIZreQLkVvM59PbgJMTR9n/MVqFmJHk/B5eC5rbXe
toNDT3LYOsO5VAS+dT+Syj2HYXwXmtr0xTcyC5mCsSqym8ONZU/p2H0oEJVTEALq
aCEEkUaolQpFRoREdmfzRWpCGr1xKDfRbbAZ4+HyH+AVeyjrrXEPK6oY4gdZPWbn
c5Dfh9qQwRPumI8GkFTWFGV30UN9zeDZLXk4FD+8u6E5Cl0hR/+ySoZ2LEMqI2nn
aIJG5uQgabtVw/0ZgekyYbox962wAjUzSO6zR4s9lBrza9Qjx1uPO13vJcwKTh+V
m8/SN1dTmts7sT8QhNzkLjoM7tIJMoJGj4/b7kteQhj6Z8yFVdMX5jKg9tN2sQ7w
EVRZvqtqaMILRzA7Dtht8S/ITKbWr6B3wuT7GZuzrKVvuZhxblnKdsC/PpVwgXcV
O8ud/L+KtUJlLtkfIIfMx/E1OdSsS6soq1JaopcMVD/TWurikHOWi/xLGEDi5vca
hsu7To/gY1mOJUOVOhi2kZ0pVoLdh0Hco+xNzMhW0SEM/8FCmKjc0Ii/bsmINeZu
SAniGOvi+lrQdfbSUljOwQ+og53/DfGMQIicML0B3JifDmgUSd8Ye07NY50T6mdS
CB9mGI0U9aTqPtjpcVhR76IV0XBJFKEgubfBY9Rm0fK+FK7LpPKyZxNhDBASuwsI
OuS/l4V3Ooqc8qoeTghLhzlyEhHwtz9xyTjjy09SWKhcye9pJRDEuBJsjjoOIa0v
r50BsV295Uho54bYZp54EK0tvJgi3LY2SpBy5rC0W9TveLrxq+atC7lG1uArPymr
x03tOnCPv5x2fmOKZbe37PxNZsckFZiJOUfWg327uXgsSxOXFtPx7G0eYxReZbrP
vYXtRudyXeKm+M7r307KilkwA/Xv7TDk+o9tKBfwcp1i3EnbPhT4VvwR88torw1v
8cSEangZF5nehVDgbpi6ffTOe0+ImVdMCBsiElhvXGfFGVTcKJU5pde4JezmKavn
1uB047zfXgwiGMqu1mr6sApeNPGPNhRvxEiw4fOx4dcWNMU1gd/rG09GPhvBTcFL
nYA1XzaVbPkH/Fi/ZxY1Putm8k90Lmzzmx6GEccNECy2jiDSjV9mwRTKMJf8rIBa
ypFsHbLYflzrF3qvVvvtwLcQ1ayAXOe4M+fGHT8fy5EF8IDRddL28AmpAubP0nfM
aQMlejWq32VTwtYT1w/Ph+pWRPxUpR4/UGLBsLo1FzwCxaGBVgBNzeosI3CchiNY
mXSsP4zq71ZEf+Pj5dPwIxT7+rSnjNKIRvrMiSpPOESkmz0fnTZWTD1teBG43w1D
JQe7WeZxaPhfDqDIxfkgoAl08tCxX6hyHvK2uMEfIBKa0Mi2Vpciy6Cae0Q9MHJp
4uubb8tsHeRDf1zeimWw1OE+OKQLF5gH4ftdVRBnBRyaWMRwywlpCZzB4Xb8/2Wn
TbOpXQyT06mPrgx2LZ+svSBlFyYUV9OucncuOokf8tXetlrR6YSOdduZSVe9d8qn
3CIxfSIrbTcQQsUC2OGWBRjvo7cFMpww7+mx8sjMgiTsU2DE9xiraVScU6GpYLmf
VXPztadZRmGcB0QWMnv4ROQUHQ0scVG157ddmWhjvVMH26oSt5v2O2fce/IHAMet
F+VnbXXIYi/IuK4CwqoDrJIZY6BzrvVtFrtWvOXTUtAXlcsn0woG4TId97ZjXMMz
Y0oPZplsUwatOtpGg980UsmRCod2Foy1tsm+9CmNSCsvfSq511UhJY4uWRV/wqOG
0kYtnFXszhglw1twAhtBJ9d30PXBSzZRQPYhLSvfv2R6QmGxd68wy+c3LGT+zHFh
56yMKdUTtpXaRXsltI7DE4Fk/aHQuGRzwk1MsMJ2DWDL+WLSZh3HlVowxhMJMmdK
woMhjrGwi0GA8NZNIQONBYk+IjwXa/pnDA6faqebZx3b5Rw880zzjy9k8nvv2e0q
7ez7kowAi0zdtROdhsqFXVFChwe1/gT+ZROEv95/kbNFwaZuhLH70p4mKBdFJv29
s9lxRTF0WCl1n7W8BnRTguVzMp4dtUBV5VyZV0XnF9kt/GZBtvIFUyziaB1hZxLi
yvj0OCVsjPTSqaKPRK5HfcxhGlx4JuCFid19b2LIJLTSuPanrHn/mnTf0/EWGWvk
DcpjA6mOoSdiqq0Qf/15jrWqdCMyb5k54uo2klhIs4/17M3hFRRrzrh9A8Q+DW3I
EWYrn69LVbyuWaEdpc8AljSMz4HNiM2yL2t9k5Cjsgkz4GQ7eLMFyCNz4RfL0Mi0
WPGUZoai3jVtbFbJtnFad/1hlnKfS2iDOE03e2duWuZIrRAamxblWOBqCTTVwH9c
SYr/gSJg+Kqi7tOGq/cecF9ETcaOLcjE+ckDaHaOKUH1jeV7B3e/v8PUFOSRrEHQ
nZDR8Uh7VjciL2k0vcuRDhVZB/j/W0IV6/2vnRkrbhBYIWVCZxJbsvWvbR5+GK6k
W1sqQwYLcLNRqjLD3ct1iafodp2ibtc/WN4K53sOuMGVNPeqBNM83yIE1FRSXBH9
k4cgzyKwDOCwnchn/vOIQo2dhVdf5TFyxG2hNNvUGNB5HhfJbgYIfNDYkL4kZ6Xq
vzIVYcHfFjkwcSWaVAIT0GxCMb6yv6fQthkOSnhZ/ln4cIb7XoO0ww8z15CEFWAc
BeNfbt5aEbHiM5MgHQN4dER8RjSUnKswlitd19QtkD86yAFgksW6+3i15/Q1EpIB
frQEdAwymEF8IZc+I48cmDP0GTsTpC+vidTkFkRERMRrVQ1iHWtuIupDbUrE/4Ao
5jnbKSG/DLiGUvPYeRfAufb21GwrRmavXkOSnjTvdcc7NRhFvvyq5K6D8sw1wCTJ
hwxng8Hs4MtNQrmRkNFBH3RempGbJ/EezDoXgPJQFB2xj44De0ISLg4nuiY2M4Ah
6czB/DE4buKx2B9Zrizn5Yl7+eoksD1xvU9qGwx248Bq5ORpeM1cL12xqkLzZWFv
zb19L2dA2jSBgWZPMWCdnvbXUA6F4Hi0Ili6EQhcbB1AxfH7b2b55CTzPSV67qHG
5Kmtg6LswbTzyml1plQcn1kkyZb+poThXEqPM7Qz/J3nhoPcTEw/gt0wye31xMAj
YfrNyXHSTpKiSif0r0VYFRVMsg9Ftw7pwEN+4O1T2Bp5hWJPnnYMFhVYwrOVGjFx
m6wb3azvLxYov2ZTlueDjDKjBIRj+5YZXSjn4gpWmBCYW8Joq9k53Kg384lAjJxP
Tc5uDs9vNnUaZq8Nl2rbIXLxzkw4GUmFVqy1MUSg+pQDBPQSyvnyXqNKRk/TM7ME
o4Eia85jlT4jdaSjq7mZG968NFadVBf6UPi9HJM+hsChYbwVxcO69opyLvDVCCLn
Skz3hXUJ3ELI8bUbu5gUpany/W2Bqlq2vGiAA3b8Zgbcom8zTwJsazdpY9hMf0pl
7u9zOqlsWIc0NVCVL5RMiX5wo3mI80JoQFdiM4uFI0F9Q/pmkMtUsK92bkwV1uBQ
4KySP/uVoeu11tWoTltI3OIS+wKnMXYtn9AFA6BSInTMt323lODJTJ+Tu7ED7pAC
nV5vQV8Hw/N5kbgkpriS1D33JgY9mOP6Tb43NujkL4Rh9h8RD5EyBxe95LwPjtOJ
UxNSS/zKxkYWstTC+rzCY3IZjAAZj5j+EsTES4xW4DUILFI9kgQVKAmJO6Xscihc
SRB7vbaZ/H86OIlf/hiOWp1ioBi9JOmBuZgmLLLGOQOGKSoLEHbF4gr61v66K7sG
KiTQbXsemIC4nUp6p5vF3SV4WgFobyMPD0bTXi07I0g6F+wQHTKgKcjmfYlFtpLL
Xs56zyLP2n7Gecdo68H84Pq6RM41Uv+YIKoXs41ZIxjbIjBX53okIqQSEyKnwYhH
danqN2+MvvLDyCxqqHUvOtB1d20sTliYXRFM42jyQa+2JhofdtJ/YlIXXzAYwFxr
tu0Fhp7r2cTvlltcOms515hngWzohdprWEBafXeqc+yYnkryP8nFxvSID9fc/a4T
W4Xmnm4GhxnGzhh3cIjc4laC/DcRFpexTWEJw4Bujz6s2n2QhVyoeSpWoY4I+3no
CNhUaZNrMMaRzlftv6RwDlUC16cBfwAE+S/4DR/cl30YeBj2CB6Rg5P3AXvea54O
CsmNTBrfokZZFy3YqBU18A3Qph37bYc+5rauX/o1O6NaPMISNjni/DJZ3SBX8rKx
2UQl1Cu6vslj2Se3hJCg7WsyRXsix68ji82GWKI0n9ulN++f11P0YgvfVsBXMnkv
C9cYsKeh2sv42KbDrUjYomAgwqwVZtcvJXY7tSJkCKHvfXJYsMLWa2Pv8KKyEv7d
fs5tRuf2K8ae2SranWaFu6j+BMP1badY8YG1yR0mLB2r5plg9IO+hDTWPPGw1yrx
Wkvkbl2vEd0tik+my4ULKVBY8QLMDUEYz0UldzbYRqsZ++bEb78VZuCMMpz+wi6W
9F+6VKtimFe/ZSaEhGvXspIE7aOe9ul5QuEmfsufoxuZBoHsQe1AzdtPK7tjmBHv
uXZ979o3E99dpBKkAnwZcllA1qef9C58hrDHW+jQEg4A+H0JlRUXg/OGxrSNa2ZW
F0zZZucqiXa6JOpPNVgCsJjQL/RXKq1tY9VCwFfOHCRroAMZAXy3SwZ0MBx9tMZE
2T4MxYIrMJya2oqGhv1lxxYNIEGCLjsFj7OrThf23aVZaQ/YptTVt8/BbGvexlYo
J89TQ6kHK7igxqYAdJ7VHSkQLQXivSwAiBpKnftjgHCJ34/YSTewCX1pdLwEtsEI
kIByoZVEFmQsbhRCppT6X85QhDUjfm40SlxrrhV4n3zRKMKYaM87aHE0EWHy5+6j
sp69J4KpJbsVSAn4xyOsmxS56UYmtMqVIVsj+oLYDe18RVK9iUQT0Sgd9O8pur3f
TUSytdrZN3xQANq1DLPnqM0Zr+Yn6FE/X9dXekEHKq8UfgIt0GAZucsC1upET9Oz
QwpWuPVeM9Z+YHYEkEOLuKV9YXR1WG332a5N1pr2TGbdFD7oHBIzJeeGPr6aShP/
HvsLlE8cIpX1Fy7dUKN+sxXA8KHC/gpPuNWYD7anUayU2GYUV/jv8Qidam11iFdE
wf+Bp1A9R6cEFkuA3pMfaztXRdI3W/xBCnB4uTLa48sQiBpT2J6zSBJW6DEfqBEv
TwoxlhZDOEOXZYBPUiKXqINzB5QuQMZtvNGXJIGKeWIxBb7aYVhPj108F+mCoKxq
oo9tKTs500oJ4c2wjVLHavw+OQ2s1ZQTkNxDukxs8Zlhx8AdkRaVmTb2Hic64bBb
GhaH4EC/3u60+kEEADo8YdjUEGe9HmV6mUpyK72comz5FPlbOqjrtJrTwAfj26OU
Ai0oqTxNqGAmnubiy7DaxvWLyxGgcE5VplAtbD2tQcOlzM3YXBhbMonieHwTUg4T
UPUEPXP2srZfLSz2NwTvd1JShUMKvupzrifcpa+rNoHsPv7XSqHQBAGU+RHVHfwl
ggSpzpFqsS33TLD4P94ku3p7enfAhVb3lecMjQepEjs3txa8rTZHs7uruCmRzVg0
ruudjYFleH/WDzXJwKapo8PWZO17iqCPH/kkG5fcpdG0qONDUFFXXulSVt+pFLn3
y2+aGoKayGDJpBhgGBYR05eSbKzel3eD4WELfdxQx8MKEvxxUuumCRUc2t6xBvnk
Vhp3aNyO6Ce7mxjQCwB9rybIRU+gTLpmmVldaYFsEc7qIfsDokmEJr7cqHbvBqzQ
YSiqsth0lUxJKmHdIrL3+yaNcDrEjDrlIW4OymNjoqA6A/qpPhgfkBcb/br1Sk65
gb1fDEHQQTM4YXE8gLSNDmBA3dZE84TX8/tYPuASququpZCgI19oQsr/AZoB5onf
Ev2RDKCMV8lxfFvf/vWBerj11mjx8SEvkNlAqgZySS+aKc8WpV4kODehEi5y3LuY
L/+PGtLfHkWoCAfvYNkmeqd6UZZP/qRm52jBllU9e7n+vEcqANNaiiQM4CncbvUv
YB4Ec96IaTAPd6JrzGCgoV9eLVDG71Q8r/0ICT+UKQ8eud9Q5lfP8ZQ7FN/KjMyb
Kw8dTIZvtWjYZXQyJi99YeL8hCzjvIS4ki9PLPuRyLpx9UNPsF1WTFARtDu5NtRE
0Fhvsi5X6znBtJlvO7CSuRQYiEyCSqoWN4FiqLnuTPPaNlzJmMzoWxSSLMhjFivB
cIldltdO3aAK14Cmyd8PNC8ozergyKs9DKKEnzzIKVb4DCPn8hmYnPCBghaPMXvX
bV+fCs/POP0qJO/5+vL4eT0gKNJZ7xEHZFgX4CeH8sYkU8y6pVqGXjg2A8+qntVw
/th6j9phLw+AFbu9VMiZRSvPNBU72to+epJd2DAX3MUohFf/H9ic7IyO1BuPxobk
u793Y7oIbuuIDIcba31NAr/WtXBFAbeP5Yv2o9BTHb8zcu9dTEGsvbQ+hCAQle/t
4vvv2CfTLaaOXZQoKVKRcbvi+qYUAtQWOGtkRT8MvP7eBpS375Fq5UyJW6ls+2J0
8A+UOHYHJ7pIkLo93CPPlMgct4li1V0UpVOqwkCvFZsNAy9C9oqphybKzEIC/twU
zBZDRiQNyPCUaCq7CjXsn9uXz5X1OZlnTTdCrcT28nu5E3VnkaZK5FwOL2bjslWM
UQ8XzeEHww8z2t7rKfMCwWnTtny/8lKZb7+iVfmBuBFkp3cDAa9j48S38f/QMvtz
ciTvWzcNIlQSXyWiiWdFGFAmqfB+cv45s3nM4sMELzv3R9SLi+6tlQWifoJ0THXH
sJkqSTGshHI3I/pZNJilcJsRAdARFa8lbCT2zBinS52+2FF9abTWJOZUuU04J50N
gbKjSVKvwug3tnoK8cAPwrI1xI+sTK4iIGZ0scJQ2ZR9WxmmPmjXPA+7ZETkHwN1
/lO+vvTX6jk8XxwnbsP3z6m3/z0OeMStDGlE1gawqdixJE4Ru6GUdQSS0WYZoyWo
ZfLI8wKpoolBjWLyPv0HyKiD80W+nzf5gpu496Nog6NSFaY0SRBEtHox1sf48RU4
4P0DTmnk4jNeo4k+v58IBJxI+gB0mWPc742FV6mmDy8p0hXeIC+hjfY1OXvJj/mv
DLLs9QHDaiIvBR4OyWi3vNEXpZUY8p0mU+T/Hm8GhnKkuju0nCHz06UFoaLxSL7f
ZUDCydc3xd8w7I4Soo9GwVMwTOU0xgKLqHfVGR7dX1kCMYssKkBizXoll3tDIrHG
t33oh1FpkYGDGkzJVIWuS65Ddd2kw2tRDlHm+cH1eVldruScBH1zCouZvXKTjYvX
BVbVRlP2uzwYPVpskJ+OvgSKijwWFyGYwPEispaCNXin3jIV8eviMhwGGwmZiDlh
13yiL/LyUtHas9clH8zWLFGlDhY/GdgJnEDjZULcRU4+yOfR+OT2hPSsFyHUpHEX
LM5OOFmmEaIc1H02tJpNd+UGmLb0f6jMoP4gvAYx2DfEb21tgTV00lS2aD1g5GMM
qCAM6EQ0354p2Sh5QAtxKMJm8Y/VPFkYC352w+VnrTjvxRbwTPpZ/e3PrcAorSSi
q7z1DEV4auQnwFLRk/N83oGcnU6YPjQ+NcKwumVz9SChHV6JcJcIAMu3soUqftnc
0LFaR4fQ8gtNBNIiKPNP1TN09BcaDcMWZ0CRAcOjH9ZJRqO7Ax69gY5fdmkdZNOm
sIX+2IYmD42dN7WJLdgZHQGoqgbT+niBM2UmbNaGAL4CHTvnueF4tE8lYyvi2kMJ
HuwsLkzT/87XKXY4qX1vm2NWWftxWZg/rJ7GzBFdfpQUKlgMnTQrNesGK18zDXb7
5IWaf7JgYSVsuFz7XEEv6uy38U+vO4FVnlKCgW4UCjMsGJR0xylJtfDpgSpQo1pb
O2scDUWOkcq+2nAjzT6j5K4dFTI/lPf/qgaAXXVACYEODp5DzPddKKKUMWfAGeci
6dB5fdD1kGddYf3aPFYkPgOFw7n04kdtVfeJ5kcLXMO9pKkgSh0lzodGCfoiK5hr
xoYNGKf9MfvNos1otUaRajC77hXmg3uLFYL3cCNO8/YW3m4fgjb3IIAUgisqbjlD
heP/cRfeMgVMMmBhIP3N/Pp4wyMW6JZTii4FaahQCYlZSEY950LMEc1vBcYFUS4O
7eLMvF3ebKAa7tEjIL6MfTGM2Sq0czLy0zsLvObPxWjIjsEbQ8F1YihHgUR3p3hL
UFOgRpb5O5l/bKZx4xpA/w/wawpx2MbkWMedt4wcYIVHp88bsCwROrVtyZl69iIi
Ro85uXTUcCHJuXoX7y73cg30Wkj7z8bdGDUJWmUQaeA0Nj33KMtGvUUFxQowVnbh
q5cSnD2ZvtFPkPIkdmDbU9U1eP/3oO1g3QULXV+vYHH4QsD2YdAoEasb/PTKP00K
2BoKySmanjy3uIgPFFztCdlOpPPT2TEj4z9ESNUMQWlbMngEjIUiTY2nFVuwFxhA
s1haQ4Gg5I1JR2xFEFESoaXG9VI/dYCxIJe0o/4l38sBHjdrYRaR0Xw8YUUTLYvP
VyWYcUJpG0b9FscjO2qp7clteL6qq3/xxiZW7KtwIvMssWOkzYIzRsbCmEbtGf2q
FnkvaH8orFDjV+FgYx57O07qkUd7CCbv7XVZ2S1JjLtc5iHr484dmfevg+orsuFk
FanjwK0lSRkWiIh72qES9TSrjVct1QEHj0EOC4jFkxI78C8tcWfmRlBqsQy1G6Oi
+0KnKj84RZ6YTyP2Xlhke2rIE1koCHvFExMpgLuDS/lQ5sTaAv9XJpQDJs+A5nQ/
96Gb2xwiSuN/ock81fy/bPo1vlxAnB2cJb04T469IJi8MUlah6MJ119ud99c+Nq1
YOd1cmdT8x9k+iT4z213lEf/QgzOcauqVlcOIXm13FrmblOvcsnsGic+LHd/UZfk
7T2gMAWKlMfrfcBs+XlF9JI+pTBT3ED0bxIm3XNihjUBe1Scd8LGv2oFNPrntZL4
mluV1zBJOTmf/3cwXZPUsKxKLTKw7b9L8vUjA+BOz8YbWfmdg3lS923D/GX4DmQ9
lYde/2oGmblRdi7e/sq2jbbWSpihGvv+Ceq/0F+NHlmoAt+a8rpVGJyt/TNhUHJc
IKz24gwwmMXTmGTd9wglnuylSFxYLuo/6ttz3idCk2wntm46kexzOK8sSlH6S+/T
2Y4zT+ZoOlJALjZtr8Vdftdjym4RzkRV46BjyE7yFkZ4coIG+PdZZK9kzs0v4mqi
u3sZq6X/Bwxzm+DhXHSRfHZKoclCDg8O47kHhs7A8T4wAFW4kN6QlN63Xvm1dKwX
NRne7HTESGXZyIo90q+6UQTVZRrxVfbXo4f62Y512UyaVfcGORHkH9IsFP6JJnfc
UFDC9oZSuUV82WBA4zeI07irVZVxI8o1GsasFBuFtx0n0pNziYUW30ELdDkZ6Fgg
G2l4+BjRnO5fcEQUmpBLKjt3MUBfJtVHdGQ8bjeUT0BhMtVSi+JQspmEsp943nNC
w/HfCsv5rV73kgVVTdulSv+UHhKGHUHqhvKs4YwQ6eftVkJMLEoJ2M6353DfVdly
YeHgTQWj+IwVC8bP1LvoQYXqu7mfLbPj1JX0hVvy2Vd40Tj9GwodPIJWhT8pWiaD
Dm54mtmu4d4O6fUppjqwgIB9MIZPh5YRYjJlnqWsySEY1LjXoWIxOSPd1bB8FkGQ
jJ0+eaZwts9ktVgy1GgGeJtHlREp1dCq4sZpw5SHSG+pFH+W4bK7WH0WfLDdaP/N
wZMF06BRrysPhgOJq/8mjDvVNd3f3u37H6wvelLBtBYUnfx+FYUJpxE1SqRF6Pvw
0l74k4BwbbUcMlh8xX1l8VKfRiNBJKWa4CPaddsxrYT4cmLqlhBGiy6ej31Tw4+H
yz5wCMyUesfiQo7RsO1Q99ZMeHVjtLQDPDNcRjEO5HeYZgc5Q/jUbBvLLlKCHkRx
C+NRjgjth82cJrP/RYDHo8PbMd5QCB20Jb3AaQzviStZbevBawnByTpuHbYZmXGk
Hz0mmi1xfnIvNrlc9oG3EF9TCdLInSx4BzO8GVMO/HA1m0FCnWn/8RY4kCh2G6mH
Dhe1BMQkkhVt+/L5AV2tmWnH0P6gxJqd7//pzVx1YXtJ0cbVkcPFyn/i0J/1Ei0o
u17FEGkZAHsgdaMLe3wZvBUeaMWGS0ZuUArfGOAqnSr4NZKs66EX520zR29HZjnZ
hcsrBTz8XYDv11biewowLabMSCGBbNiGcQAj7ORYWodnwx+fHj2nci0ZKoaehDkl
nSM6AJ0WZkqMdZF+2LekR2UhLbCLebUHoDk/y1Lfgqw6LbJNASk4rYDdLA1/2C5n
HbY3jbPSh5A0dGS3jIvvzOc7zlDx8CRCbP6elbzMNSHzhN1amaVSpw6mjPRdfmwl
sFFYaJE7VbxycvQWPYWDSsTaOZtJ6ClUrd0KITqjX3PEKxhGpvi2KXYpVAoJsJtq
JyXQKBnokJKhuB3KIn7KLqgrFY/9WEqaVxRpS7ox2C7dlRpyRrU2SuPo+0FdHnly
fP5CEOUy6WM9Hvp1ZtsAUbwYFEgr9EwyfPYT/smsOBAxo3F5YtMyAeiQZawp2qF0
sfZa3KnMoqHAQtVgHQJL08P7AuAyHDc1VdsxJjdNvbNVZNK04O9zxBfC8K1AjKzk
fQWe/mYEW3J9EqkWFLJJLxyg95FILtELkOhAFOb+WjiaPjYOS+L5Z/ofY1xPbwZV
l3UiCRty9UGZfU4cwHqgr+9qZrucSdsBYSp11Ojz54kye2Zcdo6bpsj+C2IqR+Wh
pV7Ol3m5s6i9FNJllFBh4+n/juadIeZZJem1sG1ZHOAWL4ed8YYpM9OK03ypCrxj
Ql1Ubi1zgKxhcNsKZ5+P1fok7ErLQXadgHnpSOReJ7uESFUiiwXJ9l1SLcQYEQ8k
zaN8tQA4Uk3yS2EG9+LpVy5zxryyr0aMKo3BK7d7JGlXXThyapvD62rTrdyk7xjr
YHSuNa0K7CyisuIBtTYTAGyIXpAXWR7tagYMgFO07Eaioasxte38Ei7uyWRwUgzV
s2LT18fGsKG9hlxResfzBLY2XJ1xxmz6jD6uwbVgIFJQUNGzeENJyIN18OfkmICz
aJ6fq8DQPWmFwIVQYCvOlPe2twY3ZJfdGehSlYkS9Nbl9fGNFmDkkzaK0BjaEB3j
L9Swn8aimd24T0Se1dNXaRw3x9kNXYRpxwuFFQ3mB4ZlDvH9eg63cZCzwY+RawGO
LH+0Z5NFcc5UjQqJZ+h0J84SgKXh3LBbOi915jaXn01K8Wft1KGCML/MPgBPtZSa
4dSCrqGyI+z23B/bkt71V105LYHWg5x8VD7Iny8JjMunFRY0HTwlrFYfDfzh3Hma
w+bwhiDG537g4Hm7KIQbIAVlKvKbBWdL+d6qiQpdH5ocm79imi8TgGx2mSbR1/9v
BoWOthbJWafsupIYTvIh0tTxjKw+e8e4OP+W8UtQfTR4W3YaqDqP+MLxqFu5GNLV
fCf1HOcv86kn+KkbUCvDmYpBYsC27K0vU6tKqHbx7pv1jfU1jxRRtgb2T8QfZx84
PWZXLJwdShH1/2apt/4H8CYAfJs7oEQaknxIJIq0FedTobCQSAGRkI6PV8sKvp8g
7kQU2gMcOsX6tviPWLpz4xnQwxcPZr/M3XE2isTVXxIh4nAdZgYNTELuPSpvySrl
eU3YLrVimbTr/tm2X7Gg6IbPTOjECur+pR/Bz1FjhuQvJqkXxIfDNsDU/RhAi7Tb
pNKopuT4ijEwk4kStv1LzPZtNRr3LD7Isxb/lLQmaFy1txk+ikYsoIh4L25ZzH8c
ig4xxQ3FejJBuANHUMt9LqYet3jIIY2fn4HENucllDGfZfeffa0oza+HQaqXkpKE
c6AfQTw9wpIkz8HzGKC2aYBdgr0756tyNUQ07jUFWorS7AbsmQAlEG/yzbu/XpL5
sNoROsgqn4XdBZOuQ1dyhSDmOOjN/TKurZJ3bpizVbBJVfez4d3t6IrpGm9WrmdY
azW22uIZ4xKm1K2nYS7FMXdTI7HaBKGroDzT/HiXjyArnt3aLOVUGrOQGF6XPbl4
Lsyqtt4JHPJ8XuOKt+IL+aVo99g+FeTk0gOcrj7VkntyClpK6JpXAbDFTpjLvdFU
dh+oAAzsky6fvUkv4weBBjdwyEOx5fcNFpsKmelNQLcHoa2bULIaf8/GsW0CrMxW
7A+2yccbhqWSIzSREby2PoSr1Ci3R1hnXweMeVSj3X2hyL+AdqGZuCVUvXxlrKy6
wbJQGipMonE0k4XzdBXbV5nJ7o4JKNKre0yE2Fh8LrlULfdXCWSESSKimK52mJXJ
2kG6Z3/2CDCLh80fwDaj7O2C0LP+fEwkqtEUQIjdLivyih5VVnMUGilq8Gd3T6eh
C76qdSX1h7m1qI1nBkdyrVF74F/GTKKILV4S5pvA4JCQLXaKMDZ2qTRC0u35ora8
paZ8uEzrY75xdp4NHlE+oCOcRe1rFPqSWM3wRmLxMS+RmXMXhv5svaFu7CJM/W9Q
Dyamd9Rjpdvjl93AbvAgBMcHXEXUe71Ow3SMWVGAy6uIYINwg6gU4bvGZ+WHY5Y5
3E/tGtoPwVL4jRRGT98eJNFGDmtKAIVCo0/2QuWRS/e7MVPDIMFwRlfdWqpBWOCr
X3b3ygUxyr3SXerJTGU/E4tR9R9UMTPaCmEOtxn2ooKwTfCdhQU5Yj97b6KGSKLc
oktP5VIKX8okOkHAbOiA1wb3VA9iKLhTGCIO+Nn82lkwICFparIwlAJq1ob9oWfe
2NSFmb0t55SdIbFAmXSQm235tODoHH0NQDMO2pIqclSFEzptAbSBD1bhYYFdQhpZ
+6oBLVq1Y4xRdUGq19J1DOF+Oz4aM8H6pCoTHZ6uzhgwdQE10MNRtTrjADevvlXx
st/boyhID3afhannGJfA/PXbxB2RQA74EXZL15uY759TeS93uMEO4aP6zL92DUKC
CNVvhtYZZ37fvMaWwTlRw4BZV1u6YfglGt8/xUrPq16LvIfTIYNeg/hZqeEgdpp4
nDiTyx4IaOxhh848qrTymjqh9bOvZ5pE+r03mJHb4+dUMiBoBrQe9tc/6I/VF93w
o5nrYdRCI8YZynl2TASXwohmFx1BVsclG691DgGVS3pFz12jxNvwhBFK0CyJVwtn
KqV+JQIiEwFhHABSz+Bb+VOQYuvyx/Gw8iJbtE5zQF/Gby7AylqPfr/lUR9dnRW9
7RsWEWDSUMBtzwwURncD4LrFaMFqUtZMf6HDU7hxoKWeH60zNdQdXHhdoh7pkPdh
ieNeW4i90G3Ornf+ZPkyRy+VU17BOBArgdo0lEb4mLZ5VmRUJ8wQtYZLFkBDuFHH
5QVzuE9TkX1caj3qiGRnEXM6zJWCdRGU9GGlXeJnFZesPXCUGOYS01J2Jp0oLoDB
frN4qCcP/XusffPu8YmdjqB1e9cBOy0x1g9M4/jGG/ux18im2dozxCVxfipI+Wqr
XsQ+j3nyLwlXrxVrUjU4RHvrcm9gIcQHIMsg84ISEZhr2j107E/e5oDZ102FjK/t
mllePuTjBduN+eCATtHQwbvv4I3aOjjIXaYhORVdAXz9z3D08l+CVrdOyiBIhSLg
vGquP7XKTdFLNP9CbIulE1hg0XQCM8TMh21beM4pO4MZjW9RdYWCgubrFu/5fUqB
WHeflEeW0+6iC0Vh0R4z+ylpRKXZ8h0iEpb3xvDMMXfrvKo/ZMjzzDqegN5w6Bgk
aCspWXxqpYApjjy4Jevx1tBdk904cGp4jBVbjjCy9aPZ1WwHR8egv8KdWjnSfQUm
t5batJXOE76gx9hCxSrnmO8rO68yQxur3UjjU8815cX+QUfzlmhu/Qlxln3NUz/v
ghX9g2IjQHWmLOLZuTnexAW9O1OSFrGKtm4rk2eAtXidwBJLjszd/QosnukWpn5n
XH9fmdHCplhQ/c6SByOtjfRdEm6W+1Q99fTxqj35z64exBnTWL+ERPX/2zTeoO4Q
CKs7tbHKd8a9bqsGuIAth43vqNeDd3vPJarupI1CH7hNbbgsqnUGmrqQw9JHVuk1
njbA430YcgXSOwqksOf3lgv2DhSXoI+QUqM2AcFyAhhFfawCeFZkgnTDss4yltnO
qWDk0Yfz9n+KK6Hhtda3XMi37iWqqkPIB+HAyHQjWXFydcr72vevdUPH6jAXDD7I
kCSs03SiSPI2z+4FBz0OG0qzpmHpsdXcvaODtF4h9r3tPrcN9AYP70Y/GRK0qYWq
r5Uhbf1eF+8EVC2rNbc6VrMEzD2ZspLU0oK5bfCBmox+CBfvi6v4/pLX8ZUbtPeQ
/4No+k6MM0Y8kvQmz2Ny2Xcx3Rnp8s6zGg7pl6r05dRGtmIjiMz1EuWQZC9LWDYK
wJFioXvpQWoqqfML6azDyVIKcu5cJxCjTVNdZ/ysnYKQbo22fEPf6eKZfrBEgSEP
TH0KhLn5WwtUjQpZSx1ceM2ZsDTwebIuBLScxM5cSCNdApUbYmOLTPyoOim71x6T
Q5FZl8bt5UN53ajp2W12FLvbHqi7IrEs12Og8q9P8E4BbkOiY8awznXT9Une5WgB
8j0p7H+FqrFEScHx7a6739UHfXEJ79fCOrP91CkU1cV4+zKnNszg7YoLqBdV4niI
ArgT2gYugvxjzDgDlhbp2bG+FvrV+qFYluIrjF02z7tsOQ9IyJJbOlYRrAjQCki6
GjvjftKmRu+sz6z9hyRIbWFUudAu7Br4D8L5FWGMx9U59U+Hv9XPDumdH9V0PGGn
X2hcOQhltYT+NfCQnoJskzwN17JxsKJ9tJQZz9hmtXUpJS9A+wkXEWtpa/u0fyqr
8wZS2MFz+7CKXkSUoCu7s/nnvyDCaNtvd9GvJ6EkP1W52rujlPeuLTfyjAXoudDl
5D412xbdpvXXH0bN/Rsph9zxL8HVojyqtU9vadSU9Gr+004r39/eSDoqVhzYo6LV
hI7p5rCQO59Em5ZoO5JeYRXBKcNFCdM2SUQ8Ed1jEzswH4eQVEuFwaROB0T9vdAf
1SCC1I2mdDIi5m8wHb2iYHSmOYq6otCoDRyDtQzFRM/DS73/DOhrKh9HcbjQnxpe
VBmpSepZOa1j5umCWHP6fv3PWStqKTaIaX/CdZ6daG0kIl6FSnFS7rfooMHuk9HV
vhoftiYVxUYnwInsH8cfyTx68WJU7SPPIlYaBofY95NgmtnST+XpbFa5Nbck+hDv
cPVWQIyc6b+weBA1xogi3q7mmRL0hH/4DDvsdR3gehcNObcdmoQ5/klsidIng1WE
v4g0aWUZVtKw/W2PE5GugFgzsjD13fRaQ5ur7wFL1jWB4ZoTh+1dyjOAKjtFG70e
2tSV1tSaPEBwdMR2+ayfOENvKiibReBbKh/OoswTF44lE3NelwdycNytuUQl5hvf
h8EjA+rleRMDCv5rzeLn1VsVEa+8QqatFFcyxcBcmj6cfqvY/TwVA2tEzStkSSB7
mt+OZWAk9xbY50q37DixqegLpZ1ssLAhv/vcsCnxDC3sdk9jRCDVjVJMgU3iz8gB
DYSnIrBt46UCl/72efg9tIyRakK7i9k6F1cLgRgf2CS++JlI+5kgvbv0I9BZr7fc
XLgRB/iHzQUCvjS+XeQm1YoQS33StRvFKWdiFD8zK6at3ucZVz4mTCknpwMVf3RQ
EXWfCZohc7ZzTRnsd70fYrY2TL7Y6W7h3e1m9Q3GXJf43HKIeOVfNfM50bqHXs8g
gu3qmCy73LKYFtkLhmFuPsCxqtLQTl7V3mHqW9osQhcpWmQClg3neAgCKTgab9zp
T3mP7gLs9xf+R9ZM4T3fHjXLFedJR29WVV6lwc4OvMr7xOpaKfQNeVaPA4Ejh7/u
AS34q/g5LMt660EbyevVWJwiE8XPzuz7OPzt8vLFi81st3gL3wqeINR4r+qjmeBl
MhMQwmDSZh0977aaF60G2/GN7F8mWonrRNcmaeaggGd5Usozmvl5APr6+Ft3vBEi
ItKco1J2pPLv0Lt+EeuuHQj6td53ZQBhRJrj8SntVg4mNUYtK9JlkvQCl4hQfXlz
5Y5O28zDg3/EY7vNcThFLD5+gJ3dl3BRT55t4uD4bo77Iso2PsY9fAlXBZ2H2NqQ
+X15uRQvasjKMNvX+ZOfkvJq+Q45+Lm3m2xIBYTGsxDK37dq28peE8C/VxLDM/Bq
UixQakwyYST7zxyyXbauuhjuPD6G+/DZaJBuQoCXHmvqSaHMTuTQoOzPxNpzwFaT
6wlC5eZiUjO6Ii0tB7g5XqsfwPOKNHGzikQFfENoZW3o86ufcnI48Gj4ULJkKTvx
NCJolLJ+1CSLt3T3Fxs9x/kxIJdMy484k9MZeGHQNZMht6GJvT/qcTRR9BkjF6ov
nEC2VWR3+DKVi1ZotDvgTr/IVEFwhTD9QyStxzEl6VWthLxlR0FevD6QDxtT4MAF
OtdPjdj621Bc/h/aLzBtpectbEtL+1noVPOJMv27jPVHrmefcsrFlwXj0IAWtL5X
iD+uSEI79mbmq5+1G027W4eco23drIh6Y4Wj/HSTVCm+YfBxQJdzIgQuYW21geCa
8WErfc7I6CpHV9okqUBm1Ug1UfVzTVe12MMUgo7sZ1Q9TSc5JSnQIe4sw6Jb5Z9g
fs45qwKqoD0AR1Pm4zhDPwyV/lqwmwPKOG9cAOSoM4QPh8L5vdePRnLHVVwCOM7A
vx4iDEgiKyE17wJmxQNt4Yf8SdY8k/ERjN9xJ8lHSU5wwc2TeX8/kym0OxtNa5BG
WF3uknvzuFM5DRcZfk9Y7XOpQRqSPW8pAW0NuIX6goj7zb7jBS1tD9o+IQ6Z26cD
mfXp2+IDxBrvUy5P53KchlIyFbT6gpIf777cVvrBelRPAELQ/eO/hkDLiUy+y95d
+Ewoh9jy7L2sgvsqbXanD0K5LuFfi0iejXxWsUMTZGgcbIYO5rLlQ2ljF/uxVqpA
9wWufXtmeZ9qdPyLNsxa6PXDMYv7ScmPeEEuKP9ODSUWNvncgpHUP+khhgXD13+w
3WHz4Vbu50servpqiw4IV+yprl+MfLukHuTBEmuKsSEa8nkbXXKmJtjA25K+5YdR
FFwG7gzSqt82l5IdR9Eln1inz9R0tnm2fFykhzADIKZQt0XqvERDy2NB+v1GBKhp
2nAyEt0YQM+32m57dzuHbqTR3XVxFXVOdpZrAvUM4SBGMLxQHRR4WBTmDIZWiopO
GNvNYPfmyfFmfwNxs8xx3AxcoVv07I7RBQiYezOLwlzptCDDN1Rg/MdqDIcPlFWh
WUCZikAAcwM9wB3ZQstjbyUaON9DWtTnsVZ8t0cqkY19UETBzYmP2hfyltIceNfO
paRaKh5A0QqMNvMmoZQrZuG6uS/R7fLW9tBSmBzg1+4=
`protect END_PROTECTED