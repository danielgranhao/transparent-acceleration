// fft_ip_tb.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module fft_ip_tb (
	);

	wire         fft_ip_inst_clk_bfm_clk_clk;                 // fft_ip_inst_clk_bfm:clk -> [fft_ip_inst:clk, fft_ip_inst_rst_bfm:clk, fft_ip_inst_sink_bfm:clk, fft_ip_inst_source_bfm:clk]
	wire   [1:0] fft_ip_inst_sink_bfm_conduit_sink_error;     // fft_ip_inst_sink_bfm:sig_sink_error -> fft_ip_inst:sink_error
	wire   [0:0] fft_ip_inst_sink_bfm_conduit_sink_eop;       // fft_ip_inst_sink_bfm:sig_sink_eop -> fft_ip_inst:sink_eop
	wire   [0:0] fft_ip_inst_sink_bfm_conduit_inverse;        // fft_ip_inst_sink_bfm:sig_inverse -> fft_ip_inst:inverse
	wire   [0:0] fft_ip_inst_sink_bfm_conduit_sink_sop;       // fft_ip_inst_sink_bfm:sig_sink_sop -> fft_ip_inst:sink_sop
	wire   [0:0] fft_ip_inst_sink_bfm_conduit_sink_valid;     // fft_ip_inst_sink_bfm:sig_sink_valid -> fft_ip_inst:sink_valid
	wire  [31:0] fft_ip_inst_sink_bfm_conduit_sink_real;      // fft_ip_inst_sink_bfm:sig_sink_real -> fft_ip_inst:sink_real
	wire         fft_ip_inst_sink_sink_ready;                 // fft_ip_inst:sink_ready -> fft_ip_inst_sink_bfm:sig_sink_ready
	wire  [31:0] fft_ip_inst_sink_bfm_conduit_sink_imag;      // fft_ip_inst_sink_bfm:sig_sink_imag -> fft_ip_inst:sink_imag
	wire  [18:0] fft_ip_inst_sink_bfm_conduit_fftpts_in;      // fft_ip_inst_sink_bfm:sig_fftpts_in -> fft_ip_inst:fftpts_in
	wire  [31:0] fft_ip_inst_source_source_real;              // fft_ip_inst:source_real -> fft_ip_inst_source_bfm:sig_source_real
	wire  [31:0] fft_ip_inst_source_source_imag;              // fft_ip_inst:source_imag -> fft_ip_inst_source_bfm:sig_source_imag
	wire   [0:0] fft_ip_inst_source_bfm_conduit_source_ready; // fft_ip_inst_source_bfm:sig_source_ready -> fft_ip_inst:source_ready
	wire         fft_ip_inst_source_source_sop;               // fft_ip_inst:source_sop -> fft_ip_inst_source_bfm:sig_source_sop
	wire         fft_ip_inst_source_source_eop;               // fft_ip_inst:source_eop -> fft_ip_inst_source_bfm:sig_source_eop
	wire  [18:0] fft_ip_inst_source_fftpts_out;               // fft_ip_inst:fftpts_out -> fft_ip_inst_source_bfm:sig_fftpts_out
	wire         fft_ip_inst_source_source_valid;             // fft_ip_inst:source_valid -> fft_ip_inst_source_bfm:sig_source_valid
	wire   [1:0] fft_ip_inst_source_source_error;             // fft_ip_inst:source_error -> fft_ip_inst_source_bfm:sig_source_error
	wire         fft_ip_inst_rst_bfm_reset_reset;             // fft_ip_inst_rst_bfm:reset -> [fft_ip_inst:reset_n, fft_ip_inst_sink_bfm:reset, fft_ip_inst_source_bfm:reset]

	fft_ip fft_ip_inst (
		.clk          (fft_ip_inst_clk_bfm_clk_clk),                 //    clk.clk
		.reset_n      (fft_ip_inst_rst_bfm_reset_reset),             //    rst.reset_n
		.sink_valid   (fft_ip_inst_sink_bfm_conduit_sink_valid),     //   sink.sink_valid
		.sink_ready   (fft_ip_inst_sink_sink_ready),                 //       .sink_ready
		.sink_error   (fft_ip_inst_sink_bfm_conduit_sink_error),     //       .sink_error
		.sink_sop     (fft_ip_inst_sink_bfm_conduit_sink_sop),       //       .sink_sop
		.sink_eop     (fft_ip_inst_sink_bfm_conduit_sink_eop),       //       .sink_eop
		.sink_real    (fft_ip_inst_sink_bfm_conduit_sink_real),      //       .sink_real
		.sink_imag    (fft_ip_inst_sink_bfm_conduit_sink_imag),      //       .sink_imag
		.fftpts_in    (fft_ip_inst_sink_bfm_conduit_fftpts_in),      //       .fftpts_in
		.inverse      (fft_ip_inst_sink_bfm_conduit_inverse),        //       .inverse
		.source_valid (fft_ip_inst_source_source_valid),             // source.source_valid
		.source_ready (fft_ip_inst_source_bfm_conduit_source_ready), //       .source_ready
		.source_error (fft_ip_inst_source_source_error),             //       .source_error
		.source_sop   (fft_ip_inst_source_source_sop),               //       .source_sop
		.source_eop   (fft_ip_inst_source_source_eop),               //       .source_eop
		.source_real  (fft_ip_inst_source_source_real),              //       .source_real
		.source_imag  (fft_ip_inst_source_source_imag),              //       .source_imag
		.fftpts_out   (fft_ip_inst_source_fftpts_out)                //       .fftpts_out
	);

	altera_avalon_clock_source #(
		.CLOCK_RATE (50000000),
		.CLOCK_UNIT (1)
	) fft_ip_inst_clk_bfm (
		.clk (fft_ip_inst_clk_bfm_clk_clk)  // clk.clk
	);

	altera_avalon_reset_source #(
		.ASSERT_HIGH_RESET    (0),
		.INITIAL_RESET_CYCLES (50)
	) fft_ip_inst_rst_bfm (
		.reset (fft_ip_inst_rst_bfm_reset_reset), // reset.reset_n
		.clk   (fft_ip_inst_clk_bfm_clk_clk)      //   clk.clk
	);

	altera_conduit_bfm_160_oln7wka fft_ip_inst_sink_bfm (
		.clk            (fft_ip_inst_clk_bfm_clk_clk),             //     clk.clk
		.reset          (~fft_ip_inst_rst_bfm_reset_reset),        //   reset.reset
		.sig_sink_valid (fft_ip_inst_sink_bfm_conduit_sink_valid), // conduit.sink_valid
		.sig_sink_ready (fft_ip_inst_sink_sink_ready),             //        .sink_ready
		.sig_sink_error (fft_ip_inst_sink_bfm_conduit_sink_error), //        .sink_error
		.sig_sink_sop   (fft_ip_inst_sink_bfm_conduit_sink_sop),   //        .sink_sop
		.sig_sink_eop   (fft_ip_inst_sink_bfm_conduit_sink_eop),   //        .sink_eop
		.sig_sink_real  (fft_ip_inst_sink_bfm_conduit_sink_real),  //        .sink_real
		.sig_sink_imag  (fft_ip_inst_sink_bfm_conduit_sink_imag),  //        .sink_imag
		.sig_fftpts_in  (fft_ip_inst_sink_bfm_conduit_fftpts_in),  //        .fftpts_in
		.sig_inverse    (fft_ip_inst_sink_bfm_conduit_inverse)     //        .inverse
	);

	altera_conduit_bfm_160_3fqkqha fft_ip_inst_source_bfm (
		.clk              (fft_ip_inst_clk_bfm_clk_clk),                 //     clk.clk
		.reset            (~fft_ip_inst_rst_bfm_reset_reset),            //   reset.reset
		.sig_source_valid (fft_ip_inst_source_source_valid),             // conduit.source_valid
		.sig_source_ready (fft_ip_inst_source_bfm_conduit_source_ready), //        .source_ready
		.sig_source_error (fft_ip_inst_source_source_error),             //        .source_error
		.sig_source_sop   (fft_ip_inst_source_source_sop),               //        .source_sop
		.sig_source_eop   (fft_ip_inst_source_source_eop),               //        .source_eop
		.sig_source_real  (fft_ip_inst_source_source_real),              //        .source_real
		.sig_source_imag  (fft_ip_inst_source_source_imag),              //        .source_imag
		.sig_fftpts_out   (fft_ip_inst_source_fftpts_out)                //        .fftpts_out
	);

endmodule
