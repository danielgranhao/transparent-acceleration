-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
XRqaRRUeE7C5jP6qqFhsT1uCveMmv3FgEin15iFKtnQCJ8SjuBr0OX/MyiJCdnUW
iOlH4/BKfnOA39+5vnSdPKnGRBt4KPL9gNUZ45kYfAggE6ak0rc2pMpRqbzjXxwd
V20j9P03IEiHMwtz2XAotvOTYB6zXRlQIlhnW2VYdFFnriQMQUGEzQ==
--pragma protect end_key_block
--pragma protect digest_block
3XMZw3G9yzxUIFtU013AK2qOokc=
--pragma protect end_digest_block
--pragma protect data_block
ZzS/bAQv9tT+T5dUa3fbjtX9jh6/KwmD7IqjB0NpdGrVP8O56fmIW2M1rXiueczJ
OCIX++9HmdR2VJJcHp8tqXl0o81vztM3Sbv1cC5Ewhp59lQPa4h54a6whdOJsQy8
9g0WNPNvzEjk5M4SHyAciDGVcT5WVd1TP46s67kar7tH3cwiWhKEnOqLbF1mHXR5
7+aZhX/i6ip54wEBCxTUmj4+v87ZlvGOwbLZGxxU+Otx4Uwcw7vecZGZR/26EhJ0
VNYcgi2oTPiw0UGtfF85Nhma50x3+U03pKmKrAOFtwkjUtPwWBVKq0vuY/LRrtUe
xMQsC3BdAc4SPwUchcOQbTvW1zbBi02SY9q6Hf5HJpdNgCDmLs2DQ4YgfRyV3I3d
VX29EfDZgU9FvJirIflilTrO1x9nLcYxkSQqMY/oHHe3gqUflZb2IBn6MGbcPLT2
mAuuW8ZJfXvaOzZBgFoJz2dnzxTwCQZvn12E7x6+J/hyjLpYO6YQL/P3/LrCOXD3
xbfiHEYr6CbDZ9quxpEIaHfXrV5+16Vs9Iv836RMJoNVCf5bsQbq0zAnVxazuBgg
tZ1j9cCLPK7NhXW2SHnJeezSxQQcR8jQi3XLKXm9XUH1sSHu2vmOaT9Au6wbtj1O
Co+TZHlY6yROMARMTCUoPq7memsAoAtGHz3NZOdIb4WkD5jY79WXTN/WsCioUA27
CaAoRDwdvN4VsCV0wDg6MCQIzqMLr3thFoZWAYHmvbNjPJIyjlH4/mwq+K/MUy3X
3M2U+zP6Pl8RO6+eIWum0IYJ4FNkvSetvxBeuWhNfb1zg3DYYPfYbB9NGRrkDsF8
Rn8fIfvqpybjnPdqEX16KoNGayCbQSDChzns00jtYQKML0kc+BuPNFQmb1I+HWGZ
jJ5mwHdC5gT6BIzqDBr1P3zyN2tv84c/8hOX8cW4xVomduHhaCRdPL5Co01Kb+JW
pLpdunc9IHqQQLYcSElpovhGFbvEDAYO2eMCa3ohxcu4HB3a0IuSWfXbz8eykHUO
x58Zjli4Y+5h85qJEPnyw2ztxckRkJCEF8Z4anJqVxfgHoSwulGE1D10Ytx1oZAd
CTOe3ew9LcMfUjuGX8+VpP6kNrvwapt4xkvmG69njkZsqlq6vvf+y3RdlMbtMdwM
3kE21MgSLVCddo6zoR8M3VF5TRcs3Qft6uO+ibdibgh2TJgtqJZUnI7+JqbiEkrT
j83+t70hB+Tm2wmUejtuKdnU6vPJRbdqs+NlwL4OJATwCkIkieKss7h+fyHk1AW/
7D71FkoSFSdFgQDk6VEANUpL5KSPpNT6sU2GDZg2r+/7r2SD+LnG+0SXnkLv7Qaw
YQ22htvBdcDBKKlp4SHDMGnMrPjr07+18rupIkAa7aNeBLqjR/ythSQtGwQrz2+n
TCGApcZgHU26joNV6LFOlbXmXVjqcV+HzK2LWCbG2vICwEUfsIAYy+9AB1/RLXXy
vGln7Cs8pu9j6ndPG/5iFlFTLL6Cy7m5ZyKQcz61af33meLHhT4GW6wSS/jN6vvQ
3nLIs4WN0Cr/1/ncI+dzYrBJsNmSjGWIOWBOk+cqpE4sH+bpXkMfihmvG6Cmokvs
GGSvIhHagXPYgRE3ahFTJykYzBJn+vTjNawDvLcfR23vIwv35zTl36eWTvcu/lj6
GPn7b6AvK9RedrxpIqfyEse9Pu10R0CzGQtRkegnpnBjOD0eMI7i3APELAoNOdjE
IxhFH9zFULispL80a2+uwLZx3IwskHUIYZ/g661Bth4+j6bVKzaWcHU4oSXrwpMu
TNTzUK/CremhnqC9ad8Lf/y3Dj4iEvExmzPsXo5j1KSfkTuahEcqNK30kn3qY+41
Z1wKYcDhgnjwOeNPk/NSONZdu4bnCSOeLRuUzibhg8rW7T0FPApKz/Fn9GuKfxad
z/uMvDlpEFw5eaCf4wQmd4EqoYhud0T7uQHJin5hbi2bhO61QYCigi8yb/LG8H+N
Su6ZL5wmYTBTrp5wdZVLl6EJy0o22HITmTF3vnSI1G1g4jc47caA9miwqyi5UZzZ
00bij8AtSdZeGn/tZzacnaG/lgIpX+MxGeKTDTl9wqrFLMTG5q9fQpKxzKL4hi95
OiwNKDTomH3xp5tZMHc7TWZOIWSmdqra7xdc3hjYNycikSiRVuU3O/x/L6PiXxCb
bNenkf9uYfcFiegfBzj5ekAPlDZ6ODwTJp4/WefzI40bUcyIfoFKi3iqk+5LwIgH
edtFENJifBxM4xsyPF+CsoVBd5ntZZm6xEny2t8pfNkUfHNoR6ZExVFrq8Y09ZQx
JkXus5KWuSW3pVpmvaagr/uI/F6oGwqQqrDGGsJkMXVb4jjPEA8TmAn13BWqryLK
rcWYBzFOvIfLOYeaywSx9CFbkbTVtWThlx3wHd8XtI/YwH1HEWuBCiWLAb7d6TWA
PHH5/Lzp0A4Wp2LLO41XOk9pHgSfWku1OejnQAZ0LhA8clpq4vSe/YJ03AqVmj8i
aej7vjlfGWsXuLSHnm8E1pfDreQ6AlF/5G3X4wtNROgAzZcDw++VjZGf4/SmZ6r1
Nk+tou18eiEiTtDJGMN93mVWSdUrGxuC/1H4T5yGZwdG3w9olnwMk94ae+BD7Niy
58KRigljkLUTaLSCCytCf/MzsvDVOLGj6mS6g8U3S8kQ7C7jkpNPN1juW2UlBMNr
deHuZ91erqVsjBjIVyul4aL4UW3/vdtJh643hIaOqi24FmhPmHHHzjNtN6IQTEhR
bVIgQepEmASmYrAbb6GObtCWh2ZVkWK+C+pjNtvEy4XkWr8Wll+NnrR9Bprn7qIT
Py+wWQcGizzLX4MSPzNIp/LoVyCal7gwfEydTvo7hsHjGSMDKjbRMLlaQLuCvhrl
Ws5COQtoRF6h5IFMHWKYsTK5DMqjxoVlOFoNRjgehWeVdYpRP96e2Akah8AVJn1K
0VsuE22DC4lKE5OX14kq5AC9z0PeiEjgAvYvSTXXo555gj4J7YM0ehyenRThTNcX
K3uDXoql1dfPTidiNVsH/+8GTk98dKflIUTNY7uRn3IY5erDVXLw22fTncXx1gJ+
V3SvkMWBv0nmNs3UJvtLsxs2zqclNdhUM4DLbLQW/VehrfZdAeiT/TrTIWFpo8Dd
LKUbOErL1mA6xF8MzgkcyRED+TYDGH9I1qAeCwmW05H/31fRxRaJgY9kaC/W7CCu
pTC35540D33hpAq92lJWL7E4zPzpa7Ij6Am2TeZLKoio66+jdJldGiBfh7kGs7It
6GOQBTsfbd+5QddcWQC1QAAMlLtGttMfdScizrUpWSYlj9EE89XQ3Y2FYGO3yJnS
JpaZvX4CQ/5FGm42vWzqkXexBbwHfFQTvoubo8FiFnXOwLoXZ908xqvzVRXb+6nv
sG0D+CiFEW/Z2xy72qMGuud/0NkE7teTpZcNyZaIW9Q+e1F4UXbfKAekLM41Qih+
qccQxBO71GykruER1QCrE8mxr+8xPHDqNE+jCMdOMfbGRHpWhZ+xi0xLvFM5WPDm
AtyeNm0qCNt/7OgpGJkCdPvLKSakV0assofz2p2v/8ulWTHPm4Tktq66b0IcTzX+
IVaD4burmrcbbxPDdVh8/WBTvykOsKeedRbPI8CzB9ZHU3KZhhNQXANOf/bu4RE9
UHsXXJvckaD16S/2JnPvm6ItezdBb4x2M/q3nlkwEmafCucMkPKof6BflNPw/PC/
WuD7FACUvk/rXnmsPi7BfHekkaL5w4osjGSe4wgu/DE6Sfzs4Hb69t2Qs3IH+Dde
ZpPr78gj5CvxMUZcRDk0EDIeADNWNINmSYlwx32CKh6bHOa19oIEoJUv0TpysVM7
0h/KQUlu6deqBH+DKmXKlbkfJN9+5UmCdg9cChBdF+0suVDDy4aQmtctZRx5gUKB
OEzVhbu/4LIvr7ruNoylSuPs7r+o9LMBz7Gq7+13x1h7CmI0KrixGIyBthScpS07
ejFFxxEoM4rnKBQ42ySWgEo+f5bk4QdOwSX+LBzvBmmx1CdkNF1AbOaWJdJp7aqJ
b94aCDJ1dZgh1MdcggHqHXJg2ZHxS9AZBDEAR4lQgVgE1RnmFlY0NdyrkLNx4L5e
jOCfoZPTRcvYZr87DJI4iodyL34xw1lkplQtjzXonfS9DgWIufXInbgy4TOAoEc8
dhG1slEvKxtRxJZilIfRxtE1bOk2cSyudH4jdi8FpLEHzH7vol6q9u/LoCUnVUyH
nlyeX56jQcx0tV75l3k/lEcrz+UlUFAlf6W+FHu9q8Ynoo9HIXYz7XA4c3eW6LTn
G5u5NAr1uGEHqd0xtb1pmm/KMY7JO1ZdzggxDrkdSPBKU++ShuFivv3QHXP5ZHoo
OgscF5pwu/vgBAOAHR6o4AkQp1g9NinVvjMdQxjIxxawVOUd63f0n6E0HVF9mID6
R2KHcasqf+nIwD33PmIej3q7pJy0AiAZ4NmcrH5zADKzlsZhY9CNU9Of21sFf8xi
QMYeFRHZWX9mh7i7CYyO+j0nHrkipdh4KhyiAEAKA9ilKTso0F3Why9WnT4N/yeW
5EicbwuuGGjuj8rCu798qWh0XeF7tbkw9z16aqpdJYkvqdgLbR5Ifb9ykOhF+iTv
dZ+nhGF37KIxTnDOz6aXKdHuw/ZDKlzduRyc/AnrOLNfC7yLHM7meOsPT0MrGJ84
K+yZP3luIUfurHCHwnZHYlbhb/FjLgNFoJv7GYA8qm0vkEL9v9J+tFNvG8tB3OMY
BRvdR/rIEj5t7Je8bQvBaHkzMAs/DJvuHwPCy5PZstjpWtxjKT1Kx7isfRrv8U5g
SehoVbz0VdH57aZ8oIktK+YH4y071LCdn1eEK11uKs1Z3wgENrCFr3rVS1hr0czR
skyC0BP5ajKHO2hrHK8zeHprIDwb7grIUHXbRwwJXVUh6MFuk9KzwcVsP6+3WSP5
0QgPuxNnBNLSE1Y6X6IkpoQnZx02mpBj1Rz1sjnVa0SUXZaFUT3yUcIV7/ulXVX+
jrNCE0+rs3nHuNV1EruMrRHuYXq0CM9gX62tNCdzj8mIpotCWC/j7vKGSRTn8hi8
YgAjLZM5cjLBVbGWtR2g8SL5AqAJG1XDaxNMorwcr6tQtcH5eLSbRll/vggpLMQy
ODHUX/ej6O++aVHjhtxodzL4E0hMCZ6or/KbGKjPqYVhnhMY+awmYlU+RMHtG+sa
rjfPmlZwOR+9yJKODn+9kZ3UMqp9wVelHhgC+ZEunOr64oi9ZM+AngOILOieAhsz
fUbxxf8T2L1vh2Rwt7pYgtIb4k7k5X2DE5o06XrsoD1fNgYa8DOa0KJwTs1G6EEu
TJJ5Pqd2xuCHhAwvq43C4NDJCfTsXpgOaib3Q1Z3acDAOCT1qkYNAq71yySzJMKq
b7RAmcK1azVjloX0ae95S3vgoEKm4bazwqKPOetk/0ae49oiRECgyFBAEnx0wa23
WqiREbpc56p5kirp/DYm/D4FNwQBXvw5KunqUKwibjJIe6YMWzo38dCZKEheksgX
BLzwQBSkRai3Gnx3eLgCQQvgi7/SFXEAfHNGQkf8LXRxP+YvVhmKLPy4jnFWYg+E
wK8lLWhUi5erPnD7nJr6DdJjYJ6tV3FTRDGT5CuGdHOfCKI88Le3rLcyDB4KGez8
pmCRkoNinFIiRCADqSNIrfSwCR7MRD1q7YxDu/0azPUZPjE9fMaR8R42VFwoDaB8
Hq2d6qMv8WT+A2xUdh5kcxlAEqQIU5XSDm9dTvOmjBrKrefnaQ+MoI/YAA7e9WwP
BemtO+11jLjXGzMzUSNlOsXai4yX9M+H5F4ZAYqbB9JUiMmLotyDo58l8QN7RIAZ
XEqOGX1ZglKe9V8T1E9ps1AGPhC2qWzEd9JSEeqA5FRXLiTHa3qwqyGZXQEkZi9J
uhmgg+OkrRiZRHyxVVZZ+vtwp3u10lqVdcLmdCoveX6SJsbGk85D23sA54RdU6A5
BkbvUaosGlizi8GpJT10FKuf5w63qcHinS3DU0chHBUutitd5QW3kd8uHiWIpfzF
bDpGpb8fV0DiWGa7gyy+Eq+qNubLY5N8A6Ga+L2k/O4uY6D9DJLqO4+GRkjp0eLZ
9yeeV07cW7Psy5/COoT9jB522aGBG0njO6VqQHcY+gvsPkJUU7ydrD6QCX1kUe5m
VA2IkXE2xVZYGhTaD98IaUGsncMyYpo/btVg64vzRTanCBn8WCKex/+vYn8ohs3/
FEgZ6vF4qLljeY1lZKeIlUCsjbqiSjm0y3+oHCVDbrnS09zG8onmE76MNssgt0de
+I8CgoagdfmhlEzMYd+csdf8+hOFMbpPv2HRiQcyYY0+xPaeF29r8Gchty8zTeLA
5ptXjv/wjZpQLyQTo3iypIiN0+rPYfd9oMBewQLfwjbSjErpI9dFyKujBV9TbR+J
JMO4OdqiYkKY2jHICWNMYdySoLBcsZyL1P7oFRSsRxzKFERvmzhgwV3f0XiZ4/Ic
m1UNP7r7W5XGjWUzjsRNh2vOh5V3RbSkYYXnt+4Y19VirFDbmzU+D409/MSa+BfP
7x0Vh89wMUI/0SbS2Q3O0sgXJYdRl2Jnw40JjwDCHV+PfNWUbLWhJIHPGlazdTQZ
VjeDjLloDsnFHtZlSWfRpOJu3N77JRE9o1GHXD9kVphZtLygQfj+Co7A8GshxtEB
FdIWP8z7E7z+iVniRS46mBKr4psc2z7AyR68HUHc+ahNtOZp3GVhuStY/O6tCJ4p
hhHuBVypkfH43vitCLO8cpiXLawh54NtphBkI0zIWh1ygGJs44EcIWGlrtZ3T4Mk
4E2ciuKYS3Vy9y7OjT5ZgW1mRAt7Tya/5fwxMr2G352/diE863kGyW/TMHH+w9ZJ
eoOVJC0vMDmYRAjP74InSFrCtXlR4WOeBgZ2xmhty4CgP+vlejKMfOpUrg5ekumT
5PJPO78m2PM++Hh+gb7S8+pxufPPTRR+dwixRnSYls1LK8OA44aDVaqvmQhrdSwO
v481fHRDI77IpzcPhCTzRjjUGM4B38aS1qIDARdocK189Fa0yi44jsig3tcB1zBA
2i4GW0763bdf+i8MLr8ntluyonHabzznKmYoNxS7WQum/F8hcy1oFoptoXyhkHC7
WjRLqGvqNLrFIaBZjfpt830fniuRGhdmN+TUqT1LXdIsN+dJ6Jbjl5g1bOdV1iVn
ZjJxKtzkU5H9qW/EM2GdwxpvA98W8O7s+xPK/GYloEBTzLM72RybALK+lpy7+p5M
/fE25jj5TsxQqkacrQ5/JaTDPocAOT+bJIE6Md4z7nZDzyzsWugn2qllW/uF/Oho
WJkgAGW05DjsYrQC4x3eQAZFyAymMN8robJvhcrENd+3rvdm1pQEnlu7i5n3jEwC
DTXY83MZ57qIPN16devuy4WN3oXxM86Huh5OKovcGIzB7fRqJVtMSLMCoatjE8nP
0dMXmDrWs6SS5FL7Bbv30e8l3QN42q8qCbog5X//woR+2qH7sdKxWYLewxFm/zV7
qzubiMYD1dqK+MkmnMM7txngIPYzjQzclGvBjdgMagYmL/e1fGHjmWhTj7MLfnJb
qlK7rMcQxKJiZ9BFLUIYdDJxMrtF/Nx5F6gsr32UsfdSXdEjH6lB0E2FW/6Yhbuq
LzVm3deBQa6YI0Jq+/3Ecut36yqUCdxpeQ+FeLmgO3772eM+FbH8It1gEf1ZugtQ
fE3wCJeW9R7SQrDf+jIbYr1onRa+NP8+RC34XqdjFrMvLWDSAGsO3I831td/opF2
O6707Nvdu7BVobkmqtG9qvXaJjuzgnEuSNWpseab3RqSkPvDltoB6TUa3xd5HnKJ
4h6ev7MWqD+4Ey0punqt88RCj+bw8w5q0im+EwVl5D0M60lN2jsSXjWNw1v8rcXI
6FEhg5SYMdRzjeo111FjqNOu43Gg8ZdbpcbOqTvZEb3C1jMMtH9OG8FTXqzwF/LJ
GwOUrT+wdIeYI/iA0XKFHHJ4wg/tht+WvtoxKWgj7cQYR6FGV0rudlcZroY8hnPO
ZdDNa8HjuEsahzfsPjVpubL0JK65YPW0+d+oBifCx51gJBzQqoq8s5B/hGg66bfS
cQlf0wlXqUSXsNp7Rm+7fZV/YKs+HHxh61Yx902M4YjqjMMntmkeM5DyPcDGAqR2
iz0Iu9X1BYSe8OC46+PQy4JtrcI6m/x7udym2mc/nzkZ90YXPDwKoawiOY0sT1tH
rdb/14v67PDFfHP9j1kjZjwTEimrzfEM7blyoXgqUirZo8K920nbN0rYBOBMlmyy
ipITfdM3IXqQm9ZQ2d39tm520yN5+vltevSwbpdSlCO2zkkBjcblGk4PrynidaeF
zcrst8wPd67VYBqgCB+aM+svZgqNUeC6u0B1vp70vp95EPmTlzN+6pczziP7fxK/
9Z/fQj1x8wwNBmLhU5I3PDndEncSf+SeNBUFDOofBMeLTfMsEae3iQcwQgeSEhj0
0GXQukG/Ajmo9W8qYPxaZRqx/cCd1IgifFf6p4iK7/M5ygfbKbymXn4ctV0/drmG
+f1/LpiSpnE4NHAIG0gaQka+/lNLTdMO/b5JyBLWC4gLQiTL90IWZ2aupYHvhUdP
CjcG/ybEV9IKQ3fXbuaYrxwlB19tePXMuBA8sz7qmf2WxNGlhmzM6C7PM32Z38Cj
jtwvdT/5EXSE6byByHEniTQm+IrjJhD4W2tK+jeA47k1hX+0me5yd3nzfh0JEzLt
iFKb8Q+lgRb05/alZIscOaj7mrR3XycRd4Y3qzh47BZVFAkQUPp2+K2oxYWls/Aw
BDtbYkGsGjFeeDpIZB3ou/xNQByrSkBe82Ct3q8YT+8UOv9gK2A+ZIXC0O6uF58I
47S3H89yA0kgwbTf0usS9nzjVqtUIew7kEee3QgNDgHEndUk9XSienuiCJsS0jvD
U8upDJzA6hHpNlUMFaouln/itiee4/AD3vZkvfilg2bCjK+kbIV43ZTALw82MlQf
hQ1aY7IFo1sdnT5+HlDEPfxs8srKoIbd9kgXtvBWa1VXeE4V0lESQawaRIp9QI/W
qt64OccbQNkiIOEw6TChjzZ4gv1IfV9qm/+Fx8r0+pOtn09gMAMcPQWJq52dd9d6
DFpBjhP3oLyZcDRwWbAou+hk/8sJHalEo/0Q+gr/4e2ZR8R/YY8ucONojHv/GwiV
DiV7PhJcSPZ/hpVlDohInQ5xQ4IJwnkxH/KWVbJimbO2BKgl0OSiEVxfHPtZjcsO
UpFtOxnt760p/zBZzm6ttgqgpveTFXOtmXVF6+DKiPul0szdTn8hYw37w/pZvVY0
nVdiSA0dg2O//QuusBnGkPIXRhw7GTLoeVuKIsnUik2cgrNa5jPxz0i3AYrGTFSM
yd9XpKPOK8cSPgls03LczDLfubqfjfxItREjMC3xmBw988QVQYsDQMP+NeRq7PMj
jJWmyflan+mI+KJct7J04IjNu9+rQHeJp+ttieDjU68S64Q2Tk5S3IvgaB37pv8u
jzTbil0G81e1tqJ7HigKWx29PNvbJql1fOYNBa3jzD/fEyDov+eVQIBbbpoF1OrR
82ZIc8xVE1kikriP9tKW7JWolu+/e5UgSLeQDZKyVnzrJ/K4+CAgsGbk5f8G6lWG
oAkPazIlSep4PYs3gfrVrDW65n4h2PHnO0cSCt6EvPGX4OoBXra1fT8HrERfAf2t
zLqCyfoIVhBJuwpWJntME8E/zZNqE9bkIUJeol3cxmH0I8KRI7oxvHUCfCWtjER1
Ktu7zt5AvFGvUKyVr5oUaiT1ku/tWBqGQa/4vjW6sZjHTLW5POLL6kA9sPFi0rUR
fQ3iZlgLn0UYQZGh/dG9IsdP9I2Au3R5nLwWekacgc67UvTZsG1euMJG8VUjAhBJ
ugtK2cxIXS7LSRSkb6Yixq7Hnq4Zt/xKelSjRdoXdbL7o5cjPkWE2bb7/CFKIWPv
9wkXlDGB/f5e67kLRLPxPgtSxd+7IyxjRJ/Uv0DsKTtdqZgKMb53bS02X2OkrPGk
UlSlCbEXW3WeRSyCtXQjLgg8lV+WE6F5TUeN3gxunBPZ4kLD9ErZ6f2qNtfL4inJ
tkF6iecfiMza4ZgYRq+RBHgfdA1RpFbtIypA8nrzFPz1xQYzDHzYsVov1eQm4prT
U7o5DOSEg61EGvsiL2g1hf22uYUgvV3ZgRNuCaVm4h0rmMiyf9H7YgKNe58Mt2cm
N5KtbUdKgX6RQySUQ7vZtVykj9JnqgUx3Z48RscuMCbJXg1T+BYnGQYdMETkf3GT
2+QVXjdbwdugEPEUo0p81xUoL9rGhCYx7eFCvm6lImp+0tvLtR3/SHACUupyaT7R
IRXSOeb76Q7a+YGMmJLnMsDG3JNZS6gjbTrQyBRbkfwNwU1uXzyioeHZP42W3v0Y
rdmV9LqW9oD0L33i5CVBg/HQgVw1RnmHzhZtg55pkGKK0CiscALXUqRYuQxFmHPg
uL1wU3j0HKe9RFWi4FQ+qUf670e6CBWes3qkBFlm/RHOAKs4f8C8D1aHs0FbMkyX
B7sBRs9YDzcDc4T3hB5rb77GeNDGptpE04nZhhH4N540COBNUJB0nAYbGQTJCmQI
XGKzeYJJAL0yUIpw75h+vjiV4YQGzC3KEULpwRitstO/2BvUO3MUj4lZNDTQxNWa
rjlAdT6tJX20jtoiseOwRiel/fjvR+jpObUHkk+1szCNfB2bs15G/Y1kDZpKwnkN
kB8PUcfKlltFUq++chwKsEnu61VR0wSjc+LailAn9aLOLMUPoID3BVqhBU46PFks
iHYcV8kwoCXRYtdLKB8l6roDK2yXS8r5RqOrh0mYkJllCxwHZ892oisR94tyxWGG
LP2cgceG/wwxqZZdd+mylPtvRhChyt3HmtVgLoSYHjez/qJYojcQjuJI0bLiIFhq
Mg7Au3ra+KkLVEGDtxzusaup3f96aPEce/lwH08jQML8bQ7jvEjktdsOt8bpS14I
AE1SojuYVzt061mE9BPL3DO57kiNzA5cxpx5wkMgIidw8a7+VaB4X6WMZWt2DgL2
MstHViKBNC6Wm/XllZG/eGsUJW7a+KVCyba9/tCyd+HldsnTNZYbG+OU0rYdIRVB
AVSRGnqLD+Lms0WsvLspCC9t+Kki1Xj21PUqxfi1AK8qPSDRACi40TMxp2K+3SKH
2eqGmEJfFNAKeMin8QNF7n9eUiQ5ZrdQj2BX4R2m4+up6387zw8CMvKpddXD6fz6
3Dm11qKAwQJVENQx8sYTxp9AMXPuTzEYLJgZ9pEG+JWvJh1PGpEj6ID2lYPGCOSh
x0+tP2P2t17df+jfWdv6jBn9M08m9jkzk6HwLHfdArPy5n2+7LgPyqbQ0J7+ZBQd
N+c8484iyqEay5f3gc2YGk2sdfW5L7JvWjYffDulGqKh65QzfHQ4MSbj25rQOr0E
KWeB0hAB8F2fURJoE52FO6wlz8Dcc4Aj2yoJvuSZMGqLB4mLL6ANcT0ZjYA2D/vA
UMF55mQgwEVk4+00yu/E/5iBYcIaYncJnjYCvlxMlC5NZhUAf3ah78GrSOJkjgw1
B8LSQ/T9uPHUp9H9CI2cSrKDL4FA62NICcap+POevDkQ/49+XrmDawN6EU3vfvym
o8JR39/6Jrxm9khOOouE5bwdXhv3laoQGU2ZtDthp1rpr1uhUpB2cMSgFtXfQaeS
7+4n3GY4knwUTAJk4zwR/6Mc5mZWgTBIzWoHrKnOdlUR4+gmjFLO6Ds1rKWoFR0E
Ignip9DQKTTH6tldA21oUU6XssspH7nSPwNqcqj2570fOLrRs8PhKSHUQSs4WAgu
3JsgDWyv2QyDe1J4KHJwCh9ppwb86T8pNgCBeWYTN/y0L6sOwT50qFEeK2vkYocF
Bkm8Wb5p4wBRN6EYuEY5RqxwFUC8D93a2X7OlcysJc4XPjhqc/B4BBEkCKN5b2v6
jf6e8BWHHEbPy19y5uw+jLg54NKStkZysRd1jDUAgGAvN1cJ/QFCjbWFe91YystO
sSeJFcdd1jgSrYL9uIcAb4xcBrWMKllE44QxtX4eBd4JrN7O0ETgNe7UYaCMPI+P
squHBxruxVHpO+44GooTwNQsShmW5eIglhiPDIru4b/MSBmx3zO/GS3dwOzQ9/0E
QVPpHONypfWvxkYEUcLeVLlNn3ngpBOaWyDeiT82/QDZWj7cDQAbLHfxFDamFMR0
722Epll57CT34+woU5jIDSOIi/VHFQeVPgkkD5ayvlDBZJYNXMub2GDojYVCg8eY
dVDjE7bGEi/8WvtE9CHTwoKIPFiG0IiWQlulpXQ7rqAl4Tt9LZi1RUfp88GgbQGt
rMOmn/dkLrwtg1py7bxtRdxpBDkAacW/V1ArvVU3UTOcbzi2Fudhd/Jtd9w5qNWI
FSQFRaMFgYA2HWTUGWfhx0cO3QVSpuskGt1SNa3OvwMsrIP3IjDK66AiOWdPHMp7
iw+VFvtyAVquDiB+Vdfp8vkG9dGEQJCOKyGfAbjcfEiK8COunsoilrYi3/8Mn2vw
kWo12XwIe/BQDhjBY+asoodcHuWWqMHlQENuqRcseO+uZZJwugD1LmvGQSqRQjjm
nH+4BDQtQIxfcTqG48Dlyo2K8v4AM8GO7FrdOw/t4Hrigb6Arpy+rB6SJIUtZFLT
hlyUsF/wW2sWCmLBoNuMgNVcQd/63ZF6fzQi9VCD3cVyqaTdnUqJY1/rX3jknabg
JAeuZApyLYQglcU140d2QI+IyoNmqadYX1LBTFbN2jT1HzsZQTRKeRVDBtAjVklw
SQeQzmVstOqXPowJ0rJd3eInNy7aqlgYmIujsXdYQOZLqojCQWpbgRKOgzW15aT3
Oa3muSBAkczF4tjTRb8fSWoLdc7Awm0uD2fYj+/hE3hrtZXbXzVuS2qjUCyBsNQ4
tukhrkCBWztJ947SqnN0CKTAuVGNbi5Uf5SrjBnXRzLaFK68D1z5GMlKImkoF2lf
dEqcXoHZpyOxxxidqxHsAbHT9AWDxz85YgjG+87LlgS5raeMqPbil5W+bXyMnPfE
9mVrzQcVJjWP2/jxyV+NL0vDFwYDPmMlKp/EAyFvKbF799ERdFHpmrkJFJi0LxZ/
Qr9QEdLyW0B1+aXiFynVM2vxDcfVHcsV4LW5P+LnhbiO8AOMKg8yySMC05lrc0Ym
ozwqvG1N6KxOQistf2BoAdCJQA7lW64FoCtZBh6SKHZro3gI8tcGw775I+JVQxM9
3neaViZFOrmloLocRnxQTVz4Nc2OrQQeYrdyoIMpGfDWS2mbkRARGExw7huoJ2X6
umPsfDH/Ey5wanFl5cpcQVk+OJJa5BHD8+3oh4s854Q9Zrl3JcZ01b+5gLN9dGsG
bqKEfp/YfYx0QxIg66mK1VJBBR0S3itzd+vvSAPQwOzMCSHOj22aKph1yHIta+gL
+MJH2gP0n4279Px/plUnZfBV6ZvP91N9f2bBmtEBmivs5iTzwo7XligQ6AhONkSz
MyPKQhYlbaJB7LaRosa6xTqLNjLxpAMEbl+H+M7oWSo7NR5XxsDhsRkx6780bOX9
aH/FQx7YLQuhfTjhkz65svVjBLNy/2GyyHkJsNHm8BFrlBloQzPxStAD/Rm8J74r
M6/OZMPayxnwJTHVJNouVV9p9FNWIobtZ12DOFw4v8HsE4iiVfScQdb+W3BWx9bb
TeEbaIBPY6uNnFyrkFYXlk1tLzfDymR10uI4FVJXkAeguAvssXp4JmwLRzpAH1nm
E8vfqgD1oaniHDMfhlNvn/BQekFnVbE0D7jvduHV+d6EtIRRSoU8IC8zEznWzLJt
1cWUNr/6vO1DBj2z6ZtD+tETW8h5oWDRuD1svre3c2R3r1VYNVMcBgbKcobojdCx
t2WHpJLd21WWHXVvmScaKcu8BqVOhPqdm113anqoS6fW4aCuPDIFOmg395ksuNvZ
23vV2rMzvdke0HGT5Th0St4+MDe4FYNr6yFUcmrRys0WZqQpot/bAHldRdru+eEu
a0CRDcOtf5aedu4JzouXTYcYRGFF2XtBC+FgTZvGftmsLvUUBeS9ynCFlCP4QHDM
KzlfFqUpQLc1XdvRON3j6F3kdpelRXzcep+WZvvCOa15UkqT04FDn/3VjfmwuXHk
sh+jIzOL4YJFi88tT6zFYcfqRgkGPDyI9OSq3/WXyAUqLxlzyk7bt8Onwm7pEl+2
7fFCd0Ppu/V/R5XGFGino8Q2AZTNVdpZ9l/Hll2hQ7PvRwLOUO0QThbnXVJimtdt
aLd4denwZnbWnYsgbaTIiO+2M3I5Q4TlF4w62/7nDjPd1KCuBO5iH1AYmFWkkbu8
ZQXULyBHOQ5S1w7BcmctLHzlTRZ8SbzLjVL/NFxqrEAH4OToFKr96P3Dgwk1S/nu
uo3BknhX7fYkQnIMiHW8iMzmyQbNnsH9y1nnqa+HzF7k6U6sGazhcvY0lWE5Yrot
BG1mW9pCWoIUY4RKJUCOZG15y5s0SUzG69fq07+3pJuKcM0hEkGxQGVhKj/Op8Rs
L5rucjypHPM1DQ+/PKxy9xW3zE9yB7ZZMc0AEr3QWuCcOI1/JUNqsAADGpN/KnHw
vPLvok1sdtdApWYlhi/1GBIIekEiUrGtzLS7hXZt3qMHyS9Rl9bEu/sYDscI5CBe
zTbQmAz40DaANPvq0SJN3b1aM1JqpG0cq8qO/L81dsK3rHZhvjt/0h7y1fY2P7gp
eRnFj/0UaaHsorU7+glThzkOU0BoCl1YO9/V9CwtNBOnHcHlG3dT4G87C+M3Aah8
WQRqQND1qoDfRG+Nl1jNaI526/PEO7rpl/GqbHHNl7ZLkPfEYP7m8qx3/xdH3y85
tGiIJP5StO6klFYGo51M47XXkZMCTXdWTIK/Oex4amXSKy46hKdYcUvp+vMS9Bwn
mSvMN8U9x+IqzZY6oF8ux8XaNld9EnPKr4iKar0kTNdZ3JPmtWYo6YJwsQHIJMr4
Y9YY/fpK4Td8os3S/u8vhThLJFCLf3FkXmuvrbQj6NNyIzEcXUpHvtmdwCtK+W9Y
robY79+GxLMmr98kzVxFGdHjvw+Zcuk0MIG+lhcDycYw4K3hoD5IwpNtBZKp2XQB
a+rxiT526E212Zi7dhQ7gywHHOs43ag9pmZCjnBKXwLle1anMSNmnR75RmeG12Xd
VCae74noNeUlI/jqUI4nU+ZR4Xp0idbgyoGYBD88Ml4UWKtMQYv+9wGvU4K61Ju6
lvUjCCmEI5lBXIVolIF26tS9cfMdHzXOmARjO8DyBba4sAfaXDBvC3fdSg82xN6h
mX2U6whSY2CPPVoqFB4s0ojV9yOr+iRD2AbErNBy11u6waEIEygClUkVM6oK9hKZ
BR+FY676GMAx7sHTd9wSQrxmF+Gng48+YFt27DL4nTHwW7+RdqUai6hG88B41lST
7SFKtqr6iRyo/uZoL6poQffXewLxE8rn93dQXDO/yDrgdnqhdk0/DhOLdd3p11zX
x8UN48KyUnbLVTSQrKSJX2m/LYOmtNSIRX//JlWVKh+uyh0uhToPk/jZD80DdpEt
dm7sB3aBRQXYegfUXj45YB4I/EA1jM48ixONRbwJ4MSFN8FA+/R/gRppIvb9zk8I
NN3PXFsaQJypKWpJtOL+6wGfqc6bdYoHdDqXG6mZfjhhvuVnH4f/Mp1Cjau/n3Yy
QcHFvARCm52dU/uvcu3Ty8fco2XUBejt+KgKZJGbAfXrWwIL89lRfP8uV8U/76ge
yMTtktcuzFgC78JM+SJcOyXJdrV59MSe1I2O7Hp80GZIGVpht5eBQjOpxPpzuL9v
d01zG4FAtvqWDyoybJAEL8iENfTikXGH8zzXG5qC7LreHCWEp3BUrYr9jgCBE9Cl
yI/KLM4MnNLZhDEQ66qIxhALUmzFMKfqbXZKb+4w8JZVF8sS4HEEI5wuPmjxkP0x
EXfiLWrObdqnh6Mp9dlCBnam+EsuRl8RXLEPl6tPBMWsNOiES3DKi9gNHwF2ewmq
vo1e+nk1noxgeyOp6zCHlPZK6DiZZAyWltPYYuXQEUGu379OinItFLNgFTP4W/+V
TOtxl3Xtt8R5jhTvseK8YsdOq5WYoLl9kSk/iTSBLVWjwP/gn7D2bLYsw8TuaHPM
bN2M5BXgKYJ/syB4fDwrr0GUThOj+KpBQD3uFx5Eu/3gOcA4fsr+hp413CSXLUd6
k5XqLDW933S7ZQ4cNfG/65WJMKoJP0s22aLFkCMQNvJD9CccVLrV0v7m804/ipTI
jSRNFzlyezg6mBVs40GSWessxQlR+JLuvreP9OC/LGmbbI+n7u9rFTw6I58Td0k6
Hwghd0wSX2wELuuVueInBBlEolc0BPSsxDCCL/OKv2haOQvViAtJITaRUh6AnZ2L
hKOqvTdMkvP6RCXSGVSDH45dIsgP0DepL1rB3KIS1oeImuDfyOZb0iI8WHTcAdMm
eHnKH3DvnsAg7pVDSAtvIBFWSdQdA5LbvgHavEBtDktkNzUD126hbHPG/msyn/qe
ipPi5iCRK1B7TpeJrHi9+dHZ6G8yQIN5VauJfJ19p+rzlJsWJuvCiPFZx05sgVFb
e6uBzPnazK09cfwz+t2kRvgrZp2XspZt700NkN7joM6Q6egCgSZdA9YdjnsW6pRC
HAITxN3P7cozkldxvWV/Mkmr4Rh08LQ7LnUey+AmkKtFccHUSbl/rzoA4QvgmYGd
XKAxAYzE+a0ytnows3uqGDalCbEYqlliJvFgJh9hwR2/vTkEtNtczaerqLPC+VcR
PTl1ItzGNZ4GSKT28dosUofTNLB1KqpLdGStJ7dy3S79wHjd+lDOkG56m117/Q/B
LVQ2L/jAXsPRzgIRD/kr5M4WFgYabwtyyWfoUuFLK6HzalSTqzurK6p2W1U7KDoA
sP9HZQfosYsf7JFea9q76tMbeWiGrbqGbP7WjDpt7aLaQL1ZQWD2A41fE3QyfvWY
J1iigyrZ32TWZZdjVdN5MR5vrKsx7hjDH4YVdU19kgTx5AtEOXAQKXQ54VSQB5fz
R59TB9O36+Vgu+Qsf/SiAqDkOiWyc7UG3VavFSuNMHfSjtldVicmlhwSSL4K9RcL
sHdJuc1ZYN+BGmu/V7gQgQ0c1jk0rDBXmQqTUIw8SYHLAlnHxk/jvS2U8dTXCKOK
zo6+SxdDU5bRFwJTBp5H+05LLMZM0YH0RxVMgiflHOhG6m0WYsdtkbf4PusQKzh4

--pragma protect end_data_block
--pragma protect digest_block
J+qOwtMaervyHzHPIgRE+Gdhn9E=
--pragma protect end_digest_block
--pragma protect end_protected
