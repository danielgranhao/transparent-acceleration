-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
BSFlBtFi6mkb6+FATneAH4HjUmgQs2MkNtarKUN0/mrFUx+CdI2dIlc+xDad+wRD
0BFKKvmTMA+feogqK7OA60CEkmuUNAabhs7C6hvc2Fd2WPnXg3BMClt3q45ubP+F
DblkB85weyWdCU75Q5rl/C0fwXy0REpqo5oWwFThyJ8nkxDUHJfw8w==
--pragma protect end_key_block
--pragma protect digest_block
66T/DUA72JC4o2SakNh1CbBfTvM=
--pragma protect end_digest_block
--pragma protect data_block
rBuslZ3xmnBOJMH63qgHuuAGyKh0yonfgw2COMoFtoNmAbhFKLwSJS3XhXId4SZC
TDcjt/ZkzCmMbAMYhE38Adtd3LT4RAqz8ZAOtd5ZnMj3UDZ0p06AS7Z4UOp+y9Qg
hCYCIAOIIG0oSLxaB524118EZ2o3+0pWLC6oxPc1hL34wHokE9bL3BG7SVRsvhNL
qEjlY3pdre/67OM3uthn4Ija6qZTvswzUJysVn/G1Zp/TMD7F7PBCQtClvc6iSOa
khmNOATI7Y7/D/ErGeGF8XWLa/8M8IutmnoKmNkKtfRN4pglC6uUCs/5yg6867Rv
P+MHDCEndFuA0H/2qzMR9ig2giPl9D7ThIPcpYlh6ruLbMdEmIaWHD2IU7jYR6bu
gUYciPrqzBssEDR9f2AW4iPnGIDChcDGffMz8gClR+cL4m+B/kEeAsUkjB/xqvyX
mkkteMPOiLdpIisxHcVu6tv5DnH2qetgDNJCcLTe8oNkndX8VWXQfSl0KmcfZ8dW
JWjKgqAMS5TTS4OrEt7LIVuQa3mXntnALWu3QI8sqgY2KJhSPNNNG5AZHclHFZuV
/V4Fg5yTGDegYPdBm76MDVtj0yrMopMYH+QB06WmjApfe0lBiieF6CxbLUwzhr9u
dYaaF5GUOvyLXXVXziTxgEloYCCddGO0uxevTYSmNvyP3ASBESL+WK4d9qDvRw26
BBWF+wk5hjHD1yMxihqcedfTOpxWgtk4UDNvq2mfZ2nimUhAC7kSzbt9Hdw7rdTd
HW1SNEhr4CwH1JonX+UR9Cza9Q5gM6GMnRhO70n2wyOAzpvKtDL7ASWQNE2kXIl7
aEwVJxY4EMoGiWvZ66doBmOELal8Ck1y+TXRhxeuFbeimr0N7R5GZEpkjvIUz++u
++12T0zNLeDgovTY0pR01leF+c2qsrTEUGKJReHQJJrU8/T0PFHmHLxKAT6GJHQs
SL9cyI7ItCJJmaeug225+aWkk+pZDOqf0Y2ZZbcSLwxOVEorpefqnY7j6E9tV6yF
gE+7DHLDBvx9gM2o0ZhxWlhGGzawL3xzX22U38d8Z4/f1igYiB2MCQ6onsnh3piU
Jpk5Kvnk6dGipEsHH5pyR5YHuiAWklVuPflc7eywhFCZnqjT2aclEv6Z4ev6jfwe
bjgXF5jTd1GLg9e6sGQ/f50zA2zCghkGGftJ/LT0LDDraTe069V35ncVV+XM+WfN
I9Rtmb2SpgqyBYQFqThfVIqCcJ/wBtGER5n0PF3w3qyIgV7/GoFmh4ZkZxI3ANjp
1nkj1uUVBczKa/1gM+QSXl2vUMo1d+kD3DGZIE6WkGpDkfWcE29eiM5Y7iUD9sOs
f0Y5ZTPYmffjDZKVq+excYZPzRMyZEEBC2t8+S55NTUfIk0KN/Jnn+LJsCVcQIjb
3DxbdKDFyE5QejE18VYYLAcotohEP8ZEp3fM2SlBbB+7nJK1eKwPc3dymvuqjADh
Gu8Sbp6h5NCUJ++ZFlv+JFi10mx/9fxCz620ElM7wqRsclYowPzv8IMzjuRG2pk2
S4BX+NxIss3mVSyxywjUcUTsrIjx89rf2ADEDKMzK1SBWbOAxFlIiSIXGhek2P6D
iQIaBrcYpdlo+8Y8On97mEXFPRHwnJ1mpN5t2JhF18pypbzqsDvLiTf78+ma/7BZ
awx+jDk4avALIVMXUe4YDUoG0wS+oV+P6OAtHlNw0jon97poEisaqLnmqvvQiyvj
mQGcz+AI9KN7xhFFRwjTbMX+oJb7+u+f/xI7Bv1DiOFSFCNMV09/6Z0M58qFvuY9
Mf1EwxK/0VVkqY3RpINxG8QMchtCSlBzFazKOzIG5BqlW6+A3HaF3LhKhNLFALLO
nZ1/0c3W+GJIswnKOkIDGq9Js7+aaxvJr3LvTvSUtKlBJtDa6eKeEuoZKMjK0wSA
ViF5+uhfsz3tEPABjUURT7C9TwKGqqgsU1YhOS7T5ks2QZB7NTC6PiMWfQbgtgCy
xkYkzSSDmwOL5tCac3x6VcdqjszryOUtvg/+WBZhSJOEeNqWDvLTrfeZeqA/BNbg
oYIz+Qa1bqXvtIVruB6sEH4aZ77wkdHbbs1kHY6G7hijXlRKNLfNYUP0Eq7GcLoh
579TSnDYmUI9D4qnFlUnWPNF7SZqoAdguNRfvP4cP1hW4xoN+0iVOI7m8+qg+c1P
1UNZBs14k3hXNi4/raep7+7ft8mQajVLeVGf9ODgVKdgaVFESl5J8NPZ11Vx4Sm+
QeXggzbzEsits7432IBQt+a0iJtvZCHCEIHUvFN142wu40iK0sCn5B4fRG62HDCU
Xr+efaA3XQNhuoyEnk8rFlyDx4g3vjhjcWDgjISjuqU8cLnKXHTxt6CjYpHPrHuP
g6m8RpG24Uq8lDjkQsi9l/QvqJlsoV5aMcjm0fipTpRII0mj7r2OJ9xJDZubIydj
F77J0MKbn77rbQkRoRp3nXz2epLxDr0Ksp227/8cfbayQNAXD2+yLfIKaNW91dgm
5Z8Kf3ttfENBmENc4sF3F1ZRPz4ZS3phWm+DQWdADABSHxuJKsdgPMBaddP0vxm+
2rZjY2Llwr2LOu6L/lwGvU4XDv1ImQrqk2xzzcS2kHZlluxE1OzCAU+XRS20x1Yn
YKPgRMbUJCH4nnxHIlPgnE+aVjTR4awxKu02mjz7taD2NzaIEH9DOM4JVykkUhfG
JGysekkos25C31r22uDRzo0tOKiUO0qJ4xUS5PehY48eGS03c5ajgd2MIoPre5Tj
2qmklRndlmhu+tavBUIc3r6sDmdc7QO57nPScEqVkzr5pLlsx0OxKSny4HbGTe6d
mJ0/SnBjF5FjmN/G0+KO8B818GTZKa/W23NO/wuctSNMjlgJBua0Krj064r6F/sS
oL8riuSI/kMKej9oCXeYW8+em7+yV/+e9h4PeZSfRIt3ZVO0n6zoDnqi9LlOqnmA
MvArrMYAuEd5RFV9EyszvqsCthq2OAAxGGgekIDiUopQO4CfPA1wTgCivkr0HdnY
9xq8ICMrA9tkezo0Q5vGfik/vDS9LxyJHFC2fdPV5qTgFq/pyE8W187aAEpgSEf0
n8X5zsKCFIW2SYUyH1gTFCh3fhS4Et7UAkOS/neqYe4sYKjlswdTWw866S6FkiSR
oRdLyl84m/yKAY0WuK+An9Xn8HdVOl75YuMPzahBaHnIbGYpC4w1d/YLqkMI2Hn2
6FEFDssjkmwKjxsefavuPpGbVQxlAEGWMLUhG0GiOp7m7GrlA14hjp16Wxidew+0
hXA9wiIViGF8WzzQhGoQjfpozoxeH+eTBBbdLaUHIBmEy9SqGHCO6OrzF09GiCqU
VvLYtEXPIr4TF1zB8d/gDG+awVU3JMz/jq3/G8h+0hzhvKojPBE93S888cQKW054
ajbGA5XB10zwChS3Ju43J5CNUTs3DOYoum/nbFmJvaFaYa/bYRNkYqa0bKNGAfFi
tnECG4nz5mihJJNIr85d3OFD7TqrCvynIo7OwkH3zKYrFCiI1XjMjhPXCi2WY4kt
dUx+dpHdzv3taxpb+u9X/xvSX5X+mVmJ4E0wxTIHse+MVSXCFn/SqtaEkUy428VP
Gp1Bq14RHbosokWbGTPettZFlNpGr7TBQg4/4+Zgk3ZGvjdX3SignDolzMyU1OB/
qA/09CkmuPFsiimeP8zM5HTNMPt3aYCch+ODs8nLxM6XdEem8l5dFBAELj316GCx
7H9xsMyDAZ7EJjseq/4yAbyTtgCT1o+lgYQAqUjsR633klGLJiAjruritQ/BdH5L
P977NCHkYmKbDEsDfuZOdJfvttRp5sOH+pLRAE2ey9KYYiMVlAk5DNHdCF2ZJl10
GAGPGnze5vTbmhIXL20JVhP+WLK/+9p6t3Gk5puj7+uVKX4/2LQwKBM7CIMntTcE
14y/jthZU4ot4JYiFWRGpBl1nEl6lSLOd/HPSaFs0FlhCvqDhS5CthSor2p1USzw
CklRD2HviEnOeeQDclh/nkSSqsSCItDtChT8uanMXC8Hvip7KqGV0KKG3WGuN1XH
55SFX6aTdTSLMosi9YNz7XxDzw0NjmReiPAai4yVfI099DOCHbS6Z/Q5p+1h/irB
LH5pthm53pLnGJ4bqs3YTJmPaypcaR7ApbJi6SoySL10Vfvd0V7Ii5pM4RDCME51
WV4S+pMy+X45MaLfU4YrYjjK6u6wdsTOIfYR0Mvo9L74Pfl20EuNgqtTKsUCFK24
VQlWkSsVAJ1yUIAZyaoS2sN1DNzinmTDvXPgLt6WXNyGEI57zak49er12sZncDAw
MNh5DRAGoDZrQh8XbIo+AespMvdtR6S9SPmzPo3v1M1JrFdpaXZKj9ehXX9tjjkE
OnMpUnlV3lfJYPryMM1Xl8nFWueuiU+BuaDlSvszGHU/W+DPH2gatphdVYOOj2ww
81cPFHoT66/pRaLExcz2SHfYCRHeRXE1RBokikz/FDFWTylY828noX7Vq6JPvo1y
JZZCDepz1j4HrAPFjN3xMWpVY9AJqJEdnMMcZaGs3PetwXHJ2zb6q2lzvbmmfYgI
nWx0nsGuGGXtDUqvJSACUfokFnYEIBnJd8lVhEqK+3cNlMymlXBzrSHkav0+6MdZ
cXtgznj2pGB2u6Iid1DMw3rcLhZdeSUxjS4E0LtQRFzdSMDSYpMsZo9g0BZYD0Qk
RELKOBAOYlcckXRQzBOQkaIDGPhrv3vuh+RuK4ONZ9XfmGm8mxHVm7gVkRrsj9sN
JJmgxcmOImCMqJD+MTx6pBhhxUW83kcCGAfx5c+jFY55erYWcCB7nx51w/yqin4N
Y3uoa9yN2YyqrwXOoOgyer3K5hDIjVovIzUAlISXc2EzjRe+GLEfF/w6sAhag/sf
wLaOGmKqlgTZA5NrsHAogtrqfh16ysxd+nXCrTgTb4P214uy6cUc0mjMSfz89Dq0
aIrhJNjzjWipW97JR9cXK5j1YNGRqXzsPvyp2Vay/aWqrxrS6GPCyUpWBO+/F2zV
dzW1FI/5peDSMq+CZRfc1HJl45YznqYlKXPgaLF9dG0G+ORA61u+kBkL+dE2r2WC
syoI53m6AROL3l6/rsZSfg3ePyx2NxYc0Zr6TbfNPZ0SvPvPEJsDw12m8PTeg5m9
U1APxZ3bg60zvbKYqeX/K/SBxSFRlbQXE3L8BpDl4vdJblNqx9qOpMNYmOdAjv5Y
139/jEO0aleejOuwrzy5qHIkNrZvNP8fBpASO0WxLs2cWKdhDLWpj4KK26QndERq
8eeAYDFjG1jWgRnNvHqlUT1laR2WHPtZ7p0wAr4Rod6PLR9SwfIlT5mCXKepdQwQ
AR/mq1Zaflue9u27JEVH11+GRbBYadYxX0uQ103bFSuFDdKeaXusUQfC7p6n1TdW
3VhnxaMl0NmpwK6fd19QmBd/TupZ5sP4fHdMs6hSjRgZLlvi+Ic3zjfjKEAyTkbL
dh0xa4kNZG7ncWoZz09N0sblVZZN1OhhQo4RJXxBU7wDj8ALOhHuJ/aTng8AmntP
sEqX3Q0blyOzWrFFFlLRLRN8Imr63FhzqxpxXMkeYSITD18qSN8/ILzbVXsmU9q5
Z7c72v5hvxkpJRShRtb+QtT5csoDP/rBD5zBarUjnoTSpneyGwI17nh2unL2LqxV
kYRQThZo2iJE3v3dLmtpwTgl5NT4KiZWiQFttC9pYJzw0USRe7oELj44GuWc8Ugv
2KTo8i99cChnPLIssAuWOKbg9aOWy/7JKB9WCbHyWDefzXsGeIs781myRjpQtwjR
ctcfFZGkc2QzN50IHHOn7P3KrC0RftkQOBP0ZZtuDqPcTldHvIVvQXJoDdigZCVz
n+FUHllVqoW3cx7Q9IXxNDlouXwxq+kTJQr6DMufuAbQreWi7XtrBDVcnk0AwEXk
rBy5CTt5irjAidHk/c02gKDa/tKmww5RyeOdS/z47dZaHihjbKfM6DbP2LIsvKlj
hKyhfKAEFnKTZPQgGqg8Mk4pIgcsgvYr2fTbDZ0JL+G0f/W4Cpl3BJL9q/q+b64C
xcdylKIU8z2m8yve54TlHZCQsAAaZ72FsdnPGjkFjFOZaGTvLkGVcOC4IqwmZhZ9
Bz75wW3yLxMWHLbRQ7EC8WzOqfn0wPAozCB7M+2GQ0lAIpGYN67EgY6rq26ceMT5
SD/dQe2UuIp39+9k+76vQXyavm14LzyjU3rFXahgRLio6tWsovb1mA4OH5Pxhilg
f+SukR/i3oNXMdukvTOXwFIYPcQhktlYQPYPbzO9WZ/jzE0mJAz3rWpMyeIktK/n
xXbcSPFobiaZFtaBksOnHb54oCsK3SoravuapBlZLkxJPRK7FeCg/7SWA0FPG1ue
MJjSeopKFsIbOvYvJgVqQF8VpE3a/J6Hd4O8Z9k8kD4l0yjSVS1rNbSPiu2JfQ0v
fMAEQXnVNc3SJVZWUW2pRUOI+xGjzrFmZIGTJkNcvrPyQ1WLpoByun0RkSm5Vfmi
/1x/OD2f+SLEff7eiGxHM3zLVRtrIrJ+OPncThsMtvLyFX6VJdH8oU3c7CwGrBNI
c5L3qK99UEg3qUGZgTKakLEBTH7VOBINfjsuuuEYtR6v7mGxYMQWdl7tm7Ygitmx
4oCSF9oOBHtYUUld4u7FxE1s9Tdppn7II4XDoSHeSgpn5e+jz/e0PrECi9+EtchG
ZI5kzzbQfYOO0tHLGDj4Hb5VexdH4FQXcD73nRlgkY1hTmBvkbLop+VwXczXUd4N
u0qQZYU654IRTDEsVMe1VxIx8HjDaqcTkm+2QKt8gGN8B5mwaiXl8V7Jb6Nm9fdk
jOFKYkU1CoHu/GpDgyWtlzYjhNZFT2gR9rpHGrPkY9g928MlrZQ0iZ82cFsOocyL
JQ+LkvJlTfpojNXrTb35ub9f18I/uAx5Jdh+0WZFhQPZ5MkQ/mmmrgYeiXHN+p7I
bcCvWGs5wHB123s4B9ZnumejM1Y6Vukl2ssmKW8c14hCwUjy4j4gk1zBp3Yk4bLd
QldIT9oVNk7XoNEH2TdlgF919opXGMBB/+N1Li+enPxcWdou+v0kRLkaxEQElJhS
5LN0wHERt+pqtyhCsAgAOasHAUUmN97ggc6XYRVd3nVVluUCHJxuxuBufOJLWUmr
lwIUfnIUKwsNC4MSGI4n0GI3+vE+Rn4grldWaC9SImCq1AYcFS0swudzshswHQ6P
CJe0aY+ghq2K+5cW2yChU5IiRPVo3CxQfbVhKXMbBPsRZ3vNK2p3nRTA7QImx7HQ
ACyoiFfRcBbMqsDstRa9972lLYpMldSVVKjztAC5VXuqMljTQB1gAL9AisqajwXK
a2OaNbR+g8D0SpGB/thPXRIvwlLKrhEYQIgMgXYlVsDnwqaoUtBc3qQrWt4aUTVN
9O2JOcigpt1eVWy5H/2SRe20cX678RJCo+yli9MPm/W6F/F5LLGlAL2yEvN6M+v0
J8mcaMApWexEy3z/9uj0sXIJpBVUnkT6PlAVXmIUC7pVC/KpUFoPe4gifEkEMkdk
z1VOvq+4VXk++nQ2kq1YuFVqdmDA+PbGUAKMA3zRylkVeEqcN7S9u+f9uQ0mjGPQ
hslfK06zHwhuPE1zh7RA9daAPlnwWYnDMKopB1E6t4eJ6nMBi/4CQieJJsDEFuld
VhclsqZ76otZGytAZ3Ay2DC5cqIL1vKmzMCf8XRkZVs1FNHC+3jh78tk3diLWAOw
JwQcVVANjv2vo7qb4oQiD9AG34R83tpVqMty6OlLfDVt+cxpThFyiWNJucYgPxzy
1EbFdgrTxa6MLIWKzS4qkkfhooJrf7mW05uB4z2CavB2McnMnZaY2UZYdiHMg2De
LwgS0QV67vGyXf2fs2EPsicd59yFOnirL3MWDZUNgcobwcuqulACjJHg3S5H8ee9
oPmEx1GybJipWchPzLquX+iPm9FahAkKc+mLertEqtLddPMbZleCWTa79Xz/MwrX
AWvrsnlAYgqqZ+teIAS/q/oula14UKfyBqolWlJaWw+lLd1GBNPnZDxwWBUg/9d3
6osA+iFBEkKKdd3u61JdO+UEY8yFqlR90x3GTp1lmpeau1Z4qNTOpdckWqG3DiwR
l2G0BCnpcQvKvUQ3iqmAoA62X6c7zb00MokvZFKoTQ2HpVbPdoU68Qo8Z4HdD66Q
wg+WaxBraiBItP5kHAcwaOXEbkG/9VLWuVkKY7tizUfwYKtRxyznvFlTXpPrlel7
KCqnjOTr+vqLjsubNai9OUt49nvIPQK1aqlh9oS50uHIs//oncCovh7FhKsyh8DD
kv6tvc8QXjbtlJCLEoA0xunIcdHq2AFBsXM1gJutuirAh2lijZ3BlPzIqXMhS4dV
seKU0yt491gH2H5mtPH0s3Bh+pDBA8G3abVlXBAprwHVdCrbZHUQgNS0e5KPErnu
5IIMZJ/AabzMa/J4gy/H7CTHGwKSj+m/1+ZKDpEqE1qzboaS0MKHOt7LZiNjRGU0
X3R9EpR+tuNRv5B4YIn8p5Ub234MUjyy0ogoxNEPCB8ugWXbT4UAsKi/17XnJ7iW
BOEURGxzSPpoOBP+qS5wzg9Z+/7pBCoul1Fcia61IljAYyoT450JC4be6FasZ+4v
F2OdgRILaaVVqN+Wsuno6vqJk5yxynDF24dHh7fK3eVSCeaUrSKo2Ky2lmm+Ql1q
+0TGDgNGLhg8LHRnjKU5nN3SkbAK1AF0bUo4CHKJHuXoKuSGcnrwspy9WTaDOkBH
W9OkDFltHAd5XwiTBzDL9xnGSDM+qPa8LD0V/NMplthL8Pe7ag4npMLOU1MgQd71
Ou9u6syck+v9+F10E0+B+xToI8Kwz8soXnho+tu2GjJor8SpHfagLOYZ1EeaJUJd
eHYml4lfpq1zmp++3xK9yOUJrHbZk2EV/FyvOkreuhOe/Utg38Ef+7brffeVB2Q8
9DSWYj2G6QJOONpcX4mH72HiXPk+L6aYam8jtaAHqxAdG9MMXSgxWLek6QWVnD1G
iTGnVNgdQEqbXaeQGnRXqovEjj5cteRioLhpiaYpYfPSgara+XHoOJ7KKDAaMPFS
6Nv0gZxq9+BpCr3RtxcrLz7tiZFHftcdWSF4KTOD2rH/C3J2aaO9qXoGaASWCJeH
PLpNZ35OFYYIQCK2sSE918fDIBvxPiP5qlnb2D9vXYNA23vcrU2rb36xvVgnFjHG
fWApArHLAlLhMAQaSEkuRQVWEns22s18o3nOllJn48R0G2GvlCuOSBxpQ7MCmq1c
qTvIFGT3/XxvjolPXd+1j2wgJ31hJIDasRsUDpNJxmgWNyUDZeBOTDkKC195YcEb
e7y++nRdn8wArmuBsOh/sP/L8eyPsChtlxqpbOhapoEL+4aQ7h6CBgaNz3v4Ncal
J8O3sPJe4eP/jcADZZDGI6f7FKTcAzkvi+bsqMlrtr5ujkGYLILXPioz1IVao4Q1
V6OqEKywhG8zrRhy0964QGXwuExSSrTqsWUQ/XMbnoKa60E7uMnOq/6S9oe7fQdL
fJuYkgawGcm0rofh+RreGZSWI4WjHXrG77v7Sx3mbgnrAZH4UC3frLmOHT/ztNrZ
khnAmILj73n5gveJ+y6m0ixaksCXSc+tAE+kwZvvczxuBV6qq7YG1WGwmp78ieM5
3eNdjAKYhaYax1ZRE0TltGdG/pUemH4uWDTJmQcS4bRxMUTn6PBhQuYwbSCxFKtk
7ro00JAfxizbj6no8LbcErT+C6m8PJebYx0nnJz9zsMrkQYLiS0cTJsOywptJzv8
qGJdy68PNro3HFaWigtSdzCcfmC5kV/v//gDKE4G6BrggIth6Fp21HHSvPp3IM8Z
SIhfnWOFqo2AHi7T+yyDH1/n33CfaNVztWCq6WHC14EXUZ66HAIvSSa0BteYyRmZ
xCJVgiSE9H/Y0jZgCXv36bI+v2Zm3Wlg6qwN6cvNVwwoFjk6sgy6fXybSs6sUsUt
PqfrfEs/nI7yRMWy3YO9+LY5w5Rp3+/XwuRu24HAL4HrWVjRrCsoMMldDrxTxhGl
DgLTYyFyernJwZe8kYbLCcY6msbGqUTXh73YJOoMrC1IgzVWhL0p/cdrdN4KNL4b
BaYP9LRY9LoP6rCiyiOqfNnepPTomu+1N3rJnUab/MuKZ4PPRucdEXAHa5Pyxd5q
g+nTN9xWLWMaM0FwJA59yjGhs9FgRwlQf7kPt35LQLShB8/pZ9pT8BrBp5huJfJE
NbXN/2UbwkpPgrdMBKE3Dar3buIsjCBta9eIGOHqv66h2QE1b2FUwUf4xAvttk8v
FMIRiBNH65ZGBPKP43v5Ka2C/U54MjbcBzwGcap/0v1sVhGBzKunz1WKk92tOJ1/
2LtU5HHaOU/O7ojJLYe8bKhR19K5jgKQ15CA5z6k9dmON+2whvbKFlN2gWguOFJz
dMXB/jh/MZAzHKM8SBTaKtzer2X0Cuu6AHccaCzJJvNdM/3WIoX97T+hVFdPCTHr
05pT+SaaC/rGZQv0GCdYw7Qnj6opN1gwbWCylv9Ptk6FT0GWa8U/fQ0KYeoY7j7Q
8g4bcVSYyJeW06JAwK8cs2Tg+MSeBBJGI85nrEHfPCHkPGmDc8/blzCnq9W41qjt
zml6mMD3eFExHzdj3yIsEaPC+VpeH7IePtx+yXPcUGR/ysiims2t5rlOwJ/wS3z6
zvg91xqOFD2ZEPFpyGi3jK8veHE7IWkBOY0zHg2YUKowS6V9osUezs1wCVcnhIIk
9jZB+UM1EG480i5bBx+5nvhKqy7FXqObiHiczHaBiI3GP//MhUquU3SNofKdnxiK
FXTIgKVdp2YocN/kk8kYMdJuU3BchZeXSexDeYqo0CPv06bfEC+m2klm2WswiAzR
Xu9uhXQbQILV4t28/SK/hGdLRfq+p8WuLD8PhqlvlNl0Wf1ZFMP64Lvqqnr2S8cK
B9dH4HSrrHeTtsN8IH4GXbFO65j1E3tIHlaHVO/0oeWIA0MGN4fjJX/9/GpWtxte
GLPRDurZRJnNq3tLMVDT1GCrhAaywmUkMa14cD9kQll+OM4qeGT1LCIkNOo/exyp
gSMfCA1PrHWoJTe0hd/4nt2wuGNuujh4QNKxt8Jv0ib3h2F0KH3NVipMR+Okowa0
VYyNOOX5Uztab1MBwS1ZhEZtvn37YvueqM41/Jp5RjA2ozg81LPZrDySvHuvU8n4
TbuCaOfTw3aVh20D7BN6I4pQ8b5hi31C32bITtWBeyFn9zk9NRWVgKZm71G9aUvg
/jOUj0xkYXtTC/C3ulfj7T7exNEV4AClIFTgCjn7+C3MMA6Zz5AhCb1+12TdhUS8
ew4tMkghUbk8t0sa2H57youmcA/58qACdJ+amz6/JkTsU9KSifIhPkGp+hIzWk3W
7TBai1DMuabXP0Pv7WhlXRb4xyTUyBsfzcsjQ7SustKQzkT7PVkYBR0wfjXm4oBJ
y/a6hai+AQk9luf4uKiRcx5Gbh5KaJ55oetThq+JbxN06tjJ32dH6iPlVVKh4+hu
bvGjqOSxkmJab1tR6QW99q/BSbLfCutc+mkALNX2Q+MsfyOzCvVDRkOYooIg8Cfr
Z2d0EAWszqcgmJAidnGolgyMYt9iWSYIWj8fM+A7xct+v3NNwNpu7ZLGxJmQx6Z7
1qxJGkN8fK9hI7IRwgvnNeIxjaZKXZzQljVv6n06ZPtgRzXNOtJ4Bo8bW7gtMtJh
2y6pzhvny6Tgx5RCwE895PpOJZzQ5AlgERkySxY2EdEZ6i4lUBcGRgT4hKzdw7Ld
NARHnrma4UGQo3/ByR6k6TCKcUgnzi655YqCUJ/VEosmEOJz1jBqyqe5U+QKS9mO
QOatv25b3dm5pUqCX+5p1P3nuooDYRhe4E5qOcc2FSe8QQ1K78653kPDglYY9kv3
dFfBFfefN479jqWhh/GkyT/CihOf3XSyiacjwIaaX4VoPIw2/wMbfxXJr/SMdJ/U
+KBA0I8DJcVUgi+lImT/BE3LJYj7lPJFZyUW1kpip6DZl/Mx9vviazJApt+TcQbn
9q4mSydZO8YKmNyWnyQFr1A+GZf9prb9Q3Wbw7Q394w3JYbYuO3rQv9SL2sNOOt1
GggESzoBlEcxwvxT0xaGucUqSuWYU15tDPjMylEFVBSj7kcxkMIF4ye8F6xvJedi
iziX9W+LfPPD+68J9Jnzew==
--pragma protect end_data_block
--pragma protect digest_block
GvfYrltRWcPzm06DEgcFIf2xMQ4=
--pragma protect end_digest_block
--pragma protect end_protected
