-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
gyx0kYv9oj8mEgrBBuw8JwMUD5KTxXCYWbePQeVdHbnaHCylRTjguQ8M4YAu0RSh90a0Y/vrFz1u
u4VbR4jp2i7Wvv1MQB/YoQLfwlsbfYK9aZtInHyWj7DLRPMHqzmAlrVpxrtKlOc1QBdpbezUHumd
mdFbfYXbMkEPwL6gIsu0IbqOJrLoIfUNuz7M5ZwK5PPa81IqX9Wl391/kmDAGXdYS9XbaQziJWrq
BdnYG+1jIqOyfD8HAi15uzEdWNdrqho6W/95pYbLQ/xl9RPBfQLcRfL/2uZJcXgSckHnmb11Olgb
+wJLz/fF8gDdOSPsaqEpLWbIrX7qxDk/6kf3Iw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12624)
`protect data_block
yy/5mAJ9Nj/7k0/pG2RnUr/7WS4oJQoE3kUWkYzJ6NW8mz6pRYsSW62Q+wOag33DOZJfRKCdXYlz
upE8HHeWHgqudL/H9nYhJItH/IkvP7T0YfA52U1576Ve/ecp9OUv8Jfg/4AlgdhVC3a6ruvlbP4+
cIP8b755XsBcAY1ZBz8Url5UQ8hHuow2HXlGKujmYOaf/1hDrm0QKVfkicb67cNVl8qe6D0M4AGZ
/VBoKkxblrx39Jbaj4cIFDw9eMge0EOJyCJM3scFNmPwRYASKWjt/QLISYhkcTPHpmy7theK6Jvw
tjzBE8Ru6eVV1hxMigoVJCvSsdrMKmrlGv+78t2xkFhQMjt0pp2ldEWBPoMOjxnFlf7MbdGU6avK
f/R5KkrcbeWKDASjRn0JoPpPUmSEg9MNxIzP7+hGbTM0Uo+CmHJhCauR8Pes+hirBYyCa0NRPZ+/
GLAN500Xc1fTfxW3+6SK5KEZy94SHEdErTldR56jwUkmKW1DqhtyTQ/kHLGDGy3Ey7HtH2nqXUz5
EIzAJOkZB7yLzVMdbQ1VH/p147IpjISlwUOUB5IJwAev/sq7WW9AzeL8AqjAEENEs8JSa8gkIZmX
R8+iE+tnqrEnrDhSGgiC9t3q6oAx6ad4P9E5tYC8Ls8jEQRXkY9vzAQXOaS6P8zcaR4MZOYI0hfK
DwLbYxIU6po1dJIZ9zKVkpeOs++fEYJvDWQDyX8JiGlD/36EBZzhw7j/nw1Yp7N7e1jBlPsUUxBD
xiqpQazJ8dihYdZRvSqrACyCt3ksl/lybPYtMhwFJZueyun0YFQeRtshpO9Alni25h3obzo+Bz7f
6gZhJ5c5xQsZejdFLJYlbJO31D2MSsfZPVHhjETra6ZNv9q/l7bFG7TJeWB5VIViYPr3mwCaAXMj
FUpK7g7xFz8vSo3ZCd0OMF7BSxB/wLYiy4qizwiWEa4olzOv3KepFi/cVIQBwpCgxM3qIlLr8BJg
0A11uP+RRePbRtzYTVtQsGfPZxr1VB/EjSv37oZ4A+XbMvWhX+4y5S4VEktgd7pPBiXk606vBgVr
PbsE31GurWt2o7sQ+R3Gzr+rLYO3keAcIpfdrkO5OR3jnF/lLD5RVH/eA/nYQWbnZa220wzFJ/B5
tJgzFCvSqjNrXhqfjnSPoFPQlwvka/U3dol8ESEIn1xqe3rA1xx5AzJOoR2CYdVHEY1e1HFQ+/B2
nZNeLz3v40YGU+tOmzV3O2iQfq86u9YvEWVlazAtjSi3I1rzFk/HS2vLjFVzSge+o+8jfKufVE1O
iZL0zQ0jsAtyDDXi5mQjtCf0/ACjgkBwoPFzYtWfrm86VWqv3NyB56+QcTwAOmvl1RTsgk/YW8ZZ
06Km/CvfSmB5BTkhGmxWpSMc3LMLYbPXqHACpsCGFifhIEALuA/EwTEaxxJQ2iqKolei3tN8yd5N
0bnoRTl2lGbJ7F0j3sv28mEWd4r7Aw7DL6vPVFrHOWbw2vrTtRH7GylX/zXQqhGLwZk7vq6IYQ2b
phfmpg4VUVhF7GEyOHLPRMUZGByfIBBRbkByunUpvUjb7gOoGHlBNwfEXhpjSGQ17hA5zkUJyo4V
1hDcYvsvBnmdG7TFDBu3g0cUdXUivlQvKK1I1bjpPrthMtZ6TuwT3cDqTAK+yu2N1ocq/jBlQHye
09WQC3ifodMQ5dU3mKzQ/Su+oe4KIiNo63Xa4W4sIO6CDKmj7tp9OcZV6Jx65RfA4XgZMGZgPEjE
1vUF5pg4sMd8nr4yG5vlKFarBmpj1fFnCUmezwobNIHyDBL0IVf1t8GZafQlBzaVnmDtmg2zRAnI
uH4WP7T9xzzVnAZ6HhtS7/3aDiTabbElvaa1VOat4B1NG5HXtq8OhG/FExxzVi0xxx56oWANMgJU
yZl8JZDhwfqeMhBD0YnN1mrtxZylyiNXYBy6L1omFzgmWZe20kWDkeubQk/UT8bUIWKQk2qVLgCH
1g5JyHvKT5j81cHl3ExM60GdclZp3fqB90RsZZKVUPazs2+APbyEvsvmdX+I4jkxIR6/wEHHrwAd
pX/Bwpfox68vNTAo7ea0quHlZSDypyRKnpTNUHm2A5L4Exqxrjsxh67y8O/b70uyCP+PsAyNVCGw
u1XXKkW/QXHbRpkjMq8O7pCY8rVO2ETQPcKE1zO8V9668ydV+ZQZr6X1VQWBWyN43HNXESWyyrN8
/dMKYQJN4iOlYIDGYwdaBiSUHm6V7qJtGljLr0m2Xyh659rzxxf1D7L0aPRtxXpto+wY3l6j49EV
+Bxv5OzYkWrHbVzAduJVt94d1bI+sREnYRoKBnSbrfC7nsOrD+Tk1t7ZiCp0NuBIBkM2/3g6ISf0
hSeip4gPkscQocwHTq2hBjvP74eBHZMmSdxzcm1rDDAshX95jV6DqKDvyYkMbX5SlFiBfChPnOlh
54olMZGA4bwuezt1eBIhm9Itfdgady01vaVFm6mkiLxsUdsnIYNpsUdI3fjR1M9veTOC0na4aEjz
vWIy+ecDxnUM6Uzc/VOFbMgWdxbv6rrPGkFg5+qkCDVB0KgnlKEUC0AdHEokAF1+viGrA93e0x2+
UpKt3DpBrcfn9YrTLl3Y+xeJLPkMmJPoBIIXmZdC/Dae/JnUumyIoGx1n816aP0TMkBPuqLdp5Ew
HMWilK4ycXQQnR/ZDjuaAShx+B4vahUXPfyWRnZ4faeM9nmZoMWmieqgk3UR0ojY6wY26L5ENu1U
avOS4KOg4sPEwWbaNOB1xsxvigWCGSspYvlG41sjRdHfOZj5vCIKIapHXdQP6RMEOsjcm4KmcYon
kfTuMO8lEqwHiPpHcrq7Uzh5C6ogMav+SCw/XEDS+tuJUmmIwPXVcH1wqjPWDKXWSOnFeY1AmD63
uVn4yx+RbXaW1lL26E68pvQLTvodiNYcEFk7Hr5DjqkJw/kubau3mPSvfUmq2gbqXWwclzSdx9Vw
tVeEJpHm2Bf17oMO+oNym5veoidvWQsNcj4T2Ca4VjLE7Ihps2mHn6JFjLaneUSOTuBqkXX0akrH
2u91Kdn/4uhoH9rUysxq/kZshp5f7FwNQI3K6jBBRrcfn3NQIEew0mcIQ65DdzQzNw0rBoI/Jfqx
PKx4p71PIYCcbQo6ggCvIkVoTXe11E/mRxcDl2Kb1+xm2+PIiHwpTod9cCTE1umyEz4Q/E/CqPcQ
6CnBLtRpCQ9iIT9k6qZKtHu7DuGokdfOgzT3G8g+e8MKCICTlfG8XCLyvrZdUHzu9C/3xoT64bbF
3STAYGc2VqpIP8c6Iqi3ZwCyAJHDTp+BmIVW95lYrAGAaNzlQBKW9/5YMXaPiHnh4j3Cmv/u5dg/
aCvS7c20iBml9cE8sBMYsLNXu8frl72KyuDTo2cWJQ8k0xbeUId1p4MBmMwxQQdE/IXspXyT3RGZ
+YhPGaFakBMPZtZ+e2VmXr6xEmjsRuBnuXwawLCLwFOOcqDPKntpyqP82hYkk4s5irbDhatwhQWF
ILn0ttxLeHzpAB3V1h1qL2f3o5fpnB+jHp3DH+TV+T5CP0YcN4T9dqj3BF0chWXJUQaTbMSmjCmZ
vDXg2p3/zsl0XZzGXAzhPZsVpNbg7S2DAvfLEt4SMiQLDQDBJ5otbpRQCXNfQt5jJDhR+MiQ0TuF
gnDx9m2JqijMZKRiF2cnQ+KYpIDFvPr7milUXMSSEbyeYjw7jpl3pHPdtY8iQONcJV11beWUIjeC
TJY0cw71RPib/9hRGNgfZROU+x55HNwDxHwVYiVdDoW0xxZyjQ4AlIGq74D6Eg7S3EBWYPpUP/Nz
2/UzyvOgAqz5B32SpXC4mlrrqJ4h1rqNcCLwzr9Kb3fLLDuqVnxVLQgqkMR6hpPuzXPm36xIU/eI
w0ga3CU9jp+AEHAjz+torpeGgGrQWxHn4I2xXSB7h5jBHukOoUEWN8n/QwJXL2/0XSEEc94YM2tB
PZp2r3Tz0tLertgel1X9NbVlb+LPIJKmPtZsyAZdwZPS8049OuMSXuqfImG73tB0jwFeMc8LqBmw
cd8i77yQVgzGyC1wMuw4uwyDYcu/mESNRdCE3kM0eKN2aDNTqYc9OUUcVawpj0R8il/oJgRYe6Z/
oa0woDwLSeYVmHK6vWb4loII0yXAZBiXOoGEIeNZB4ESlNCCGoqAedVhllMLsLlyqXrqa3ibrfhj
VDbXzg1EcOFP7l1KcpBAVCVH15Bpu8g2FPQyDLe6M8EHZKJfNtszN8Q/qlmFnZdwCRATljnt8Soz
c3U8bUkk6Qe8U5Gu3DY9ZioJhM3CIE776XYwHu2SQynghDDDcZeZ+besctn8ktsWLnj51emp9U3h
rFPBe+OpcRU5R1qkoYCzMDQwNA2wERw5kN/r2G7faN1gGmhIKzgGUWk/+uTM3K4U22HqCmKmoViv
iI23SERwHxY6qAZ5ntwJGro2SCdnfx6Di7eSbm4RbBM21soNSQ21nnI6tK2rImLJOHZjS+6E+lOU
rrBz0PefbjCM/xEiBztI0oD7TWOAlzFErG7LZSLF4So9zqgZTwQ83V77DqjIPuFoskiK0TQFlalg
S+auJPKduC1Hr5wmUkQaYBB3VLwmT2CzFkwkgKO72R1CsJY0ydXJl7M2tO8zhsqwwIuY+ZyTkfYD
9mUGhR1q7DkzEtgLASb6hiG4IdtZO+aVE0ydVtvXH5GuTPieE9fRFJ/Q5T17VNLahHpI5qp/0xdm
mxnNVHVfqGxeCEWL08u5NDiJKTqHGco3E7HWXCmtxYz1DhBQnoqQ3dZgSbnTlOxvY10fpfpNlj6r
6JjreyVH1BMTZcA+GIckVwD7dFwYErdKdy15oGUZpkNvypl03Cmy9rwJKUhuLA/t44MR9Jy6u+Wk
G4EX0sB7acQ/D/ZPeZn3dj2T2jCtTYmHQblRj+mK9HPKY/EVp4pNpz3c7SNlAH03UoA8zOQrZYAV
LflDeDPatozWEgLPV/seGH7vVRGIPiKM/xuEAOZTKPNWVp6snOylXCbwQpLRC3Wa5orMI8vZim6F
ZChSISQKLlZ8N16gxafY1wlW0oU5OhYoHTt68ixZ5gjKBbxd/6JAQpkSINcIaCSnMZR5yANhZICe
lDBrhq1G89gMU1uNwDCNXncTmFQljprJO5ADjE8+fMFIQSbLygacTuAAXnJB0AxxXF+Ac/59+SkP
U2aFCvPuNftvYBekzOLqbEE83//N8M5iSLPAtDrhLRCyA4Esh9FWx3+NmdLvyoUlT/xFuvzwHtcm
4QPXjE8qsK/LMGJQVIt35RQhY/r9m/U5GkJ42kJzG6p1PSYoj/IEABcdoRRG0rJJvcz4l63EmBHm
95pQzNUasocz1oYqz1pn+9c/0mSZtok2tyqD3d4yxMeCzpSdiHpjcRojcRjkAGOvuiMWblHT2ujn
DP+bt0V+ZMCltXRcSVm217qD2Gtw7BQhXw2A7yBj5X3924sCp8kQHF6OcTaW7I+z3vrAisegKsCt
ESrBeIHxCkpuJaPWHGFOfjywBMrGsov5YbKTA4A0I7Tg1uUCky5L89E8cV9qsp26rNyxGUEiM29A
R+kAj3a+OPlZjEmT6jDpW03VOJyUjEo31K6wVDkz0WIBoimEKvTJtWod0awnGqm7Ery6Mwsq471d
SQcCORdjdcgmiGh80SmIN5cPvj+KPhEeMKFgcl/WyRTvog+W+c0Z/FMq2vRpc/7I0BhHEiONb99s
Vl7SvmydjwRxWqrMY01uAwivHn/YZASY6/PB98wUcN93DIEUIaTSHn11yy1M1NLmWs1syfYF/V7v
EyYpuF5cNPM36DEC3QO8Yewyz+ASTWhIqa1ZT1CfG/85msQwt3i5zMjaIGQIExCApTLXnknPfDbg
toACpTll6YuX1p0J3o5/NFSNsJ35jQ1wY+a/JJjPkxa2GxYRpDGm8UCG305tN6HZkI8tbQWjTuwd
WRCehixfWEj6K3Vip4LfUbWgt7YSepm2RDmONF6gSmZQ0Ivanz5dNrqxNLX/BP4RFfR20G/8v1jV
WQvhwE+9ct+TNJsGeBSc2bxFxj2bq0c1pUSthkNLGAtLkFR6n4m5EJzwo1Crb+sHamQUWkOkLqZt
pdPi+U584AphJFIoLwpSA/iBBD5LA09SR/rR0JUdnkbIdLeN9H/RR7kt/GJe6/vhDPTYTKEwlYIR
+/Zl/gUotNTWbLs5HCpOlc/jvlfaume4aoLlyGHZ3kW+mMCbI+O6xfuPWDMosrFnnaerP5tHqM3F
NkpDINgk8iFZimi4x4sjAKSZtjZ0BcQt3+AoWjvXhVupNNgTKWBpOz9A3hlmghETlO1/B+HsBqvb
hFMLPPyuantURzN9QUJfw16jM3UaGXvkpmb76g3W8j9v/1DQeLB5HM4+vRCQs733JKSQOjTfewy3
yY4Sz2ZAgcQKF2V8Uqa4dWSSSl/CsHgqfuNaUYLgOfHhzrKCf7drip1W6/7ANhhhV0S2viNvB6hb
u8NECa0oShcnA2VV1wxuibKdxSWhu551hU788nAoqrGflHzqZAvgWGMndTgBWFZBz5wkynRMNc9K
YloPcDkuAKduEc9nOKVxVboJ2tz3XFveERyWZ6s5ek9QpOUUiuA2Ykj6bvGBPzH9Md/JfMMLZEeJ
WqYEZu2sb3BQHuvjJ8bLq3d0vSOFCpnpQdH8hlzSaJr5r/BAvsn19p9NX/czuewsfey1dArzZYUA
fGrJAo7MPiF5Y+v4B1fc1CSJ+H7HjDUbP8CE1/meGuhO5xy1dG3S/xIcIMDErSlFN7awOdBw6rtT
DDPKk3pIcnu7ZNssNXZCWinQwI0yvEdXRV36XruELwIufm7E0NmJ3V6E9Qx0vZvUeyG+74ixx9Iy
kAUy3QWFv2EhbqUPpJCYloQxk+JnXM7AjpCl9sSgVJEpN3uYyhCKbH7Od1nh5xHBc1JvnqUxKr1h
GEddqeTUsf5XRUTHeCwR07NY/uTBJ8w/OXBA8//Zv2+ouwlTKqOh17e9vQWyZ+ySnyP0i4KBUd9H
qA8seGXgzdwEcOjnVYKiLAmu9uDWJpchX2sDlmLEgF7QdZSYhZ/lH55PHrLil1EOB/xpyVVoeb0q
CH9xxBxtSA2lxDgvcZ/DVhIRe8lNWte9TdFndcMjdAB0y1QYeAbUvi3u5kHDpF20mQ+8Xls3F9qT
e5R2qhITT8DNYLkUpaF+f47uxWAhhjQh9x2QwMts1PbU1tuLhrkowHKQxEAHory03NP4icRZo55S
ox/dG8Y+TSwMaKawO6xTT46adCBw7P0A7bZ2unViBTi6oBk/tzGSOLBI2ZP+Oh42WWkzYDCh27Bp
L7YIbE+fyPaSh+U+Khj1WJqYUR+z+emBUsif/XwwIb5aHMENOilehg/bIKoc8HXDjokL30YfP6nW
4wZRv9sHR68l3BP+qArDncV+hai14jzyrupdJxXkkYDAT8r01u3M0Ib1angcPRVZ7RRXnqE227hg
Zpoz3MC8mz9yzfwJK+DV1jyTaro5hmHkaoGuAtP0CWNanZ5bsgQOtEO+vXucDOC0UmZrzQZsXksV
G0w6CE0ydPMEYfRhncFFz6B5ZPZIlGQE9vmG7/wAPgsNiaAjYWJJvt1ERiX59oCUfomOFQQJ6QUA
pMsboyqvHIMoa6nuCDmIiRXybHLUWhRF5hWBkF41y95YjwCVK4P+YJLJxaofp3wjHVtl+X8EjbNM
jWwshL2VjR2hDAckEQAH5WrSV5IVVcypNJNaOs7XLgclGBEL5vCfK3VnZaMToWXPooENU8B9nyuO
PwL3smju61uzr3zFj3t9XjGFhIRVZeKuYelmYWgOXmm+O918ihKE4T4n34hnTYlr4D1tfeRnUUYJ
bDhpBUQP46DWbUiW7EzqjZCy0QVfEBG2OlA5kIOvKiD2t5ANBtuHl6xed7MgUdlUhT7hi5p5yuq/
1VYWSGyjwygSXEkrm6nEFHMbm7Xq29UG6ofwFVpHxWGU8WV1ImRCmqaJxYbBe7HzSH8/V2tgojdS
Or5xeLpDmH1htnFtaaDjEQcsgZSBebCDJV7I100uY495LmtlS9Yhx0F7y373crzpDANOJVnyoVBZ
F9D1ngN1eflFoTpgf4a/0dDcFwBssLleCTdKbysZt1Trx9hSHFzktIUAA8MUB8RGHO5ar+S7WX9R
9HznwRJrfoxvWMaNmWi0MtiHd7P3VpWsOuioXfBCiZGoEHnj9Obgh9k2kYCpvSdld2RtSA/NiUu4
A44vKWvkjrsZpAml0JfMXnj1VyO0pgQ5Xk3FBQV+8X7GVMPwNpLjiZ7VpyaL1eW2CErnmNwWCUNB
8hSxHxnm82A+w9UOa0xYUfwLv9YYwpP5M6damWfXey1FqLC43zZSe6RAZzqrSOUaSwh8L1NrCoCS
ZM3IDBHQuctNrFGKRIQUbl9rnhHHIa/rcgj8SwDnPsfm7tNTmUxk9UewWZ3660H1zV7UsjGVFKso
nXpML9hK9ODBZ99gbVvZQOu0K9GalNwoTnvp4SzhorApZkXyYM66vzJ7yqw7fQLV+QrJpiBHu7Ov
2DcoQtiweHvzBzE5Btz/uKij0PhsUljK+ENOgNvz55TJVYi4tEY8u8rD0xI5Lshvd8VaOfK04RSc
5O9/ll1Mc3/IZ9R6xYjGffTfm7j+M3U/TTkt2STenBe7hqNAMwcIDcwyaGqikGOt4/0tz0So0Q/L
cZjKUSB/hcQrRGBMtkb5ZsCdtxX7TFf+vCk7apFXDxZmyDkMxLnlZjDW31PL8N38ecBVAnrey8Je
iEPiZC4onKO5DFDu8xVzXGG384nMqSXz2ioQUQbzA827d0ls9xTn+pvdSd82jCoxkXQwrwhdjv4w
ajFh879Gsg7wqzGXRF22RS2cwfOZoE4uthIFksW7vZ1uhZv10Wq6HK15bl0eNtd43CIGyMQ+e/s1
mM8HUPcxvB2akSIkIUcDv/7G+qCGq/A2RfX5w8baRNSW3Nhi9b7ybrKr4ns0H707touvHnxuapwl
2/QaQ2joH4kJrxM8RReyY3gkwjhHVHWQ2mp7+HJ+pzodxRfflgg/zdBx7R4ADeB6CAXAkYSQwM4R
75x9MRSLmcoKqAShZ1O48Q77rjtS+z++YNyOM8F8CNdqDDDVayCXTzYs7ZOMW94leJDXTN4036wm
+UqUdAQwgytDfHG+/hwRWCIlr5x2dxZuqcVcvgwJsIUlfSrKlhnZnyP9QNSO3lWRjK7GHVHrsYV6
ndKlPg7ErCEWmRQcRdCYlJbU+iBi3V6jk3Z6s8k1tS6WVdpZImCioGNm0BNTYPvqKRmE6gU0QtM/
c8a76Mv2gT+jus4OF/iEaKJ2HDrFhWu/eAsW9YK1ozXWdtaSZPi8ltL+XhZYGkQs2CEGh+ZaCoh7
UvucVbBjTCs/YNtg286B9ENO4Dfj6ctEQMRHr4RXijAfe/61IsxY0JDPttxvya8kz2GTjLlVn8a2
LtlUtGrpqfz6nhLjOM3msSOkpV7+g+ODv4qNzMaulJF4a9gvxP6iyjCBi9pB8F1u/1sOGZbusmX7
SfYDqVcYjl21zSAmwd1IzEiC3s343AZnlWhLWfXbltB7R+SBQ673XJAQDSIuQbO5R59W1Tcqy8xT
8f8CBX3vsBvKqQrGgqvN4E2VBnUWBGVv+1kSBINu40UQwiGnW1KgV6I2CjjIHM6V7oMklEv9N2o4
ZumvNZzTkhcDWY36WN7/iGfH3wVXJJdzDsUFusdebVoruvuPLse62m1O9FwHDA+cGIcNh1UIMSvb
3aD7qCjQ7WMjJACKAKlJQdde1mZgKQ6r7lvA4CBJNfMhY48uU1j38s0TkGkzC9x8Dbuzxugz825z
6bkJrtc7/hi8oVFiQr5UUk8xJ8e88NfoLbZX9cobqeHqu7vJXypyzMrHQvlD0J6jcjHfGsW4hFW+
vox6jrWj1Mn/pkzNzXB/Gs4tmiobvCXQj6W1PV0BD4oOn/YhpoChIVYokC0zyTrY3qHZbPyvhQv2
HYMdb04bod/3j/vxclGBqHqlfhi5XUpvJCBvwdySllnKI2LnelRTOuP+F64vpN806BrYtM0xpEUT
BBNWIEb5fuYHwcIZqma8znL9MAANxx17nRbUwtyoemSXNQ9+FUcZ12jgovtMWPXKNRnmn67klXx1
6vGCeDjZpjmRcgmtVA4tV0Z6MeBY0rl34YV4rk7y+rtZnRnzzLLiF7PH72BUpQYkzEQXhjaCs+W+
X3c5RVWuDXCDB7k8HTEIggBh5o79Gxu8ysBXyJlX5g1k/0n+OJTvDQlwaedWK7jL8065lVWPymIW
P8DTRR78TtpN3qsIrk+1JvESRzCka4CEkIPa9GDC2Ti63i/8vv/p6xs8/GDfCSUp618pYw/og5s4
MwGsm9yz+bylZpJFOK6B4jraHV1PARJPSS+mljSRK21QzUyVX8igDJrvZiAgG+kYY5lfVllM2BYD
+ndWh6g1N3P/2BoLiDnzkH964spEr59ZpAuqUZ0XMtHQ1c1ORMnCh0aAImh0vQvUIvZ8LvZKabW6
jq4jg62S9jI6J6L2hTcOUD7KYQIHD3r6Lp7qsqYbVZeQ2erV//USSCz1Yd1imv7uLYpAI3+HmRj3
5aZ9cTf0qD2lMHUwfa8GpcbdqrultUus8B1AtsmajcRwD9K0sWIOuuLHqk1rDb2qZkMQsRZA0/L/
0IaP9oXKaCnBX4g4Emh/fFiXHizNUv2jrzb2vVpxI9Qt/YD+yb8TpKQMpcNg4xKjG7HRAH8E3C8m
00bM4/a3ssvh+PMES9KjtfrTYCzW1fJ2Rlf2QuQTY1pEwsuf6LdRdRasBjdSNKkbGcl/X1hGZ6Ga
q1erLgDJciCFJ7o2yHJPnbPz4uuzM/bxjZawW/aE5fUGJHkGem4Ndl6JsdDdttBXzn7X62VB8lVC
hu4nh3nlJezyA0AQEhwq5WdEaxQrTfkDslBPfLsevXo0iKeks9Q/zr/mqfRrzoBAjTi0G27Fp/Ie
j3OYQWndGfN0F8Q63/YMw+8XTQhCHB9/c+mMURIn3USpe05e9nigytlgJkpmCmqIzWP2XWnHO59p
6aAfLM7XuVQblITE/CvKoXL/m/GtQpR3hMOYMB7SLonZzr4tgsm49XpDGLWxY0ZkdRwWHvlGoqFt
jqdYVinaS8sKb+wAJCVDabbXpptRJoYJvnsPcXPbxFvZxRTEo5BWUnfTXBJWsB2/UE81XiLjXMjM
fLTBJOfKa2+wbYnThxKNY2oD1RtCXOynpEB7fkvFvDxgZNxPcy7KNqIt18maoNhAzw3KhuwT62oM
jeSksAp2M6c5z8pEbjcWU7F+RQiMVDf2BexqvPRfu7SY2a261qEmRyXgDN8JsvzjnL52a41s2KRg
i5dW5ZYDD76cYqY9E22GJ8Yp6B+dpDp5vv5Xefhy28tpXvCBEsXPOdXS35MOIF/C7ijelok8i5ar
xRDnYW80nUfEnRYsZ+PpvVblKPV1D5f0SpEcX0OocsyMuBAH5IyelKWGRiTLQbnOxZ9wtkAUnBPY
BQ5oDj1IUJiB+OMjFHyvb8IlJwBEqDYKC41TBX3KjD2eOapJw1B87ZTM9i43XxXtFPJd/lRE5YKN
foFonAMkpLkjh+IKRuljeWsh9lYPeTA/lzHFPIjqMYOXs7C0nmPj11/huTLLEFx+mL7POng8odf7
nY81WR2h7UeM+g+PaRwOvIF5NlYVWNZCWkYlrVpdgrK0Nx+joUyL8N5Pq9E4OnKjotTUDAXFZZEF
oX6NrF7NEFTe5WeyxIp/87AeubsrbIJpxGpKA1fT9/zlv5kujepi1fPT38qY6MsyuGFm2LZJZ+fY
J5tL66/cwpsKN7IaSuY563dI5VObesDnHMhXSdr15uDIg79XihYH7UED9BsVC7w2Vh6ium4dncMu
SMo6zmJIrUqbdYoa3NThENbZKkUjndEBlkiFUbBzQAzwGPBT3bWS15D0as6UmJc39sO5r42HtSXL
eUaea9KCwvGqK/Gcj38JdeyFAUzCgSdl57ADECLPWqX22s89NTGqOTq7Spwr98U/QGJGKLJ8XY7S
OREFXGTLdipA2pz4tFZaBsXkm8is4cQL+rL77maSpcyx7tXKY1JKC8P6CofHon7+JcS401JlhiMQ
28o02BajgjmDxGRFm1DoDsTp+7IpTwLb7Nm49AjGDjOgcZxRdXAGFyakfPfrIeoAMEJNGi0nMNGE
U5Udw6GOINLCYFItw3A9bRdK2lz1HHpEnhZ0vKOVbaWA1QjrxIU1EugONpt216lb5e4BfVnSvD50
G+yHLd5QQwJPMCZBKUzlcyH0Rao0hZZKgjQHp395kjQtaAopvFakGZexgSlI30UkLZVQYUQxMTec
Q8xa2GyvcHxmgGb8gJprNoPgt+ifFDB3qfuzv0UMz3P2KYNjflbRqXr8LgAQuhPGhxB0Zf/mBsOi
aC/7VHNgPM4qZnZKkIrFcVEpDB5hiFYjPE+3hFkutLbNp7B0lE/cPkxz80C64Qc+BgjhPpLllxQo
m5u8d+UH1zjiqV6J0m2uVHiLODMJ7Euujj1ZYnhnNlgRvxKNgOXJtcG/CfgpjfjfGSnO+0Qk7ldP
pVNg4SZ8fr+biUfFbx9URipkS/jpaTyL+B5j471nghBhTHEF6QMzAWAcW21GBFn8CI2jY5j+D3tC
Tx7o2gFi8Md2lFhxKqTklVrkVc/ZhRA/5w3Yc/ewKi360lVf5jy2N0rVGWbTjOjWMJdqyFtHXGiK
TTaBJ6Yxib7rKJ9oAPIX7ST+AOnuMoD2/FD85MQLEuVuWBCRsp0IW9LUyoNRfXkQAVWSKhMINduf
C+OBe03xyoLgy4Rt6fU0jLtylL6GsAsNmHvKs3zQulPnmrSac6NsVrmjgDVyuvZc5AQizLVFfQVF
RagwbQ3yVJFjm+Ib6eXjjLHrpAenGuddcBv/X4J+vxNtn/HfS8Bt225mmeqKUPRnmQ1Oo9ncrVYb
msgtRMhVsZIZ3qAOkpqvDXsHEwmbGGwkUA0G6A0SR05YjFScorswGPV2SenwD+K407Bct5yK0WtB
aFdUdmMVaWnp0W+cyPqy7ZrXSI2WqcmOxsXW2kchfOWIZ4tEPkMxe1NM9o6XMOaMlF93bXfRxTg7
9yE6lHx7lyowv8zNt5NTKW1F2+SBhz0iFKLZeIl6QDb4BLmWO4JL+D6qvUP4fm777TcD3OIU0tx4
ymRWFh5sRt/xDLcgFPwI2h7VklSiYW+rdz6bEwVbcl0ZacADCDZ1xug004QJLuLpHV4MIwm1c+h0
vVbLssZiwI6AuMnlmO3+yP/UWyPcuUMTTwVyPtAGq2AJJDjHWsXRylssuCXitgIhwY2bzR9kwya4
FABcAiXvXR37A7SbU1Ztns+PX4oT4yBbcFcO9w6dvVgMQP/FVfvCSpSNaiQcSpRRnhEe7JT7kVYW
6oXNw5E4IntWQuZK5bh8rFLheu5BZ3IueAXwDZ9eLs6T5ZKDZSumAxIaQT371ZWQtkjy++bf3u4A
szy1K9OXxY9YmY7WxYyDFl4SOIjJwe12Axjv2TyIZY+RH1wdmS60LGV+rxIR+9uY5NgVnvNAaZi6
EnPj5cftyUfhmtOJ3W1hwaIsr995YydmZPONDE47xplmAWV4RIcehwEb7gUQG0ZZCTuXinXuI9Ut
7PuRBDtQ90dDHShwHguGM+YfzzQOXCgXrebca6avHA5oxqLX5YdMCcn3Ig5rSlvMazsc8eU/n4tg
uhZGkOHxAWi/lYL7Ss9/YF7GNkmkVK7vDQsRLFm2QSakTrcTGYGSRfZkxNkMyIWQ4bgU9jCx3pfi
XbSlltdJ812WSnw1Aq4dt4VsAv856h3ZL0LTCN6aNWG64jxAj6CJef2GTm5xJv0drNFPLUCesJ8K
Xm/d1Pefup27lP9x0HkC5DmEeTq8jaXpvzD4otUXCwXQ3sV4dfNNfc7tqMZPoawlorp4parxz/lh
scZG2Uty7Pnbs2vB3Jykweh+ar/o7OsjP5luUn4EOIKGlHcnh8bBIC7N3VWdnWBM7xFRK8WyjCcZ
PsIeJYdns4ikpgxtyqZI52xrcvUV/iiRQLKPzb/4Ku+Rzfu0nyQo1a9md8gJlDcBdArM6ooAARLE
GBU8vOfO7oIz9rzQ1pH6CQfPw4rL1xo7sDq3Cy6H/ZZCpwdJbuLwtcuKOmImP9yY+QAOe4XJoM3J
rdB1XuQjZYBHsPyys4MntY5QvaTSh2yjXg2tgwGnjsbPcn4XQ5Wv5JZtb5DTPsBYXr7r2r8XybWX
ojF4WHHElMBiZ6hQuUxGP0l2XIFRwyDW3bRWUJ9gvfucOtwpUVl6t2exsStEZloa9wYZWL1PaJHj
IQi3qzmqbAn0kB/vdsm1c4yxTU+PD6T97DzGzqEc9bc4dEMsLJ3JBAZCNPEjR5OXWEgdSSSFafxZ
LkZ6fENMs+Qz4RiLIT0IJp0jaF2Doz7rK9hTQEPYBBgL2P04ZrgRSjqDqyHLq1Rg7Kh9CdO7xj2L
Y3xJ+oROnEOacoP27qpjNUtWZiKErKTDXJMEHB90S7qEPg/oeOHJ8cE0N3ulIyOryUPmFo8+KVR4
LSzmiOLat7/PB2hgyx0z3DDTRio40X2y6HNKR1bYRspIuPh+VET4+ENg+JNtcni1oEH0+iAMToOB
TG8N7ibu1/BmNk10JB1hJjzlZOFY0vkR6SEaN8NmMjscuG/bnB2rbSMVrUxoELp0ToYO/jTm2Xlq
edMZS2a6XzDCH80B6TTEQX3n5BQbOOdn1GlPL4sdbu9/xlwvHGK8yIK2Nv/YNxDFEwC4treJ1YWR
zp8jvILh77RBfUgyp+Rx5KqSa9qMhF6fYYeKnDX5BkDueLlu6jxhSugRiJEiKHFDBuzUrKkqK8fb
88D2tDi46d2sSjFYOWJC6PibsDbiBte0ttlAgWXq67G+APq/Uxtp6A+BDTmpkb8/sRa3lR9jZyIb
krIy5HckA3ODPm9wn6JK5qEdpWNV+yUWjfuITmSBiDkZok96VBcGx3571/7WT/yL/t3Wm8ulHYrF
HSupTZhkSmibVYaqND3V/HIlZIXWFeiNuoyDTQnr0L/9opKIS9WBaLw2ADBxWjoKDWq/xsCXoXpW
+BMAWgBqePjfgsjfZ/gHleg/ssPHu13WVjU+hpCOJbzkzX4/QB0Hynalg/WUsa7gORbWWOtIOOZO
aII/3w6kwCDQZWc7VtJmJVNKgRVGKGqTDxgUqeJq60IwMenp+bhoKtdJq7UEezQvYupQ2qPX5eKx
mKUwPQqwAGwFSuQXJx0Y3lKrSGrYOSNy5zGFrIN+OZq4aFkmZE1yTAmh6jnmoizaasdXDs+YNEek
5KUcKJPzly8NxxAfNONERbbBUQYy8h0bROvGr649twel2PW6eEgHgKz7ABHS4qoFhvyHwZupM7Y1
7rKLxHwAmIDISY6Km5z+gTiPePoicW5FM2ciJI/NAyW05bELbL0VYp76DvjBEd2m1LAQ0vlZDOxn
f50kMTUxmTEcFQSlF8GaUnc49q7vikFnTahUsAYfj1JLOjcCV+3WUN2RkiWBivWiWQQ3tUlgDJIX
bMZ/MdYOJ00yBzJatzs+bjuuOUhYKe9wpVpt2PV4iab94GiP7zp2nk/5t4fmYwRKcBFjWd3fugAZ
WKH51sb/SN6JnJJnbI08T7qgfOUC3bL8WMs4ATpPIw5ITSV699TzFG46eZBlgAexUdvdz/+vHugg
+M/+5VObwo0xjm2lPI4firJL9x4xHrFbnXIW77SBXjUdrBJ8NnnYYo2plkzJJ8aA2Hf8Yxi88sD8
x6jQroqaz2vhFpM8Q2YzfvK0VbHHjJ9VAulWENj/sSCEwUSOYBtYVheC/VNFo3Dgl+jqrFLrCsUi
7QUqO5MdIc/K3TPGQWu4+jppAlKqR3FPOWaEnE8WCBqmGSSU6EqL3U604mQ/mqqZQYFH5EjnX+Q+
5M1lc+fzqWo1Dsnl7hmJU//3F0fJCngwAj7U9AVYQsU5fJleNT7pYjg4CneLsp2U53AE1mbDUaX4
U4Xtp++jNyP+v4k/DqNXX9Dl3XbzmxT7heCU56EsRDjfyFaf4YHbBw702RAlPnpgajDxQWyPLBrZ
w2xxq1f6kMXYWhTIW4Ab0ECxYPwya7YdQDEoDlKyWcju6glXKLKHAvMpKvDhGadppAisf4rbnr0n
OwoCzBANcochXYowbIwAVF4ucdQyDNyvqD6r4cQWjzRYyPZwkPpxXcALJE+domsp3s2tgkKH87IL
qQIvYLdEnf3nCpEdc3BgLWG8zEulFXL/EzcdvCFiZma1IcBzOQ22XMz/Cx2pwtOBT7+1BU2mDC8r
Qd7L/V4R4NC5UNpzmTFQ2xc+Q/DHro2yQxE3l6PbOY7v5lKRspyy3gjLv9r4JN/+ZQii/RzhAAYD
8NvyIr1KIno+MMGL4uqZ429tLz9WQW5Rd+IOwp8SXJRX5w+c3cqMjk9wJyPQKKDYgG0/RkfMmNCW
t/47Ku+U+fOFoxAPOc/QIpQalttwzLn735tmckGReF6on40OgjyEDXLvRemNULkxUgEsNa/WcqNi
bON5s0YUC40mpUucdHZZLhr76wg77VcDFa5oSB5cfOlKlTaZfK/q5RSI2cTyV0PpOL6mCGtylm3L
38c+uf3sD8AzR0W4S0wnzsLcbUakPxb8v+gVK0K6wNwb1XMVf9scQUkGEf5zmSO00OVFt1i8/dox
utST/r2Wo9b1+sLPBgfg6u3zYvKE27FA+OryHDqPNHFNpE51Qjmsr+k6U6etF7Fxm/cwrK4Opq6g
sVKmLTCYhLDK5z5Vdtn230IbLzv6Y0MM5/6wPIW18jphBWWQQ0/3eXEDXZWLprOXSocu6STr2NrO
ns4YG/kTBjic3rYyl7Z2WCjdVekF7xKwFFjj
`protect end_protected
