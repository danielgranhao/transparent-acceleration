-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Grx5Tycn4wSNWMbX8Eyiw72t9T9eJWHLtLEcgSfGMbLQa/nDAjRisHsiyl68NvJRNsGofuc6/xnk
BpKghh2UhMCekiqzvV6OI4szCuzkEgpf1JS9zwXPmWjJo1cxie1HoCBScgdGUEafjHvf8HdUoBai
Un2bzLWDWDheFujrjj1/LaEo7/bMZaaMVElEstaGH7UCB7sxqWKAdUQwVmwANIfNbVe3UXPYWwMq
GXMuTzvkSfomY96JzjlNkEFknI1iCc+1gLER8BG9zzGYmRv0+UQI9kpKpYAOFYO3AV2mzLZTKLOi
aQ6EAXt4eSBNVvRgzo/7XC+ldWtOqa8RAN9wPg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13600)
`protect data_block
DjPVgtOeQufNfoW4Yj+Y7N3w17em1vrqOp/czWNkfg/fUI631mt7ANVAVsiIWj+cizwMSUz7FIHA
2m6cMmiirbXMjFRY8/B/zkNms8dxyNu/KfT/Es4CzEh2sR9+gCO0EVb46oN5kB3s6oVu3ANHYyau
wtS9fUVnTyCkZeqv4CQmFXpxlpretQmVVgbhcxcH4wIFiSRUW7rDeMOXxhC3/zOOIvQyKm0pLfFW
3/Srhz44ssZOLsUjkggw5EKp1PMA0jawvnjIeN849Ye6DwSjscUzaXKjNwvofgqnDDDNab1Fyl/T
NJl5FnaqBKup11c1XnoCXOx0U/H+lAEctO5bEx8SceWWiHhBL0Iy6FGn8lDDX5D9qJZIZjpV3FO6
Kew9Skl5D/yNg2rEJeXuOQIOa/n8OOYpxZA7qDBBtQHwdmjYdhsqpzE4ZUphbUNdJtxPiQOjR+Wz
ylnrLiWk4KxkdjJcpTfLL5ZyNXPEtRZf1UDlQ4nDO6I0YBYH+b+X5f717aY9U88IdchlmLcBLltY
enOPxLt2vhhspBQLstjnE754e2dZHMmM5hbcE0QzJXbL80CepQnPoiu/FX/91uwBfhWuKQOOphKX
Fko8o/e0W7vGe03mWDEO6RTk/mE74Lk0RXroBMeKlhLnSsykU7UdjGMPq/UOxZ6oe87WPLAuvfXS
8L5aiIuuUzhmLKNFsKppYjEvDNtyIBT09+OhmLJ0VvMrhRsrUCMDvQPz/fJE28KdwZgEimIILaO+
9fl4v8teFX55DSZDYBDyAKVF9OT0B5/dBhlFyuOoMUypIR3R/sns7qcWDEWur4wSvWw0AmxYc6v8
whXOjl8rkD7ObSFFNCvKHXa+F1NvVScOWzdDTC2uiWFRZYMxRzCkOGzxVGMVcNtUjjZ4mYtXI22h
YlGoQaOqwiFfUBNaOBmezm1s7HgmQtbxUICnkOjy/N3rlfpv0W/Qzbl9WDLGCNA5rz5gOY3RA/U1
EAgsCNKjSVn+GEC9Pd6rgPJQI7DmiyyQdmx/a15vSC2Wxi+nHe/EKfyeOFSLGdcc5BDeV+epdV5L
qKojQi86vBYZMslgGO2kgi4qapilhToqx+Q5/Gta4F4Gc1AgMTFKG9/mTbW71rWH+DcZXvXNml8u
i70S5fYVkU0fEGEI3CI6zjPkrGHSS5uxiukJ6XZFYQ73i8ngKqaoDQZlktLUDnbwvW47obG2rszv
v768KIOvKn/39GATMg/Zdr2NeE9yIL07juyqfLwXirxTfYf4I+I/1Hh1wfsrZBQsSI4Xp9JlNztp
8DcI2hwCCJoGIvEM5I8haJJL1rPoJsYJCcnzAGbYf3Jh1+SMf4kji9mJKOyuYzSFixvdOdHFa/5L
bbD2XZ/vhxzNEJOIyEifCLOxQaGuI/U+xzzemSSDdDfhbnUY28eRuTeLozax43xDBSvepwv1JdPQ
3gWobCsbsorUfHunfz2LmI1kzXFGWaInt/ZHlEW9sXyBNp9IvqzRHJg4SvskekQfbY9iJZYo/MC6
+KioRJEqkWu7VDcYUmw44wNwQHyu/Ph0S9Wcd6UypSIiDBh+GtihbVsOWI6bJIt8ciVhridlvktr
dIcEQX/vf/jmDKdo9nzxX7QKTusJt5i/WBsK8uk7+IoeuQ7LmGvnE1IH6BkjEZAMaNojY27v1iEQ
UiZX12Ni6ufqsyMjkZF2NPBGLUSvHFxfNGSllsGHW7RDKxKkN/HEZNAtBlRwAi3zbpfoNR3LXm6Q
d0Rdisaj0RmzzUHYv8wcGCtuPWj5tO+8njDTkDRsnOuG2+NFvbogWlAvCoTsNT15sMpUkuSV0GXn
9BtFPNRuI5+2VEZCFh627zP1MuR6tPCd1W/4VadZ1rPenEDcfZL8/8hEEtij/TY/QwJ0wvYpwWSk
LiDAYCnlbYarGo3TTGE92ZnzIE06PMR9KQHV657OjPNd5kdBgTVge977/OM9xbDTX5TeJnJFf0x/
r+zfWBrPgJZvGC+EzNP0OrlL/KaE6sOyAPBIxNgKkty3HuZwtdbe9EoUB8IaKkVV2AxXwY9RG73C
rqvTq8zLjy6rSLYSpSrZnJ6BmoCEN8nkDlCTJ/DE9X1CCTTHz5YFlV0QvZzPBs4HRGL2vuWiW7vU
M5PumTvymVRQJcWO8VcTV9UiIDQF7DGfH1foKOCEV2hJiB9FqIByAiMrb4UyMCaTFV95zs1kT6fJ
yQUPCGogCOehFoSk+lsfX7363BDEdBl0hmRq6IwD12pjMU0KS2YS0YzCYj8YQ0BPln0cI55qrzyG
gONPlSVHAFSn0TOE6Lqrp5565/u4KNZ0TnzMrbjolXmom0mPAX58ZZ02jwhOWUp7MPEa3CfNXJ+3
EmAso9v2QC9wglhjSgY1ZdAyX2RJ/X3vVDzxrKRJpoO4kAMtjCL5NobpSUyWwykMkCtpRrl/FaMy
YOArLn9PezXJmgRhpeMMGPnj1UqTfkKaOHaaUsi1ImjN5CuuQ2wuDGDqtpRO0FATnDGZ7jJGzv+/
lauBWnYEt/v+rjv3QGoKQao04NJiA11nbRxdxaIi3LzZw0bF1x5xBhDRuvN/6JSKY8tQ6hVaDkk4
YeyQdp880fh8n0IH/ISZN2JVL431veGMev++F6e6YgK0LN6ULYeRcA7nhLFIJzGFRhZT9NQXJhEb
+CSbiTs5RqDJJvSRhEsmH7YZeCRJtvc1oWJ185w6fDW9Bk2K2hC2A7S5Pt1ZCyyXIIV8z3NwclNK
d+2I5asfjSNcFJyNgY7Pk8VU3txuCmzxUPhH4oZpocf5i4qvRAddsgWBaqhBKRA4s9JHHA+c/j8W
PbYE01hxL/P8E3exn3S35YoBcuW1WgaxhtADa0zQB+mbO1Oqm9wK9M2Ym3+2+U69KW8+RoKX8JYv
YMz6zF2ybksnse9uc5Ii1vFRm7nYgVpaVSA0MO2Ds65GGNi6bYo0lLX9i6zblGHPgzNLsj6Liwmz
BhJolflW8ShrQVz1wzGOMWIuVCuAc7nAD1pp7bWz2cQdd4M+p/SDPS9ZkeuRMgLDAdvjBgdZ+ezF
ocdExNbbUDzFqEO8s43ukstXBu23z5RhKB+3Vac6j/P7RZdX0HFGmEZ07dcwGTEjJ9sTW6xgvyZn
qYhMTF7shXh4Ti/9Jn5kq75d5np46za7nP04hdWn74EvRjtDN7Yi+CeMd6DxzyxutaAgknBW2qSS
rSS8kVDY2hmtuw4PlXPvJ65ku+FMusfJLfKR3RN6eUs78J5/qWAJxI6oENlytTsCDTTWnUs71dWI
q5WxDgs7Z2VRrRHJ2WriUdaQAd6esJVTx4qBT57XgHmY8dDmYtBfz8npldNc41D5RaO+7HPFXb3/
7ITs2OZoPQs5Klbb0GOlE1P0Nqc63NU1mYcS1AnnFXwGAS1tSsETaE+KG7BT0acWZ0C7VI4v5H/s
/i3+cNGy1ezEQd+Mu/Hhs5SuEG0KueAdnqPkPzZYco2ciZ8miLDlTOmB0RF4COrh6KjlaRfTsZbd
eXqldnadCchI5/hLH3M4lm5i5r1uTSh2dKzbINcxNf4/A5JMPEP4JQVhLnfLUK/NRp9h5324MOUl
VXmUtYAnxMgH5tLPdNKgyP7x62Ip2PdnbNuCojr07bROq6LQtoRjZxJORjzPkaEVumWg5bt8BJ8o
IAcz/BKynb5yq3hbseTdevfiX34c3K3/6qjavQwlfa4A1YwFGDsGHtfpSTgcgxPlbSzcPWYvgrBI
HoXOOf+KZl+BhPaWo3VL9aXIMhIrBHJNksixoHDK3KgJ7tmTNXQYsAOGPVqsSHlh4pnRMpU0ot6p
rgdqrifsLNKG/FJ2ZmJXg17A5RzRgn4LeSD3N5+hEGZU6FYZTMabTgdVkDObw47R+hZCfJ9ueMjG
5I8sPtt90TbbDw+tsWCrWJFRLs0TO8zYkRdlEF4uVbYOagZjUg8VRQMsGT0a9ipQbH13L3XH6X42
ceMUn/Nf1z/xD/KNIWn2npOaI8q4fB9Cbsv8z1uBsUIse7Lj90CYeANoQdiP5ewZbh8ZSeV9qf5k
4DzO2dWbisAMwsOEB4GudaXqf7kUInVbDQdB+UQ6Z1ub90vulBod3VGCLX+fSopxEubOfoMMA1+S
tG/mp09G2hQv84+l9SKtaUeOebI8KvH7Go8FK8gZwQvio2HrusaiTVnLPVGj7o+Ru+JI+z22OZ5x
wEL1UEL9Zi5INXLbRqgHPblEjJNZnoHtct8dEjHiXhoaGOvXutVhC2SIpDhLKurZayBZhLVbPP/E
cimvDktMpyfC+SM62u6h56EFP1UwKub/nOgJSCxWGPCStf+2rKgVbW2avk0etGAZ1azjEwIyXeEZ
26mH8K4HyJ/+eb9nArHF8uCGm+a+dqmKItZdYbdEbeoUVAhM+MufNO+0OD3+MWtjp3ImJEJq84kJ
vhFLqrRtyBSWjPcQut6TG76JGwrm6/LFo5ooAr8vPRpCdhhKdgEWArYIgw3w7SEtukNsxDxTJsFK
HK1Ssv97n5ryMVJBhdziv4+fThypRbUOQKRiniyClwsmzP7gURUINARCaejLKqNFZdT253SCzs8w
DbDYjgCuq9Z7ze7PZSnw2gdN7EG5jHpd1WKXF/BJ5jw8pm8xXxNuz0l5afw72JtwFRaF9HMJK+Pk
3as4Sygjp21WjHQU8d1Uuo4O5hgk+p7mHjTigb/aq4A2I4Dywn6xTSSBoz69IvU9ndkZ1IRj6Xuy
Kg8R1TlDrVEcpmf1iPi2uCLSvencQjxYwa/y8zCoEb+5TJSDDOBREvFWkMUb7xiSrwS79Ni8m4Sh
ewOBR/XHOz6pWRjRLNYDrvP5n5Lfv0AgC0uVNc6yaBDm9utarZszmvqhpE1o2Ms5BQx7tYS0ft8O
9LrtJNWuk3yaPacldzLRIGxPp6RvFvZpLk43IM+MDnEuDIN2ABjAicaCr21utPUgA9SjnNsBiShG
VXc/nEfb37eRJW9iLXho5CMqAlJQ0C0jDkWkRpDDh4hEFI08ujgeVdHGfcM93EMmjOQ881KhWDIG
hLefCB1deQt7fjK7zGt4kddNW66QH5+BHD/hbcPFh+Q4qDtqBSgKFdBxjbi98oRpo8Vqgr4prbpw
JSBB+dbgTh204a544O4F5Gj8bePVVoxfrDoTMFRIJJJyeibD8ceEP56oATiydpNEpMNKnqrcef7h
2VuYKaA1yHlP6tMpe+hoWB0JmB1HKUfG2c7GE1OdG0mwtv94sEUCfBX/ysILD4JP/zMmw9oBMw9l
vLMKb2b/tq08BsH2Vdpk2NG/cUXcVTm6Icu/81LEn5c6SvXJKoSAWoEJFrr1ibRbt6syVW586DW7
t4Gz/kS1CnQPDOlAgNUn4t9R8JDbTHO9azFW+c8jsJ+ZllY+eDIfhjBnB+UFFsd9sJ8rVqy4u2xu
NMEjXrQofYCS+Emy/J5eo/eawU/6ZnA2cYePovBm5JIrdYQ5+dfsz+Ww5VhyeUzTo9ar90fFZm5X
2wZod6oWmGTBDFZITjlc4I86t1hZNJO954N59NJgPrE0pHSL7q5ugsMulQ7JdZnEqWz9XS+UQmqg
VkNsXeWdXTn6P1t0z8FMUlXEXdcqWz7gECp9Vn1wQdY2VNe74GX9pjpPfguY9sJSANaVCr+hTsPM
+3icN0ZRB5h6Tjhfk33LzHNNKej1ZkDYbGauqVE9WffwLHCQ490u04FvK/QqiLfzn19ZEMjXARnR
kF3r1aJAj1R/1cCXm+HoB186F5OVrx816npf7v4AQhKFJ6gla3Zzc9nRHlEmpgTLZ8zJzilNkleD
dEjVPzWyzjxmnJBmfG8SA99Vi/MZ/7lsEBZKDOtN4IiRTafsObPBVl4K1HwSfXJwlHMdPb3UYeS9
fMVfLzoDd0RxXR0U3bsVXnqJHP9Nndds+Qt47LPgc98XkcwNXnwFVGbRfuRZTf9Y836cJogfYl1N
OpzaSoNPRcD5OwpVJdQOglVAV8ltYm042+VGIyBmFQ7np+KddiVnAF39qBYOaHsHy+1YpDp/2xRB
mUeX9ZxZ/UPkQEkKsOsr/e0/CDq2DwUxfGlEiw3jwiQpfTz7p/As15rx2t82fZ2juRY1KV9iMwt1
8PXek0q1kL0uOeDe1t0p4TnTj8bdaTDt5kFyw1Bu3qeenoVTTkRzmQ/72UTNFOo816hABzhjCQT6
EBytWYlSnKBO2e/ibGTx11HDXDC2Ls1gpmYwgreP6rO0ADc786yxkcNjOk+E59hS8zWLwWg37fMx
Lw+ro5HNkt6N5E7vku8NAUfoXzdGKiK4O34yxYz2OsL6+oquA25MXS3UpGXeR7IKQr3VQbTcj92e
EfFmmWkUoBPPthxqEwsmc3RnOOOXQORsAAB85o1f/4P7Nte8S+EK1wWN5NX5HYi+TCOWYKK++Cte
9jMLS7Yr7hZRmMFpCH8bV71iPTRyvxYP5jCgI668O7V+QqSHMP1LU2a5T0cF5fwrj6hJp6TL3TWo
ICudqx6I+tfhNqrcUUjRfB2gX0NjZe7UWql7aktzdGpuGWSlGfIPAiImv8DJ1F0CM4YvqKkdoiQB
StOH1VZ1ThOFS0xA3b8LupMyZ6X2u4w/8uFBeRXrrmAu3y40R2uE4b/GxvAUzo5no2UAdd5L1p7O
jm8QRnoYGERVK7uenyYCXvlnwDc3t+hnZab6+EB22mhYkT/i7tCKtx0ViKFFrzfDdrJ8bB0TmpZT
1MjG17mS5TiyOaKOf0QVxM3W7IS4mzdKha3KTdsXFMGuHRG9InfpQUtfKWdB11RKlSYtGhdGlKo3
25tBRFXBz7KfKZ61AZojxvFU9laej+36cyFZgMxE2TFTtAPJMSvUGz7gg/7okUuKu5+x8gwBii5v
xUZJFpXFavTvETo0MScfcUqiJB89YjxP7p6tMBzTf9yQ7otS1exYq/RMEVTJSSXQFcyeYdM7x+it
U4fxeHh8x9lp1vCof0aHf9NDLNuGA9aCJUvItcU8QeNYjKwMRJiVNi/5lNMca7IXj/QQF8KcoJit
MV0a8B+jMTP3eB9Rz+15mn3ewZAXVDx2V+lXqpzsQIVExw6EIhTkh4WPk6mixil3FOShvH4Udyg5
Q7jCLYpqZJC2o8ySncx5dHoItXQJXW+CdMGdc9f71NToMoGyW2FF9IQ0XITHlg6+HPBEwx8ODivt
epzdKXJSfYTIk9Ne3/0rrR3Yhm1wtcqh70N7bHjNXBVRJH+EG8FkV+8A38sT5ClI0Ud2lZDJKMAD
LZsaxcFqrH7qurKOz30VAdGsF6W6WQhxE7P3btvRfWJoET7NudQJYSUw1iJa3iaTl1XQByEhLX9I
ogYvolwm92Gp4ErNcVDcpx5KESyT2PeMQGTnEhi8sQH/z4q49kbttBqLFcl+Gj5tsgkWxoKKSRo3
rbpfXXBgQxGjgAzo3+Vs6i1+5p3sXKLjO58nKHe3CRCt5Lbx6+j9SXWmRa7+VZ6o5e+gb8/zJ8ta
WescnbFqtOaN6r5HB85gLfJph5mGOgKcn/eZk/9M9F2Yb7zKdp+V1crCliuhk3iodQuqjwt2Ul3s
qGNZNOGInqw2sLUwPMq2MiZsP9IiR2lxTKwcMd14fJWJMbcw823noTp4ZHCRI9uLJQSmxTZd2k81
w7xC5K1xjWhiGHU8FrhtPX9gzoDzA6HfpepfDgSKRavJTZB6GD/QqIi2BoBtAnELcH5ex2QMf/Jv
2MqCHcxExK0dc/WMtA//FUTjDnYM8DvE8XnTVjcMckuOSzWRk3B4c1SaIl9dhv4oJ3esFXls64Mg
z3WZIUsVYEbAYKFQBrGrqb8Q8iMzNh00xofflnMVF2HZ0SE+LNjPY/aM2Nz6K297jZ+dHDHWWNq2
FVmT6spyDb5GLJPlhBgKLqDfW5ohQq/lmH3+mgoJIhQ7dJMVtetQiC5b0C/FmXVU7lBv+Inab1KX
/oXP1Yz83gbk5K4U+UuG2csnko66msFTCK7cDe9w7mwwHSueOQZJl4GeN+k4NQh50GyabK3YAlxi
H8nC9sR3GmRt14nvqSnASVOybkWP6NDn2cCtuYFZlCsYBI5uGgF/U59RAwlB3sbckfvenchFuHdJ
085cuzwiLIEy9aqotKCh4i4eJZEzAtZUGJWxXZ8B7CPmqArJIZTEGYTiN2OLbY2/TuoGefP0sXU4
xVo+qpBDFknGgcj+7PgJgi+hAhAnd9gc4j/qiDDcANQdpAoaXVvZm3+i47XuYoh8P+A4PiL57qGi
1hYPrt31obD59kFDGGqafoyH4kcHt/1m6yR6ZzUpeMNFEepEi9yxfemC6I5FJIpy8znnz1TnAT3y
yikv6R9EerrV9DylHVjxvNlKNCtzUVqNY+1yJo/0+QXflSuYBQIomUODVesy60XQFf7uRHF20yj9
2SAB/EfC3GzPqj9Zh+qIkDisFYmn1esBj+Vn8NL7zlj2sOBoGVIIec/LsTuj/rpttpIWKvNsZEkw
gtkf+pa7OgDMP41QESL4rR+yxDR06mVk8zdgnZNpCS7hxA+V6Sm2TwCa1XbB+GAzViFS+7l2CTAt
IDkEl6KVsYLMbWgS4qHoue3mhDv4RT6yAaINFDaojH2tkNtS26IXx2wWSQ4LfQvMZFcAAH9KLvpA
2DP/lBH1+qIReiCarrPfbNpPy4pifguP8ULOupC4/XV40AloZy4xO8wCbWQtCLn6FY0v6pXoctih
QC0CSU82JuX2zi2QWZ7R1s8KLoXfe9B67ATAIu9vzw75v1KwGLAOaiwI3MhEdZp5lXeHNzo1fNZW
u1BpVDBbm+SM36GdD9lPgaVS/UkOYCfIW9/6lYOPcqrxz66+8e7lOaE27R+kNVF/ljDF1qFH6GeR
PaOXRxaiLb6ViEUGvi6CenrHEmDAU4hyI1UyN8C1b+KIZpNLAO2bxJ393VM0fmqXLW+T+Gg1qgCw
fRkj5oT6IRbVgCwynWGJPbHidNPir5FgFmD8VHPaONkBAwYVh2sQ6/llgELQLWYXEVLNVR1u+89B
3O5ohyGH3OkggTXuxdcGo+FvKLKXKHWJj3he1gPGoCWjrVp8AHlp+OqPJSHXpV6VWz7eHYND0e+f
ij0C6WOzVo3HIE8dgNLSUpSt+aQsbAcg9J3uqjqRGy1sgZufs5dmFD2fHGye6JEdI57+hehduoDl
jbVNeEEFXh0OGU+jWf9dM8HDXYgcvtlNhj4uIOHkP7IlS6yUPhY9ztmVUfH60cT6gsNNJipJWX/A
yaoXanZFWAu9piQHj5UDpLKcAZSgC5cMRi7JNNBTPUwLWpR4oMuyRycvLjSF9zYWZ/5SgOBa3kOA
8STb69YKBJOhR7kRYVcievFqcg9hspOxeJrGAM52GE65xlikuTEiRAty7UauTsBSYevwQvdZGbwi
YQO1CkrW21bm9DcZzCm2nBCj+Df8Y7+n1loofvDCjxZtE0Ks4zyrFqTY1iAlB+q3PfFjDRlaVOOH
2PdzCjZehWav3HRgAPjWzdD7vrfNKHdRYghWDDoNa3AIptZTkgIrPPRqZa4+o9XQ5BJqCZuhaFvJ
4KA4s8H4XOsfrZX3GoTF1ZtAgM+OPIlsXPGjox9ANXbiWFOW92hgW8LgHF8YP5ySBC8vORhxocCU
dVjQI1rrRSuDgCCqGGJmuG4qWNZohu8fiGloA9NMrIkxNm4o2ql1vJdovgUjM11DUEEsL5DO45ak
Ckdz9nyx5vpzZ/kYqtuKz5tN3MPE1dajogm08RZE2oyf3B0Kufiv61Y3RWQ7xuVUocAsH4DjAGGL
hPUcuylX6ncCKDQnFGoEd9Te16sFXlUxKYhuXaZWKzIsvEOUBDslEV4yFPU61eFIszD9PzIfSS4S
HS1ztixehJG0n9t6eHeb5h1QOWIFDGNKMIBG3P73UpW9LAKBuPj+WZ6Ok5qLjx/q6fBf+FB9ooZT
cjI6JBT2gwolxPD2Hwa7gxbDdbft0St39OHPc3LcdLrgHxTzOM0BDad7TKErUJIH3g2/0moCFpuV
lGZVg081iPSmYvTUiyNDgx6BE/0X0SkqC5AERdRh0G2bX7hvQJLnX6mOpYYjQQ+rmUxlOEi5GP8B
1jKBPakxZBUi0DaOTRkxPPYeoiM/Hjg3ZlOwdc2GYEbhg4bWvWlJqNLK4QzsPBSvSEBClXo/K2QF
qj9coin7Ua4L2tFuF0kr8nF36P4PRvA2nCYVEdgdaC6wacKN8EmtcQ0B5HGDufmnw87X1zbKXFAR
SQTY67ZSFx0zVLE5wi5PdcfyHjcDNrPnp0z0aqSQda6W8Q/F7iYi5SLzxejPbgdy/GO73TDlzSiw
Z8UCuF6zkaCqkYDos6jPGgbSjCld8cZTx7App0gk7oXvX3RlL4kial6vL5MyZ35NjPuHvEHG2bg4
eBe06r8VNWIVq65QNsuOFeDAfrnSI52BKlbGyEqKy+ZxM8+gW2PsNJKAOxCGlscHT340+nj6uHda
JuclI1tVzlm1UxDExt3+6asZgqkoBszs1/gMVcmwBUUHpqPknZQ2+ViyP39rBjTWbdn1ncQhxCmj
HUkOiR8zLTuf4EQtgunHWbFrGo7mRNZ8vu+HY4wiAlpwF65u6I/VRGHu/u9dVtU9fvuVdqXNzSy3
IGI2iY5q35phnbe0G8JXJZ9kE2SfmfIJ5LVC1sJG20Q8cWaA3DO3Y7XN6jjHa3A0ZCL1cRUt2eIy
+Y+jojm3yApybnEL9mJ2MugZkgLjasCTQ9pzUCZL4UECenvEIE7Ki22rY1AYClVovHuGo830Qv03
kGkQ/LZmB1mnuDdQmN+5HoIrzihgzRBD/vrSr+XEBnJ6p86na57vlHloVwlnukrPnad5676zN2A+
zDRWWSKS44FHk7ZegprDrx6iR6tfq7i7odKdjF3snUhCCHUJMfDQv4w2IQDhHEaX5d3glnBxG0NQ
2GGII/jhY86VHaNRB3xDno09wl/QBkDrxzI0fpwhm7xBgkLsTfiB3nh9j9/DVO5y8gsOMn0FaPXl
OcvvFT//JJTVXDln3zhcnkqH82YaqTRxP4QS4ztAwGXfEGbMa1ugrINCMr7ZuU1Rfna2hKpHNADD
zL8SNsGQulH4IA6finpekbByOFksVAkEIBS5GH5NZQM+qmvDnGqNbB8zEK8fuYcRsRxn1Bk2IJuB
qm20MSItX79BqnpgKQBOYxSECRS1U0FzDbGLzP6MbY3/6Z+36QuwcC50QQQ78qdZopuU8JO6Ba5C
49vNq5N6g2+1nybGIPi3a72Ay2ZOm10K0ZF+2w9xA3HELigsdR7h90xMirplHF31jadVVSlwI1Dq
1+ScWqKzDx8awh2/KI+Ho1CQs/O6t+ob7jhES8Fu2vNPKAKau/mrgKSsEuyGicg28GD4VNECVKw9
RH7AdztHfemY+TRJ2MZoDHoYb58OV4CWsMxUclQ39IN3Dq+6+/58eOa3sY3DUj8v2/LJ4Ey5M7mz
CE3eoKkJb76ynTYfKZwm3FSlhwHKtVZyWT7UspdCNhTb9G50AlOpPcE/umgiGI2DC2kRBNEtiSOy
jSXnMsORXxYUr3oaByYAsBRniUIBibkRppiQVZxI+IY/VfoktRQ5a25kebriU9JdR8JmsnhpFniY
UDRChJLD1jxQP6DW6/6PqFobq6lMyO096TALUddktIEeqGCqWGtOWSvi2yeHas3gIOp7sJvxaMFi
JlDSK7w/gqGLbGzTQUldbOlPJtfqfg2IZtFKk4ogXyeqmWxS+YXGJOhHsgG5XaURRF9T0SjZ9Gb+
j5DVKEvOHmnBZ0tw/8cWkj6FWJA0CHkJmXoIlHytI4lJ4ym8c3Bweo19Jo8WrA1ZtqOFz3Ti3GwZ
cSiNd+et29HIyohRhbgtuhOw+21TupaUGCTS1f75+FFicYgb3v5JWQasVvVyQdRNbSktFt/TXOiJ
/IU8AgBGQwhGFwnpAlKPHlsGMUsuCIfnNFiCPss6m4eGLdVyK5+/UUv+4i4OmDIcLF2Jum6URokC
o0zOcNk+SvVYUm/8KH8fWSZFTko0t+iHDxxQYh6Qe3gMy+rcJc1JKm817NwceRDCzwhSmJr8LVjm
ud81PFBtcnbBCAMEDTn0zdhjRlrzfLeZLCRitwyLo9eF7B11dLsI1sWDDNwe76P1lNwemOGiEPon
PQLGnkCUHiI4bK3KdzHx4HsrxX4rhVqTY6SfpmZGOMxs1fyeI1nL+CX1Wu1pSA0u56YJ+iKImCGm
6FWDjfyM/rUZcn1ag+ZF+IlA94IlpbLvf9OXTOeKrW2Pik7Gv9dG3Lz3MLaQYPzy/tK2eVha6QdZ
bP5RPBSsQTPeOne/IZhCsS9eIKpCldYORmJNXL7rW8FeRsYSHykKwceRzAzUq3M3Lz2S+OCQZdoD
ycu8iEJdrdrTIxj3opUXE4smg+80zYLAYgF/ztRcfCL1EK2Zx38HY+w2s4/UFSpRifp0hcTECt8b
/rEZRpzzJlGsNBGYaZhgxKg+/LfaCGLl0vynMgmnyL7kIgLtPV/vqVxzvmdsttTI+CTT4qcYLCux
uu8svAkX8Aqf8sR0NFJ6nT3hL2NcLW/IWQIOeQD5Xyj4kf3hJyLIps0vyaTDHe2NnTJlPAISMXVh
I59gO1Fa8xKfRI7ebb81123DhulQz/WyIXMrQQj+Hk5ZiicN3ijxD+70Fq6L0W0xSKqwW2uaI1Y7
bDUF/AlSK6yhZJ69w6eGd0pEAjD2i4tJU00jtMADji0Zn1TisJy8tqG7Mbn8OD4fKhCUic2r6aRO
POdeskre0ZSsWg3ncpg/lNXCP4ttMb21ZfHqmjhTm6Q6lmwqYGQ0ag+rI2hdbr/1aJQCCXY6PlIo
4/yHZZ71tslFHmbRqHs2+0Aaqp/3pX9n0CuA+l+v8SgmB2upE0OCKH2VwZEKp+uJ+3MK1CVOEEYw
yLee1BVksOl3ciwRGyhnnDEb/Z8Vd1uFR0xk5RfXjE0WkDHKY6YpnQA1gLsEg+4dCw5xELL0ykMG
JYHZICpA7imsP5wC2jW9e+WTjCwUmx9D8/CyjfRR5puXioTO4jOKw0rVYI6INyFg9C6eUcLNoC8q
Ae9SdjGyl4D3KWlI5nZfhb1xDwHcX62CvSXZ/aoJQ/LBqYHJ4Pwr7hS5zsxYUcsk4dTlzwvi4vQ6
TkWYrYcADGYK9EsyXCBrooM6kJyZsEp/uhrJeP673bjsuRYCRth/u565VhXdTinYP6P3T7Rs5eaI
zaE061KukPdy7ZBZH5x+zHdZ/b7zERJKj9iLgbQPlIW8qUo0CNCIo7ouXhuH8jPD6GX3TCbJ1GMG
H3IB1qTXSwwlNsiaG0gBTTH9pzgLSggAgObS30SP0l1v1bOC1RXfQ+TcyIEBHBMJdGukR3Wsc6d1
4qA1mgMzXWPJX/pGxwjaAeiy3MJmQKtAKp1tdTNxr5ke2RWxWXC1/LM3GGgOTJTQTKm98pdanXo/
sToHP8anzrnDuyhukZfdrDdf1ZzIFLx+47MbCE0fz/0TsfZM25omcp3SUaDStDyX3WK7ICtcW70A
E/tAEic9/PcyBlMD9tHdHAlkK8jDJ9qpqCL4aSjncZMxcScMZMK7RHhlf71iYvtlmmdJi1vKKkNj
2vAUc4IK883mwa3jzPsVPmk7b2NEq4zxeA0bBvceYlTzE7XerdkTM99XZAueEf1E8Y56JZRsXNb3
6sW6gHM4aDM+oj9XfSW4kOx3Q6mJzU1kC1dWsUtihqK2fFolg0CCu9IZ0L36fFrxAQYhDAegOFK4
AjSbBhPgI46Dx/mHazHo68i1RN9bHu8OjnUKp13he1FKG9KxPGKnlmGNR9NhIEuKIQipSXkwAuQP
QSwgxt5rOUAg+l7l5WD8yFci3gLOS/vjJhm1K6h0+ZS11Ra+7bc9UiWPMKjF4uhnIgXqiKNy3KeH
VpOMJyQcjyOBIaxG5GeWa9ylYRla0098oT2NB+uNV2Pp7bFCeO4boQlYvwyuhiymKvh+g+y2Sgr3
PY8BjY/lzJSdKZkIc820sEww07Eih/231vEGo+p2PW4vNvngjH57bwOLdRSDsC2UPW71DWvpCzjE
k49zn0JQgvNIZcPBTCQDOjthO45V0/a25REZC/vyRv2qpmnY6rVHcB3n8SLqc9X1EQzVyTQZF3Wt
yUbPuL0gWZSz5ZqQkUckFnXOZYa1rowBfWP1aMERs7g57UnB7z5JaUOOCagtlBJNU9xrXxp/PttG
v9PKrPMAOlIHjyxuM9VusN2k+h9lseJGVElSIwzfZVsS/b6DLDsTbaQkhG6e7qayBQqwVgOasle5
16RXvI/mrcX1KGxPxmevNwlV8oTw4ytqLmeuM0rFpGE+CXCvqhv5yxLkMG/fyFXHyMbuA4J5eLuk
nwIfqP5ahgCj2wVgu6avyRIwk85dheqnxw0rJAQFKVjZURDgkh9gYxeus2IIOq8w9ec+efkdNXoA
n4kL2cN/d/20+ZpdoRQUvDD/tJ5Ob9fmG+oZQIOfJm+UqmTXso+Tuah3mmDEUYf6fmVZYSXS8nmu
KnuP+scx5rR0wj2wkwWrs+TakY0ggJj4BNM58JN26iFXCGZs/KghMtHhawQceEN/9agDAvOTOYUB
3eIVMz/Sz7qcUVU0AOUijCRsFifYAO/3xuCUO4h69A/hLi7zYE4FXKoEDATmWStugeueXmI4+WSf
ZLuKa9BwPO+z+S+IGNSbzKGEXb9BaQbRAI2b5BT2MaXzLAq4Ay3WuegmEtPD8/ljTrXXmFD+To1H
ND/1Jo8R6zHFQmuwK98MmIfXo1mDpJ6o0Ta6Eir/a8mpoUoapEndmI6COAQG7QEi//HSYdfD7uQT
8EyyCoyknkEZ4PyVy6QkdfFArbWyG1sbO6AeFULJJAUARD19nF+w2RHNDYma3NQfu1HlG0BC3nSP
7MKI2fw1A5sgS09LVhvhhWJyFp4K28YgBwT4oAnAlNxgt+YZx6cKKZMzN96pPJvYkXM7Us6NE0Ll
Z8r6fDXxgp8f4vakHlm4+tJ0QV/HK4stJwV3HyOxOqC5YMHRk3qxW8JZ3+grdw7VNASB4KJKHaG9
4/7nHtcG+vnq0IobLjczvJys8e2lMYe/KiGwotetA/FmQBPj2v6L4DH60Cn9UArw3PT875gKa+4/
64cemQQKTW/wkf6HQl7wK/G1n75PwXgh5Wo2MxzP2ki52wfzGopRWp4aAErPQlcSvDIjR+VYCQRK
hkyN5jo99JzQiFD5NGeqEwJh4j/1NPUJwHDM4wvgFYkujGRp4ECJggsVkXxuAAAJwU+oYfvrZwnA
BFS2Rxbdxcbt4P0+2MmBz4CxrpWBx3NWp2yQ4gHa5NxjJYItHZuOuO37JDoy4XkemTZT8ywgbFuO
jKwnaA0u+6KeYmPH4Mn7fRkDpUBbgX6HLKiGUZWiiVQ5LjAn3WSmR5nVD+lytDfGbwrWUa19QoE/
4pfyViUt8sl40+PDN06Gb6Ue8uP6nxwbbZnHm8e56pqhvOCoEwbowXVFVSYc/cgTWpWmdEnQhDl5
yOOUm98tarhXg3FijRjeT2UHh/AcxekKYNMQwha9kOO6TXzP6O/b2kC6GGHeoZnw55/SAyhlwf/P
FigE5HbSXMEjPBFyTesbF31/zbqR62HKj4BlsvXZT40DzLQ9z67/CLuGOtJOKB/SbLXM0BdzFX/k
/zK27svTPKQYNKtlRJRK6V0pp+DRfgra4570rj96hJHOenfc+5OWr0jyMDszrfTeuRnGJ4ibZtte
xmBBdT4z1ZWOrHrJczLNRKWu9iwrgAhDl5dFxHWj6wnAjzYVDt8j8+ffiRp7pbGurr4DPdLXO3S/
r2476qzK+p1rGVYvEQa/XryLOkQWtNhmC4OxvHcPmvr6wplG5YJcj81TCzNCRuLy0tWbC3Pz3aQ6
+o3A9qwlSo2yMs2N5m5oj1/HoO5L0/NNWDW9XP8lkTLFCRmesyW/KlPkiH+BR8hJaF9BgcNMAQb5
MXWRQizDZYpHjZIkKxo1Zh0IcYXbSeTZA9JhGx2OXYwN1B8BpDWXDjcXmim+w9BGSFzIeM5j/F54
w5acMkcIgagvyhWk/ZfEIt6ktfUCZGYScq7W9k/K4oe7TgfAxas1OP08bGdqzA3B54mm4BAt+zcO
aFf3/OqwCsCQD33Avg/sJ+ageJfnGOGuvCsm3WNn7+d5ZLigmffde5f3w1meAZLA8E4+tA9/nyaa
65VvOnEVlnZt/kYcXoti6Yump1ripSR7NXI4wpEDtzQZl70yz0kKSEeR08l2QXBVFbIZBY+gLVVZ
Dt3dhASzSF1FlUu8H/isCT7QrEZBOM3p+XhGDDYxAIa69RTPS/gXthmhTWg4DxhDd+ZB7tIlm/s0
oEul1/xNPi5gv1fGY6zyzbnO+/h6ODYYsS5rBErva8ErWCIgiFpnhv4XR4Vd40xKei8uRZBr8wZj
4r6BprkNdydTcXC7ldmnJJPrhjl/SQJmunzyGBDYylci8zdJuTsnma6FjWWg9bfZOkWA3GxP2Ck5
iI6jDgA4AY1TAFSwzzWNpZKIQa7ZmBQbydQL0PlyL4n+Ib11toqY7/lxJ5xfJ2dCirY91SoECdG6
LzeuPIs07hq68ROEzVfOMIEXAyLTbWlfggITSZSz7Ztc7KIhSOGzRQAJnNqZHFY6ZuwptcVb50HC
Kx3Yj5XLSNTRm9fqCPXI43LJItaxJH+sG+mV319SITC30eFfLFfy1Vs4TRydwi/TrBMD3F6HO3Qj
1fIWMyv6LjgDbD5O1nV3cA9878DRsAeAPW38yAHG9FmEZVuXyVC5M9SKtlvJOiwIP+ACy8ULhFz0
LOGQ9g6VXJ752nQ9aR8urDI343b5r0ZFHads87toN9bt5ztfZfQYp+MB63V8SpWqR4iwOnjzniV4
8CVsfqO7A41VQKRcp3Ku39oET4hVS8YryvrOff6HvkjwrTACIwyGNpsWjfplg3c4kyc98Ml5YKft
G3JNPJz49u6q+eI/dBUPbspX1b04Vafs/Gg3xbqHjSRyhd4bQ9fjMgz4tj19O7PlAcRBs1OCVKCJ
frpv9TJaLo09QSRR084TgEHF1MuA6kJen+U254WGtfJn9qx53D0E9wowoUeNeZPpvqZZEkNlIfpl
yBI1CzLPkBXLNe6Vj4tSbynxTzUWzFIt6YxzP5ZthazvBa24CNFm7xi7yWf4JqNu/73SiP7c6hOA
DGRM51RAmn12pIAeZN1PG8GlBcLjdeSxbzZLX4kiE+YE5IW5vhOSpJdIEabeHUshUrwYs6OWQuJZ
j40jU59vCBE/MSmoTdPpcTFGmkJDMyi/FH2geDNa0gMRvY5P32pc+X7RUaOVUyh8DXjnARZJNjLM
g15TRpXQILo+SgH0hUqhFVvC4Ix9MAgsFAxpOD0XJ0UijmfKyrJWlUxDm5d35f0skLMWZOJWOWOm
KZygeoybJirqoPhmWKvByIHLdblAbse84LA78x7HLgZzfpd3bX8p/7FJHgVphaKvuK7ul+ZlotaP
jC4LR1csoLzpXqNYXu8YZxYH/0Y6pDHxc/iD2+/olLRor08Q1o/t6BCS/S39HcqeFFAE5FNTNBqw
LMinFdrFIJeNHDxbtgUVKNIy/IeEpPvciVyCuqXnITPi1PVF35wQASePlQADODclr+AXOvjJD42m
LJh5xAEzXUS9iBTPq0F2IRnrCwRqxbKRxkLb257M4sxCiKv0QZfxyF2wPCmBu2Fp1d2avujtkvHb
HFdSiFitRpRWjXbXc0uAE4lhi7LOBfqiid4fDr/Z1gv8j7k0H2cWohixj5WHxuu/lobz9x7qSaQ5
yYnnJJXeAb3ZZebRB4VpCBYCYQetV5oa9HkEfHrylIwTH4HXeFzvEU+lfzRhIHUOrHf2DbCURDoq
GYYeywjcq+HjIxXQT3xcuVpfR9+6UaisHYVKZ4KGQBnyZrroPkg277WFJnLFedw9GysD55I1TTyX
ic5evWZTgEhyUlU9kJc+jloVt6k0dg0EFcio7LUcZXZVP6YnWLyU/X4fpRIAoYEz1NjShe8PP05l
kJP5Ib7kyz7nDgITcM21z7cX8q+KZrI4jw17BDUJVLbDfp9ruPS8weKTEpYsZ5YUsCMyNtsw8/w1
RuDH1qR3F7l9pn0gzSqTg2JZiEfgaAqC5+pQ7uBn9sXjh6w+rnIUzRQ2+sYBN6xlsVbgwyLI9P17
1dnb1H0+ALG2oSbqwJIJMjgSkFUAk5xHe86hHo0cW/Cmvw==
`protect end_protected
