-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iMFEC+85kjYM4QGt+GmLgWYjdZF/0JHRvtUjBXqVfh2EwoDOXcwEvN66UjkFQRYIof8DBUn74fh+
F+L8CDfZOnrTU5gLGvqKg1VWS1Lge87k28t6dpaeRkdReBjXc8iGSmofUepCjDHg/0aswwWb2G4z
XF7HixETm1BOXtfI+De8j/sYO1E1Ko0PstsqokAVbmsoAvUnNT13ExUP+10aloX1ipNa9xNcA5vc
Jn8FZV/RHoK2q1hmybyq0ftEtYeCbnuyi4rPRoeBOvfWAmW77GvCs1bsB09kJ6vHjh6gmcpqWmcR
O906MzCR+640iNA2mxjaQ9c9HuC5LzsdO3BxXw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 42000)
`protect data_block
/RvXAmTvda5DfH9rhs/yBVgM1tAd3rENbGpPhUlFawf3zIjwzqICsXEKk8HzXnD+R3Bm4yal2lgj
pY1IYLuMooxcvPBQX28mrR/P8uqEktEL9zRBSGsl5TyZMvNn4YOJ7o2Kq7XxflHEnP+wa+Xz1jUi
spb+1UpQ3BmSRWS7RxBv38jD2bo2xi+IA+ohxJgHT5XQqmX24hPLRhXTC7AijHBkk/fhO+rxUdBr
30/GlD33wgM4VxrOVCxnwkGFFQxLUhNBEtbu+fRWpawttMppqWD0zA3OXq3Z19I04Hxkx4WSCVc4
1kSUnmZdRLSi9UkTQAoOewJIJK4mvWyu6nnwYEsdkoaS5gJt/2/gX/K2NrY/X/8ElhdqrHIb+ghy
RWJyQWxjchoaGfVO9paCbGtF4+0jLkTcjR2pQZv06lD8RzrObg2WQbQg2jX+iyIovXdVf+mm3cPV
D24vptwo4MC7L0RuJKrwI3lfUBGgSTJwtXCHXpwoelRj8N0BmF/6hKNUfjJCeS4dhwZEDQ+7IgYq
F9AU88jOfCajd5qWZegs6b1tAlkq0LYcy9oYHbiWjuKKcmUGuxL0t6SdNi9nhOPXimNatKwXRlUr
9aE5A1iqCrhOfT3TlWqFt3RzxqOtguzFtA3Z0W5Atb7dG+/TRjpLaxegGUc/9x4ES0YT5DS/0Hsv
YHoJftbZ1LFNI3HlfkiHrgHYrWtfQYEVwlXhPD/QLEM76i8XNZzD4zZ1BcLvr2nikO6/6U/+hdIC
BnpOr1NP4mdwq1XJQLKzUHhEpRTNBGs7EQ/xS5ZbBwPMG+gp3UHhNBMVPv/OdiELOJV4ICMpG6yD
OkeF3XFtVmr7aZA5nasWTq1Gc0vUdukA4owMKMujWS4/kXpnSSQK58RKZ565GRxa4RioYEDINHgu
kOEH/IfJ3Ig86whqbHe5T3cqOVuSU8SG6PHh7NCTaJ9PcZILWioo0r01FdIF3SNZgwwQU0tMVcJI
Mdt4wYjMAbolQp/H9HSPs0BNV1/mG1lN4knbw7wEZcK3UfJk9z4xildqBR5tvYD3N5ofPAadMILW
MVnGKCp/otLQfpiyEkZ6r9ma56YUysRjEVWXGI0Q4I1YR2LNpCwlHrpI1tv9P+XbPE4ss5zrBQ6j
7qEqUGaeHxhGXzQuDir5LjVYC8/eEChAcu9zj+tNUnIJe8mOhLnZuspHXdMD7kByUOrwBlUALDkM
a/zOoksT78tmmVn+I5SfHLvsIXfvAhs53uRNLaP4xFv/ZJswSTapppI9bcPDGBkHkdGuiHmjaD3U
SW5ijl4nCaqgUomGOzpF6cs6a82aKwyLIeXpzbUhlQAuAXlONZmUGzHDy7ws7bXMhvDsJjWJYtmw
c7CdXPMP/PIiq6Czeva4G913/8a84skGNOl4IvWpkfP3zLNGgMr/nUFp9Je3f2icTiCQdV2+Rwu2
tnh4CwiaCW1xOJrjshh9KTEqEX1ZgflvVzw1KGa9IMLOVx8oVxkwoAr5DTXeXe49HV024kRENbkk
/Cnv3/kzQXIH8bMbf0wHhOwJrrxpykZdp6x8ap3bqm8bRVSUjTqejzuhPYpebtYWwkowBEH48NQ+
I19X3kZ35TahyiBY25xLFbYs4GrVptibhF38VPxXtuZWEITpMIZfDqBKG99wBfHXnhI5SWJ+7bAq
Zg9apw+abHZqMWlH/Qg+7EylOGW+b5mSy1QkCEqSno97qLB2BFFfL1x15GBGwqaC+5TaHUQc466u
CcYqyr6X8Hdugis8QF/v50PpgHVFBfQzfYZS3fHgZhyy50CLBdVrhgwGyrFASClSuyq1boyCrEY/
R3MWJ5pYvPFMSLfVRKNB8y/xJMht+6oicASpYrY1XVNeDkhDb3zeZvGib137mOl6KYACh7Hfx7pQ
T6dUacgsT2jQOVbkV4zmkPXfQH4X+nhMEZJkQJBAzzr1PDytf62d6KozGIiSoC6zAnbwZju7kSQg
/F0hDjUPBr5avxhLAekm7W+57JJBlrtd7XMPPoKg4kmwYG8xwGUl2VjfYzEUhpQxMG1chJNwhrvI
oR845/8VcuIv63NPgFcz/j8olNtnCNnDlkSqwJbrSoZjEhbt5qqTgZMufzt/I+GPxxSc1Nox275B
wJje6p2VDXPkqCcaEFX9mi2ngOWnJ66Q2l6pZKuNn9P5jorV+U8KBTN8qN/N/xkY320Dia9yeEeJ
7LpuFVvWtxg3Vz/t7b1AbtdmQWB6C9ap7Nea52j4SUREqZKF2T0/26siXwDOfExBviDm3NgcFP0T
QFhluGPn57KIv8uGXFv5Xx+kUSrzFbY2O8oMUvmAD2FTJHBFNNzaU8KXOpWeK+1rNSUuqJnhaT8f
KCDCFU6J6b991h2omyG6+D/Uy5e9jLG2wt2eVdwt2OjhUlgntVyrsuHWzpeGX0lInGjWrMsGt3mI
Hl8ubimjGlYkOnB9pnyp4tapIQoOerQK34vUSpJ6FgzVJ9+lfFnmGJuCdvLs+/WT6EBfvXN8jUzz
Bpl0ppLZbRafJJxxviBvDdjRzSTX0+FUfFaeVGG/UxbUxd5HSqLS/J9a19PbveW8AogTMATXPv0f
EX37wInt+s9bulbn0wYmA/CLLA0mKEtgRzuSzJUDDH1xIeebuwSrkdGCUxsIFR+6/mW5uBRrK52Y
/Bm56Xhs27GKdaiXweg447SScEnZXumTM1v25HXUWlixZV8a/2AIgpPlIyvzd6hvyF0cHUsnR9vh
soAdQtyHOhTahN8ujc+XeB7IiSYeZaXTuMOqMin07ouGhLLMGuy69F9/8yK+uspuqSqZYJ1glYH4
4o2tR1pRAqYl6WGCq/ACzzlWbaa7QPXzYy2BL0LXpMOvUnbUA4toxUSCwE5fWB0UXnDElWscn/3B
Z3/i+WEXM9e42CwJclf0WWIw7pTtv3wSltUPDukzusz0zakJkPbG0ruL3CGSrj0SxPEW6JQCK+ci
YRuKzFb+jtkTwlDJf4x8hfwAoaOGqWCIeIgxgO/Q0prXCuaWx+SzbUQVSCSnRSciEjGAMgXgSzuN
v6WvgwkzduyZcn+ho6RLxr6f19QZ8tfMhr+Pwa+ejtZwm0q2tyXu6i3fXZtF+gBezxOKyQkAi+8+
TZvSKx+IUiu+zPtNEbWWz0wMtenkOhjI/u8/SvJwYywcP8t0U8e3KPf0XCWMMkId6UFG6ngx2Lwq
PoLpwagMt2AOsQlBjWdmb+PhFPgJPb1ttfeWliZmcd7u4cQNId5nxN1YFi7ixuh346jVq4g9W2ov
f254QiEeUMemFPA7YNC4wdPQHYw//KDOLizurY07YG+TsHvm9Vc8ubZaAkkjsX28diEZrGoaI4My
q4U8HRzHDxNvsDGy0dsl5c3c37JXmVaeK4FxzPXwK6EbvDA4ecYxmvtRo8RbJkEJnLzZuEvkamBZ
dx9mtThgEWzfno+dMZVh87Udk2HJCNGOOwwoZkLAguR7D7gsE9LDGt3I0WjWoAgaVYkTYkwFitF3
oAxwDC6H227fl1UEMhAjbXaWkxXtq3ot9qv9xBCsn4co1iuWV4iTOw/rhVmGmnNyNofudOZJ3F5I
9GZF/DjozsxysxPM6fX7MtS9eVpp6+ihehx83Q3CBpYUb1TZ6wIhRh99KMto8pJLMmIMw0iVSv7C
fwN9yLZ1uTrN4DKTG9pn7qCtaDrnST0tbFuk3/6UQFndvLhr0qNGB+k26v5bO1/HMv19//3oyIch
Dbmwn/Y0hVb6NZCVPyI9JwOY4JhYQgtZniEYqopKbBxjZKUDlx0c3zppxav5mD0+MBTsBQr6UC6+
e6cSNYHxGEaFkwe9AzEF3bsnhxMTfznoDiXTHHlULlbVcqePoihcgME6PGYrcoFGPSmDnT1mJ+7Y
+pueOh8sl7YdZPDv22RrpaqDhRBYgE8RSwAIWj+EL7jrK7HSkKuPXCFLG010fJSpiGGl6mKi1ldc
cH0w7tpRDNvE0vUetPi/l0eEj/ZDIRm0WAuYuFRoZEpWuBu2ft1BsBDvlcu536DERHk2hGHG3f9a
90TpC6KMKKUt3ytiu3QwsNHp9d6LPgXxXP+Ciq6vQWH6hdTGQLsTBI6L7ngQIQemH8kHeoLkzyBY
2ZSlkuv3VTaWWXGl+1RSoKstWkaK/BBDL0apLTio1CSdYYhOAK3n4zfYF9gqt5Wp/KAPTyEoe9Oo
HqOmjP4+xFAffG0EaT8jzs0Kt88Jp4w/++NwB+DiPxZxD/YM34eC56vDPRzC9Kp1e/J3on4RpVen
Vj3/oToD+PdJHgSnc/bcYy+QokPy9vTytqidjS5TS8kugeWHKrldeZTCBSWdHb9VA5jtOvUZntBs
ucft0LPEaNrnSQc4noqfbSBDhooY598tqiFQeQI9amJnhJHW7hDGyJgRUYuCzeNhElMmxPDA1X2E
/C2SK0X5v9RbMicoDOOEMl0su9Y1wbOZS8zVO+kTwrgRd87wmb+cP/JStAQK2zvE96Z27DPn8Blc
3XwTu6LSxOqmOj97wpe4Cdvf1RCv0itSzE0wtiyZFyOOKJoh/SYvzgMMTvWWr3oXr/qvuI9k4Pbw
cIcRGS/QXKSCWSInuA+eygSSJ3r2rAB833gfVUzVKcMCCEo8/Akaouald5hwIpGDhePy/Th2IUqm
dT77nDBqC9pJK1oMry5ivWshbqeiUyKw2FZTSHq4QSY5Ny/TP+skDTaJ8FEiU7i7zbhqoamAAGDr
mW7cUBePgDeX6UYF7Zuz6ekVlNmsIL6j9OT2QGITIog3lAXljMCxndJ5VbdSG7cXSkLHGIXUN+0h
+Un6m9Cd0x3cOpb/UxmuGzSDQTexli24NwLMlHKpPpzcPzxO06/isDGm3vFC2UZIA6OFqAeCC2Jn
y0B5Vtwcse6d4oU0WP2vZhyIVQ0WoXEgD6H9YWpcT7zhjoUYYzu3TQOEdIxBpMYOXpXj9uyBgv2K
JUKLD8f/57oBcCrfJQBu8JMrL34+Wcs7hCixMnfUnqlY+CEPGhzQxjXlDuo1UVZfa7WpZVN/IiF7
80eDchu0Vwu2cLPKlfNtTljZkQsCPR2DWUYnR3l8VaU+G+1tD7ZRKmNykFXHmbLJIvx0M3n50k+U
Ww9nyCp/647ztm9FfDf9blRuM6ItJxz7QGRHiXU0DtFxwyJ+PFPITZGKlb4waVsO+kHqsUifTzJr
idj6ds0PwRjYpL5Jc3kKx53XoJk7ob77AWDQxYkHHRRHSTdPq8R7Ui3tnm/HzkVbPKGmdmRsu4pz
35xZcLwuQR3nyCKMTbDPtVzGZaLC1gMmN8Xt4ylH9PG8zbcx3+RjOn2lYjxmgRLDhVB7bShkMhMA
ztZgCRKByFaFsE/DsCVjQhVny/QzvlbjyoGTETiAZ03dY70fHhqahh71r4JzNXUcduvz55CzdQxA
m75deQW/WSCS6XzEdXJ21oq9ibSoxXUTh6ABchc1l5gRkZxaNzPTly9fo1FVh/NAce2rDStoa1D0
oNthPff1wZSC+A18TJcirzoUQmvs5gFB2qWFNZztJSEow8kIAEa9dG404+Eoen+pFE642HTqEirx
ILx/L+rBPzf50Tvke98/nzlh8unNPim5bkRp2OxuCOm5yzcXt5yRrxpPWQZ81GmUbOxRVppL+4Ck
AC8KWCjnEvzF5//sKQ1v25HAZgcr4x1AD57PrUznnzkw4Uo62dHwKApdHoCzkQCSTa3hTQa/o2DB
Ol1r1jXwt1W1G5VrMs458NGrrsW80pXjhG9ouWWzs1TUdRQ1Polv5wF3w5zhd8Nm9SPvrx+9MBBJ
a8pz+6IpufQ/8199Oz17DYJYx6rC2gVok6b8NpB5MZPW4E8oDJHTaD5P8BagIexIwYw5HqmczmvG
xj60QwvnpAPwPw2jBaMuzQZ0HTDaTpt8eCx9GtMYeQOZEM+qgxo9YjkCy9b/e28HPhGVo73jeiHw
tUizM1KA8yKaMzJFQcr+yjcGyfydrGVpHN/ByV1cqvvZcWVMWUKFMSxrpiBp7ZvR1X1uNtRmR+vG
uTpX07JGaqKAscmSo/WgBywFyGBxHvK6sugNxjb3a0TLO4wHtqYjNU14wf2q8pEijZh9MXG/uAsb
P+Iq2n5xOPQ2NgYSlbt1GiPmo4A8q1b36CUwg9MLgDSIh/tGK35UGUUp4p7+cAiaiEfoupJGWIFF
E+XQGY5o3bXMRWDnn1b2/umSbwlFxMi+hW2TK9bT7P0cRwrguU4Mxtsr27TpEBC9Kc+Pjhqmf68y
c+X+cSiWHP82LKEJnA7RRkSOdzkwl2dYowSQX71J8+XoBCNqRoJjZNb412AQIfPlB216xAOZASLs
8nyyF6OZLoE44IgDk2xkGXux5Q/7g5xh3iGLc7R5qgYP2UIjG/q5v0GuU/15qY93qik62FLf+0im
mmBJ4EsMjkAmT+ibft3+VrOELmsBFmhX9Vt3hilwX96O/RYe2Dh786Gm05euQ8OH5aI35XlNEtpl
eHY/nKvgys3idd2oofRBSLCeLQnPM++MfqxZeymgNqxnyzPoXse3hFBIAu7nFHnlRApVhVA0tCjF
nVlP1xAoZMyDhcczH6TSBLv+8itRx2jAbt8I8QZQMXKWx8ZorWwaWxP7AtZRt7XJ1xKu8IFmRsSK
eEWTgOC8iC6kLbV78J2KwqWFPXdAGTgpqPMq++DA91A7GkDwFkPJHYKdJmCLht75mGD1M1hzOmtY
FozaiDdTk0af7lkGC6uyOQo5QGUyEoc5XbleErUzavUeR5PO6Se2OIp11eHwKh1aZ67wB6RhKW4W
Wby3g/9Nnzv6RUq3Klm2bnRPXfmbWrf9B0nLfHf5LR021THXuCFGVuSpLlWkF9dTZ/I+dyKDpkfR
kcSKweWQyBqd/FVTWW03g2eoLiGWFMu4QKna0E7EfAC/FfCcNOUS0FMxIDlT0iA+CVImdYmJxEAm
FVrKUfSM/mK1E6y7xfZhbRcQZ/OOXeF3A9IO5NwwX82Q47W+Lq3VkirKqUyjLf2/s2H+YMxOBmT4
4F3L1EwD7a9fNk3nlX3yHaVmkN0cRbPJGg2iNPpiDelaPrUHwZDcBmG7Hd3pcEz77p2KZmHN0W5A
OpywSgWGC+KNZPlBmLO1J233ODotOdfDyMZiaeftCOP7CmRe5sRrWj7Fuq+Ub3bJ0qGXQekqzg4D
ugBERfYVPCw9fE/orVrqNo6IHYCkMAYm6FD1jJj74KMFMipWSxUiYkr1PUcNtDCq3vsKnNLUD+xA
l9X+YSDj/meZ7R34T/k07OP6dCgP04HmLWWUrcWd336GW5ajh/07vRAYgfKAaDxFBWIVi+Ee/urH
edwk4aChnymhicLHwfklak3n1S0A4DQD5da9TNDgUZJTR0UZY1RJ37oYsA4js7B0vjwky9/t3AKh
X2Av21liCiQtylMjCqF3HjX5HMu+K5NFfkCfLlycsCOsv++61dhJrit/QeujtbFTfyM0r2OYsUcV
Tr/FNET8ZofMPZKJs15352ug6hpPjaIK3dA9HOChiHiSQ6uvvCgawdY7/f5gIxhW9pNmc96ieEd2
6MyfckuHmDhWKoRboj3hIAhN1S2UoyAD/ooq2GmEikOEMJ8l5oycAmDmWgI7ktvwOMZRClpIOaUG
HmKElnalOa2pO3d03A0vtjTwZlPLX3qi1cEttYA+gPlfxgMECPZN3PZFDTIA2KdVH2bbnKfrY2AK
0m+UxUxdCk0XqKScYimU9rcXcMyHI+Wqbu0Zg2wqIKsLH5EOctuNwuO+zbr4cGOEuwR4LbLuWNcD
+cDQV/qjNj+GwW6LBhhiYQUALxGVRkELlNVsHa7iKii9l0DVncodTSIT+xH+PsnzZKutdX/ei9fF
r3q66W3uSppmQgtngD+fgVL8FpT86uF+zeQFslI7E+Q87LKYbK34/gFlBZ/5+06EhDHWl3w0JWuA
d5mWXDpMhDbv7jcldopB7qwRzEJh+XcQI9yLPMKOAPGz5ugNUV5Ep1eBj2w1XCcbLWoYIUy5FGDk
88qhrIWfaGpEu3zTeqs7aTDzXudcHOtBZgMsbVbfXR3XnI4UqOISS8c8mHs9pJBbf6xhyNBfAIZF
9zu0mLPfBenAWf/32gmDrcWB1vaWE8ZUw93AxI705decbNfSS3opatPfw0pPUQEgRJUz9rrlXsLJ
XABLaBfvLxZZeTQQHNQxfPLqdTfDi7hT+9DKebaaJXzUyXGtRSvek3pA2ygPPpjDMYqza11hFi3p
Axuq8rBcWTE/V9CPi6jOazuw6+erNlObcpSZBTASRk6wFEhK4mVmTHQzI/9paLjMUPw7WsU91tuK
udsYFMSpSAjXyjVToxHg2kVSyAU3lXuycdXsh2N7mdmW6GnT/oZ3/y438eY2IAysiRwF2WNPDXS5
svblY8KYb+OJ1ETRrauOBiqxAFOONTjPyRibMzZWTHzAIcaIpsZArRGKHmK4B3daWZ7bKw/N7jW5
O7XTB/kZinOXPAJZsUdUay2/OxIgtvNnLNfUQNzEAxkxpdLd7z840D51lHknn203GfK5adCOpfd8
uAvfq7BDLzKd+Bh4kfKEEyz0yHeu29ZF/yM+7vQxzRNr4A5JD3EX7szO2Q1ImfzPPP1Vex/8WxQs
HHO1ocfITIJS6tghXUARsDLldVc5F5853UGArNClyijfT+ZabLDsU5ZCrLHMpM1y1heKJW3P/r5v
Sb7Nza4AKbmPOUDwlzJRo9XCdWgfEnR2UV6OnQS5XJGszOpYr0IuSVvzCKgJ96Vj4d+an2DfsuR9
9EmTThCkQs/zOKlb/zN00YLv7Pj/JWCIQ1Q4A5Sd9rPW8tq/k+PrKtG4A0wCTU3eAB3PMVa7rSlO
T6zWL6qcumCOWG0LcUPrtBy80D/0zggvQbTi6M8lRfliMrWqwBDvIw0rmNnqMkmant/sl903OvlK
654lMhCMQ/HH4NQpDYL2YnPBu0fI7EGn0qkyOJ7L3geO4zAxJ0GbbRSgpan6DpEkvsrFDrzxi/9W
xilWQqR8Kvv91XbUdO5i/vkiGR7BA7Y1IicL7Hnaql1oW7FJMwCvOjiTI87EEpFmFaYNE8Np8Uvg
Q7NNsZiZAbybu9Va0k/UVsY3RZZpv+777kESFDmsOndoVn0y0JUD3C87xdl6u9y7E2CitfiUN4hR
LGJXerdaiUjlz5ld+nsmaL0iphHhcCBCw65K+0+0aaJ+6CiPhn+Gjowxwvna5pn+DwMX1PsN8ayY
xKfeVXqmvA44ylnkDjYoDgiaBbwiXyrD9EbzNzz/51GijDokR3gbJjZwRDPX53GQppNKOzNThPbC
EoufLdDxaLZDwla8xa1UNF/IpL7WFDkAm1GqPyoaNBsOgVM/hjKXUDx/dp690BJ8aIHB5A0WG47l
oYM8gwYZJYC+HvfX9syR3ABLf08aQmLfuA7Z7qDoj7yyyoJEoz8+4VZh3EpxJLjsTV36tQPnsE11
JuU/le1i2Ps/611NrVzhJDQEyrVQS+YfKl1dEWkZyPLez6WN1/844iLR4ccV41OTiAtGS9f0ry7m
6PzpUz8gUipxTpfO/jMbYySBL6VZZTfxcvqdolrsGtStSrfjceD4gk2sCxx5w9p3+E63KJ/3j7UN
ck+RJe6Z9Rz4ltr8Ywp+rYgQUavxzvLBTodOGnd4ajld44aq380WIc+BDGlWZVoVvQRqL6Q6bRtY
wctNUzvwDBmSMLz3D14YwZh8ybbMN0r92kl0N5jLAuxu/3W13hJ3r7Zxz7BoZrSxkVzo7iG1dIF8
Qji1v9YFyLfbB20cMbM4X/AVAzpEIwmc1Fjb+17FX6nvhyT0WRFvRxuMUPSY4QRAfWRhoQT5MPQR
27k4RVRGKalEh2XjVt9PUgQSz8FAHJlcZYV6lUDR8+uYV9/5U/RmjowiGVaAyPoNThVzr/0g+aHj
n0o6TZ9YrkEOB0QhQQZEvvq7k1YIvMo5hJ6w1g6DwevaJdm/P3UnU4YRMZTVNcX7C1wbUzsXVqHz
30fZbSa7KnSv4cP8Kde5cOsKutIqh1z8cdOlncgT3w1z3uYDtq3nOOGWMHfJPaCWVsPBMthVeKZ0
7JYsUynabIH1jYYMzaa4+EClRgWWaedrTlTvjYkF0mMWwgCwi30g0OtXl2343kGigzg/2qclH48a
tXJUncUkNUk156pE0m0uq8GLse4QPHZtqDftAjAefH1iChRVOs0UKbpnGOqGnnc2BigOj8d+tAUL
fMzCjOeg+r6mTcfM4qWIg10JS/+9EvmAZw30IE017n/3lLnH+4Fdsm6hGXBTb4kybj5DH/llJfVJ
7oRSLIV/I0HXVFlgPnBHhUzlXptOEmdChBnx8DKvVEwECLnLGXCGFpwSsM/r6ptkSz/Qdd5OScOV
N/LjdLQDfQPXSTyB9LAsVH+ZTOJ6PvuqRlSAY6wnW1xVKTQRqf/2HRz0fvNCvJp/whBnzFhstyBE
OZGdkEPnfnWxqyNW4/s/V6tNTr7ADW0gb8cqb5P4D7xPk6XU4sysppXQ9fbsiIhJmZN5NIcr7Ypr
a34+P4P0BK6Q0M63hn8sWiY1fN3eeksG+9a5qPjRpMn1yom0lfw1dxXHw1ovSP6puMlBLgquatQn
zaidi4HFHTAOMusaFMQJsuIQPnfuwmXazTSA/8hMUzCE3AvJoI0GJSGNYMG7kBayeH6kz8oQgN1O
sl3lSa8w4b1/zwbn1ohvIoRy8PajdHRh1k2xLUqanVXDPwsrYuMdzVQWc5Q9YDRQbTtVtyk1tenZ
Cug300is/d5ZaieiUm8hGu6sZ4qRcxxbrlFf6ogvpe0MU/+GjlRRgzDGcnRUpNTTKVHbSKs2WoWN
s91LBl87c9U69SAjvYYxWtQCQTy7rUGD5czEy1UP7gFVc7PO7scScVzt/BnRDuFXflOvfO5gelVq
EOc/ezURZY7aZMKKMaah98+rdoC3cWE2pxjpf5G6b35N0tebLrv7lKayPxEDG4vfC4RA7FyHs2en
vGR7XLMNPEjS6JiyvrWcSNaftVXwqMNKBLg/bGWrqYADUhW7a5onefdptbnTJe/ceyIDhL3qhxDL
g5tNfj9/cEAmw5vl0Xabjnm+w0A3AgJxjmWX2MUjBbR2xqc6TVU8aPD1zwlqSMt8bpo5GfYcCxYl
5AGDBGILsXNqYz1MA1+gBJHr6M0mdfcOdtgqFifTUBPSei6sHM3AX0W7vD+rxntrS2X7IQhYYLPv
6meAMd8uZ4OL7L/K/uqr8eZwXNDSrcSOX9zH02f5LRlJke4OG2g4Lt1OV93ETNh466XCBs/F8pu7
bNpw+t5yg4YHNyHLBiGRg87Vp0tlCq48jCEPgufn5fbRF/oci037JmxbgeMiXl5jMmyAmqm+bulW
fYychvYQOO9qFyZdZa215JEalbKCffam2tlyBX0fJiwX24L35vtrmQZLNdXJkDtSaXT3BCW3xJv9
/bdykHb6tUb/v+2phNj7ulXLD10xinLjWzuQ/OMgIvl49DWdI2Pv/Na+P8SpBM3i6GQAPd0pVk9I
iQnsDbi8HRoqUQjbukLNnNH/GcyjOFKGXPNtxAXXYUZbVf/6g+vuels3A/utl7/GPZrANCS7Miw2
TJ+F4cPuJeiLU5lWokYQwS1sqlsxut8r/NKJHm40Y4kWqm0Hn/Rwb742PZ5BgYnclBAaBUMxha/3
Lic7xOztX+PPRLd3xJRUNiwR79Xpu8Pu72gDIAClvmZo9MoVn0PrHlHYHou2/f+WyhYjENIytiNI
8PyI2f8WT6lN1LrVc9a715V01+3b68Xzx2m0hnpAwCb+XscnyfC53onBnmvCpq0YIaJVW0xFn+yc
OvYSFaqwBOwSUT0x026rQ/IUTnkdaUHRkPjDVVzQb9137kJaOxzql0jKXl5R0F1kmLSfp05VUhW7
lD++dHGdQUQ8A8bcFpgI96a+tMhffV7GM7vx7UGs+daLzT9EiJfcogoT2CaQR7x6+5QHE9/6/G8J
o769QBsbNLMpmZvW2TZSeJagg483C7C1mRnbiPzLr3USSwDvhfARXX03hiUEqFNuQZewlIygdzBY
EbIm37xyWedGIWozC+CH6AxuYFpDYETfdkNekh4YMr6eR6q+vbBlTGh+9fAR/V3mkEgz+5HTmTLQ
XM5+BHbI7rFtMHzZMoxF+htnrENMBCADo0nWnM1xaq3h8UbfjZO1TZiaMbcYMi30IzW/4tz6WxQq
V+RclLAqSWqMJAR0u0rbmlQUn2jtM/jidR54jdTmu9BRpvT6VWieHDBA+cUqMMkBD3mqND+vDa11
KFW9cFt29tPUw5CzyetTxcMn5xyP0+gvuvewB7HIpXp3Pmpc6faA/CmxK6RpADeLNfrkr6zcf4Ol
z+GzkgW7QF3BT6o+5voeUuYCgCJb9cUV6HN8x384xteN73iNqS5p+qnJhsk26uJ+CWoJdh+8ULkM
cgg4nDPcwDTP3FZXoR8aI/zDbW8Dzbh/nTQEm0WQxjCPYK5wbzdlPnHbO+hCjkK60+G9iO8BnxjC
tcKOr+GOnRmlUk92cPTX9vmgrQwHCx3A3cVyyBUCWqMgDy7TCvG4tT8QiQeIQ0yqz+i/lfBb6oGl
fV9wAKalIu929Pczf3WM80CFYeaOdV7qCiGjGdCGmuQ1zwC/IBYwdE2oWKQz4atH2h39XOt2ww9W
tCafWkZanUlZnaCtUjTAmDhSI3XHB1phH3sL9KCzbA5T76PMBJUKkMmgmPLi7rHqI+HsrPKaWMNP
BKtoIuc6/0ll1WuLdytNyFseqWdSPxx6fNp7mQHZrmwd49yL2bsCUuij0yLdw/HnLdGa2xaVwM/0
w3p5UbK/wYp1SvemcgokcU+ixIG5fJ6mytga1B0ci0fAV48SYeHOMiPoLOKwJxk+/Kmry4u8ohuF
PMWlAIOkCk1T7Ef5takqjfI/9bftw+uAot7T2CuI16LWRi0odj0lLbnbor1oCnPrSnma+Ik2A4+3
ElgqHDLT5RDGWRg6p9AG1naqya6TrbrH5NeBRgaLfCocVOAkCWFmDrvcwsfFSGWjEBzLjVIkk9Rl
0GVULMQOxKTWd6nm0YxqwZhz38u8ysZ/LM7H3PSV42sPQ1ac7Dbu196q5NLsFKWD1/YaJqUNKw44
sJrhu1XVi3GGSa5unY0rzb9l4aZU3OKPco+eMM7DJNRT+lRipYCPDmtnwmuiRvm40V6GuTvES0hD
jtYqGbS37l6oh8TPvaTUzpMdyxMOQgseh1EZVe4D72f6O616h3whchjAJGErPUQAPhrEnkXe9DB0
imv0CkCOGGwInGxP787DFtSuDN1JCmx7GSeSc/aUPwyXx0xktcaRyuh/rFEqSI6r+q0QuDhKe5Tm
Q1Vs5HSV0cNxLjNNymZhjSjxhDfaNCCbBLwOHsv7jxAFfr9psOUGzHYvkkJVcJD0g6zUlBJxOSFp
Gyhjg2gye4DTTSi5VlnVFDNKqVIIo5l5wMoBgW8B2vPS1Lc/cxtlleEV6Y+BHTrTscQt+mecbrl/
lSINKGUxiKR2/LbQ497fbwJLZ8+/6ImWCPJCsoRe0wEgL9CtQOcdjVtZh/7sf2fbAqCT6n9Tvt9U
8ijV7l1tPeXJmeqnuGOrKWfHaw2lqTOxw2GKWHcsc4BFp5OPM+HJm228uXw7Sl6KjPiwsX9fnJ6w
igOkvfoEDYz7Id5WqRNCCHaa6bCHWZsBzP6RC7Ev5HsVrnnyTYmxORwsS8QPeT76rUStrihcboAl
tLEbMV6nXT27USSfDS/Xvqirm6hFlrDgDFw1084zixiQwI/FhWvsSxaz2QPoPQ03jGsAJM5hEut3
n4/VScFJu5rMzsBcM9l1NbEDU4iowxFJp0hunpyZuP82xhk8jDzdj0jaak+Mc83Bvhh+d/vVeNVH
lD0U5WyDQ+Z5iectG/YY3YcvxE6N7nQPajbOOzUiESq6AUI2+ugExlkAyV/VqT1hbYMwiOKqJ+d9
XR9+8Y597Ej0xZ6zprvtsNJao1E8OeuKCqNDRmAeoEmh+JnK1z44BlzGMrPtlpQHbB3iISSTgf/c
2Btrb76BD+gD0cs3DJZ2pc7CUz38yHkl0sANGR0X0vJagETOSpFXqutQdxLHKeRqH8iWerBed3YT
wkCUBh1dsmWBQZLMIodr2sEV7EOJGeqajH0EUhCjyldB3cFe3yBFkI02FzB0FgQPT1KYC1lV04pI
JAtDiZn2kX/x1p1moMsgf9zyWM7A8I22/DqtyCm+sMWEcngQCqLrTE3ate1xgeevAD2vVWdJi6sX
xxPaY2Rjq9HTKUTPMDGyvEM0QYvJqGcGlsx7OUl00IGOdcR9DV33cIxWCCyVO9QALVZPyh6C+eDl
mdLtIJI16NcC4mBP9mrrKDL66I38hrQOpqTA0yCn14yX0UhAAILx5gcJNEz6dKG11Z7QDY28ur3K
/a2XMfNxdLuN73/qduo8kXV2KxSli92JiddossCCJ2sGJegMBiYGm1Dzm1a7ve3Wh1/AqHxyjaFj
o78n/MQyMRH6ioeyY75p6T/JZM/4fW+wK9DE5miGQWl9fmr/0VWwJ/x5IZIa6fsilI9CPndHmqHy
Xw2vBE6AzstHrPOhaFfGkn7i/io4EQwySfmERkcZQTPVWriCW09q+EwGPUDKJpJaN88M9YjEiwa/
kluusGgokOAyR22WIekAQUa6VsTCJip5spRqVKeK90JzvumqysabaR0WxhlU53RMIvK0FH28XFxq
qrXORzX6yNFg+yT21qJbsdU+T0LdrI0/5UBu3IKeP9qakUREip3is8HMWcuSaF4vK5wRbDeVYwlB
2gIyRrBcYYMBkgiQiLWXlGUVQxRWHq55fAg32x6grr00LsZwOKpJzKL0jNpvTfdB9PCdT3xqijGA
Wqa7yIGhXxENxAmMzQZW5wJVdUM/1svRshnp+Q8rKWVfAd/mN/iPTa8hYP01Fb5ANSrsTNKpfIUZ
mnXKxBE5yvcRBdfOH1qTWaHuAUFTSPSe9cfo0cNWOQZMv2EAwc4Rc5SQ+d/bBa+Nno18rF2rnhC8
z2qBElzA73YlshOjw1HO5YRwXaA3IK9qtuBmczRFkoh751DpUJ6xhb6sK8si+fc1wUFQa63tB39c
N04rG8TNo8zrp9dGZ6KaVIXY+zC+yXouKO4vpEV/9P6LzHZUD/yVhTyB10+hLk6gKjDqWBOdPJHO
feAc+jHmQ7t6VjearCrXdU84obemONVAr1nb+62kBHRt6kpMx+A/OSbgcId2auw6hYrhdAYGTu6K
5fut6jdW1p98KY0B/LBYo15mqzz5brp/GInG6uofPlDZf7XsFT5I3S9yqMpj5ce/in+AGWjEPCqh
2dkzEtFwyKacOQUgl+3y9M1DoSxiWUBoN6YgN8AIL79nKC5LHbFOQHAkY+zs0AdkO916QFk46cYT
lEaofXD3AyTv71tvNIaF6EzL59fJDpWpQDbX1r06wCis1kyw4vtKfuR5aUEUWSb1WtilHkf2RbeB
bylEToUE5JbVERYfOxmIi7P6polnJcO4iLnb8OntwCsx6ih74RjpSyO8stBOqA71jLYW6cybj2HO
SvN90t3AkI3BMatn4x+ZoDVAHDfqIV4EGqQsClEAoC3T8pIZmIcNI8hPtHg2yrke2S7LHXK++LLc
s9k3x/VvBLDDE/uKTuH1w/NjWKA5Krio3le3kqozrSYnyOT7o64PkeBIpxvCtUX0+Xo9X9035sm8
W96HyzfLEEjUz+0XhVvNlcMWsCdsH7n3x0/rlZcPtwyFM50EXqc6JUetzM1p2+PlwEz2wUSNRJ3V
6345MnU7Qmtm+UR0+2IlI1P5h9NBYY8g+EmhRNXErzhM62f5s4Vyrqh1gl+4Z00vrdtA9NOCffWK
PYERt5BsLhTRQ5zhGR3azcWc3UM5Kfaj5ADDXH4RuIJMDXBJpufdF8e3Iup0BumNIjRqIN/G4RHV
xORgQ1E4vsoKNc/AvkK8u/7qiBJkMWhN2YQQ5i4VOmBmt2OE+SZ8Gsst4mAT3+096DwXOIB9KnZV
71nmlWA6DPIyTkh31WLSAoYS6qYPUzaA99ABlvqSfYR9KaOnTm+aTu0IUA4hpOwX0JptXV6YOuJr
d9qjkN10tLKstHBWf5LNp445QUf72F2jlzAcmwHnq4zEWcbBasB4kr1yNfYPsD1Xhnwq8+5jcgyr
qMHTgATSzzJ3KH3Ex+rdQaQyLoWYFzt5z9yu6kXw+K/zur2dizuqk3iXqrwWHYwJVU5AP65zSMMz
xjeKZ/vqgLk2hozBnW4a2g8RAtv0VddUylilEtDG5pmfPfff/5mlN0PvX+u5S5r3svJzJljeflRe
3WfVS5gV0sU8l4zh1gAlneGQzz3NweYcsNeay+xNsI10hGKFcgqLNlssc48kkLucN3L40o1300qz
V6OTX5sCTtFwaX9cmQE8MnqdUfokIufGMHwGz8+YkNqplw7EZ1USprO9EeCcUlgFUGUKNgus6wlt
9CLscygS8aiCPwINRgnCMcvTqZbTeD/NXNY6XRFba/vtoyOc7ayV0WqtBu2HWsg5b74MuN6Mtthm
G/eLphNs5Vzb4P9Amqr+B6SljiM283CON60qnhFd6rfaugq6kjZNLOXaikgCOnfWadR71bchiv19
60OpaifEXn1nveErpMDDcpLzJ6URGLeUd+vJRJjjjMCk9XnfLez8PHt3/2J+EVgbQSbmhJKD86oi
PHCWcbENL1PcGwK6yZlaobfq1TEofkOXjHDdRnV960qw6MnTtZ3klZjaGIcCwEZPkpey2kVlZVaH
24QzQWuB5kjbKGQ560d82b1RYHZ5+m8rGcHG5Em9Ep0gXjJhPuhY6fdCiTA07+xd9FMyxArEZwXU
lvVD2OpjkVPacdReD4aR8ZkRmwBOgGJU/2HBVP8UtSqmclLhMr1G/+ZPzlSbQZKYjoCfayup3391
4Kh5cAOb6SYtOICuo5URrF5LVmXhYFC1Vyo7axbWjVzR1iTKJ7pYeQ1OFm08667CO/5XKjzjPLYE
bCraBkRtucqvUb0St2jElXF9+70wwiTENAgiGJGCXyI5uThm0tyT50IQj1Duj3e3D+teR6LUjcKs
89HIUwPqdgtwHfo+j22yRh6xnHO0zKEU2pqb4In9yC4Ru/tkesjYhxl+f2xWuyI9xbKP/9NVV7OK
hzpkY3LyJFXFOwd1EdcI8cBLA1DWbMBchos95L1p476HVJhIrpBDKPqyHhyJGn+YuUmZrsKuZQgR
z6QErjg8XAOlK7ZE+kZUwk5zthgIqlrWj9WHtcuLb0Us94MCxfuZQP2qpGC+ihdDpsoI0vadz0j8
0XV6pxBFf1gj98HJCPBe2YJi4EdaWIGt7JduqYIc7DAPlDUltsZ4Z3Iqcf8i2Y3yJRZcfQpDTWLI
QPCGHLeF/XxMtBiwdezmqqyWVzqtj4UZJPQWZrq8bL8jxe7aTBTb/qoxNx7iC9I7L1a/UAN8E4pl
wtlAVAcjBD//MMGxOtcPwm9lbilFTE4l/PkkX2JtM7qhH1LXTlajR0P+CB9JhdTiIBSuAjPkJUhW
bOXJwnCwafSlzLNJpKT2sZqHyHHwsQFYHUYD3CZUGcSM/mX+wHzFX10YQogBQaSKhwhup5CugSPG
sgfwcUqCtL78q7m5F9IC23Gg3qkeNU2Cy4Nlex+QR+N738hK9NAMeuthYZMtafevKGtI5k3MwjO0
EE9feSU1EwNbcWYc/wP4ZP80x8ETOjmSvFWX6UaYPsbU7/hcQYcmBDXQA0EI4VVGnNSJyFRCvrzy
lyCNIdCmDAeoBCekUCRvFPhDGWNFHZ1phgF0+P08ILfx7tO1ScgieT8qPhvdF2j4yKy8M7evALAZ
b+1M1ykLnVS/3Xi4EuWJWgqCnDT8ATUTk8qbgY0i61QiOretOOnQbSR+ig52ODuiN9rN6TDXpQFZ
ffDyxpPLNDXkQpGGOhjez/S8IcYCIMqL3nte+CmGz67P3B8LuNCCLIpgMHfCR2UeCDB3gW8VI/tf
KQ02DzG0dLJYxUWcwnHaQ3FL+J3Pd9tBcTOhzWlsJt1LdB6jyQug+F0YCXhBdHWBgV/SBCSUgXBN
B62SPlaHBLTEC0Qy0KNc7mQtjjJFTDLZ/Xk9mh/vlKyeFkb/QjX1rkB7SLw45t3x+6rwqB7g6YTX
npK9wdObGSnpN4lMpOn0sreCDQZ+A0w+795CLoNnIJXRJxEGz8vpyMUlop9MIeis+jaQMG5I6m6h
Xxzc7e7wtN+8Pay1u07l9Rqt+GjBk8kN7PF1qdC/0siJ7ECRzj6dsZZs1mDXCMAofJ1DlsjFceeT
egDABof8IRMjM6jJFgQUAupa9zwcxVvOfrQKmIU1C8RXA/5BQxMnOEVBKxUg39k/FTLRcpPqVQaz
9ttORd/slGtYQ8paOT8TLjkDdgpGnin3U94dw+E5/dk61YI1E6u2qBiAj8+GD5DwWxIZiXB2gbq7
r+cu2hXCrbv8QJ2kP2xWTael5/VWqct2HTOzat2ZrX+E1rqGJd198B0IN6u219tgOAsZ8CEKONL3
oRgVITeT5DgJuVrlapxCHM028d0A19xWiCtr6gpYRvcZFNQ6Ma+ZBFxEj/hVzFXj5nghMDhNWb0D
gAPADd9LUehdvpUfE/aacz6g76Y1WxDiNhKS1x0eyApo4QA0DU5Yi2cD05PXpdPmbV9wAiSj1/Pz
cWiax2KpFF9MU4lw7RprABk0dtlau6EGckTzk0lAu7StUmzb7Gp8JOLpjp30R8L3BkIYhxfS5u1j
i+kUktki7iDeuNI7wBhhsbcoZKCNjKWYIBMvro4Z/TVEAEZYoE0Fxl01gF1q+R5i1xeB8dYzQrTX
Sz9cnMkb0BCQ0vmWmNs3u5DKSUSDSvpEsAOQV4oxs+GnbJAOfmcNSSMaUmyf8JACCcQBSQxUJYVr
Mqr26URIvlQlRW7ycMBMw+uheHz982wn40v1aLdeFr5q8ZtL+pKimiqFbnJf5hb+60SYAI5rMGry
kpteR/mhRSLJM/8j8M22OHMVTkwpfOn+VO8K6kz8Qomxf28OtQ5BMCg2x5z1AiZG67Mohu9xIy0H
5Iztqce+npkavZLWJe1YedJBhzewVvKbzCpvhf7YmeJx8FFjiRCaxmGhJ6JjK/0z6f2hYyC8aoBF
itlsu3mBRmocrGkm3OoIfgXQ6KVkStAQdnwrIb4+b2JqyBTRqZ4gnDXGJeVLKS0lwsaJk4f6rwJQ
/2yOh31MsAIg7NSPhUF6aTn4jb2kjaWp3vPX3EZPBrJ9EwgncDdoMtgRxr17dL4bqlEo1Gbh4drs
iOfs8X6bZ8Ixn3Tov7wEYPxIV+XxwUbmBKSPW3O97ob2Fb4XhhaJeEziD1lsxRd12vXpxe7jB2fd
DcBZHJffatYdv6I7cdegS1SsDf3Z20gCS1svgwd9YihXkZ7fWwk54flUprqUYyy4fEO5XlJM6gSL
+hLFihOMcH3x9kM2JeyTIm5b+7e6L1W9VN0CnL/l9HiuMW+BZjRIloloHbDTdfqddl3+mAEDttsH
PyX0iXd1c/ZEepjSPQQvCv8bovnrnsaCwcp+RZIV0qcUJPqua0HiSmhmeyCuAOtjksgwWXJDeVvN
l1xL5RrQVN31DrqNOxIglgrOLEer3fQ7Q3RsdTQqm59VF4fKzlUFD95Z6T6f1QqILlnVz1BZSXkv
erxq8wYoPJj9ZIDNQ7DZcK0Sqo76TRYcM8U3WM+WOvIxJ+tOyXNFRby5JsumFaEd7ltEI0skSrIn
PFTIjL68hXI201i9p2PdeOxN0mTgVz+YDOqC4/pmuegZmhsxHC84dXFfdu1fNglhR5TBcxB2Ifju
RsQn+qBfe3BD5W7iijBYTiyA/ucTlomVTmhtcebv3W+s5iWatJEGqGj81Gp85kPaT9uAvgBVmY5r
t7pGW8dleY6bQ9W8mrzZAO/zVGah04RT1SFBEHNiSWHFPXB5yU8Smmg+6UyLm0SKSgWoL1ES4Sbv
+Hidt4FqwMX+1Qb3kqaQp6a29poaVRw3ivz608Fq1VYVGESSaorIGrVRJ1d8adpawUzMqTQML5WU
3UTXYgMkNY3hzExlBMqn7hEJKq7qMaGwrXBn2w7KTIYkHLiQSk6DfKtBOotSukqHF1BmUSKekgdO
0d0z4t6mD749uzK/BC5kKqkCeTXRA1Av2BjJ6q8B6TjOb8swOO0BQ7N44Vx3kLWtWSwqxWiEswpE
u9bNY58nqCK62RI846uYaONOlXSaHJi3yiUi228wZSfbb5cofgf7N0xVbITQyGFxCTsnZ/0NEeh0
D55lpTU2mz/IgVHLSY1/PlRF0Md0//XfHh9uBGARhdjPm+nuwnzLEpIqYh30YCyb3E3/AAcKqI2a
VOz8AB0zfTuAZurcSinnDsn0sGS2LnMO0LtHY7FU/kyZ1NbLLGBpz4MsggzhgJzDwCDHEbfjrzia
/x5L6pogMYtWa6cQeu6zu81fHo+f2OOn51v9F5Q4/wtyJQPOjfxdrSn4iQOcMvj4R7YGr9dJqnb8
s1WskzQ+f2swG0t5CcFnp9C9AQnRp6CJsPLVu7tW1247ITBquTrnL9RR/8sUQwvy56oPY90U1T37
fCRBRFkyyTu+8IDiPiwY7xb4/u48rhASCNwCHlGeA11rnxqZiVTXpLcbPiMJZF5d0Y5Fd+Pa75vj
M9u31kzExDL19B38Q0dGK02Jdaue2SKNpBNyT+8IQ66Oah+0lZxsh7ht+t3fb8ZUe7SrDlMfP6Th
QpTT3K27X5Kb6SooL3HOC1bEdRM6LvvvydbCXxgax3EuuVrzKaZ/sQpc3ecv+GW/AyoL4U+F1Gjm
2JWAX3XzG28vNazpY6RrkcUk9waUTtk8Aa0apZ4FqYGlVcJsbUj3bPWYAWrJXNltuhRlJaDnhkBc
yAsK3daMSddQ/ZyzjzNnONMFDr74rI5ZyroueM55agioQkPY5GLs8bJWtnEN/E0hAT89JsZ5b2Qc
iSlyF3AacaTXiKjdywpOKX09yqwZYHh10OXLWq6UU2LuzEOjecMzPDxO340cPZFJwb+efZ8hurf4
9HKRHH+J+YJn3gfJXdoEFSMMWQaoc6bo2KTlsr/grDWMGz0VaBzdfN7qGQb8An2MKmla0WI+olwM
TlIJsZvUXan4THJ6UYlRKv7P7F6GXbI3833OesoB4XokakCqkfB0tQngOy9qFxAU9Aq/9nQqFlwC
fF/0RhwyI/Fl02vEYkj4TBf8eiQ5BqKMXDqZMcD/8zDj9MdKSje5KB97GHob535b0O3XHDR+EclE
I2IJnu29SvR4M6jrgXVCu6qzWjPFiFfLxKoi6osHTktGZaPhVj4gcXxhktldNszHYE35VVLRc8Nr
E9oJmEoJvqLHfnJs8oHmf+jEpQmbOdPHv2UVoRiN7YfehTdklDogPFe+9ZZDl1zpRihnvdNNaM82
ZX7HQvyRaoY0YwF6sq2f5eotZLd5Kav/NHpGhTvLYsTnBTvGSbkOk1qzv2Z40vpj59oeQFVDAPxF
1gNOYkQczxbqDfxEXwcBnFaobWaKuK4ttP5Dj/DA9j0PkTDNzrdXtlvEn1BAElqItVGXSXmDiMST
a8412qBWG3T9+Z/TwhuvF/G1R/XWRL5sz2zkXXDuJOImWAjWgZobuTHbhu+7jMvEUKF6SetN38en
a9xDl9TOXrwY6/kMIu8yiWyrWH3tbTrloEBYgb0v0pNimj+njJd1//TC1ZSrQid0G1FSU4tts4l4
OqHgZixzJezmz2JkL6BSlrSPH0jOn2GBAqhCwv9eE8PqgrxfEB8XV6VakRN/SMHRBQvj023xeHlW
SZF1v+/82yLLN3Fjb7MLz79APx6vVp7pD8kGpjK4XYqXRAF+HHVFR4gV9nDTDRSvP0X/kGe2J9XA
Q2vXRvVFHbrS/Nq6MG0UFy8TzWJ4IBCTmFb86CvEM1xeGuVdfq3L8EJb7+QNxBK4k/R8K6ZXsza5
qai9CVtFXoOWu0ejusgwMKWqzs0YLZiCqNb4cda2jddXkcbYKihyLGuZQ0dKurhC5L3h03wJu5wf
AgZdwqu1Q4BF35g1ufnERugsNrE4bw/yUFmqZdfKec8RaOSuLmN0jTy9btKA4IroKe1YHE0W9jMw
hTrkUIxpWEFUTXnz3qXXyXNr28tpfQ8B1gVIIBUTUuvOXZCa+/f1fke1N3GK4M1ieXaNRIYxeunu
srPK51UEBdwmHqhVaD+3ihseM0n/zCeSyxOwNomiyb4SsYZGTN8W+hWlRdOozbiRyqbj+8Xr1vge
BZv2nuJEiu8NEpkVmhD1kS+aJLHGAu20LBzSjfE8YW9ETpqajaSegUcE9PIh0x5IighNdjU3jrYZ
7pSIIJuOXMw4ayqUr47Iy4UuoLVAUWtLF9T7p6ZWS7J49SoflCCWrVbaGiLpSwbdt8sI2fSL7Fpl
wwUPLYOJXvmn7X3s36gNkw6hcdebXoArz81ZwkVxdjbRU/RyOyx3TR8Km7ykcTPLr+8nwz5DevVx
6sTdPyf3jtxKBomkVVnwlisoU/iDkGosdhN1XaGl/w0m1WhEhklAgSiOcRgxGAx3WfQxtL98K9Ul
IDvBDgh/8O7mUJVT6f8vLVY1lckM6emwOXxdrjKMl3oTjZ3Y2sSxHrFRz+O7QXnbF0H3P8eqNCbZ
3pxjZrApZWFWPL/ObZHhj15nV7wml7bX4dR3sP8+Jcx0TvwliE2zdT84F32+Ia7EZEVCIH172ZXu
rqwWLN2Pf8BueDw8vkrlZGHVINLtOMuyc6BbpuQ8mkTEpSgDpRdS2Ywyi9bCRjVibwKX/TYoBaGB
bPYzmJfOgW8gMTZ8O/NRfBFEnSksGMjioCdOA7JsD9mYyap3hevvVJbZQrFoiE2KC4wSAyQPGIxI
ZBLXKBwigFdfUcMV+vGwQHRfU2SrKP0071s1Ici0/8aKi/Fv18c/vtL3I3EfbCpGuP7Ke6k+aeZI
4/2+5UdOD7j21GfIO5wvqhkqI6GpLATXecXhTVCtBgnldSYelGVK606Zs5t9kfgGH6/ryE0dbWio
0/TDWzj25l9SQrevAjSjsNdCBsSE9Ybeci4epz850yGuz+Iq7dNg3m2aUc6ZXU6ObHLy+4aejeON
0TYFFimJHaKgNJVrNSS22JZACN5DeTLkR9YtjlHfOO+PxBL+Gb3Co0Pdo99iK0Ph+Viw4gBssalG
S6IPAtW0lvrW6YrdWh2nZ5CeymdEaj280YOCmYbOQLzpkF+TQHZ+Jj6lxCM7xYpjPg9pXO9SGY3h
SbwYMc0cL/lstU/1VEgp1dhlDGALxPYYKGYIEqDCcIljIvb4dd8Hr3nUyhTnZs7W/GSsvSFSU0d/
aGn67/Kwa2xNy8jYsDWYXPUbupER9kLu6JquF5PKQcuB4geZjvNG88QqkAm3mduamVSvtgrCM1Lv
bhW10IOyfKwOkBe1kEuOptG1abvWu4/iB2Ik2j2nbTMQdP8jXSLGSDxnaSEiTd9XzU7UYPhRcVHc
WrgmFJpXGUKxp5H6VlpsWlPgao0DeeyinC41ZkVxP+nXDFO7wPTcZf36HiKoVFiSaC7cL5JCE7BO
/12sTJuGUV1z7XUb2/9ikNxccllqseu9icILtu0CDDeZnw2ZaDCMN0VOMAGuUMxR6WKjl6x86K6Q
43TJlS3J99taHTUGTPZi9kHo17et2EwhcctZz18UFtnzx9tHa/hOAo5evrF2jWmYhO2hxLcrOcK4
K/xEOYf2GzuSfI80bLDWzPkum5SYFdlLSHbRPRnBCqnsI84hT94C1U7bpZYTHiGF2K7550HjKKHO
YlrA5xJddrZcBkf6eVQmS2/E4+G5PC6IkeO8FCb3muINehjF6qUiAhOnL2TmCZd7sL69SIrUzEeO
g9TT7COyvQUSIJq1E4WncUrwwLDBEJhPC7hw7OMBDGRtBCJ31ruVxMtaNDAUbT9oXgW7nFeM2FRQ
zBbh8ZAX3H2Zkxveis3XEVgwfcQ8NFbjusyORtIAiXfEMQgkFYrY8YzcT2IZO9xV435AXCnryM/0
+MOF09hzlIfwXHpYaIzq/3F8Jf8iD0tKU/T9bfkxqCxzBf6Chz4Q8bRilSF93ugr66r5oAhPvOoA
OyeKTbz3gRJC5ek/3HcXvDiSCc9DoyVAT0qPEHlln6Q6flgXR97/kPWpERCz2zprdRKzfvPUJCqw
XiyPWxkhKzpb3oFcHk/YQJFIHZ9QWQV0KW0PUhAdtdwwPltSnI53P2Yy30sFXmuQRAMxHl7NZB0k
7da+qeOD2dKhCEQnKJYxz19YXydUCxr6koa6jqT1CIk/16+EPJGKWiaSrRJQdL9S3QEn+UpGTaVH
mw3RUheAfJvtJRguoaq8YS71jyZCPKOAih7BbzfxtbDBQt3wH+/L6L51taQpjCZtcpvOVv+NN2HH
MT1SR2BZhzPi6xhjRoX+7nNdsBS1z8n5A/srKXOQrxEB5cWDIybG1T/cw5VwVriGVuX7RvQcWRHw
2AG+l1zsmet9xjHj3KqTvMMI5ZlP+xA3KbXZSyaJJhwjbFTbTTrx2HDjrJFuZvnVGehi1EgeeERC
NBh76wMU/e/l/GO0x/cZm9Woj3dY9Yz2439nWA1RLy9i1TkBnF9c64iqfmiAZ1fjHXYz6NqjG3if
GPgDNkAq18EdturpcpDHMO0eF5FMe1XvR81IMAQSuBFIAsoVYRhnD9CqfNmynmoMwc8EFXLozX5/
xLH/8VpXciwgRtyacoxJz1zLUWuyKMXjKxuw88/ydpqIVo1H5MEzhapDvlq3KJQnM2zfcNA3ZaR5
sQyYe+C7rdeBwvRQhnedYvn9l0+o0bmQDkMqHHs9VjazDEvu+28lS8lMGrzSRppZueY77moJGo1/
w2YELLgy2mSAz1oieuoQEWWOu3O9tR9E3tWf0sAm+DPSrMQNCXwWGKVkJINI/zxsEybS35KVpc/g
CNNW/bKiHnMsW6XYEJ+1I4RknScZkPikoVSUcmeEnW1uBcm1fWIGv+P04biw6aV9wKpzHWLKI0Zw
TG5DozCREHOI+L/ZAQTpML/27i8KFiWkBk4uHojV1ymXzBncDbfvPj+Mofs/YpDm8PnA0zmqBAxT
U73ZkqdQ0WqIJjd9XRSiPn6o0L5AaqJy8z9fJtxjKoLvYedkvSZMHLoaa3GvbQuxD8Oj7JaYSjHM
SV6DaixytDBwxjuZo5XAPR8dVhu0xz5La60ERxhoAm7RO61QZwofYTtMe9ih3D6+AGSpi0E4N6bk
HJAJsRaAPPiRCpbyvjsgTIcC+v5siX9F2fEvUca2HJXHtcN6six9QE/c/ZvHPvPCwkwrChr4ISaB
ubsXvu7ADOOr2jiC4sclHTqSqxQSAFVtR/DwtVs2m7civLMTfVd0kBLjZzN1OQcYMHaQrkSIdSvR
ZF2g4moP/d7sOFNEWl+xPa4Mbt+SzeVluP8cS4pkJllfFmqLxqoQ4jtkmI88EN6rAzK+GPW0iJal
OLfy16S0oNpiTdNyWf/uUA0DpVptP5llXP87/BVqd2Xa2Swnowwl9oi98uN/R2Go6JcNvsFX3hCm
JrnWqfWffY5IPYEy7DhVY+Ow+Lmj9OV33EUVQCCe7Phe+QZ1OqVbyUcksumRdPKoRT/3czb0M26b
0r7dZFKbwHP+tFjzIo++I/5DsWsvEM4v4v29xg0sObipRUXlda0uhRri/dIZGerWWIZNDvIxREZ9
xd+qfQfa/gdfJ7cRYfancPt+bD/5XMlJUG0mfWYvcZRLcbhWRoowRGmYM38+93tpNs5RUIGTBiH/
kDc1pgeB1fhVnSgoM5l2bTVr+OOGlD9be/sppkoKVRqrTNNGEsgjdHv5YC6hjZRl+fNqqM00OS1c
g4SiI3R3YzvTbV9kiN8hvRh5MB5S9xd/tItWwZZzmvnJqPTcy1OGDYg3fA3tdAB8tUoHn3t4PuY4
WAdVOcLKWwLcgPS4cx1nTAxUqG77T7g7ltZpvEdOsXRJEGk3p9v3rh2vmL6DiW9p4xQYElJSIpZB
0IdgelEhD18xXWhH/k225Ir7omD3klPi16Kgpu2HnADwlTLif57mlpq+SnWWq45iyjjMMfDTQCoq
xjIRumFeapBEOGjeJCZvJJfgEbhUPx7t962QeU+fNAVfQ3wZ5K8u9B0oXHNXn6NRL66NmXCs94XR
8KeWLddoQ8dYmRrelCZ182cery0xlZlszTXXPoR37JhkthmMW/SlQH2GTONM47RDmnjtTFgqYyv8
PIE/+xmPsWQ9qx5CWE/6G0Y23Yf6oPP0yCnkWLaxHg1U5VFb0FL07lZAuAPjuKupgJclUBwf6LNV
KRlbChARGeHO3D0zov6RavhGiw2n5UM2eGsNRODcfdgw3d74OPimA2PLDh6KBm2s9DVhdXqyIBpF
cwZ2KaH43ckyM2S8WAt1yWypcKASuTv3vh1u+3nSZ5PgsXfrRxapxhFvQh13DNjMeZtLVcoclc21
MQPnWKvG0gzWHmcTDVuhIPFpUdm/webgNxHUUYpZZV1OssqGG0HyZBCAWpjAkr1Vm0hZkhzS1hWK
4ZzhsSbcaTGuCUoRdCmAuZU9pBsgegIiw2ziS5uqK+rnzFGu7nOQxNURbG5QmNwxZAGegCDHydsD
QjLE4+XIBjjnxODtHRv4IyAO5gQN3NjxozoMahRSTc3pKHHfZEmtSuzQbcftnieOURbiwP+av1sY
zLBRyJ8juUHzY9/qV+KeRQuSShLgQVisw+44+sbQMs4faYC1o/FLOhY+OyEFx/rkAkOYYdpmGaCd
mZQKP8IQF5clB3vdABI1G9hItGQfSM4jSqf4F/XiEaKOAVXXaWix2lODIQ135ri4DI9pUCFJD5wo
WkwxpDG3eYOKZ7jXuDpCfSKCo4Xc7op7jH9LJEHIWx1Y3oPrSGiZrcEIqQZvDQOKfesCeXeV53IH
2+Swa+XHzuZRZHv52QyzhwnmprdLvR3ijdf8UyAuzDMsgRoVs6KVCY1fWJUFajuEh/O675YFBtg8
ocVLXIK+F8SgAPxg4NYnXudUJyfC+2I1j6pziL3dp+VV3Sv+62NUuNtZFNXH5Kk18bNlaAu6Z61L
Kxay4WCuqmRoXqQ1tEJCBYo3U/esYclAoNfDvT2bNeDfUfoIMN2lrw+UMFZh7bCt4k2DBMHNea/6
L5j0B/X5hbKQ1l2nIPXIJEYaSib0GTvoEop1UufuurTZmJ86dj4fU0ho7Y3fcCN8HzJAsMtw8HEh
l5S84Mlo5lgFMpo0bz+HJlYzYfFTT1ehzeyVW7+Q9SjYkRFKJ3Mu94qQeQk4LezXVUCaZGTUWGlv
NhR/DHtgvDf9xESm7S3bn3LoJOiuUJ4IW74Dl8rN2dGrODPNOM6d3L+tpoZ9opZoSInQbDPKo7CH
RX1P4wIxranphAfHzOhWX6TidOL8TPEMnDF99HLwsl4m31FTpXdsmK0CNPOt3PIPHvtzEPTFMEF1
FTnqz8n/6qve/JJl/+gywz6JT1hvQZWVC4C9GC5C5bE1zsgzgwvF0Spkqxb31fGippcvRkQMtYCv
u8BmQfYb2p0dn/zQwOZ+p2TgaMvwYHMiSEmcrC0asHtbcWRPemO7Y4xs6fiY094Jo4/p9yQaQIFS
CmE/DKXO0W9aOf8/a73kWjUYhFfsDliAUGpsDw5RuiszGV9r0eufOOUAxbA7sSks46wqiOZc84G1
Kp4pqaKtQ9qOP50mMZZw0lk3Qdd9yfFD37eP1T8Md4vbxvViS6o+AA6rn8fco4+nRVhQ2KBUGq4C
DIDG3OtpZNAyGuWUP/4Taow9XpZpT9oUGqZ6MPnSrpH9xV2mOL6lne/r+l/18s4dlb4nvXpb7AYT
5KwYCfMHL6nW+XRGVw7aFssaPuXOoxZqssMfPciR/7YE/BcUcg6Cg7xjvUxJ0aqRYBV/7R4Tetg7
4iGCL4jaS+QeIzVXKwD1+Dsq+Qmt/DLyWh3d9aEQSgYJYlxTez644KpFLIEPTZ2PCsSAYrcKpL8l
tlBVfjq6lyID5QaifyOrfealv+YJU1WUgLBazE9q4VhN+N6SKVS/IsBCK9BX8Sr4vS8CQ551SNZA
Bs69QW0mqLjPrJC+GfUuHMDFmnHgcTi3NKn7XsufGzHNhbz0WfqqsyyK2+7PVgHy9tuwjwBtX0F9
E4zINnKyo6hek1cQ1/3gE1YjS1rcQztCUO5XMuwrOsAKS9uaPQN/kA86T0j9hPuICUMHePKpgUs6
Vnk8WUEAMuZbyd7vlVUXZH8w/ngrEyotBGCFExUKt/jLjP/t/jau6DoRl0uhAtNoHGHI9OKVt7Fj
hMDXikDHNl3FESJgCswTo6fK3OI15rZe/+un//tFjcvSeQ3Axl9xZB0hD0LV/lc8/BdLExHi2KSg
OyXs/aMk5blaAGiJMfK2fbJGkAxeu7DUj/asGlcXXqCYo4X4NNZ585GRqy64OPpOH1MprA5nKqcG
m/Xf6sfQztzntEEURfZRHdUzx4II2otARvbapPt99n77DRxaB5F5lvINrfte0fNE58wUaqYpSNmC
wxaY/7GHC+psOt+S2pm1gtDbzkxArNnQN4GByKz8ZysNh29Zvu1/bX23w3bDZes1ChdRMDfB+xr8
P8aqG1YHCcvzswW/oDofFEeQSXeh0RN4+xWIXZcbK+X1Jahsoa2hCCb1EVwhD0viXvQHqntrJOWQ
kbHMAk/6dyg+Qr8HB3hT4DkSMtE4sjK3RkWh2jzHSIQ4Ns9OnJnZ1yUM6Hs9yB0acDOhyjrJrW3w
fx9X+TwfKA0qnRDi3089tAat5QMlG4rUHyVMpHw8/+SHZ8840vluHsc0poC/vo7orHWUXKvtXoe/
6H3UmHVbStTR9K2SGDSsNqy3knzaZjFJiM8aR3fCuZC0g0LFF+ajKZKWFMUJf6/hqSRATvx8aPni
3F8cFX6NVSIRfccAFhu0gKfIExz2h3r4c1I6Mte4g4kbiULMfp6j6NS81Z3K2Tif0G8dvq46kEgy
PnJUUmYDVCYelPLIg8Kl38zpSbKECC9Pf+81S4aRzsY1LVzBS6bRjyrJcvdvREdwS7gb+xfxwlSH
rY+co0w0dCrj9OYp44t++aoZU2BiWkGxx64YtclLkEuMKZhaQUrHHW8sMItyq0Bnx1iuGOYz2ZET
qHKG4tIfLSWPJIUiLEeCBX6SMGPQQpiAkGdEVSRLQ9ZlnNcrbImcIe64K1Zz+Q9+DlbxX9+kwlO3
7x97qm9mM0IQo97gvSGWj0Tzw2t3H9E3vK56sqDwdhFwscpKZezzKzk2xb/vuC1iHtNy7E9IIYPf
AyQwM11+fne3mRWe6jfrRaC8/Ma4nTXDzKjPscUE7tpfUQfCqZw4WmVzgZpcNcjchL/I/5bA77Ky
tC3mt3FkHN/kST+WJpXn54afQhVzMc1dslThxROK1kINTguLADUlg1UgE0mvIzQk1smd9/Awpkzw
HRI3y08HddsXf2hJa+30UbM3zdC+VWDHx249tpP3QLfLui6xe7zy6T7YjgqCKVe4Ydz49lnkoII7
4mdAYqXZjXXWBwbreY/VOPoANyvbcuNjiYKTY77vbx158hwZO95BbiNOhXIuSlokTZ2DcvEn6vZQ
8buOyGc2XfgzQqyYcNJWLElemN2AdYYbbc1XlyYbKHw+rUpJNitPDjEnKTMUqaFV5MLzZ7GoxLQb
/otGlBuU6cDhZDeytIkEyY0j00c5SMR1ufwRBsa2rvWp7e7y4byAs8Tp9ddMxj2/vJLyT7vOiAjj
l2IJfFAWMhE8fkYwQXfX2s7sxSl1NXo854fU5AmGNh2R4hX0jsJUZxHpIj3X8+i1Ez9KtUM4GiLF
une+NVobABMd2GGHjwXH9FwdxS8VCHnDxv7kSHMOCmp6+4L7rTM4FMVDL3TaUFWDZd/b9TNRkOa5
CU9iX9YdxV8sO0eGGbB7gfSuoV1i2m2klHHu6JrJUngrddmnezu/s2uvqCoanYekmJjOmZgfj56f
+2KTYgNpLqBit8i8YW1ZtPXYNJ7Maxwng61B+BbFwux2hzHnkF7cVGGmwZ+yGguhvN4LNRJGRM1b
JrSvqPBdGpNU6GUet7cbQq3u2dIwnLge10Syp0BAdNCInWSOu5Lb7OxD/GQQWNqtKNs0zfZh1nCr
1gHOs9f6VlR7+0kEVUuPX2KHlmt0ab74eGcjoFbOrm7Jd3PezRoxJBO5Q0CloInQh68jEzsVKYEo
4AyOfp+eZQTyVFSIwJXw6yCaMp2BhE9BWv52stG8J/K0QjWccmLsHIn+ilYLBSSe28XdazcoWvYB
ECNUSwqVu6WreHkA6o4iYhrJn6a71ea304t6cudjd5CoboeBkeYS8wXl/tI/+WoMD6iTrhYMiGM2
jBQQg8XytJK3Loob87z6O0g58X+t4FfPt0o6eSwjzS9WLTTrpHLvXCn01LRfT1ZE4GhjDz5SS+zo
3rrlDOS5lj/GJnRWKWdXX8SahlVz5ZAZUm6dxl3jYFiF6cTh0DpJ31mE8uFBsNF+QQmoiNcWTPpi
yQ1ote7d61U2jAGRpG1s1afl7QCyfD7z0xZPeSxMF4V0I0iwMgXp0HyCH0egORJ5SzT0i+OW/fhW
SUNSnAdgVViW3+h1ZqCCZ9yWBwiqt5KO5Z8TK0DBMO54CwJ3O6FSs6J5+9kCiLW6ZO6b2hmDTjXd
otqjxmkrSlnZ+rtW/SPY5OvHvmeTR7eIsIrQ4Av4np139KrD2V/CIwUXGguWXNM1ydEpH84VP7Gg
1lgKgUF7bDRbn4hWG/GDvrMtnvVkVHnikwij5k1gDNL8Bz7Fh8flCLVnEOZD0DPF/XxaflDmoYS1
Jj948pTCFt4yC79rKLdTNcz3pJrl4lh3SDoMrAdhikyfHOLwfoMOGASGKjdZO1TaB6pXFbKMiQrz
kKFvjI9JotJTixBf6Zzqx7l0IN3VIBjSYe/QOUUvCNHHU8/zZTN3c+K8iQtkJfeyFJxIigkzuCm2
XV6582lWhltpgzRj9yZC/84UBxAxLeTz+HGB+e/gqAHRuhS2icWMo8ATf4ldgaiKINXA8th4j42K
s7PWrSyi645JxD/qTWvOkgiHLhuRwBXTvwBsRQWLNfePoCoVtlYo06dHDKR6Cbe6c+4CLJpFXO+k
qp8pHKttXyCKoH8v1JagKdkccQezpJfPpmgHnWtH1BOZg/uvX4CEHnfdfBvQQtY8Qe5YrsMq9R0N
fsSNvPNFP0fGSKwtcBOEElO3wJRqlEQa0mzmuxrz0khdX5NW0UgRwOGfcxaEvliULalXyzVybey4
FQBWP2fYnucXlXq9BVM6Qxu71QinXRpeQamOjMhpIbw2UQ9blTtWbD6xgi6DwY0bE9gWHFUahaIh
mhP0pxb5/R9a8nedQU+LDvQjjVEX9jkqiixfBJCMErKSD8si/tllV2xnZzFLjyPKXsw7YWdfw+cj
+iVe0dowlXXN5zr+nuVCn7wjj8Nx9YzHvxJo8+rgQ5AOTupEN05TgqSimJxIkKBubZyOapQTz8eN
vEcD2rexOUaPJiJS6RKhOlLNbpywy8pDFILM8L73kDwiiQ8PQrdmLKQNfJRYVhd4ctPLmrYBm/vw
XMOtLWfcEGrUjg+N8mtrYl7xRM3OcFfpqTH2uhZe3yNdStq4gnogDpbLV8SUJYfeAYpI+lUaghpy
iyH7bzw+KqbuvG6BLG+PJBbZQQ8dQhmKwTOxfP6w1l0kb4DPq6nCOJUFoqfIj+zKreggXmsBH37b
nkDQJ+qz317p61aZED3s6AHbZQwo7PTn9/udEyEsaeNKcR73c3ZuB194jVwsG+Tunt6vDoP03eWm
hjpIcucVWUK+eFpy1RqRGhApZIwZUj1MUNgLcRk7Muzj1akN2vXG1fIyJnR3KrIRb9qhjDdlRxXD
diMQOkUUeSXovZVIJX4ACydMJOD841/QrCyPnJMb9pONeblm/QBQQH6wu+uqCXs8MkzP0Ec+B07/
Rk3bfTWdt1ad4yEvjMpWHQobqN9jbWWDaZxLBlEbPuAz4cKLwVpfPQsjKDuOCYVDOspVvn6QGEle
7pVlUMS28QEjWs3dBol2A5k4GeA/wX/5MQGQ+SoqSKuRcIAQ16Bjf2v4d3FO1galCeZusROJDyI9
1xTbgTXY2im7Ah80dF3DuBy2l5/5RtajLG+nrRsbYdExqO1mnCnJ4mLd7Fb/hnRG+69qzohOXGY6
e9ytSUr38tZGzZzcOKFjUMYTVa00CaJdBtiJjFOepMni85F15LNBVFOYWqZROMXi8IawRH+2r3Od
bkq4gZpCLEhVqR96Tka7Er8W/8xw9yasugvcQLnBuuUPnTIYs0/lFHvDTwO+CACFkx4o3OLfFk6E
iJ7w0mSSrwM+bi+MxQXUvPDbU6o+P2gN0G/sSOhqWg8ueSicNwKkN3aMZZ3fRlPBezPs1fUmoU6g
aKGqU0s07bJZfL59dNlv40TXwKF4+JUbjTcRfOzH7uiPvE4A+tTwt+jqkhbCBV0S7glEexWjC7Qr
lw9+gAHby5g8z3VBULhRL1AWujptcgI2o4ffRyf2aDWdRdi/GO+RkPM2Yn56gV66J2BrwJ3ybjME
cYfxMyNFW3kZCXTHmzKCYeQjVZw2TnTVWwGORM0ThVTHQQ81LWPPXGSJcb0bnDlHmaV7FjqFpY7c
ovnLpSxDnN+Zc/VeJBkB1OgyPKOhj7k69LuTOjq3vfQz7xDAFVSPQbzrWICYAzJ3azUuLafuT5BD
6QCdOSR6JbowDmQGg/zuBdeGaXJbO3JaT6A5CPpr0MtJ27woKMyHpJly7iCCVsMtJwB8xN49+2+M
PV9L+IQMRGiHAOpNu9CGWZJ69J8LYn95zs5Hr8efrF+yJuWXYHNUMawLCoI7PlmPzcXmKJjX1ISz
oWUR2Yp8Uj3F8kpm920+XyDyzZiC8ANlOZ1BtCKRkB749aDwYdOwWLLFTf6koJRm9yZ9evkVvdj+
aEerHAw1V3YDwVOkpcq3sJkI80dVaIhXdwPmpz54LFOR76h5/ILUuxbai+LDkltu5lgB5qbOgL65
+QsAgGc256lPg7zZU9cHyzLHUHiaB7MQ7GD0sq+8iuqMjP9uYwSjqi+xO7PSB20TCHt22frnnjVi
67C7JxpNEPtKu7klxca0JSMFHNA1VofzRuMsWeav4IK4n41aeR7oGfoUk2vonK92JCSNn0hDlEl3
ASY4FP6h8GyezknK9EXGswjC4+OuurPGfFZrAI4Ym/107dss64NG+clRy38+BfERk6u0i073j0zJ
EfqI7eaAyMFTo4Pc9gPu0fCR6IRiYKbxnCc2B6h3TJGl5tBndvmQkRB5JR6kzLnk7EXyKMcKCJEJ
6EclIHloeddMZpEkH3xYBc6e0D9Qw1mpxJ2ZWE6vTfXPBfAFWKM8J1lEI8UzYu2oOZiqs1Ze1pJp
+hqgMQvkcm9cBJw7cpi08Z31KjNHvTHxPVt3IUWXv8HxIUKgaLwzraWlbUApmxO4lEBe+c2qElCr
nLGEiqek5eWUdgUyipsckWqy/Sn6WyGl/9zBWu0R70Rq4qRKgR/L96prHCSi60+EzmUcN9NjxEdh
CBhmnwIYqYwIEIxMhxADg4qa1WS7M0T/YqER0m2tk0Lfb9WawXs+tr+shwW7UXZ4xku9laHcqIFD
0oKx0saEcCEzoJyzsJC6eyMXNUZwdDdxXyi8sSNHTm86smX9VKw4bMugd39Cou/L1ni/b/PWsMRF
8/QJg87ixE9KzYh7f1h1R/WTONbep8pCKn5GrT3Isq4D3dsbkmJysXNCdvjd6iH9ZECMJZO+H1tr
etRfMAAxQaq9TNQmL/x15AXb/EI7yen+MV1dzgh0IUN+Hx8z3/2+v9MkmXvC5hu+SJePO4tNH3SM
KD5aK/JKPb7NH1bTLYf4z2UDBM8XDP44PBUgiAAyA2YSxWE7LlUOaMHH5rAk5bCAGOygV6RgnOXv
ihOKH03nc1tHQ68trXwZfIlU0fwPSB8XFPbMbD5dnK/x4bSPCLnQK3mebdvqKdme0MYlTlYW292P
QcRB0EjWpvfIE+RLYT7BQNd2N+v2Vp+bbDtFaK70J20FC9MA709WV57zCv/YMQs9IFwlFew435Hr
DQG1gA7Zuh9kHveWFeOnz4PAaO2iuKJHvJd/cXLpdreDAWZPKiqJPCpwZHoC32hrVKCXXEAT6C6N
m0//gKW/L2n3wUEo9NQfLiJlajuDquK7iW7cq/DPgjqhKGmUbw5xDI0jqzEa7KZzuCdmbnk8xM1Q
Efa0p4zLSPWLLDy1uiwj72LQo7cdDAunrFKFaR37ett14lbZ5iHtLaEL8pQ1W4uZi8dEmou4lmLV
w1UvmW8/kx18t7JKN/8OHYj5TH9qj9swKjaajXK3b5Wma4rje/CVKdsJApEdBaZGgkOzieSALjDA
OnysbpdBsQoLdEqcF94V7zb5PtFkelK0PzxmhbiJNc+nm4PPl04twOP1u87CY/fI/NynunzXaFro
LMJZPUp9UqqgW3lZXgiS++C7RLgQLTyfJt7F4lKlPGpTwiimcDH34R7TCbqHpt0lBZgALlITdYBM
RANgiLoeR5mno4BoOl+6WWDxImoBIZIg5Lw8M76NCaTXYwv0hzslzqWLyY9fiJcEJn7jZ7x/bcl/
AXGzgn0DOH/B941AdBUZ4Zd8SQ+MRU9RD3mmjTiQkueD5uf/G79xQ+K4ntzCv8MGLtLm/GWrY2BW
FeKSqaljjIE7jVRrMkeXE02QHuti/D1v8aaempJdTietjjQ3SoWy5MMcTmTBI1Pr0ZPsEor5CPId
6jDNQ5WThS+3CcaY589hdwlbsT4lo+Cd+wslQohkLIFoqIMChzM5ebaP5ULlbW5RlBr6yy1gqpCd
czeYfBrIM2vMxMWtd1z4BjkSH6AFNTWCVa1mbYnKvgTg9IFvLPfibgiqesEH9n+VW22q4P0Spt53
AAIYDawxj2GkJkO7u7QUNEd3KXUiuE3gW//hapMxUHBOeT6uoSvDkpCiqt1Pm/kg81RzQaKqZhuD
gmMKTm7cI/hDvpbCEKL24T2dcVdVX9eaTMlzCLtDMijGKqi1NlVmjrxhKWSe91DuauaSfzb6RipK
bygQC0SS+vSNn/eP1PWs8/EQu4mI0MgfeZ+ezyY5my+wYHDVuo+D1X9UTgjQYOrYNwPyoHLX5oD5
JIQct1o0PeKcNs3k6zHX/sVcrRDoC2KrqFdp2NfS7C44c9Eut/Bl8bI2BM+aFmGGPMyqYTj06r1v
jMDL12HfWFJHFS/PeYfyHKwpgy2HDhg+RWaFYxCYlhNdGwZEzEUYyznK0zOQNjFCldVbH+VBnwOr
DiXzZClvazkY8UIUpV6MyFp0MK7Y9zoX2Y4X8kMP/B4oNRKVh7Ij8wShHuDw5eRe0kdbWOd8f3YD
O/iY+8kRUEHuLZdN6EJDKKZoZ9AIyLWtxPQgpR1IptO4pcc9B9dm9EnwjPVXyIedzdKLOXns+fqP
4uiUzzB9R2uhwcjNHLPY8wslQJSmujjhU8jLjlHyDLypmH+/hqbz5xgMMj0vOHmN8Yxtufaba5lh
556eJOnGLdblr6X0VaZdsquuQUrT9QyiBcTU81iVD5UuBSUl4peLeFuD2octKUl0PIJoc5PyztrM
Tkztw2lYdSqyRjvBU3pliTRpv6DuWB1LRw0LUt4fxj6izEt3J8NCjPzxt/lYaDFAn5KCjDn2d3gq
wD56tUyVu5ujhd1RXP3mxM7ch1DKs04LP7ghF1OJWGiiz5ltvS4CKhJ59KexunhHMV6thhO+bdvl
3snfg/tWJGQfPa+9ZpfejwO+M/oGI61RoYN9OeGIoQlefxfI+AX4ijtwarQK/yA1m1HssI7z8m6P
4IT8/3FNKlS6rgupWPg9+MvjJKkkMhPKQhfYoFh33xKg7RjHRiSiM9EmnsQKCBCY2SCTF0uyNAg8
J7mYVP8Gi2vxSxfkmGqV8nAhdgqtFt84MuCqED+gx8IqRhXyhqonwJymOzcLnRD5RkdtQRManaXH
tsOeOn23M/034cdIZp4+0M3OFjmK0BPIOGkmASaC1wWrrVZ0e9H1CY10JIW5Ci+r+GEmZEabPLGE
ncetOT7AmPi1qBcR+ejjIJXPJx1Mc1H6+AfS2m+fckeuzHKzmKoL1NJmCTCh7MM3PAOPX8j4WBF+
domUIvBqcvN18VXPhiJOd2L6cIG8KI16kIau4sh0jeiasY4W516+lGAipomXHfcqitBscjubr/sU
HEZV+rqlg8rmISGWMhPdYZtUmOwK0lROLQ7nNhjnPxCeQyC478O+g9uNVqKyrDUv1pjm/Pp4eZRJ
9xVRK50rCFzYbN3Z7zxfTW9fbPsYUQEBeFDXVNSWik0n3a861qui8toae2YiMerFg0Gidk+L+PBS
4/6lzT8O3/Y9Psy9X4mx7LGU8sBPv63VsoWovn4ILWKY80ciucoLn2VuDa9qycTbOOUwTPEkU7GE
2HPNdMyYARpo8IvSW53y5KxAUk66+3eza20OfvRHtTC5cvMgHIy4znBJqbodniMo/buRhFB902w3
CHAHVOU66untqbE+1VMXjsrsyISEI9lTIJWm/Cueo3mihsXPcWUqJXnldrsBi+HCMqrVgUlrvUFT
+KVD69emckTNBvfx4+3LsQuU+JZaEw5ryBDlEl1gaX/sXuyLEPsizBjU/fAR0ALq8CRVoO1/7diq
6FAUEMKdEP8V9XZgbho0TV1BPWKK9/HN2kQiF0cauJ4hQhvvMj/oPpfm0m6vYdW002Q65zl6x15v
yMbF97iTE5X89Z7JZlrAaj9A7Kdt/DtBzGYR2CeKfy0kSvxbuqaMnbJ2q3gYnbUxuDewMZ9YZax7
YyEH7at/nbH9t88qeJEA32Oo74vhQhJM2F5CvCCwPF5G3Dcy8YuBeJ8Z5XsbqL7foxvbfCpSrsrn
9YIHLnT6FjX/FwIxetv38ZYMcXhenlQLJjx4wGqg7txUZa1vvfzEFGGyuoY0WIv+XgFcQYSIRonE
GLZnjxBX0qe/4iISxRolNBCkeeSPek1G4d9eCm394kTEnHTOdDpInXMWPdobGTTdmcV3aDzGCf/s
s7l3wgWRj9dsTcOBlKWllVBgq2FjwGuHzSfoQCloAeOollhUK9MJL1QsI+uBN1MCsx2Q45LrkdD+
El87WBN7fv53RIZDyQWAbWfjYGEA0YeWYnPMfxydDBbYeaDDvRTvOjjrwmA3MLDrMpMgB52/X5oO
SG6Ww8fctYVSdycLTiVOO1EYVQKW6wBMdtVqIQ4E5t49NuTQIFE2cmhntTllwg/E9nWwqs02vldD
D5ybxShgetm7HG2RcYcN1ISgaj/UwB0OW4lhubf6ygD3VYkjJV/eqlEgsDqdo9/u/jSU4C5bPTez
kQeNaMc5DkDwkg1uDPuEk9FdT0bV70EOQMX7G5fz7BRA7QGmSvy5VCbN/TKSvE3ZLyY5JI0UqT1D
VV5bMBIWlonXwixRb9c/H6rD4g50LKuWQO4heobwNKyXWp70EZMyr1QHJPeEwRiyQ85djzuWCl9D
iSjLvFPHrVcALe60QnlOM0Usv4WocmI1I+gmmXJQcLSlRc9SJyzVI/r+0pCdRpXDku+7xv+0C0ys
4P+SI8La42WjS8VjCSq0qXzL6/RB1/5IzeyzIN5CdAKdX7/Zw/cC+/4TPZgwNGrDprXnLg6ROuvB
M8JGQm6jAHiQN1uOl8WbN6JoqjkffPVbGy0IkIpysj3FOMX0/c3AO/2xcEpC8SBkEBFejEBjCOut
m9jdYN0pW8c2V4NvV9swQf945bLWk/STB1Nr/hHM3NnnyNi7/rNE2W9ECx0ECUz2/iz1QG0HxBs1
Ru6kue7tPv8rpaWa5zUFdN0PmPUeEqWh1YdVbCq0+1etvciAxlwJBTDQpnq/xp4fG/s4ibLile5X
8YYKulRXkuBOZV9ifiM1ncHFTbK1qJvXAVA1cE2oXW2PnrMxgNV/pGf4aBDRC2Bmx8J361RqQEla
Yz/gQCAjNPRLdY6R7YEZ6qYtKAlnJcnsANEQiOhCTmKPcTkMpfCG6CiPkugn8ztZJxESKKK4f8Hm
xkOmIyPGY7yJ7w1YQ9CgsrXJ+q0+QqxGJf8aY/3qQOx56L1QdjMmlmVdW+8e72LpGQjzgjGCExOH
Ni1MD8Oc+GfMRpg9BF7Zzc0tB4HQfWmFG1Up4yFWTSmU0Y4jymo/Dh1xGeEexvbr0WBIi4iQeJVB
jp2d2s0O7VZaDo2PNYH6wzU3h67zGbWATl/eyzyBau/aDlxIaK2gIq5UumaLx2clG5LqPH7N8ZmZ
f3kH95pcFe00QU4yQRp+bmrY6zrphFAVA9fMLJkWNfGFSCcgSOD0x6FpQul4EQG0eQRu8PC9rnRs
6iynVCLottKTinmXCnT9mli2WepI5lmR4Q9rOl6wyPZTRQcNs3a6mi5/2CUKRucOP+xHyLtqkdG6
sfPFaqvIW8w+sak4PFxjNt+inmRGKQhxdXx7c1CQlXviTwbcGKBsDqZzdApxRZlE6iB2F6dyKhW7
GOVKNdNR8z92KwGF6ZptqMMWBWf2AyR91VL9S3NfNdIs3pQWvyFOnplOXFh6fYAUIKdCT8qpSMrU
fLFobv+hwvv8ZK7GisNCEv6kAJKatPBvKfKJlSRy2JJZ+2JzQvR/dgZiPFrP8iKRsWQDEAGIr4Cw
W0WIJjUhcV9pf7+BnsTfikJg9rZizwxJnnWauIc5yy8zEMRwbJIxL6ch/qdNV/OHcbw+niIsxlI7
xrclYmfALySAZ6zV8FkkKndSPfyHSZPJO0b+pcfboyDkQyK734Z+3dn/CvmGucZJzi66iR6ez+ej
fDWyKeLfbEH3bDsKD22XNme6RnTNDr0LlSvPENQmWwPCmiTKm3cxLvHlIn7wwAcCDENNdKrunIaC
83JU6eWuQVXf4xTEMRJb0h2pFdKpX7RjxgN5pY+Me57lYfv/Sl7tJdzR8Fz5R/7jtvlyX3VDDDmi
MzWSGtq1Tn58tsQmr89OQYMZP5HLAkNSt7LwPLZ/OuJsLKYRt1yqrgK9A4BfY7z+lw8IbJ4MAOen
X7E+PCwOfInfoSqlBEp6lYEhcDQByd/GC+ux6YXxxsNItrN7LPDRBVQQnND/FFd3ldeGdG+4Gx6c
PJ7xz8GConhFqEmQ45ZqRLHlwzv1ouJ/9YGX2UiEjaTmfOoHsvf1q6Da6itv7sIy+6PtIu/bjXI0
yeqX8JzIPsvgRVYLLucCQd88CzGqLs2MPKoCQ2GsIeHh5u5o1YZB/Y/KBYOprTH/wn5lOIkTfkci
1L7UjrsaRxJMYgqIcNbbfhBC+L+GFVaYFvhk5uAOX11+1jhHgd14k+Ga6+/6mVYkyRDtHywWsexm
qctqaNMDrwG1SYx7bLfWZZ2uQ0/+j/ZmlJlQ6Pnl4yofqHm1BnmyPiqZo2QAfjfeoJPiNVUIOVKA
nvo6NwLjPVMa0GhtjyxysaPZAWzEu2/6d+mF9NSdXC1IXyj6B/nNmPJ5/3A2QOUbGS9lR/0aoAxO
dF9Z1s37LSjxsHjwQgeLfmIYjK1zNmekjcS1NZ2GaZfKmiCP+SxeEWNSyPTN7V+y5r55RWJ8Bg6N
x9xYtj6bqSqj//bZ9tQe2dzWsAeagnhWaLp5OcjphRYY75/2fs5S/2VrHUAcSHw8cMVcRjn1oawT
jXI5xPIgR9xqMYlC7QysV2HgF9i7hD93X5CmduspoNvXV57EPD9YM92AJjLV1P0vZJ9xn6kWCXSD
LlygyDwdLwgPvZmOJzqs5KgDjpKzuiwJQ/Ud5RtZSDN39tXu5LzNqB2Mwx67UNi1fyUF+093c3ke
eT7wAawHZU/uhfPxKn2pDSh0iVwYzYdnhPuyn5l8Dkj7nIB+Rhas70SxJHs1VCs/G0IDZ7rs+6l4
9Up0cmb9sckzsLSQlybuJt7iacM1bpBYSS4i/cZvW1DZQzqRP7re5YVTY7J+8RNSrdmiolOcLC2E
A/JRWzo6eBqnTuRXd+R02qAzIyb2lFBQiQ+ykrcmuzr21xT+XsnGrdtEphZ0KdqWsKEgSi+VGpip
65rP4CFJEix/XKL7vvRcoSKEBTMe/sXqAk7e3j8bcV2jL5rDZFtt589SYAe0Aoq118iLS34Sil+m
/pPJTohnvKBjQqBTSr04jZ02Sc5UCImdcCiQU9UZWJlB4YE7OEQcMVkiSJsf6JoRc4Y+oihI/wVd
UkoW9bnMQ059FFpw5jU2WaBdDdIR0sOj6fcJRjJsqx5LqExEZRS63SUZhqEP/7qjGvMl7eGbdxu2
/PsaDhbFCdoJMseH+mASipg+/7Ubufg0s8FukcFJu+3xtiEnP9m6IlcUAh57ZibYKhUqv9ZOkWJl
gfCMjEXh4Tnfwb1H1vcb91XiZ3ULhpHia5BqGYqnF0Q2wc0N6hvZZ+mFS8jJ6H3qEJkGZjKDqWEb
vY2gJXjmCw1c8DB33KC6YNnGtyQvn775q+IdFfusnWK+W4XWjnhn7WNWta/B/gxADHuCJJcaKcs+
BISf3i881xLL0Z3Jml8dFYe9MJv2FeiH0oSScHEOJG/0bXBRtI2Unr15SgO3Jm99FIeJfOHw+AJb
y7gEbjKT8Ihjf9mN4ibmdndsQ9MaBphvwA+C8MuI6xUKnm9D60jtKNn4MUht6Z46jqfPbvg+kkN9
EHaNABinE0OKTU7j+kxIRfF8Tan4A/V+6j8ujTgTyZ6eClU6xo2c9eDAFKcfTtzEJK/DdP1yCkgE
mf+ceIuGU04qG7oiJbv9vPEL2qlP1Qjur5fdVWZQOViuWZcpUQSSIPc6TyTmJMQ3bfRTGNob174P
Ns79oL6Am/7BqQG/ffraXcvgEWiA0s8jrIC/grIQ6ZvXI2/bbpb69HDroQeBd6HRw7NaqN3wECfA
C796Wzm07eE6hSJJQV3Dmy3xayzfYkyK6UjejQqk9Nls8F+y6AJAA0Vv3yiodBLCL7Po1mGRzYC5
tGTikNyagxKe1bT6ivEkxXfOq1jWgPK2kvP9a7UVEixHfvAzz1NznAEnH5/W3UkAqkDhSyuP139J
m/xx9162Kou6Mh17JtcERhsOzzCLUAQCSNQkrczdwAT7RvbHkI8hkUKhpLaggBaLLUEsN9pqJiDg
G0ZBdFfWL3gc63Omnt9tXbixzMQvrQJJ/il2GL4t2AJmqFDT3awpqxPn5OHfqiuGzzZJvvNW1qNl
gciE9Qj92c40ags6hXGYHNr8XGbQwwix9Tkmvhtsbtd4mkJZs19vxsJdeeZGHCroNS5dLjAzVhNX
qvnm/98qDv+rtSN+yeQQMdXBozCxfdN4yorS6ahB4bOTISzhQZo3dLGv6uRSLaxF9vfiKrSA6Fxb
vfiv4IimAjpxhV4ELia3Z4wca62iTiKy8qWAADbyvv7vSzqdiOvNFOTDOAfpHQpzVnrr2TUnoMwY
uCnriFU65RDZhaUlePwKnOfxJk+QcUVSpIKT2IK2HyMN4CBHqi/M0rEV47hLPoZ29qk+zw9RrxKz
KmZFlvsWBdNefiQmIkRsCdEEpQKkjq1Vf3lMj9b5xzCnsxyEJ0T5SHDbhefBNbeZeEz2jOc1aJ3u
JD+Q3yHjOZwJDvfwqmbbiLba85VBrISMk5d3PjyYyBhsaqMdrkxPZQTOvh8ZVIBWYLaX/L6DuZT8
yhsE6CJWK6n3vL0E8ZsWSYWvivCJwbd3HWh+5U7kvC0YXOz0GiHq4kaMClQ8C63y2sVnXggNRCul
+7k3MsMUNiuFH+ldkg0wR0Z3akUyy906kzVDgGl4mDNqf4JrO7xIGeimVyTni54/5Dh+bjYi0Yl2
2cm46JynoWPKrWfw+WHPM3IQ7N/gCtFbavMY3p+MYdDWCoyoTBaytz36qsqXLhv/y16U0D/ZzkhE
FdUz2gbZ7h006VyiT1n4i/lFREdh8PEChWM+SNz4f1W5Sw+x3ggELgIJfrhaKxg1j+OmTBooyVXq
wAQtqnzFJXQOV9gkpnkKW5Sj0soS3NidTHt5SbLxDRvHX49JTCOnoiNhg9SohKS3Z4r+Hok5Z58I
mX53z9KyAR7OZp1VjcQAZZS9DuiFN7UBr2B0iY5jRaOsigVw5234QYvNJsGYeTw2rpSgbv/BJXao
KiQVcC5V3EwvUpOPR1GS7NJZVssgDgJgkiWevbR6PS1Y6XVvnEGk8/vo637OgIaPE09in9dDvLyU
Yi9bZbET6V0kDXV4wMJVOuJyWcfG0au3jUqUnFVmyf6yPcRZGuTxkGdDk9wgPIEwv0X5Hl1gDSNE
qbZLwmqO0RfOgQ59H36oCNUK5zIWxF2p39rYBsB7UZsDm1q8slf5n1wwSck9XpyNdWfp/5CZis1d
noxTePyXDo/gWVJrGl0tV6DBC8v1wFfZcvIef9UR1cbQQiQKkOVpUL0WOn9pxr0xECIvWvglIww3
aAiLF4HY6tTYi069lhHhuiAW5XVElldncB41vou4J2I6zeqQKaSQZen+8p0rTnlu0H88x+7jR/ND
kqA2rwtpA8xvmPFWCd2Zrty0Hq5EdMDoLpORl9tkFLCHFKs55OGX+ph6qjA9FIaTR1wo92WHww0z
5MGYQLkNovZ2endk3HZVT9eh/aVh7rHviUSuld4KTysRgxPJ841v1/VqB/k6zNygH0AjC0xe7JRo
hmOKkmZxAaPt8SZg+kU3cAjYYx90Yp0ReXYDfU4PY1x9+O6ZVeJbk0ogOhMcD+618uFVqkKem3EH
uAW/BHvqRvHFfmyjiWHu0Ral4XqjD/sFpUBPiCJClf5nrlLUxETdrAlHp9Nlx/SgATkIgAcdp0yy
csjgquDYtNhzmY3WESpV0MB/ntE561zx7aFjwZ2lfwy6GRqTPyie1Tj7FZGvhRSioKYDqt47PYQl
b6EE3Q9OJkKe8WsPzXiNEHP8t7pNU+QM8YrpG3O0bZbtb54mxXoUMu2HgmSlJLDNQrMxpwE5g0xQ
KbMeP4McEyoU/l4HAvg4gm5gf2h5/LOq3Hx6lOX0P98A9YJWzFfAIkj6DwmLAhgIVhzpq6MoOFO9
jDiphGqbOjfpLiy58Momyei3KI8dXaIM+iLVJ1qmsbKH9uQdpyUlT3eP62IyZsMhJf6cTpUj+nBI
gOHTAR9Kx+dOqIoSMUHJSLYzSzczvlQxoN1MTMHesJLobOw8l+ketx3CbqKnUArtRTy4Y5icJiVK
PlXJGS4764lHNBZQf25yN3Skdu7FyIonDa54mtuI0/WbPGxH8Ror7on0OAfe3hco2W2b4lSDmRsJ
T5IZkJNPS+bmfIuYZxL6zHFUk9dH5uCVeS27rdPzLD+59EpVVGAaZ4HavonAR0QFR3Ws4svmBdxM
l5+SSf8/JzgL7qZqILSAgj8SlYJn2DTsX5bfinHcCGK4jaqwpXAPgd9+OHNOmXHv4+Exbd5liIha
6nG8cfH6ocJmeQnVM8BEzG3Y1a6b0toOv2PWhllk1CqgJoaKnMKPLFT4cLSy8h+xC97vUXx0p8EJ
BrH37tt1perVi6kHa9KGhZgSL53HwGDe6BAwPwcmIYonzk1h12PlERGB95/TOxcJ081zeEonbbfT
2cX/u7dpHOyAdDpmLM15lKaGbcrmC6OvzPUXFiUSRMkOanTXjj7Y3hamlVIfoKfzZYB1aAZbfi6s
tFYG9Odtdk3+Z8YxlfoFygPsBFxBbPijC3xMWljv2+UZhRLy7wKAPBBavbBMaokPX3KA5gl27d8Y
rkppCsXAVt3zIFArxyd1ydPWRkGBA9SgG5JpvqyXiG/p8/XxqDRVV4h1vr/7fIHOZ3pQJYm8uf6S
6l17cG4BL5vYC64bGGVKIXqihLrWXlYazI8W+MKCEEcnciRSWzeQOesU/WVVi82E8Tpwozy4mtiv
u6rC6QcDUgSP1kw5ignAc/exgUD20Jz1tQtXTWvuPs07NsleO2AReG4irW7jDDYOAABgM/T+LZ0T
BP1eClFfKeS/NOXIQp3gRqLMaSAr+cQEUH9GhyslTjn8x84TKF4e+GJyRItZWbNVNenkYzyH4d/g
YIZ7SUMQFmeRTxuWGGG/CZX/lTxchi6pnAMq7DGAjuwmWlY62azaDBvfAqRl1VWyINRd/xOh6eFm
PfSph1GowVgZGtKyZ2gTqWSbVMGj/D2EBMpsXybTGLzeWQ5qp5Vw3FBjc79nkZxWD5JA48iJWmtp
tMo6514JxTzpLj0kdboU0MLrXdDr6J/cabl2MH9kwlInkZN8IeoWPU70Vb0MAJv2YJif6nRRXAy8
cCvyq6ygrMWRYKzpWrnHQK95rKDOayicEWJ57l09zstnrldx0z51/uVsTzwXqRTPhwVqqkjiOccB
xjvYDIkPw2medjEIVQw2BvtezCSj5fjPFklVH8KdTnldTv5K5dLxv8EhIaqpEF5j6+bJ/Qest0mP
vMyXoBTvoiBNGMdnPG68BmXDWZ+rIFbOJYLKwbTRv1pWPQJmheQy5PX0fzOpT+U3M9gRap+AYj3z
GLq9xtC/ko9PW087D96CeRNBJB0YYZ9s2+2sK4GcEVYh9MLOCpqkV804WV9+U/xqh9dtT9LSL7bz
1trua0QsXv9CEbgDj+X8KG5ydZo8cbnRKwFApxtpd1iCchQan4SA52Fo5fHKOUA3YzSiDeGCH1wm
q+o7wZejV91xnRigQdIjdisF9T72kfmneYEyjnPylUQ6Fkl7Y9aObz3czqIIPBfwx3m33VtP4HJU
ihgDzFOIAi7F4DjYBD93Cy/iUfc7pItHkaWMBYk/lVPT9d+40X69p7OJkYbVmxy0BKh1nOzjpLcV
PeJqB7t/fFebdut4drutUBjzD7XjMfI6wcBSi5aLgKBjgLWGmvZsr+CAgyhrmbCqM5+oJ4OYakJN
dIiCCqkPqeKPqC1NfnwGeq8jWR/R+BVhkvprkmF6XKEcSeBPHG0WdhgD3LxwXp8xV4M+xZzO3HJh
ztNNEdHyJBbDqLZeBfZk8hHdxArU1ynOu2gn7HZyM5uKU0T224CjfXoPq+ClgMqowN4HNnv2ZQYR
xzYZy3AIAj9bKXbCM/eCd4DMO1r45zorGZRTtPUXBJDAx2y+8uRGEuOCjZ4SWzGuHaxnqGcvqlPY
yGcn8MJ9SZXyu0H0DL9miLZ022wlo5PrJT2w/JpygY8/K7JJzPuQkIRGT7pH+235ktx2h0o7PrIC
tMAKTY5qL2po1iVSElRH6yLHxg0+YfyJm8+XnuyoAebJUoHerY8oh0Ytfmy05YN0FJ2F+1iKHz1Q
nhbWq7dEZvj5KiwQvRfutB3t7nAbjOmcP+vzdz7UCm5oChbF/sMogGc2jUtRUObMSHgH9myk8hAy
NRWa0OXNtJsw3JuodpkczdXPfr1/cTS0v47so2XKgqykCPRPItrpCsmVRjNzghZnulEYKGkUTfO7
6d/av6x96LmY8jpGwfvCWbWA9oaNe0NYc4ocVyMQklO99B8WdLahWvOQj7Wf9F4gXii+17knvkP7
25Xd8Jmdmlyh87cvuSgeka9TVjrCoiAPKcg0v/pMoNUipTQg/8zU4EiJqfJBJehjZTEDh8MP3Jdk
yOmO+8JFJaX3/XbUdqMtr6Hcei9ekRqzbjMKAEmI5kb38TS5K2ybPWKvTA+/ja69y9QomQB7qjTo
kLYnYG0/JZABziPMrIR5A7fPnbIcKr+KgNEVV6oz8B1iDIpVX8eP4rOg1ZfPKcDBF4lwmrRXt3GD
sDLr5dW+1CvUaQRTLTvDdh7zlLL8V/Kt1WfAXargYTBpdEN++i7i5vY0IiZlC752bqZjWVTG3LIB
aXNhCQGHw0O+48mijYUskhUSNsCG0Lo2SvIEGxVZBYFIoXmBEwh6VhGJtyOf12OEpdVUIv+k+qn/
6feyKo3MNkkJgeiybH6lhW4/44JZGAZwHzuRids8CQcucACaJDS42NSZUNaYvH80LFaeLi0owhTP
KyTKodp5D+4AhKLeuD0w3vHfHFaXBz79VPjwkgYKF1PpdpFugCCqgMunKLdBkxXA6lwNcJPY80LY
9JsztvPe6AEoErTtRHIJubPBN4pqLJ2Wbr26lE42WZoRmOuyzWhzB7TlUD+NC6G5IatntV5K7bdI
zi1q9V278/xiv/6k3XQLRg9Wzp9jmhmhglPAT6x+LX9qG2oPx8/7jOd7I0nIaswKniqnXXMUKPnu
iWi0KBw41rsxois/CckAKyy9DnjG/b1N42O5qRpOnIl5KEqVnee9HL67yuo7zHEq4RFR3ZAawAq/
0nPA5ne1JfhZriMnMvhohcO+uCtYdNnDvSXvhJEgPRPa/3ByG856pQZisYPz9Lfh7maZTG/g0lEM
m9fUAkppz4EFaqtGwk00Kp76vSyBstp+SU9IBUVlkiosZ7bjSCT2+m5ywFF2y9sAYE5Sq/fBGg6M
ao6yXXTEo/tP7dNKd49gu79xHsoRL+CeZgT54lkVoAcT0CyapezwUDU89o4P6P+Mo4Fgt8dvLIqZ
FrTbHEJyDhT+26IGrFCJyyilUimKgJDQDtA0OB4FzgAFOZ0a80OKogVDcnAzI3CAr/JfzTAb5v89
WaQRHEiUeQaOa1LcJ+SYN7b97DKZQJDbBX9Q8WqVUKW2w3WpDf5G6S5PdlCBpi1p8CtN2qzbDxrK
3hdZbgcOm5Yr4MN5j+BxL4GGGC300R1UPrKFtjcKEX04Z72YLClDoSIEQkqgbDpzAKmHtO3cU/Ep
SqBYiVVRlLHH1Dlq14E11t46Q+lbksu7ETMrnoF5UMqZ13d7zHaKIz5MneOU64gaVxY9GPHJUn0Z
u1W+5efDhrIXe3mcOKLgSVc1ALM8X8grD5VOR/KyVNQhbL+2tGYB0LGCnrurDaMOVITodwh7mMxr
o4ZkLWOeMWFLxHWmNIqjKFIbtn58GzO2tOqja9i9yELNeWQruoYhM4IuFmIkB9cxjFs7AEJsaO0S
UcECjdQCIdu12SlrbE+kI5lNa44sS9FMWf/aMbecOnpkQ5HqRKooSlrIzreLib5iXzOFO57qzVOl
XcfK4Dg8pdhWfm9A5lz0R0XjhRDeqboaH72Poe/zaNRqmAfoqRFgUY4ce5WMqtRzW1mRK51kJI1k
EqWnPX8JFgEEKDEUwdaRmw6uYocXpHJkf9lGHqzYei4Tgg+HV5T+EPF2F6vI84nJd/bvGQZfQzqP
6QgkJlSJFEuKmQE47gJwFnNXyqwOcrrQFXDA+B0zJJW+WvqpbQoRh3iKRArXOSUaH+jAfCbAyerI
LSpssk5WcHk7npACmrl8bdSEW2rGlIGzreU8LCDj3vgUMkWdUtPvHw5zh4slF4IsvV2A+Fj863B6
f7nEdtgji7iZ5J+jKUz/VFza1bBynnsFYxoho++dh1dWtbK9jdTKIF0S8DMrZWn703WMGDPQrXc0
qsCjUbl10o6/ukO8/rhgI7BSlsZsyEMtSwWGxOFXxatXAhgvD7skjW4TVQMNLukEkQAWNxMSjG72
0BuW31euCh1eGeWw0+Je1+s04NkosaSdz8CTcoPbOMQM4jFamhQab4M/nWstsoCus3YUo+EIM8Om
kSV1UzhzxRwJaDkAkpPRNytBS6S6NetX1Dd8QhBf9Opip+W5c3LtSYVlZ3as/crbYeRwedySTY+Y
yU7kvzxriR4RFbGo9mAEguZYgsTKuCX6HHu/OmrcBGfaJjWBrhhR0GT29y0YAQrlc83RgLl905tZ
49HpbezGNe/bzF4w6Eg99Qub2eqOmuDOXmZdXqKdaLZ0dL/PPoBtlncPDvVKM+ua+9eHzDrMIJjy
b/13T+jObV9eOdnQVq1dJ1ccyIV5ApCyCjTa7RPNzBKVVXFPhM1EQPtspX4IHw4ed8sGsQjsdWQx
rRG9IHegiPO8KfbprdsYJ9B1OSiUkENgSyafwn59SdgVDlGQt7YK6YdSSVWfDQKa21aiEj15pETD
Gfm338jZ0DYlRhNS/MzVJPOJLeuSFdASJhQoq4VgUqFcOyV11asLN11OmdLdFQ8phWgWaZPD9JdA
aYg61M8SgBA9FxFuzEso8sChtriLyTxh7++tUnWXV8Dftr12RkCr/bZQOncvPgK6U47moW9Q9RTe
eRs+EAaM7oKF5ZJAGebu807+w7E1CLzthBGXaLGB8IBafl2QTKNGdAdvL3MRl0NeINyDI9wbV2re
UkOwAkXxZLyzo+0Es7f60ttlla5OTEbAUCRu8Zf/bkJTwYajw4JczK4/QNkBufhaVi2Yi4fc643o
DvNmp33q9+RE55yayzqGwwdkY6J8BOTMHLBUjCnh85/fdv0rkD3Ep2229NrLZYaLFjV9Nt8ejpba
eAEwAzCLedpwtKdawVRK81oxaKNwraEy5AUiCEgDaKwkG1vNkc1CF7xPYapAqOQeBLudOcPCc/WN
FfX2LcKnxqvFbTWYz8zeL3z6D8gLvv7FhMT5GZ1YlWYs4KW32QGN7Ja1o3A1HWVGiDkLojNsXjMI
SDsRm4OlDYQMNMiXRNFYEMwhzI8mdESw64hPnB+3Bcd3KlDsx6MmMVobi12ZGp2u87klbbjUxjPG
qAQt03oQNwvRqh+nC/fSJTICzTVjjB12KTts1eeP/CatuCihMQurbNEPCLr6Mz36nKC+hHhyzXDA
PocwSljwG4LxNa6wDBsFgrvXr9RJn9u2pW7SWmH/9Nf0w7zt3Zj6LasAqe33eX1z58SVmrNNSz5a
Rq1isyLsejZM9quM4tISNgrjQzNkOwM+OsOOGYuUFUY+0RU3FYI7jPs2LkBCZoUWjkvw16eFug+a
zp39MC7iASKxI0FRpdH93xNotvBMu4ul4TvI5VDoht4x7I7IhApwakswRdJI4m4MkQ674lu9kkIR
jwK9fpCd2HIm4hsKL/t0O3RvfKFhQrJy0jym26B5P0wLMAidLlzBdz7Cjgp9m5OVhjNuslDjWw31
gDmqjWahEIirKZ60UpdaeXXPduxVWUKaYJIkOibG9H8Hyk2D62/XvHPn0HFpm0EKLHETxDsrlnk4
VIegfQpX0nMgSFIwWQLIBrV5u9SM0BDdlJShn7wiR0/YOd6B/ihFhW5PwP8vm4BD4133FsHo5AO5
1lhEGO+0jgpyPVZEU2s+QF7qYzVpykl8RLCuwg4iOeR4pWeeaB7xeYP9dprTtIRuIu8LXhlDOgVt
HtlIWiFLl1tl4WiWRrLiBd63v/r9wB/YlHnhsH3bplVrk5/WPvNc3qhmIx1OK4H9sD0V4cOfyBke
CdbRpr3EcWmur+uI0W6f6RoRzGWWD+zHVBFLEwjM/Y3lZvkWdcqxJh80iQwXyw90MkpYy2oESbQc
bz+vofhzNXswQl+V1qu7KaRCM8TikHczNrSroh/t5bFYQaWkyfr5Xf6ELhtThokz8WYliMwHnvuR
Z+PwgN99Qqo2YF2zLk2tYWT5vZLCgBi39NEaEloOPUZB/k0OoC+hwEG5kluveJj22TV+kIMBswuC
zM0z05kzbtAbHGezCC8ETnvtGjVYh2YW1L9Hc9HuMD2O/6ZDwxK8geYT1z5mju91n1luCA2LR/+C
kw2/XlanuK3v+kUzlcxxx340K6tm0e9phGNsbgTqJq6YGfBC+WtX2DUDyVIEHgrE5EICW03B6FXC
DmYtLFf8pmFuvtqGt69adm16+Ad0D78POak+sXA+DSfrEjQhD48t2bxIXSqQA9FfukfD7L+MVI75
prc21bRbBc+PvYGX2JIMSzCqx57S0lBh4k7+Keh1uxW2LF17Wp74GfHsnbraQPqc6xCUAk4yzggp
y4Za9/hkOjmy+VilNB+o18kbvBAS2Kon8sJ8foeA2HHRzVTancZEgr9V6oChL3s7tf+YqWWW7APm
XMwlp+a/ID5W+4Msc+8fn7wd5RGaMx+VVlKq3NzdM4183poecmYIATwotZBJwOh8DKTGpzvFmdGC
YQYvU7Srg4yByTMGGzOnx4tXaFGZGnvXqytSZa+WgMnjYLQddu6AsCugvbuhVM4Viwvgq4ah9Zqp
YvqE9pbn6fL7aFHBike4l/bP+WVUH4bBOXm1Zgqf+wumBDcDvAxK5Dz+cQ54nKpoq0V6RwCnr+6N
yb0D8n5lf+rGpMyyTMvPpqTl2rgz398lHdsJce0u35/1d/mM7fCfxCyGhBNmjY8ILUdd7t1oPKFe
LYQ8v1oFSH79pIyw+yjUVxPSPnF2JyQ6EkBnv+07wz5J7R6vvykMnypySEeffUhssRlU1/b0KsZ6
+L7tmp4ixfYX3vC3o44in6XFvOYKEAyK34JcSplDojkFagzm6c6vcrIQ1EaQjaUeenJzl8ey2lYN
hzkbE7RExnCmL8iSqHCqGozVSEkFSdxpjeEHerTH7MjsQRy1bwsprGH3+6/+OXAVwbSWhjOO5jV0
A9wKaPNf76jSy6DNFvBV6BwegzKPeqS9flvgiJd4llMRR5/loGVBHq9/CM+LCnrxS2dpdwz7xRgv
TaN6mE3yglbYE7WfLSMlTmI6iOHZiS0qVl6nCJ7a+3kOf7N1LwZ4AqnHErMhsl+o6etzuFarX5/4
Vq6EHiDGtZlS/hgBpJ2NLUE9B5Kj6lyKpWDPp8sOuHfUio4jA6JcfjplJ4n2wN39CqxHR6SVylFg
onahsyWVmkCTelalgrNDFYbnINrZJoyu8CklSbFLHF4jj+Lq0sXPZW0K54q0yukumlDJBz6oicxv
pSpQxE0Sf135gGe6Gz0WQ+awL3JfILOXNZn0ESPnFOaObonMJ4E2eaw6C0jhdeNJnozLSVhRb6Lu
+XhZ+PYITlgdaOlBNtxrWYWkcQ9W2GJ0gCQ6W+bb89v+uZd8cHpQTYhLl/h+jAQ47jcZ8uVnIBkx
xnIJX9m9YaxD76/9G3vfnvuut3Xr5mkFgXUFKyvyRU7KsPjjPh+2YWY7vhuvq1QzF3rctqf/yjm5
irxNUjQqsiLkuza+im4iaZ/4Ydz3/8bkZyQ0c1F0uYbpzXJlH8S/CWMlI7grKOyy6GUOBMc9v28C
l/kl/1cQyNMDRKWryCnMvd3vk4omFeGuS4UiDDh9d7K/D6cQEmcdlAf9B0Dm08kaSms9RUaGYNCY
dNocOEE/f2x5dRk9KChfX6zHBtbXydauDL+RtyWFdRMG7GC8+VVF5vOVn8tUXDYMDOlAZCwkqOHO
VfmcSSM8yPoR2U67M5v2gVVrXkSHrixqBVpDDo7eDb+aiq3pAaEgP8dzssoNEe6mQBKV9EkklpgQ
HwaQ1kIpcB47GZw+Yn94TAmgTtJFkBjBr7XVicqvlatMhLAR33maci9MQx/pxMy9VOFnsu4CkZrv
CbYo0lbGAIFzU2FFBtQnimkJ18UgaFbum2z1Og6k199pQgvqIt3/egfEVsyvim2SYPwbbG9HnAKX
rhYtIFHgMIGCAGPbOWGZPpci9qGzVTIjnRTAJzpBqaYQ08BNeCRQgTeWC9b7iYjiHHn96ineVwkx
Lq3l1y0Tyw8UWsvA06S+jxmc5kjAplgvxtOAK/+xHhBzC3XlJZyPeSOlHZfK73A9T8lUMZFIgRK6
NV48+B6dvpcszgm8ZzmlA/WAScPn/kUGWofuhWgbMqmDhFJad2Xk9Io9ndvAPC/DljKu9JUzWuBA
Jp9MPx4p+EVsnKG/BwJSOaN9dXr7nglHCTKITHBxxYi9sYlCtieX794YHKFLGCuOHQfydcjAJ8Cn
a0DO+lzLxJI9ZpFE1x7ITnIpUzK1/sjv2VA6XzvHJfLI7hESEdBCbEcnM1noK+D7qKLf1+w4jf3c
j4yx/XAcfxtTHR0yeLK17yyTG4XYY7VKpfsx0bitKy/Sqk/GpI+HkFIQO/vP4fvF736Qz2rDbI85
RALaW8+9kGFUdttILY2kWsgRG1wtDGvK9FGvbSRFLbvOQjcs7VrzO/vEjlBqdQP+Baj3Bnq9nIfc
MxpLutsWooy/MVtmQq+ehh+ua+7zkEw7AjXGLQAVT1E1a6aQeZdwy3zt9bZA4d1h0T+U2U3tXaiD
L0Eg6n45BPGR/aplZeDdkyQUSLIZ0jdaIe+PD1qgaBsJfJZr089p7ub5+0rdeovDKXkXi9HvXd3B
9+M9xvXCCFSa94ejjS+PmbYdNq5WeDL23ka2tF6s+ZmQU4r1E+/1FB5Qt4JeLdbtTAmjjq1V49HY
P+lfcwpvQHHZO5YU0+w94M1sE88il6P+zb8wj6e0jOF49JnlbbI6I7SWgN5dEgTX22CFR8JC5Yuc
UyoD4dGh/T6uf3hBav5pJfhUbeG0K5/SLRY66J3t3XjXmkOb1odG6o7mSIotkcbcgIGKc+ayZRMR
ueASGoer6ze8RDbqLsT09SutGatpHCtD6Oaf8XIQXgiS8WnCCwwYA+APJHY4iirqOrBXBgujaGrT
QEI3nC1+7dDNC+gYi1QtlawYYGU+kiMhFewt/m8iaJez9aVg/wKBqgCGWjS4pJjeEidXwYeqrKBJ
8bKweHiMI2Ult/kcVh8CogjwvrI/J0G7GbBHgZ8MSJ9LcADqkYpntQsYNJHbvtDYuFtR1q8bQdb+
iH1uC7XPElUaLhCYxWmjLaYoDd0sTo/fbCG9aazkAx9uVsJfhSk9H2FQwz4W232BZo5yhv7UaO0M
jotLMPIQ9PNgi3c0PBPXfYDAi7WKP1TZOv7+gL9DgmGVzyKIXpKAXn65LzFG3OROzv/EiW9um5UV
FJcHhBirfJ4ODMppwBGW7IqaBE6FelS5squOqTmgOK9ooW767puSvpweCQSlB27FWjFhwP+PCSTl
9CTiO1ROIQg6T8/BLhUF5qW8vJIcnFtyXkrMBESK1X0A+sUYRs8D2uihkAHWXCBfqOXWnQ+hn26+
Rm7g1lp7/QDkVrIdjpGacBZnS8fruqgeQAfmnNjfDlHBG4Px0GAeZQmfF6NpeQaqf6Vo1kKnLewM
cidskRFSnEySs/kzmW0pmy2wWcKvCWg5+Vo5cyNt9s9QJwUqXYxfo+gcrKn5a5vmsNLCRY3F7c97
6Ftotv/rKLoyuidaEOtyHdWvBAAa/l4k71rW22A9Tptug0m7RKyV4idMlm1KJ2ruGIWhopmXpaR1
5Ip0Sh20+8uO38NZxeZT7MHcRZuiDqCj4XemfMryZVRZBTJHGt4K20Tf/O8jCoPmpJJRrqTgSPpu
JMAXB9pEQ1Mj/0b7kvpq7X3jcfjosa+I7z0QosLm7wSBmUjT9oRtKYrKe6me9epeR71ri0mGEk2o
gxTRNRFMNjZDuXGClHi2vhs7eQVPSbiV+6GjMZ1n1NBY4zRVLODhWUHzF6+ZeA8Zl0Br17ELHyAD
ROZA6/NN6y45UpN1euYT/EZ9SsqI3gLwpyWIYYI1SQYjl8ZDrV22+SoGyyzdUrS+tSABL5bcWiZt
aqUYbvaQHHY1m9PNrGG+8BQtgsnoTKM/AcNId/oRuHMsGAWUjyChz2DRme/Be7axcckCSDR0+GaZ
b7LFLgSxGzjjSPMAVIQ9ZqJQ9bv7vvk+vN/M+jRgLaN67KAU8KOOEsdOY2x8ciS12baY3DgE/A1f
4Y/Yk08hVub3/QgD21iXVs2ehgkZogzBEi9bue/LV5VIii5bW6WfEOPBwhmSqLKqlT/G1G5itC7Z
0I0lGu/pvFnESDmHjZqoF5f/AftNoFAptL5qLO6v93Nhln0A0EzJzYd1wraXadxrDM2ypgkaouJq
ZlsLRgYohUUu86falee9JviJsPUbYXpv7J/+Jvk+fqYwwKkZLD9PO8lJNVKYRlgYxTRnrkfae6pG
3uFmvFVlZK5iRF2xR4OPJ/I6cx8atp+RwG9PuGdcC/vkzYghNQxgYlscxzhW3YdKYWariFsi+nbh
0CZ+AUxf2pO9CIAD7yUB6HKCcWRcJ+xDWAEfiyQd+YeUzPUCeB4FCfpos2MF5iP4HTnxEBoAI2RV
QdaQyhCuL+6pWCieqECZHqhl8steBnJt4b2zgEzPPoJaFQS7lSVzyXDACYLYMS7kZ/Vx84Lhwx39
zirXuDB7SUDDE1rPIS3lR/rqxNcou4YePHGt3dLd+NTKTnToGO43o5m4zNlBcPSAA9ORLp/uphRV
i6pTaZD5gRUlpKFYdQpSumhECoOwDxLg9LDowMZzTh7hrIfaofQxmuGpV8JkKZzsKjr6Zj9oXlrc
+3AlhzeCR+16xJt6qqOKZmB44QZbZVX1wcmveXCv60zZZZ1y857X6wP7NSzabFzbfINDAbqHH+gb
K6158lMELcg78ves1kYXRiCCoQv5jvOsn7mJyjsC7zXCfQRyvU4HoV19tcsQ4bwvCJXX0LBI8E1A
n+l/gSMInaItuEiEBi8TlvSvxb+o7Ap4bYpydCZju13yfCaHtVr2YybcJhxhjFDDEcgG3TPhNTQt
gCM6lJvhdHQasor4BBcQcFHQtQsiujBs/6FpUyXbLqmiXOkjZvrn1yvwsqyG8V9C+7YfvWRCGwsx
JXGuvskWSsAql0/8wY4HfK6Sh3Z74jmyMULFkv54N3utevNw1uhit4Jb51AZvbE0EF0eE/AeDZuR
BrKi2gno5CLkMKprvxLozOj7qLnDnDCFmCBDIz3E9QwbptyayxVdnqJntoKHhI3OPX4GP8E/F2yf
Is4TqVCW0kuHTAcVf1ju7enSfiqg/Zlo5CFmZ2oao9x6pNQHFyNwQ/TJvmh9Z3fTy6kQ+uoaoS5U
NQ+CS8MXZ6BRpw62j6aWm/nDnVToiVmQkpwZC4qB+inFaLWE1umkb2taNQmzlaL8HonEchQO8E/t
CjAmNNk9TBYqeuUYj0IdLiC78q5WJjv3KPNN2sM1bvdJAZDwB/aHSi3LOCP2Y7wll3t5iDtKottT
6XNpOkEvwYbCSXwV1AY9pQX6RJz6rlBSxYQYU/Q+FgMKPTc7xtRV5afGsJFak0ZOZv9LbN2UrKmx
KSs+tcJhjTLla87D+jdYhj6nWDgb8/fUbq+hdOWmlHBSNE/XsTQgZv/Q85ZtuRf5k62lsQSgxPjJ
Tx4opwiY3vXsPp+Afeva7apeixMXyiAYrDAgiLDJYwacJZXzgnEXwlEIwD7lGA/GXsXmw6bxHCeY
mb1eaBhf8DAB0g8kKwxbp9vcxwK4MK0fLkAWECl6k3Mels7Inww779mpoWMia4p6I22k0zkadBYz
5j26t4DTMbwo4/djOAxd3uHT/bhimrXSdvGOeEo35MvipKqw4wd4P9xF4uNHvgf088u47BTtZHlj
RwWi4Pz78ZaoXVNsKPH5VNtQFIT90Z1uFC1lq4nCQa1B+e7ZYccDefTQVCeifa1nHF+7bWMaSMCu
ti5mjltGGNBFjLvqw1aP7ntlYAfP/hPxYD6gIigCw0ZbD+rWI3gWA1/9PtASzebIFCCtew+unsQW
Ybxwt1LHwfp1lwYGKVTNZaa+hXx7lJakR85lEyXfGj0iRrOwi1xUrfGsE/0ywPGdKXhHU8l9Z54C
i5KKsskEIgVjvymNlAczYsfcf7SyYSnQ0y9dRRj6Q5LNBzEkVKXBy5wFX/d9XszP7kM4KU5wAJkd
SHunj5cK/kkNOkibda/GYTdAWlbFJsiGVL0TdR8CwPr2aNMgkZi66HSRhjVDnUK04OU+shN48rHD
cZAObpwZaJqOUnt3cIRxF2sg/YmpbMemEzUXk/4XL/3qFU3tbkfHYZeLkgxr6jlxqKE43qWQHXuB
/2NQ4elcg2enrJME/R2v0cF55RfHy0EhvmTs+BJkG6ASGA4b80OpTfRMDqLonJ/ghvHI7dtsk7Qi
c5C69JEyeZqQzZ5GXrizGXX2BCbmuD3ftCWE2jYLX4J0GFvXg4Dbc5A/fqI7ujbivpaHBZUsEa6m
a8SZdxgC5RAVxKNaVIMVqN2ROc1Xnm8UDO9ctc6VNfnh8TeCZAHxLKECKJkcSHEuVpLwLohyhqJp
RTYYEnusASAGyYMsEKbq1TgEf+GC6RhKuXPkfNfkQ61WItWB7hlPdhjqFP4Iq/o3wJRgLQ3wR76z
PUF/i7c7DNNTT38cRj02GHoBTywl4H5fM44/42RaCd1pCoEG3v7ulq/HyxPh396CW9RjCvkmMsZo
Jgbb7AbfPTTza2sELT4E0CfW4iarwx2LVh0NtbNE9ZjuY/xCJucHO81WCWidQn07AbRpLOnTE1gM
4oO2kyySH7N8r00w6uthBvJyCa06dQQWH840OKcLO/H4smYKmVpNhmmzZzHIo4yO1kHci0Mo9mpg
WeI7CFB/ER2IwB51njW9hI1AYGRMMzzW7nXM+qhGy7G0PAoXGMvAgnjXiPCb+DZf
`protect end_protected
