-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
h0TZ5iABhYefvki2faYctWwLudkvAaZRFkdfpTXL2qPlE806pkhGUm4eC685sDZa
2PzHTg+gzA6OiyQGBSAX5mr9r56KJ47ddkN2QeBFSK14YcbPgK21PBXHTXqBRdny
oLu3vcKNEsaWNyxbpDxFVgrcEw8Sg/16zdAHOWOStIw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5041)

`protect DATA_BLOCK
c+IvMT76CQwAwnvFmRfeWnFiPGylcoegWNPV26I9UTQ7E72QKXOVbaj5kAuP7Fnw
cIFx8PCWLAFhV6yH3o27eRAuhO4GvDbDz5BOm9jQcS7z/tGbnx6SSFBMgWN4zqUW
C56PhkrAloSU6gFLmDppUPlHzYqgpct4IOLGlW7ZyasEd9KrkPuw5Ijb/i/bIVuM
wSEYqc3iykyv5ud01u9r6IVNUg53mvRoWZwcS7kZ5paT3U8EkVhYJ4adTw0Wr3QI
J4k8CfwZkj1D/2XzCCx8yH7nwJvVjIvXnyBItyH2bdURXY31KR3GEoP8VKnw2COo
baijXupK68dPJaHyEDOlfmfNLysUijE37lJfcZA3Nr66dNrfSMm5Kxn7FrQ96ewi
yttYcshoE6pX4Mmx26DPEPks/AZJEkxbEMloskPgCt5CBMRD3rCimVC/JCr6T+am
Dt5w5KKBOOe8HB2kROLibkONFaf8PZUyImWoFzxFt26KgatqEo3bGsssquw/8O7Q
iXFPFGVilAJSHZaqsygSNYA1thMJVpHsZkujxD5MAkgcJ5PI97dNePQe3gPv3RpX
2esttgnzHcKCD7uF6GH8CblDlGS/nBxNlgoEBJNc3ss+pcb450IqHqjnuBDYPtSn
XZKlnj2KzwB5nTIfgNzx3Y1LT5qS48WpCxvn+UPB948rpqjmadym+jku9HFhCGnp
4uS1PrF98kynkrkUG+FdYCmaIgCAGUyk/r3UcySHtdupUCZDM1tJY1ESCyUjdxX7
8wNqazPyZdtWHEEa8S36bf/soCLdQFtTIr/Qsi+ad/PfESGOtlN1W4pjISe0GqS5
GLvSPLck2XgeoGj80sjiScycVORE24HwM93ObwH6WunSqgbc8bKSydq3CHGpNfKH
feZG6MRGIgDe9oPRsRENMju1AhLlIzC5NUOo2cB3CymOmdv6FHPHJlEz+1N5M2Bv
dKerBPC5dyJjV1X0fFc2TvcgS9HffN6mDy1WKJhSzEz3RPChLkFw0wHna/fZ0LS8
sa3usrpAGSl8/vKlsjJReLnMmkEIxwPFCp/wm9Owin7/Vk2Si8sJ+C2FuORCVZnM
w/3ruzJ6B5SHygok5A3+sbn+EK/uQ/anrSogPxNjbdYo8I1HJo/Mn7lvGyLSFj0k
rFBV5Ia9rZGbdWw1FMJ1hoQpqgyD9FOnH1iqxxUqHg1x6qBVqF8jHtWXe1H/l7Ms
cACmuFXGQFdx9TnPNqpCpMuIP1hHAbY0DyO9uOXbpSLwEZZ9Nj+9TWyLG6IHj5So
Npc1f6pupBRZUI6zi6Cy2hqw/XKsJWe6HdsZFUFkveqLFXD/SQJsAmDbLuWkCisz
jA8ZodOanQ22Y3B93MS6NgcW9dwaX/OKhWq9comWwnBivvJJhoNGRFX42+ai4Da4
V2p3mI41TBe/b40wC+gq5EUhrPZdmnmjwDZ02c9+eLSLwnWoI2YPHPf/XQrYrBow
mzqHwyAqjiSNO719SPRFJGZib3SBlkyFJFTijmwt3eLYKwa+FmL0L0LKKNM1gvxO
yMtvXPsASCzGVwE3cm8J/iYASiXZ5svsWz4z49c99wp76Ixdw+pJm712EeABAdUV
20gmcTZBA64cdjOpQcGxJvD41Jjevm/qpxNd6aKV28gymggWrAks2gDaTfUknGD3
BOA03tf9v4MZ/WOlni5QVfwq7TXZr5OySpJuA1tYB89nFHSN6H4WsRuA9M0hTjtV
vQYv10bk1CfT641ByhCnRmoUiPkgIDrelCxc0YiePpKQcB56hhzv30Pcw5WBPA1k
NOzbA/N8Edsq3qWmtLLzg63Y46DVI9fTnN7MoXyVMujESQwssxhixPP3+IRvwgM6
jTF+yPJ4joboAFhj9u2wWpvFVjqjPLdaVBgZGRdGopA3RhHA/9zKaYc4sjnCvpws
ZdmvDiq8PeTw3xiDPeIfFlsQSUXPv0xKETCnveUCQWRbSXl9f8tV9jbhWy6T6AdK
K2fWGR6MagElkZ8WH8d9yAQcEQWVUKTQH9yVg8Ypo+47H9MhOtFEIlqbF9ya0wfk
cYhAJ8goALuW+DLVMJrHfSPI0ddvhgJd4+snogfdphzB42K2SksvI0iQ5vYiQpyj
cY7uBZPvzjfCYXnXdYjbiI3L6Aw9VGcIm9gw1iympxSpqjsCKir8ofD7WX34CtUO
Hxzf0zXFT5cDxI/GbkJJB40U9lnWtQOFpZGKXVcKjCtU6c/ZwV/F7PGFQtZ4nYeq
6UhEUMM10RG9uSPJrOXQ8j9UEfTHZjBtHaCvWoHahuZOAdsfzkSXzWPdJRSyvIQk
rXZlc6nvY/F7OeJPscdclkuQOikb+cGoIAWY8A8uy/XScMQOTZzQPMaq2KIjoaeS
H9oeVjhN+z71xnXs/6kAf2GQZvs3qI38okkMtmoHUIS+xbmVSUqCKuOFEFQ7OUPp
2j2odHwd7mdJ5TW5t+UlhWgH3TdNUI13SzZxXK6mTpZtW0ueLk251hHEeDCgdojU
FPlLxQBhuslX1UAuG1LEAgLN9Z8Iv1MAwmZL5YqkRSZCgtSToUgN9GgDTHzHdsMd
hcCBcq5R4xxCY6pm0BLN1b43xgGLGF2ltNE3sFj7aVJ8Ksg7AxIqT4UMzfoYfZWa
BY8Ltlmvd8wo/LcwXa/GL92YEZvN3cJEEJQKaTNKWG8u7QGbflos+up1pUANiQs8
WVU9CgVGWebzidNLLsYcQzu/Pi8I5y+hpG1saVMh3JHeXa9NCILxM4BSK+EbUyMR
mHFHD9L7cdJyMmbpVOo49Dr3je/6lVJ2d4C/MhDxm6VzhB5sTZEUA1sCP+ya3EfB
z+TcgPj473eGPU8FrWcOcERzrrgs90ynpiJjCjA7G5rtf74vkf4bFJ8oAAlD6Usb
+KCOvADr1DGetY19qzjyM/WP0pElWYz3mEbZlSzroIe9EA/WFqKX/GEiFIXZG3ss
opJB1CBxvfCpPnuZdvkSxtsdxw+O2Kh1sl8cFI6xRG3mhIQ2u9MIudRLDPWp1S7u
kZtPn9g1s4sCvBQbQmnecd9riVwEbcNQJ8K4YN/ODeJqj84JuACpfyLqAkTHmQGN
iZoedRPSvwhaj2fqGpCQj7+4Vz5fQIQnzqtelKKcgpVdWUYdG7HmncMIzRvvjbfQ
ZsxZnkqORJgQkidRprRoUC4bAFT5y+NMlwEOcBEom9NqP/qhG5dWLZMQwUNs0eOh
TLoO+47ZC1xWHkRw3fGprHfhCIHcYj8LIKuaD22bRjDMGMb4msmv5nrvfjssbK/t
gY1dO86/HqcdiCqRM04picf62JXW1PzeEyzhdVUa3sp3f/a3/jt5IkPT8fNiXM5G
uaCk1BjL7/3hksx3sQegi0MkKqzNzaU/1VBuhTeZDliO16meqOYEAoBpjCNB5Q95
1BfGlM0nu33XnXpQfk1kh6zgJCSdhBkYDndqM2AC22Z1XAPiJ9wOHNwFQ6E3+PCH
hhmPlJTHHCm1avRQ05XdCXlp6dPyjI1BPyiAji5W83ZMGzLAZImyMPnTUZqVnaGN
h1UklMWTuyYQzV2PrVmH6hFsyn8V9ot1IzdCrp6ysDivTl2QGsZy9mA9hpcwSnG+
d48ualZI2Yb0GoL+ShGJDb/xPxSqvz0iuWWxAmlDzosDtTEyT7JWQ95NpIeP9Vb2
afCRJw2D88A+RI5ZdEzZXdKy1gs1mBKOmEL/At+0CXfLAIBkS0VNdDDMLIBo1rBo
mhxVSKhowIMqYQIXUsggKtUsfcSCMSCT0Ygl9Nk3ng5+eXsETqlsNki2Cp1rICzz
KJu6ZWHbxPQzmPnKfRmGPp/YFuJJCmnzaanw9+ZcPJ46ptyIEKIKCS/7vaGo3YVf
jSZcZThjDMYEweWrpat2y6kFFIP4ewuDvzD8fBIecY2pNtZ4OxRlbe/tkGfvsLPj
KmaC91tVzwKzAgZRA2LIXQDnSoiGxrd0bM1E+C78I2rxwcTvWRoCYPS649hM5VvZ
/J/e7so6QAoVlIDQ9eT6Bg1tOSfm+d5yPcUjA5ZUEkTQ5kwTwi86VHk50B4udQus
OSzNFSqXSYlRTqu5JKue2HpTTxyDf+evRxz8j6lOG/GM01dEPRgLOUvyGw2bYsCi
dFuht/Y4YKxYOPa1M9zMZCgmyxlC2wVxNci/mld7Fg7btwS+gZVIfhemC4aiw6HB
KTdU09h98TI/ptvbQyfPYFJeOwfcrnuP5gOSs8j2LWHp/DqGaa51Pu19HXH45O5l
Zbc/tYaL85PeGJOsT68DPSOtA+lsz3vmFSzj1RX/GoMIMsada83jsTd2F9wHhwVI
XWOuRz+6ijQcAa7hRcDITSDbRNKfve+mojLhzXkSGWqQh3LX2sZ4evNospEdEAk2
L3cTUrDTFMXOTZunZrx8GpCdrkCc9847xhsLDpi9TB1yDyoypc18e7/TOWfgvsj9
HBMvN5m/PWcYGQGQC/gzbdDn60x4NewJFafRP12x1RSIf9XDVP9DD7l+/WxcGiCZ
7jnf4FvQVx8D7zv72W3hITMo0agWyeWnC9OhlAC4CbljlUATuQJbNDViRJ7kk3Zb
X4ZUAHynobWGFCr919YVX3d1boyifR2nSR/t4NR19sKcyjI6nlgjPV3dcK4UUHvg
j2PQIqiWiJSjaB3oiSoDjMMNMtFwuZFu5kPATXf6EP8jYx32zzRGTmkGUeQDqvE8
0b2vX+Mho0hG3YwsccXfnxQzICbGhmFZjNpuZ62I4cAKz/Pb4136ddv6LBtammUx
yRPENXCfZIXukqqItdxkqBvY3Updjw7XqnBcUh5OxBLdtrLIrZ5uUkF6aHuXK7MA
WQ+XIGxFVxg0XpuUfVqfPtLMtz3exutMWt7ebdhlAGnSJMYcECpsFJhL84kBhVxi
YKaXOKSVMKI4ZNEUSMEpFrqqtoaORwYRsVY7JeUaTAnym2UHxwK1l2VUX1ErLrLz
WW3ZL+fwg+5YRToCoobVVKuoFxHL1C0hlqyQZLaEUs8OG+1ZlL2lCMLQBPdlHR2j
Tfry33Bygxg8xwV4NQ+wTl+pKsAfzC4leLHyV4pIjq8hWUrpHpY3j4YS8yK8wbi6
Zysm82ClekcWhzRjJOBBLXnf2pajCV7/FHZRRbulqBcOrajdzOqmW/badYS0twjr
wzSJ1p3A8en0Vt1j+poU9v1A93VAbwq7mEAGP/DFADsTnAtXeplgFsI0bLVyE2Jh
4OVwP0SFhPuD/7JyAhZCPjJu9y15ricXF2vJXaoBbDuvRRDKzw0qdJX+EgMu2iUz
J+yfhjrr5IZBT23btIwSw3III6B7XvWveK5YufwdbazGBV+qTxDmy2uPrWz9UH/y
IvZ2uur7Hb1aytQbdKAt5jjdV+g6E/dhoztP34RCwnlkN0qCouCjxDT7QMpxmRBS
9RfJGIl5XLnKYB4+R5oewrTmbPIcdoeckNP8EOH0KWdpC161VIvZ7pXNWPjY4H6M
mSi3WDooJW0fTo7Pxmht86DTT514B0dHSioGw6K3w2t8HfxwGI7nndKt2WKO+Yfx
WOSqo9+MzLmzfHqLfBG1G2kct5DQNe+0GXAcsqCcLk6XLsHM/v6bHw8wNKHQOS5b
r/ifYx2zYfb1kzn4cR77xNwCxSGC16X6UxCDDfQmiJWsblWmR1hS9qKv1HZEMVUS
/voWPfmuKBP/KWM0Tfc/dQjI1l5w6DqxwWGo54m+TxLQz8E8TmTHscVCQrPGxYSC
PUBY4cLo+mAySneAzODaIRfYBUF5BmfSuyT8VBJc7LC22mj9wVMoxN7aCoNkOaQL
jQpDFcVCwIyoOt7Y0y8xcEo+4MzFWKIQ1il0Ma6LkGXzVPqHYL9uvyly1LVH9OHk
xz8QTYY0jFoFxqdufW5PLRj2tT/Wg21f88XQA6wZoTwNvVpQgEP26bzLVuPNukPr
F3sUpEiWRbu6MHuhmk9+xBtAdLEn627TS84MeAzVIydBSQpYDHeDXBnlDUqThjHM
d1pWgDXLSGNOCuR0EtVBIJY+Xp6NAbglmhdlcO93rKEH6Fob78+zt6EGGgK4Hf0z
35J27RE9pcfFxM7AVwdFbl5g12qQhSizKbxwAlzuwzU5j60reo767BRP0tqiczlg
J007rweZyMcl8Tv/6uu6dL+j+s8c++W8jqgNEFwjm54Hvb3cFMisnI+7Gb6vnria
P/sJlKuIv7zoS2QH1TP7OUnqvAOjcauMd87bf38duL4S3ExVwXp9tVrNOgWIyy/6
IiZD3lHEbO1ELFm4acLMUn/9h97FhCPyUxYTervv4dAHYIYp5WW9LieH+ZNrSTZP
UypVPKCJRrtgQEKl+KskgDBPecFSELd5Q3dQTwzWzTikwnpyxw5HWjH4muTC9kbe
pXN1WrIgsNkqg4sWaR0qe2rW+XKRbTmxjNKLCtt/81nD62t/EVMFKIR0i8/X5x5b
0PMoZOtPg3fUTWQWmvapSDuiBNBKybKKhtl0FoGRESwKIJcANvxoTCoolIhkeG7m
cyxySETVPePz0UmeCdXAq5GB8dtABesBp1a2eJ/xmNTlnCGJOTekw8zPSSKOIQct
854SaP62oVsc8HrX0/OergQNtAFZjs6ybUo+nLvMHzbpo2b7PL5Mz+oCfFGCR0wG
3+5MIaWjuvxbJWRC9b8ru+SX0t7mdz6SyHDxS8HEXgSEItg3y8buxpOZUuycXEwZ
wU0pKinUPQapqKu9YNEHWKL8UnstOfZpHEjr7phyXIP7tRFKyCSE8PhL3PIdupv3
tkb/eStDpVquZxpAz0kvYzSa7vHEvnzT6Yg2PZ8tO7o=
`protect END_PROTECTED