-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
gEODrYnOXN2yxMG0F4wdrDP+1aHpSv/jaEAm3yPpWGgZMsQFIw2E9ztJXZ+rcnU1
smEE6mEEpYX/6s4cvuYaU1po18yLFLozP+kEqwmID2XCQb45L19l4mQHcDLeOcNf
O5jNTrpi286/rWUgEVEBXjNWRQdTMnWSpap2vSFz76g=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 6869)

`protect DATA_BLOCK
+Rezpqi13LsHXSKGdl6KtDMTQBgN99nedN73579vXwM2fKP/2qNf+c5xjxavMpHa
q5GKNTKY0g3va10LtUG0erldCgL3NnzsZZdtckzkMaKqBswIHbGnSfvMQTuHA93g
X9CIH68Y2aku2g0wcT6DRar4n8tKYKU68+VZ94YAg0z5/WNyouTYIAMBrTyIZhts
vl+P7xzO5oe+wmbPyNpXCip/R2uCR/PtPWU//jYkQCs/c3M5UkaK5dYkvq4ZM2K4
+IMI4nDj6OLSGVSIsoGMsVIhinW/945fmHSyuY1sa+/Pn7dEDKt1SSVxuQiypQfD
UxAJhuZFadGqdIjKZes00AXEoR+159K6/zivF/5HNSijltH0ib1/lGHEJHGpkD19
HdKJ668ficw4r6Cu4hBQBEHao6xA5OpGyIuE7u/d4vG4egpnJPm/A7SCpu/dlIH1
MWc8jJAXr/YIkOmriuIldHOLkKFLM/+AVDWnnZeMFwSzedOmVAwjMwK29RtVo6Jm
4nowBaY9Ff9JUJT0cGeV9dqXbGaH4M67wOg3A1n3c0pPrJwSaXLzF3yejTcuLjrW
IJMUVEV+O6UCXL6d08p/a6sVocRRJZmG8tyMVrIrceK0TsnPtwFfy3pV7rZcXhnX
+5RN9GdF0ivpeGmb8+AZOzCGy4JDuO2aaCtjpNFF1crQOiCIzKTjHyHznALe9WOu
Lzr3pBz9KEWv/BKIIpWlNwOi035asbr8WEzDFcxQ6Pt2ajhwzOIfWFrJ4xYhPgM9
j8rXKGyDv8flL5mTecF/KqE1pvBM9A1QeBgY6IZ9bgHofxnkZGAgJiuRNhGI3Xtb
CNo3icBYR4ODGyjgkKg5mS1Gq8XG+ZsS8vSLVuZC7sDmXOE98gWBGEhiOaVr7y8f
lunU8HmIrwl3sRfEg+VLGaDHpEgDmw4rjwoE4G/maxCTGlaTJBMkHH/TdGT2Hxl6
8NZTrlzjYfEOb0ReUxmvJCvxrebXSkyDwuLqPUPf/M51UnOcUOlnOgFJycT8T07M
YGVXGcK/X+9rJgo9jH+JQ18hXH7PqPqj7SZFtw7fBqt0e/PUUuuol6i6fEk9ymPb
nCNjWVlVzmmK75YqvS4/wl1m1IWoc6gsSlUL+B2zvk1DftEr5fKk7gDsD59RTolR
AXvnVsCkorREJ9rvwr+7KsK7yMjXVWd7c79n6jCp8rsR9oApgYtWQUyG+1XdUIKC
OjJah3iqSCIeA0DXDbaz1axAWxY7yOPQd5giba7HnrY7sW8eaNzvh8BXJ9pcKcDA
tFDRDOAgqI77+2FFHHy46G/Wg8axm5Zv32suo/PuAIOJSJN6Fc+6Ixr6PeqJDsae
ELGOb8ZlzhvW4NfK29QCHFk2jEFyNAAThqWDtzz1RhdX4YcE+MfhwfDAjdKLd2Hz
CuHpSF3KxPSm8PSWUXA8pcYr29LelfAab1dRn2PgHtEVP06bANfoRaWWkxuMXLlT
NrD/w/iJhUAaaDPz53ab2VselfPtTJDF/Idb2MqEqDEUYCUuwsDULy8c78tX5KG5
x0dMp02KQrPpp32bwNlEMTlbeYmoGvaoRciPtGCnRulcdjLZNyCD35odxE3u6PpA
e6pGtk6/z90iTTjGrEzcTAOQwCXfpyUZSimVBH0XQFYRgkymSeJS1Ysv3E8eFrMW
1ScoJQYBiGnbxUN321JIJv1Gb9jgFhgP26PUG5zkm+CLIn9l1fyQmxO4yjXbPTmF
g2MbH7IbFJLfDjmK8AuRKZs+Ha0Y0B0nOWS5IAYmMxfDLBU430oaquVk7PANhhd7
g+NIHCLX4UXXiVKDa99i+dxZlutkMthNVYp+d10aQu98bIXVarAWXCFHBEFlyCKs
mjhWfhGUbraEokXFV70ZZh6iptHYl1gINKATy8itxR2wA3krXKHGdKNL7ye4DT5f
sD36RH79qjyaq9iR1xpxbHFw9NBinvS3OB4+fcyT0nqME085eCLiRYhbYa5sT1Vm
cnhREab+3RUvXASkwOTTly2iD91o63Ybeg3MQ7PxJSa54MVGb3751I+CItKKMPwd
bqh1jtjXLkOyjAcJsvcbVeSUCYkMpAxC0ph9zE5cXFEA74KDaTt3kI7+RBtENJBU
++GJ/pdEqCqf3fg9YgxE2ROT2d8WkNaF+aZenLL2j47ElH71UVJbX9a2mWCugX8T
7SeDsr/9EUfbXsEKZwC0P6JYMIWdQN6Z5eVfVsJ8M8RWY+t++fbQJRwFbqAQ+E2S
F4UgNgxxfb2LcbnSPN+coqc3vI5d7qI2VxvqoATt3lOS2cvkfQqC0uWeIHF0jZ4K
VbY8gPcMS2BbA3oEvv2sKO29PrmPT9TEmUbI9eT8vIHTByXbFgL0wAhkYggAwSwG
AnIdJUNExxExwaMKEk1f+v9SqhVwJQmtDme6ZCrJOCq0Ee+4O/Qqg2+llCp87zgQ
jKjh5qCuE5Bd0WD7RvNGNb65iEH4d+4sTtptkz2FiAJI7PwX8u970bciNTatNaDU
ZnGH4zkbxS2DeRpFgSqIKAAFFT92YsYl/xRbo7jBqSfiGzII2ujJN0eLh3fs3MH5
yGbKwirxlO3RV+K1fLZLyeNFsVcWX4qBCcv/WnWS1Ur7BPfhN2O6yTdlsQuVhVBT
gLWDOBvobdsrIRUKGgxHpEQVgVo1NvkJZEYnPJ1OfEJDejSsgeCid634HkbzTLGt
RlM2YUAsdjZSewzoGPR0YsXn7menz2grw57sF3kUyu2NaJOwe4+pvBAoP+dhVuN6
2gYHJOo2jItWBvEhLavQIWYkced8isBftZHDr+8XXcFsTi5nrgqZMTAzsHpN2soN
4LyjwXl5Uuh89BrAnP1nKO4+dDS6eh1G4PCNkRspIRHKHMelhihH36vrmtiRpVPc
X8xAC/l/1Fe8E7TBRvMaBzISfD6aqWa0HT/T38qRaqt5pDEJUCiZkv9RRwqKKkxD
SDlWybRBfyTNEkg+uBURKjfaMs6bs5e7JHYGXb9fJ5AMCaZ16RDKoAU4I1B6Fkr6
2I/1sJxFZ/BWACA1UMUtsU8dlUwH63SgotJLlwXe4Yct/fUlsvUdKhmvL3d43Tq0
SPUued3vlYVQHTWfqCE3UuWGAI2MaMu/yReMPhPP4hsOoAwZ6sncTD2Be55hcU8G
qw6XQra8dI1Zu/h6Un0EMl2a0FRPx4CGTDlNzeZWrSrhRqjgX6Qlb7dIrWt0GlGS
nHyjGNsG1oqreCjbwV8vFIiASWHpFQ8Gimtv+Zy73bxWLmmQuobonaymt8LrPGxz
MqzVtks43nbFlocwrIpcIVs3GCA341kIs7YXT9nfY+L5WcsCHzMcIjBOO3hq5+FE
OFVXNVgRqRHK7FS/MyWuBnAEfqjMf5+q9QLlnQvOagKLk/mhep5vV5xvaqoiG7LV
h6VltHo3K+doV13We3FeFte4A+Ry4+9zS6sDDmh9XWk2Vp+xHkkacLx3vS34aGYU
UiNFWTt8CF03kM1/HirrmoJoSpVNMK7Z9KTRlIUbOl4FVn66fY0pc36k4zjgUdil
Jlc/D3yc7OhnaTGU1yETGYZW13P1s2wV+aH8bENXBpY+BBXF7ZIjCNJ90DfpSJr5
4folQFVT+pv8P6/IOqOeimAOFx1r3drNTumyFgcB5wKbSNAI2OZ+lDty20CAj66+
yYcPEcJEYj7FsuXsBbkK5X94KQQBHB0RSS/XARWUdweRcNWA5NgW4BmqyYmeUkdf
kqsU0C7vjX9RBH1D5b2GsgzAK7oiqDHtcJiwChVZyKG5/WICLlT60MLIEqXsvmNc
9qeHCu1gG51zz324hqpDvkbCpNu6HYDj+Tjtb72RKrqiZs+Rpy4hRGwqg9mbCVPd
UHGBmsbgWXGuwLMbGEUKzHzhaeBqDvOhbd7qzMWF6OGr3cbg7onMcYXZQM6OLZXa
7mF/7ZtuqA4yma0ydYRvL8e6vsh98hC+7Oy5ubC+99uIWxRkeKveO2/2yj5Fm8rv
zYhiXm4WArcFFJq3hCY/dQXURR+e1qkhvPptIGKj3sL1dShRh8+XmgwZSt5wVSv0
sIv62cKRQvDZ2dJta8IiNESioOGlkuJILcE4fLIIiKnNPU52GXQZqiDKcp8zjREH
dM344ZWhtNLejGK8cT0xcfdrq/rFeVheVXCynoqMfMYsbp0STDI5eo1G9J/un/dp
RhnuJ+BgmRKZY0Z3WDrQpdugCBba3Bv8i/3LX/AbBaut/M534+kAFP8Ygv2Obo/u
xKj7cR4l+c39+wm+uR7R0Kq+BxcybzSExUBOizl4KbpZyBUx+ML2dy5NckDu6h5a
tjmjFPGRBqm81vGnNqfOk1KbJ7i0B4EppFmJf6B9iccmpZw6Epq+SOdneRzJbYzB
H01/HND9Zbc6P1XA5uoRRJJhRgKez7/PBU1dwZo3mkm0ucQFvRNFttSm47hjmJKs
xVcstHviR9ok9+K7HU7AkwTW17wWSBe/luQ+EvJ5hd3RKaBYAMJ59aHkwTzyNn/D
4JMe3G2mcf1zvqbd2Gqmy1tOF7mBVvhuSfbDwtecihlPUGqgC3Sl+mEZNX8u7W+p
+o+X5I04k+g65AOTLf2zloBHvxududy7bmWFUInDcLEMJm9PgZktNbfL13ciH3dG
fZXl6QDJJSDvqvVbrGT2MBU/KLMLtwv+gc7UJFnqnPa/iRAroHPG61YVVpP5tgIe
Vbvoxsq+AXMXi2gFEtjIcmAgWKGm5FTZYzgcK0csry7fzH35mksJtW4Fel7E8oVD
9b8EWspiOWEtrUMnM8VlVGX/77yRps+sKCDO4lxF5Cgp8k3MGxza64DN0H8Mrz6t
nHqGzhLnHuhlYylMACMPKePNPqaOu6QbU1D8kMupNIy0LUJfUWHiC1jD4RnuA1LG
pEfhMKHAMgATWbsAMwbfeAhqk6x/fXZPaDFnZSMnY0A9217dQDfKHbkjJmacWEMh
aUmpFvZoZVTg8Ru0eeuuSISpZ8Gn2myHGDzuOcia0glYAKUTqGupqpH+4it0Lpdn
/IWCinAtsBslgM1jE264uYzw0pXT+s8gHTqnn5ObAwkSd4qOd2vgVNbF4nuLplTm
OPvf99VhU2Ew+xV088IBIn3NCN1fsXUScuN0P9uDUWaUWLBARfLndBB3G3mQ9x2N
5tFluL2bRW9n/wsGZk/q+T7TtBzv9qRFpFiHQN/A3Ise4se+oxYKqs5Mw9jsC4uN
p1gVAv1UL34H57lUwb3QAkHB0ka2LAe9TswyT5NFQx6cXj+senNOCvM6hLIp2Y3L
ZPdr6ikRoCPYnjwq3/0cRfv2CxcOSXSwOk5x1pmsvAvzNzDd2ZdlamS6VThcu6k4
ic9UT545A6+/s66fRKJdByVyjTvcz8s0l0rTXU8KcgBO5agW0zmbhC+1sU4/i0Z4
h/iB1oH+PR8W5wYCFZZcy/fRqpDgkemGC6/vg9QtyqTp59hbv5ALHnm0cDghMUUf
usl+sABnGDf5LWlBQRLpIi/zt4mgwfTQrLXGI4+K7jKerUUBTf2f8EaMmLW+Gfgg
3PRQy7Lz4bioeWfUSAH6FDn9S6DgTzKzbVaByGui/xJ1sYgOCHlJmvjynNASK3OY
4pkhjkUzVRl9Ikx+OEasaSCzdv3FN+DNo1bI1UBU3EmDpZ/TitAwpNjVhnb0zxIv
yXeQFD/VMKavkIp6Yjg7xUJWggiKI0xDd3NcP0zZWRToIg4qG2C3YqDIl3yuHvU8
Iu2hdQ23tAkFrrYVU5r0CBP78yVVq37dT/mTS2GttMfQj2snJWmPdAFExI/NUWGt
3zZdziH36UC9mVlHtDO+G6SC/nH0OEIvFC9xs7/LPAP1xEE+xGadIg4lGnloMtFk
e38a2ZDuG2ntQtOahKx5lSHmjokNxaYBQ2B3BhWGsMqSuZrERxIbZI9E9E+e+3WT
Rh2FdRBh+oS2Wn1bpvZdb7wIA8JwX35ptoZAEqTnvz1NpmVdo2Flyozqva7CsMtd
uuSdy9NuhjJ2vxqG6Aw4GtpX9oXp1Zkmhf6uy5ieYBowprBvdW/rni20ilidq3sT
lrw+18ZEG/Yy2lXqT5ZcBxji9dyV6Yyx94UIR0iLdchimU8YpNom55TyxvT4oEUY
ZToUxKFdyFdL8vG46pja5ZaV7E9lGBIs60iLRWuBXDrtXsxwR5mg6iuDyxsea1QV
CVCoQ6p4lEbfd6+nipW3OSxGOhJYnHC2KnjM7iuTGREzB348ifk73ZqadrnU8+XY
OXgo/4ZTtCoHZLB7OSahab0F2c2FpXL4x6x7RTk+QGyGqZT5nmAvPg3TBB7WK8Oa
+8ky15VQ6i4LXA4vnkzQjCtAXxGn3Zfwah6uVSDrBhyNKGMdtf1blKf1rao1+puQ
zQ8PQLKHXR8cOEDNWFqTpY/fF8vlYy27ADEMITkxeRlkkPfEZKVFFxepcYIyG2vI
y+uIVGKSxdo2hoTu71rGRbX6u31tz7Xt0DybXSYty6fQq0bqpYyYFDYg4C9thlcI
a/C4KLG75kkOf8FOucTV/bpbMOXeAvdS9vZYLQ1lbqQOV7zS6cew27UVxPLzO25y
na7VqCh5hQDeaFzCMn/XOTJ6xdOgPmg5srfZYes55kVbr91mGkerDP9sXmzDplgP
pSUUjmo7a62hhjs1FFbuPybgUqtWUwstqDh1uChuORLqA3l1kpdTVH21afn5jYVh
2KzfteN+DmDbtcH7Eqgy8LC5/hcxPdIncRYQZVZxez1GkiTVg9S1J0GQXxxX5sC9
OBjCqqz8uTTxygsEPaCaaaL5Sh/plyFzqJuJ4SK9BQejfWbGiRT11qC3aFrjenaG
ngH47rjDj5Zm3552Rr4mhxLJfNJnQeV2WTMj03XTUkTnzEzkQLC6BNLLYUwCpGnk
4xwOAWUuX/Zk2LwbltMKdIXEquY0sT+32fOWtTr/5Op9fWG+qLwEnel77dQk0V3O
+xw5uIab5IWKUVggzkdikVlHKA+MGcnwjmMFTAhdklx1Q5+yq931LdHpFY/BiXpX
ZlgXzGeXOhralsIhho1SjRj2aBTABJTMAfgfgip/+0Q0ukQ+r14/QDWNdvbadAtV
B0RJ/IjIHJZMwxQHw0EZOZkzAfs2iuD5S1Ayhy+SGAqrueZOUssl1m5QO9NJ4CVm
vutEiHdOoJcnuKnlEARbTHHLC4bUTOidSWoaJldsp98H/dAWJEc3xtYEmdkKVL2e
sRpmJmFo7pgQ06L2qYmD2aIQkq3XnhZ48WKvJxTu38EY3PL3StejnK3l2UrJVIDH
euxXSOdAdUs+dmVpJV5E8ejxlw0Kk2sOd83B2DTUNXS+2sc9X7D/rtHBqwmkqB8d
kIkrerS2oqXdT8ZiKdoIaZSDoB6nOIxckvH8hHt0frnOeyNB/Wjr5YMr5szpu+He
TIgkKpQ/PNZ8N4b6mqSfvE6aV7Ec8aZbqmi9L/Bx2owC9hQg2akhgZRxr8OMoY+r
S8yJuwqUFXBQZ8f6Y73dcdA4hIvdA8FEHzwmG7JtRtvAUxf0kuhGkKGUaadq8KlK
YoDMBJBCd7KTG/oLCT8VuRsaS4qrMhFK9VwSnSWId7I3TY3xRmA9pai0AfLRcFv4
TNV2MM2L8SMEQ6WKG5LnYgWBkU8ryNczBr+/uJeWNsOR4DC7cwJNzvDCBBBeGDaD
65zkG7Hf4B+teJ3gqieAyZLaz10HbepUP6t2bAUw4m+IEAb2/AcvEcCjqLKhDiAH
HS3iugEycWwjdSjPI4lc2ECs2PSbUW0sj60rA5Lj6Iudju7sdRv9VIdMQmaiL0js
ijXm5QMlocYwJzs3P3pT3RFh1uewOY/plaZTfQhTaHjveFM6z4shNMqK4EWtT91s
crjA2Ws9J7s1ovG2cPj+NQM68UD8r3o133CEnqcZPSiOwoPl1f0O+iI3KHs7l2zp
ioead18qHh/7+0sjA3gPkp9tetbaBp3oOVrPER++rdzvrcSHzABta0Y7yClGSGsl
/4Wu0PecMH97SkQ+mjAXS5tt5D8oZIhCecpgv4kDiuqGLnEz2w8t5uwWyP2JrzEp
5Yoi5uYGUNcKAbvMcGY2w6Ziog278ENkvO5y8C7p6qSdB9A1gJXHcXA0S2siubfv
EQ879NomTO9ANqX2nHmgxB7oAnem4vYCViYIiLW/o3j3EloZXM6cUkwfvuLninzM
QwOByibXEFFIT24qQ2pFyPmlgDZUXYzvVta3Cr0KEJdBr+4thmcvpNCHmmyk+x/F
1P1KVztw0L/N9DzX8hw1f31YsxTvGUeAuONj1p1iOFzSeJ42gEG1ChZpGyG3va1b
oKpbtPqD6ohsy2QuV8Ya9VfWSan7s+huy8NCR69G3i0vQLKM14Ay4ooFNEcmAbgz
XRyAsWNY4rCtgxqoeaP9kKenMt5iNRl5BwopLyA5tKE5rXNhsCgf5LPEb47JCC0x
NVWonAl5QMdHjrGzoqdea5BbWeFFtGwx0/AS9zzsK7NsqwD1KPR0dBjmkDu48p3q
XJ7zH4Wuz3rTweyn4p9ZvmFjhbYSb4GhdM34xVL4B8DbszDyp8JENfIQVrHHN1PU
7wjwrvVdqQJUz3JRm7ZSdERS22bvE8galI6KsjZhLbvh3xgabsE5eenQmEg0cX8u
QrC4uzf5+5o7j9TJ5hs74RZPTLF94EfDhFvb5ibWZV4tESDkXm9SipZs4VbtsH5U
AVXcOv9zy71KVgNT4bvZO/0Qanb2dBashdhMiUy9seicz4vQf31RZoCq79U5o2Tg
gx6D85ZyYNU+ApeG2/sgI5cvXdcUWRDluj/CYR7fZYNOc6U8CoOBZRZKR2ILxPjk
lG+eGwbgA9O5tGCJ0sUnYrViWafENBb2RqjLMps8jlJd91xbmjUUL0fmrYLYpSiO
fO383rtI531W2aCpy+y+fwn5ojy1s8KbTPLSWVH49LACpBBo/17PF7XjVQz+oqdk
KeRz8n3DJ03omTJ8lavgWH30zyiUGVvi6sx7hBFDaVQrM1mdmbYpv+ar3Ac9BzcZ
G52yo4J+eJNiu3wUMYrYmoYuPsOOqQGRQaaZDU0grwo1LvkOZVsiIPZRI0koQ+fL
7xy/dHP21nU6th7Yr1fF7OwHfx88IYkHcNjmfwX/tOlYkvXmtMQUlpU1ARO5zk0P
G8XvpyGrNohT5GsNC7GXbP++oolMMfHklEfVH6orqh23oRHvV8VobolhvssN8oYR
jere4ZU4HJDfXEUWNUEoLZgiCygxgcmSJ323fDqHE7E=
`protect END_PROTECTED