-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ZI/Lws0M4gF02ZdVL/6pFAsgRoHnd9G1kkSPrhA/T9H23vfT0wZhwWn4J/LqKQso
xqVbLafCmJZZZS648ADKPXpiWhMroKVITl+lWPM459WGdvTXzTTsByV8S+JKLTf1
iFp/SDJrOnM8K7UyFXUppDoUi+ZRceu1V0CFF0mX+vr48P/BEQagkg==
--pragma protect end_key_block
--pragma protect digest_block
QfA6cPnSRbq2rXl8oiUehFHj888=
--pragma protect end_digest_block
--pragma protect data_block
FSG4wotyum+4v7xx3WkMVLJBfeyxwjL9KS+fZByFrXA0HZgy3XRwvlKcowaWje/c
awc8s6Lxgk/NeBL6pEKSdOExIJ96d+BAUv0hnYXtg5LnTQRHxLoG8m8zQF9S3Up2
DwEzhYNDMkcqmbnslX+31IcY37H65AqWQi6DLlUQJxHJezceTAnyWK+v2EViffAz
6oBru306R7VUFcOhnzO5C3Q87tW3hPYsIMB6g/rv4i8A9xw4dobjyy8Nl+u5/JkZ
tq51hCiKhmygLv8T3BYsCMITGR/5zoFdQ2sldtNvl8V6YbnEWnFWLlcLDFhyi8Z7
1+Dk/fSfxesoRJ7kZvsk3pNFVNMi3cNSfUyqwLwIKRFYHGpy1emvCvL6scGG75wu
bU8RQosJ2SOGjzHp4poT/MZeVYwY6f1QCjyA5HSvNkIzQhcfLhPi57uGLWc4rBNN
D/9rGIzoBI3aY0OWsaB+i8HlhlHKy0CWIPrOLu/A2Xi8zHTV3+SDWPacCuZ1eiSS
j6EdvA3tpNo3T2KKc/z0JuIdjG6TthkANRWVTsLiZTKoV1Nepn9GJbHG2KvdAHvw
9K3Fyiy7Q0pIGYUrK2OEhKfBUTF3ivQ5QATJoZkraDZLdpMBW1OBx4H4AGeYSdKy
6eLveQy6okJOMLdb3xZJCs/jOJGqKjVlKsYlYit0cTT+JPVpGjZTEarnYIfy5zx+
E0fKm6ySn4rrjVA3ybI7lTrsk3dc+mICJa028dkgxQ3rnq9ee7VqXAj38fbkf/4D
ptwIJSVNG9LoyOJc86hDuFUXcD4MgkwVhYNkTypEh9223KmkacPeUDxlFik3h3wm
AIXoa4h5i/zt7vSPzVcr9ruJgcASnqnVqB1jHWo0SnYYS/x4knEgtTI4kQVILMVr
EX60iaD5LrJ9SzlFTSnmw/wzj/2wHge7yR9pMxao7dUI5aYZ97aP00xYhh6vCi64
jATziTt9wR+r1f6UV8wdfUhtoczBM3QBt1Q33DyLslEOsnkTMurc0yam3ly9WCMF
Wp7KI8a8uAcfuEpLHLlypmqUUvr2aGhoZXGZuAN+fLQIbBBZxaXVihQyaSitTv9w
u/f/if5BWDokQ9vvmdQLkDWCiOEfKKM2vPc+M5ZKDzYS7HYXAZbtcluAdxhZ2MRZ
z6WYdjQwV8B93adzsCLSKL+D5flehp9Jw/mW2rEN7GIJcBsDXYQWxRUPUKu0FtdH
kPvDiBnCKsT20q7A30Ry/oMqyQA3JM9rr+kVXCqoRALkeVaF975WQfP5PZKrehCn
rchem23C+Wi3KCJSKkfxuv+iUp3LKlCZu+89YqWae5BX2KnnbEfWRhzja/wH1WTX
AaPL9HOWKVrWbvrXhvzWPaC5H8m3g6kS2Rjq4xvMpiwNau+qwotbYUsBRWN6IKbu
b7KHgQJBtu9fz3n+YGi9Fv2BvrTeKc/6SnGINOe9cSVx+zlmE6xTOz0UPnFR4f2S
cs7kkPqoz9nOm2KS4XqFvDxEUxLymPE16DyHBDmR57xV3ryZNXRr3B6eAhz3zZOj
4aM6sCzPmy2fZ7gO+D0mFRHKJazp9CSrsN3YonR7aElUzjUaXCmBM5OAX3Dr9nP8
FkvYy/UnsDSwtSf3MVNhQAePjFmTxaNXzXvKVmORN6FlkIFehyIrmHrJ6bulw5Qn
XPy2p5qyrY2IExLDAum3cuD8yQTsO2r2x7/r7738933MxAvNXnQrppiJmWkjtoTA
ub9F/CsqTsWAGgjgY6uYfk0Tcs4jJw7AlLyVdMKYS2Ow52lITTP+vZFTRMX9A3sN
iP8L7A5i2ytw76sLnOSAbmndGC9UNg9PYPdypb0GzZkw2YPZk8DDWNu4NbCNWAcU
w/+fcRB5lroX5Wj2EPM7NlsJh7MeR1z5S48PCAtJzSCi/MM+/C5EpI307IyCXmzJ
lA6yLTTBt8sRVyMT5gXaTBnx4PdSQ2QvoYgw/PV8gXm4kviFeDl+n6bbInRGPI0Z
krNerUIltMpn+jMeiRUCKe0/3Lt3VxjpNIOAM0730vW66d9u9lMJ178Org7B6GRW
F59Cp1x1CrgK3pcIPbowtT/8wPTgcohrC9xWRvGxhceMejxZM36e1ZvSbBD3flMd
cAd6CldPx+rL6s1kPisz7NT4EIYrf5NC+bLnARUhW6lRe45CDIvCG0180L/UxltW
3ugWBYs4vSh6/KykDVpiKvZWkWCdS8B02JRO4FIcFmu8gqLS+HagurVMRymb2CVJ
3Z7R5QXgX1QRzg/uPgrkEkRJPk8tkiem4Dx6hIW5qtboDrFL+cnDFvDO1ZlU0fs9
Q0Dp8t9K5nojuH0AcAn8jgU4UXxd7nCgeNBl1jUB9UPyyQT+ibK2gwDBEWFjG6PT
BnJdC2QejBb+iytmvo97tsZqp3vLJDYlSAqeb1su2LUo3JGLyA33OrE/WsYEd5nr
FOBhVGY+toM7Du2OqHU5l6Qm1HHmfgO7gz5V3yPHZ3H4NozmuevIMKufEq8Th+v6
AIyjat3Dl3A/iefK+OxpHf5TQtAb3Q6/Rr0f30Mxp4KEAjIUsy7H+5r+gHMa+bqk
pU1RmI9zuZS7c9XbyNW82L+toj7KM8WSOCwmsc8pZWbnKD5KS1+xOX8TPqNQGiFH
V5ehpvr4qLlvjtLkYhUQa7bu5aqzCjvreZjEKAVZ0pfeNkFSr6lP9qtFUA0nzIVc
LR/TinD/StEhnZSjW1iD1+9CKvDJ8xqzWuNKbRevOrd74iZd+Tmmlc3LobD0ALLh
f/grfTX7+CjcD9AEHEz4ZGq1buKRDPsSIKNxlaxY55H0aMsnYvyc7ccii8qTtbGZ
KlDJ00eMbWEk5bvwpDk6Fm0csluRWmLuXEl5udj90rfcTr4mkxCD0eK4dI3P9pqG
ylmHGHy58f4SprJNHQHRjVfiDBkaV2z8UPdsgTs3jFCWYaowQklDqLIGSoMgUole
x5E8qTJ+xyX19kVxnP6FXRxSbQvp2/lHWCoaq+iEeF/GmbhqmZIRDBgv5E82xaMo
5/FAz2J8J0f/cyHHRmReaMw5wySOvCpTIHi9DxnTB8tC5BlJ1w0XogGr7yXeKQan
chOJe/mR5/huBsK8UCOny7UBjPMvotYrETyL21KfhVNLeGSzTg+Gst7ZyH6AbsYR
JdceOlPuFrTS5yo/MY6j0XmaozawjAyuJ2kptECJHwUeOFYiJQdfC15f3U36nO7g
bARVTZTMketUUI8pYQB1e3dN1TxjzirN4dE8+R2Bjo4Ko2xfLTDXhCbj/cp/QDmh
7uy8MNh4fIyk9MC9bAwqkiugiOpxvRta3f8/JMU+b6DUZizW9fBlZUBkZgT6P1q3
UnZ/o4z1Ajkm+gKU8XuMrS+YAV4p66RcY2ITLOqKe98i39hKc2aoYPBi8aeKPRmL
XR8yHu0DdPmDmf3kzqNLD2FnMGhduIxkkLJ7DV/2fW0UZsJgc5LuAxJUT5Bfk4qq
fsPbxvYX0hPOPWhdMmr9rdejD78WHC1DG6ufCNlf3mtYhNBw0CAK6sgapridCMq2
MlfbIkPpxtMnOEvNENBX3FsW1ryv+5AIS3w2DolnA/hnnhc9EGpKEKgcAXaWZMcH
0njAeJoekgfArzrUcCyNHPhU0EC1C//6UwsikQjWOYk5UtCF6T/D1NAuMsju4Dxh
ZJZ4uTKKbcApQdfMXa3UXAbnix0KcpFUixE0hj6Khkest04RHf3Bz+Q90mP5oljn
voncDmc2lb5iGb11T/09XyxMaA1diGliHmPfoQyYnNCZHdRq/pYZ26siAfGJd0s4
23OgOVZKLtvUet7UbPaC+m53lJwHZI89VLVHblUSM6eNBoU2iG34/TOmy2t+BMMU
KJzlH8nhvpca8w2/mHDRct17Ebsuhbj4Ez4oPSOYYAS+f/uB6+fmRrs9OgLsRcS3
OmDAuruGs54LgNkC/gyv2sQSnMfdDSFP86/vb/60pKnvzojgAyb1q4dMA81b5OKr
Wn5EnZD86pTteDMHOpp+v1jYpjG5aHJHD+Dw5DKverARTcGSlAY61vEErP3JH3qt
AeJMiW8Kl0UrIj6sTCE8nqKpeF4KMGxaKVudELn4F5eWOqCUGdiNLpnWa0Xsv9Lr
TuuA4oOQVyrcdQAxJeA8NsY9ym5FpgKg7K/oStL/N3vE7TuchSoDyToIige2lu19
TgQNw32EkJ538IWLTstAJtMM7hEHNEv1o/bgTwLm7HHTEqFrBmCtMPCJ1IqCbHZU
QkHNAs2yXvfWQn/JpCIXVl5U2vBC0T1VcuyUHL5xEmuJ/IXOV6SIK3BUPWI+/v4s
8vC6vHqzXoGbg9KbMTaE5HeU6s6p/bx3JF2a/MVB7KC0SGcEMGUREUccKcwq9yuW
u5iQwSDpvFKeWaf/L7oR1xJh4n4iTSmSC4L51seyGyeDABVR+pAqvXapUyQpjyYZ
9NLPjvjJSEVz2T8Uk45A9QrH/6q04GcVzQnJAh3fK6DRMbZuzp0qwFAuc+ArwW+b
E3Y6WpF5pk6uwJH3sJoBRugKdr9RMhOv6/LHtvdN6qfOLq5SDTlEjBPkTA5VhEkC
wM1kIuvWC7g5jTazK0LUV950qMCyfpe/j9yJAh/CX7AAR9hFcG3vEFPtaAO2vmm4
uXls83EqGSEnhEwQ4vnl56fXWV/LVfW8J3hd3KrcmmPL8wsvihxgXTciNYS8r2qg
TbnrksuaVPj05oNg5yazF9ZGFHjZ7orfFHlHrJ7yi3HkLKmYzUaAyIvHnlVJDqDN
OmIjssvY7aOxiYdcUnSbdIb7JqYtjCxLtzenJp2643nWb1hbxqx4e2EbyatCDhNB
+RbRbbbAqETszQ0iLJwaqyUt0e2jcLvLtI76bUTL/FKQQnOdGkWQaOZmvLjIZoPo
2//GcR7Id/rLI30Rlh68rdzgbGDq0la5pL62nBFOIV25IRd3X8G3NaBUSV72ehTL
BxUtMJ8ROayYpNpePKdvw9FSSUflqRnAG602UTJdHLOI5hPZQMGDYwzUIMwo1d/u
mbxT1jrbc0p6KbOaUZAneV7NKAjA6ixSohCyb0i021fN2Lg732dqWWiApM7161Tw
sfNn7yjsOw6jN450zSZok2MRpqGSBk2BhYBzk0WitBoXJbe/TdoMhO6xsp7aTZ48
E6pNYxwoWg8lQ8fa863SVYAY9YjeDp09JU0vKh3q+tWkFSa6PPwy+vdmu9pzRZ9N
wNqLDikhpw9zCrexH9nfFer6y8q47wqrcBHon8E4avw4mD3tmeAicYcSxRVzZ0UC
4YDY6bIquwghIUpPs1y6yLptiHqrN9SCQ9yZJrwAxCsI+uz57Dh+InTRvM/ZnGoD
ucnJ+dXWkDO3by8DMGtJdwHAEan3pZg1vCkq4EcYp5Oz9ouXTjklDMwQkIhJLBim
Ns9tDd0QMOaw7yCrzCQ6uXwB70oZiH9+lTMLD57s0nWmOED+ew6G2Yi91vvrSZTC
cuadST4iud+8JYMUF8JlbOY9dxGjAfgC52+o0yQoH4WxkUiJGrmZYhuXF0F99j8j
pbzJt7tQzLeqBXixOU3NoHrizBRlMDAMcKU4gAR/ZC+hhmG+qxjYil+ppWxSTery
7W7Yes9bN7hwP0WBgiVrYh00A2GRrAXM/eYqYRUGGc8PT9tHZKpV35PkqztO4cuJ
rYHmWDyjK69H8D3Gsq02s+SCmjGX8mo/J1/jHHhSNG4eQ/Wu7mwY3akBZnWK1i5B
GxpWWSaaC7wcXAXIAw8NiDUZ09yYbmskqUvhKUKMAqTndnmcBFUz+i0LFA1hswNZ
qeEoNO3Y8B4X9gSruQWlZiCW6pgnOU9Ds3WzOrVC2yWR/YfqsbIqVzQdQu/yEQCH
RB7sr95unqt7Otfeso7Ij2zE8vgmlAJFur56bkIisMo4Gz7mVnG7nlxPlnBQYJ/s
gEt9KDY3xhcJj/+qC4YSqxRihxWm3yleAxecC9sNqjLetnzvGFRP0tUQWoKVFxD1
UnjgOCgcej+HgGm4TUY96GZC44bGTW++LNQ2PD55etFFWHUMjo7LZOG5PkhpEzZf
BN3Xjg5ajfU7Sy7HxLzrUPasJVA5Mbn8qVuBT0PvzgEsaHbk01tjTfYkSIXUpTbe
8dGfQ8x9Muwv/mQKcgGwOieYPLoCje4bRknC4H7WsiA1jJpJ7bBJmQw9RP6gqOkl
Ng/npCSo5Z8RtU4TT3biEiWojPWLRoXsrduuiaNtxK6h1e6LDp5Re+21xGnOuVj4
J2suUbnHSV4O92mP4w3YU++/rowSMw/njDeT/mPHTRtToG6NuZB2Sdwp3RM7nai9
4L9hXFLAzm49szjHEA+GnWA6RkPks33IuudxIE8ve7yJFkvdt1VzNKKgK0TO25FV
/IvTwHkHqgzT7GaOaxVBx75J5XsGkiA7hjOWlOkH7m2d8BBMxJCWoSB3kavMKfV5
/c9/zzVnRP3ZUj49BE7yc28uzjrxw5Y03Ivuxxq5NEqHo3lJEXLaXvZHD/uS2ngl
+Xax04iRYa236+PpS7V26yWioUXXmMHbpR8Yse3O1Erxd0pc8ychlmTA8gg6W+aZ
l0k+ZFdr/mbEKJLxlwCuIIX55FxKlHGjyF2/vhjnWFccbChKjC14L/rskqVCLJ+x
4GDqhFm97BxQsiaGuPfOhhCXxA7cUJ2HU2VgPKRlv7/R92ZLNTPq6CBk/Im6mihW
lGVazaoN0aUMNCRyRnvMmOvNC772b3rFhlaM2qf9iLkhdyFyuG6ivCCRcsU6Oxu8
k0RRMsqAROQHiuV5YjdpLiyBnEh7zKL+GISq2A1VL04tqEZnrmQy5U6aTW3HPWUX
InLFWb0w0a8FgwR1S/GT6KZeap1pISO5ZaVXmz5R7J7GedmKh6bSPtYZSaF7Y6Nl
L2434WToE6STDKLp2/PJUD/tICvU4N7tHC+Ert02uXO+ZbGhvl/pSjBKE4Pl2Z8X
54V/+7sf76ClTxRZUXv9X2krC60linE+O6uV2MRjT7YOUGB/Un4UkZYsQOOCAMV+
ykpO60Hr1FjUDXJrabc/g3Ko91tDJXDQI1fXw4ciQpDg+mL5psh6HO8JHXvXfvnr
z6bg9vBq5s+MvhVXmMFOZRRRtxhhfxbTylcqwPzQ+JfkvmIh1zt5juAvL++c5gBc
f+tDi8Q7NvFEPHbW6j/t8e4InCbm8eZUHsykPASvilhY+XHMTaFwenT6NmilblsX
RrK1P6EcslmSIL2AqyKGiDSkkrdjTg5SqLWGR0eJL4emWAi2LoK10UiBr6y9pcnp
TMRpy8UsRARrzckuYq30QNRTqqkIKIXIkIqKvndOQL86bCDKoyENAkFzMCdiyWLY
gaxc1n/Ii5TfEpKd3wpmwxsCtazZKxVjgf3eYcuK8TcXualOrFMzkeUk0o0sbENF
UJUpAVl8bOYuPWK80jyDj1SC51wGOEQRrx20fiYyNIbd1wuo1jfhpXNJpaYulNPw
R8b0gWrdN2UJyRNwEwi8Mbc9JtInGwCwZgWWDq5C8UU3Kh7OTn5GwxMkdJX6jCw1
q7e4NVUP+YmQ8/4R6TiZmksg2pR+knUx85OTHQw3YCA+PAwEVv2XY8tnj02Qkufy
OvN/63lb25Wvf+Fd/DwjmrUCx18zd0KRjmpNM/R848rGRYhuMAzEOxpft4OdsKzc
gEw9CovcvE9/hzzXXCoGMsHgw1+ct/t0ZWNc0ptwQrWBKDAjgt/Mxx0kivGlXeUw
0+vGklzOqbzQXqb3FoH0OMm/fqsE1MDAgWLuAGCFbEHjyuSauDREC4bthnrNr9IB
wsBzUVZAU+XNRTDd2PGSXjsNe6jtUkZ5XCANQJawkPWNbjvDghpgxZ9OGnS+cgYJ
9eEhWWB5VxJI7ArGFL1XXNIrMe0/A42dDiKLY+iTNiACR9ZtaqJZeQn7ozPepVcj
eZqCXXG8k+Js2X3ar99dz53SPgI2XNBOraL0j3kyQvYiE8g3Qs/oq9+D3azruovi
MquBslKi5o44BFkWZ3oDqMa17mFgqGhX9w3ILGQOgsDLpwNA09l99vHfdWWDbXsK
QtC+RZSrcvSvZDIfS46Y/HT0rIpXQf8T0iKBPZGHKzqCxEQTPcatlOORt5Gepo9a
TV1kpCoDvRvbRSj7thmYFSRnw86sUHtOH0TLVjKpNNBZUly6tdV7RMbg/iCLZ+tK
PnqVF9h22p68U5UoBwzg0+TkOHvfU0Evs9CEWENRlpyEiHk+y3FNF+Q8uLa8L27H
FekazH34DF9QP6v1BNZ9EW1qCRcJL1ARS75idS4D+N5AtQupvX+HpeRzHR1KPMy3
Vk0OQ8gLIlWziYUl0qcIKPq/9EfOgDKROHPvOBc5PYgzRbUpx8vsYR8ttgG0Kj3t
5nigvg7Oic8rlFhaoXcWmaYXBNmEqxnN8lmGdyLSyzPIyQij+4aWv2OR9KQq6TBg
Hlbu5VUkC+87itODlue1Cjgl5gkQVOsupTfoWXAXsi4jgpQBAGhvBFkn+lPIqeDB
AcXtRViqSnC+mXcKr5Bd1N2zpofEAIDZEv/7ZXIr7XtDX1y9/xfsc85/IdmKVOB8
K4MAF6zwSHR6mT5nBrZVQJoSWW80xJYVINJ0j+nkdHBFmAmo6HUkoYl1lV2bpMnR
3TRilcAH0wBF20oq1WF9YnBgdhWOL/uG9yM5PKP0UaLnhLqldq92ZlN3PRehsQyD
NR62ilD7D7kVacMnWfYzx0RkGiEh5fk+/n9lBEmr6VgNvJ1IYdKiSak7HEx80XjT
wa2Y8WcvN47rEWFPgrtHEwNdyRlZrBK6eY6ZB6Ht9msx70g1lChATlp043Fa5Ery
EjGz5q2rFiJ1vtBackn+QqSzQM2cQ/uB025+hg2rcenKEPEfodmcAmlgxHT7p91Y
oMf4YOueLLVhAhkW6foacjT4XhkJsDKsGVQm3v17eXJ7XeNa+zePEM21nE5llfED
dFZSFb8MD3G5m2kN2Vcmcrt5ay4ZTya3JoKt4A+bjlEOyBGbUeY+nu7SAqW4CuAP
08/oK/MzgVHmG57IBh64pMB8Ne1gO9MA//79/+aJKUVKVenfDUIM76/N01RnjRJ3
sA/ukytotsX3/sC+ABcIU3MvxrsYruL2qYROnNmJwQItefl/dYBSFDqZyMugA5IF
mo4XAGABG6zTZD+yie8QBMAd/otTjioNddxn2/RkHeQZsSXx6qZrktVaq0UbJhpn
EKVhlp/20JpR+bE6eWYwP3RNrwJf6I7LWhKeePMEOP4dlM9o7rQ2hYtlzBfq8MCl
x2uG3XjL0mbR002OtRCdnPeC8EB9kspZ6d0XKIR/Ctpp/XLMflPWxsydI0SMrAJb
4Pm137WNPpcsB/O9o1GrxuEulx8lksKAjnIapfPk5l7tnw1/GOC0CaEJWIcAhknj
beJFbakZRdtfZcX/OCfEoVcOqVpxeGz5LDGn4rF5EWk7A1DqtFGLBdIOvjJK/LuZ
Udkwx2UvFfLQyQI/tfp0E0a5TKLwkUzglWr6gCid8DYCtb8d17dxQI5vAgmOr0ff
Sm5twA3ohwl3xWMzsYPWu/z3ChuKxUi5dUfS8dXkKk1oW7ztjvhgvqBz1PAiUeWd
ljtf27nJdeIpi6MMd01Qrhiyeu/wbKDP8ZmBXRP5Dy2GqVjbCHhR+nz/dgNuJHu/
/IY7ybUNUmOM7mzwk4P7FHRzKH2teGDQq7qhdA+sio4GPV1hVUqMaDIJqDm576s6
7jp8OTr2ADmO4xTM8bRyLPD8MiVP2D+tcELI1kxJmmLJytjP3HcV8vj2y+VL6mLu
d1lyor3V/5tzLHWGNkqta/bHufkSdI4uVId1Fk7b0DZzov9GZxFb3KBiodTo3gRD
9jEiBK8OSlt8H7wmQc+H8Zo61yRnejeavAXTG3vJ17wSM3nimquFmC1mk04J+9Uz
9VHLIPCzkd1I9QboHQ5PSUvWWXoR0WMlAzaU96H/kEvTxiPiDF83atrBrPLHJJjC
3Fx5zPug3rQf1+0HuM4QHu9zRTmuDg0BBOUphgcR7k54mqjttCXy5rUyiGnIlp6a
TOIZzXh9P4VrseaJ4XQmHBEYmsTg5kAiGiI4oxgyYzeViG1KOG7F0X6i7HDsAE5p
KD7pzPcgONWFWD02YOzBdSofuAJygeqr2BbE/1/p9LAKceKk9Z20DZFHpbmaOWT2
DtpEL0yeYfX/Dg0DVVhxQktHpWEkzmL2WT0fvg1aj9GZE+IJSYYIMwbV+i6FDyXB
IDNpZzt65VOgpl8bqkEL9akyy/+FX32S/pyxSEXt3b90H4Vsy1gTsEqXiiXlYr5v
VHfU0ZmSiepzgtUmb7G4lAXzaKi1n6YCSjfHtWAi8Zv9dp/aGhjm2LgvP9iymRmn
qYjlJKRreAWNCGTvkc++OkkYfvkQyxvDbfR1K7PuNBq8NBSb+s76V9q/b/FXuJV+
yRzI/3tIztm+HmHFovJ2QAxGyaP6HoO88saRE35SPYykm0Y3XzmXvWGpI5hi5GW9
eXCTqmA/7zf9GBnFejWDdYUKlgO6XD/gK1py81Loygfh1zz3z15mo8AKAfd2ih8/
wdTSSpZe4WHWMSqgGmoxUtc2mWCb286+E76qWcuera/GY6aKmyH8pswIZQkiLOGq
ASg2Fizg6c0LcyP/NYA7ac4plJQVFgzyKlFAs4ady4Vq03o9UzM32rxSMH8r/GjT
0+jfDxvjq226BY8r7PKxBN8O7wJ4x2k/62tos3i3zJctoih4rj1PEc667MJZM2Yv
zFbxzYRW95WfVoxWGk71+sU0avLC9ZkcqzR0RaSWBB0kPIlkAW+ph73mCel5qaeI
KQv0STuM6c8sCIIyD+QWZMbs6sPjglBuhAwOoT3n892D1Q7EmtiV49U2RRe9E30R
+WD/aNDntQMPrhR7Y0m+izKAnfAMcS/dMgd27fVPCTmMK4DkYGG8ISEsnk8HbbPt
0Lgri7m+cdFAPKLLgYg/WoZtQIVKPNejd6EJmie34EZUApb67e8rPn0a1iWyapsD
tbdNURvDsW2TzxESOgUbO0lIW0WsH+NFBfdkWlKWeGw4gzySt4TdPlHXol2p/yl5
5a0MWQfPC9Eyuh+r6K4BvAG/ANO/PnhjMvcHB6BbZXegF2RDvt2F4MEh9Xjpb6Fx
wxyobkQAaFmC5Ry4wVpoM0k9R+I4J9gVmqn3JM4RfAm4MNVaCr4NQE5iuhAWVWH5
pcULfueHN0c2WWPwnAk2yyQzS+g5ywcFxOBg2vCkfUMI8xUSBxC5aNjZbjqK/B0z
LgrKwfc6TuNnGK0BF78RFigHzNovloAGXbav+soOYixE5TV3mTWLkd9QOx5dDVzr
mvHAZZBjmQFOHxSp4ofMVCm4wKAPjsZaEgycuzgiwZH4swjziBTorxzsfu7O9Ifu
Eu2feahFss+RJs3L0SI9tTUY1gRDbmyxZ5QufFi+GvQXhu3pRF/7RHlvbQmy2537
wX3KfaAD9WeDIkP+YbV9r+zgK5BMst0Dlx4R8D/Cb99rm1GlIV7CI/dNJuVn0T+F
HeakAMNHQZnR/QEZbnHlXhuFTzMJuJgBoh9V6PRkqKI+2WKOPJZ3064nVlx1nhHm
lRnpVszWMyA1MmJyoFobNdx21QHgwDKtMtO1D+/nIruHLGbAb/G4ZxBSuLYcPT3m
EMn+8JURCown64xoHjbP4nKsf6RAd0eEvmEYQ7+7AgLLPFpbGRUF5Ke04sFIk2IM
+ybgZDqd65xUHbS2HRcvQqHMMHSLr2zElDRijGwKEe3e7hsqH46gehHd8vqQKAq8
Ot+SiH5IA98s4cDXzBOUm1tka18xKFGmBgxOiRnYh0YNRQxBF4SSiDO8zGQD/U/e
pjV24TIXFKGLL1FQBYRevcim1ea5dHKVUTq9Cy/5bNcVQn4JxBpqcdvi3jucLjEO
zA4n5gzpIPXiACTgwxah7+rJuG21oFyGF7q+gco7qV8QL9XJ3u6jVtqmwjYSYcfr
SyL5qBzo7UBVgixzN8zjMVMPwPaAimpCg1wKFUGx81VlFnVqvzux2AHHHpvFA3PK
P8N6opkMpZBI2b3nph01EYQlVUp5VffGJBvDuV8Ca8Dg4V5kyePNPdd5d1eJh/fU
EoF2GiywGZaCVOYQwKPjrZ90y+ApS/4rqNswg6r6hutADab1ckQbZP7AsWnE8Bmt
5e63P46j6MFW5hIehH4dPztpMzibXp3xKHM4dHm2VXBZvfd0tXb7Pw+W3TLx/fyP
yMOtv7vyNV+BXNs4/puIm20nU1sM2LQYAPndgXD7fqwXCxPkbBX+vQywT3X+wVF8
tlLfCpoPXxhEnGmqIn53+HkjCEsKgALJ1s3xpCj+IRsobJ5U0eZ2Jw7ORVObth8m
bffYpurveVm/3r4OYnLo3wQHWMc7EgXTuXkvltEUgWeJZNQdM2thSNY/shBs1oST
AW9NaFkCr9wno7b9JNLQ9/8sbhVvuUBHbs9MUCTbW7S9KdiJFzcBkRaMalZ3tnLF
tHSSmu5lTkOVmMHsfGxFjogogJGKjO28SvZ090kFhiklA/awYZHoca5mOn+HSehC
VC110tDBqkxUM/79VMIleTCLIfN3w/RLFPymML5wImo0QogRCYAn7lOrTShTdYuj
LguP/2nzkShtFv0M0v8C2iBcr+YB0B15/hSOcXbFviibC4tRe1JJJ3JDjuTuel/w
bCyT072na50Spv34+kggb/3R3unuaHn9qdxfOZhDvqck9ThY33yCLderOdNnQZmR
XE/4YajlIHJbt08PHbjqzxrTfJDV/6zQNvAYqr4Z8JxF/0WCp+t9K2mXPHR5Ft9r
J4wW9PfsNqNNndo/RPZoLnbbozMfG5Tamw4jn7mI41L5nbK1O0DQmLV019H+Ffh+
bM3WFvS1ut+vQz7Z5lxOTo400zg224dizlI7nStEedOruafZCFoZtBXrNDCmS5xm
5YtP0z0tWaeM9SQjReh6EDZ860XnUizH1x0aWcMuR6ZlCM1pDnoyOa4GUc2ANjY/
34+MEIuOqjUoz3iyXG0wUsHABncXYnaY9b3ETRvXGrLXe/p5RPdCr+W/YotzlnVu
aUGIXkEKspPvIcVR4TsNdLi5oq9KyJYORK69iwVYGvG+J+wAFLz66VD8x6Sd+XVO
O/J9bzoa9BuHzv6krS887Ovf2CWxunzvBgA5saAsKMmy4s/fjuMYVTLUtB2r0Xkj
P0TnddbJgrCSWih6y1AytZ0/61m4hSULCWvp2MPTSvHeBn8nHkkC3mPu8Oh66u7i
EdfORP0DY60jCeaJ5gRpyxxltDg4pxQTw4Hz4IkmY5V/RjH6InWxb/DPf5EVUkDj
5Mr4UsUGfouoDWdV0aqc44kstcCArJOP1hPYyKPaJM2PxgkSDe+rPaTqSW/Rmj9p
yw/qGfxXE9ycsevAUBtkJCxUsOUptFLZpraExuPRV7zYNFUuxNLi9AHZD189DhrJ
5jDFChTBeyY6AGXlL+LKQ6eBP7QdT/1ypcjHe8VcE97Kgvv2h4+R5z9bt2leCPjh
T6uH5JHiTfR2H5G4XBMv612o/n60gxXZ6lYvM6vfEkSjHUGoO7UwbvwaNFn08rZt
Jvrqi0Xf7iPANv3qMj5w8j4YHT1IGJ0JHWxaR/k6mc9ltFePti11+rj5abquEy5e
SAScMkmyCFNOfC3YLJ3VP/PaMj9KEPgDG7zcRg66wdSnkh6wIowSA6WxxnWf2AwU
WEPOd40i7t3IwYuj6SUDfEaGH/behJjYqzmmIM1ch40C89LO40JsG+qgQQMSH1bH
1KBFphp146KK+2YOROH/PphrBZUuZqBMXgCl80Mm2jUsh+SQRwiFXJPFm0EP8zxS
OZTeOK80lVmbRil6dg+gHwHqHx4/4ecAciCQm1gT/8z/jq0vanpgCydMVsWbvgOx
Ltt740r/utJcDBYtRRiMJoyaqWmbqjPXMnwF2y7RcG9sfZo781GQJn+6BnGaP57g
Bh0a9aq9q2q4b6UrRqaHKU5s0N62OcZz5oJaoNqkNWnIryxc72E88uJrqFONpKtQ
RAtJkAqknWfY0Lus+plZprCiXNOtLxMXI1YkYHsa8yahuTskPHEOP7oGRj+Fm8eK
HXF8ws/jkKYn/4R6MOlNXAM4JF0Vp4YeztxF0sdV9SnEd2DX/c+p0iqdmELMC3Nw
cVdkauudqcrhQPrWgutOyySwxGE0Qh3gF+x03KRT9W/wkkdVrhrRe+DlAlZv6dsh
47wnNT9BsWRO3fU7rQaILAAdTy9L3jVUCZAVyt3q+JYPqdH3wPCVU8X/ad60fuzh
FJTeAzVRhaXp+tsvz8q98cYI+X4Xxrec3iVswR5Q6yG2ngWhOEC50GJPXqlvlVhx
0xBPYknpuXZ+mSy62mmYkzithLvSlnx5/59RetuViUnsSrH2z/gAFW6iMw9UtLxL
JDlD2siEZNjIZcWYL6aqx5b1/AHHBsngiHvMAFWnQZAz/zDik8OTGTvVtrT04aRb
VCFIL8XaVdd2Npy1VYi54xBnIIy2+4MZiJo1swCV9U2FiDIpUKc+ZqnT6OjXFN/s
Gh9IQPdnv26N3rgGBpLkMczcSrc+uaTnsVeLT4YLpuAZ1l1XDtZGayWDU4MybhOQ
3F3M0lnuvGR0mwgOuYVgvNJqnq3SL8lTvJYHmBd96lj2fjoT1/zb589xdBcg5x7i
hgrzu4r77BrfkrdaulyTyrAdmlqSl8pkvxIMZmoUTNHi0DdrDKk1vPPrOOiEhi4M
X7t9jzsK0RSbGuh4pgtyn3zamfQj9UrlBBDKhI0QOiIDfKPRCCfo/6AQTLvdmhA4
uKP1Y2+JMVBDQ0eF4Mzck24CE8c6ei+iTZRhpaToD/BUtUEnoQ7qjy/hhagxKJRh
xboRcEjvM8OBZ4sHH1RYldU6BsmDduVpGPfovv5XBSKgT80UGhCOy2Tg4tyDeiuW
LrITMsf48/Xrfmkc3X4586you+5Bdtfav2XDcX1N1gxxkSPMq63iMlR5ZKYgMvrN
QU1iKKQWG4KViQhIi3lITPIKC8q/xa2Hk83eb2mipxSP3hjUxR1yCiyI4PAwtZlp
vIvSvcBStZMUhwvZtfiOeNWCF84qljO06Y3NTIPTvmfNAdj88ncXj4wER4vak1LH
+CDsS2uZPX+HPL98d4badpJuhdZFFtJPP1XRj0N1TTsUukYpVqUAj5aGXMDAnTov
sCWjce9llrMQxyZUmlROpWgpmaX5VCmKNHKfpaNlsv1BqzziiczjGIcqlQwBs5o+
nrxItgxujznCaQeE8LgVzG8gLdPl902AxOPCMUo0S5LnWnXfai25f9tj7C1T9zGO
KzPvjqHWtPAfj4YnEkMFv433s3x3d8b8WSEjRz4OPTnWDyH8vbKc1bBbAww6YBzU
2vkVgX1KGthxz7vb0bCow2HOuH4UxPaYFEa4MXgyV0IAylBgeKhl6LVJlr7QWnk/
oGJVRZhv+k3aRN/IiSNKBr1MOj62K0bPUjmt6VLKHa/ZU3UgXHRP7gocMO7C7rdc
GSEF68l6dwpnmPXqTf2B5+WIY6cry6OEs9/f5n1U9Re8TjLD/VQ9trNl3i8UaRRv
ihEuuBliYUULNCkkP4RYZKIF8V5gD21kkj5VV/tr3aZY00OLI0d9/8QIfRXT1nwj
SqIzz+XpvM/LyJ6+B4YynE8iVSVaBjZ9peAvNzLLR/39CuVvBIIKV2x4JtHeq5Fn
h9//LZmted2geYTwM2zw27zrwhLbuGH56PaVFqr4Dtlhfgt3Jm++jHur+Wbieo2x
jRmFX3beHm1SeIzoJ4FHpEcRlW25k3x89O+Syjq6QmTApkJRXpcxm66f45S1YqkA
QMG+FxMvNB4bgZ7Mv8/n+qiwxJtoUc7YJRxyZtvb0elMPnUC/eaVcxHbZuLErC2x
ZAUZSDstOweKpPw3bp4BUMChKt6ZqYGoqPuyhz9Zv/pK/TdSrNx/EYxmpZSuBhSo
y4rwjUhYGpCr9fqxp41h/J2w3KHTXYyHkkip0benwSPHGkBKqcGxpvEobOSXem1a
hLNWXCJzA417XwvEOJ4GSLAVw9kk5DTw7QrRS1tA5EWkB3ydXtfTWKZ+pQ+SwfYj
tcmN/KHZDj7fWnXLHkWSxonMk6/p2wwMVgOJdsZp+0kAJ3IF+7X0QYd8QQR4WkQf
CVWNInwZ8NVhoUKIO5gp/IGI7mmIMh27HShrki8Lcuj88ZTcENmF4iQJIxxM5VxO
7gCDA4SylNF8B/nvPEyVnsnmO9uFdzrbiaJwbq87Fs6mpZJhgUdX5LwP32jVktBX
cMi05Dxb3ovkINumLNDKYXNXD0OwAyKtmuJzSmYgWqBUaULSATa+Atz6QHcdyBPu
14XbPgEuylRciIvjtjELgM2YMIPytoryEsizq4C1u+GDDFxK0GndXcBpCIwjj6bJ
E7EQySLVnrjUdGzlCIOdwarxxxUDiW8smVw5Ui6Nd0j6fmEPPoXykBJ0R9ubth5X
up33jTG4717WKUW2GmtPKawHE1EZ9FAWeHR9Eu215cxgJOL2NHhHBcd4/SnCI5AV
48FVfIeUsvru1R61MfIsXher1qQCP1f3R0EOvz5/i1MbqqfgcXUOhO/QHmVU4X9o
etPDECUQ6f1UgsFV+MsNxX4K/H9jJpbK/Lsk7XLILZg3+3rMK/SSmH9Vjjjjdk4s
A2myrO0CU+CeqB2FiwsbtkZx9ArBxBWtLdtFLJHrDfYTReyRiwGTYPprG0G+tHux
rRKXhzySMqTQHkRE3Wn+DUrq3w0E0TDuXLplt7yqWOjUCj3FdjEkLc0FjpdG9zS+
LCOanBUd5Rwq6RARVFmg8IwRJI+RBdsywjAHYzTBd+ESz26BxIaibIXPWvZgBYBE
ONozLRomdL+YE0JIh/PHzk1MqfG5LqBN25gpmknHII4AK5oohtN3V2X9j+Tq6FON
jLoUU7zawHohbmHCnRi808ZFf0jQt1o/oabFUNq7i/TvAX3mSg7iCCRjGIx3JECf
1TnJQCpyoVhHvXIYUv3GHP/ai+1M51TiCGewaJufZ2JFoNx3+GiJwUn27PTimfDS
B56iEXLAw9ELR3ncV3uGqnJ71knD9PHuqQqNXK2eNHXx4iRVnHY4BTxEobsqa3YK
tmpZ+ilud1LV2xlkIHHoUMrM7s2PRHSSftK/qp2tAg10F/4ysugHlC7RuGPgcAe0
ur3xzrQW3dLHXlopO4e+ZEYxKTRQUGejvyKJ0TrsoN5zIyMR+To4n8HNZG6EtJd+
eLe4JO8rQkDLU5xn60vWiaZMWnh6N/m7rLwE2YsVlQ3u/GVySrmEHIQEUuZxkHSA
w3aNT0anJkwbSN5ymlJ/rXWCgSJk/Mk6B6xL1yDZdkyvmZCux1DYZBDGPnVjqO4K
OUGvstiq/zDEjw+A5OJLtV3B6fQBU4B+seUC0EjzzseCd42ptNjWH40C4LQ7fFTO
T8E0ja+gXVFyveP0u7K+5wZKGubf6Ykkv1z4n80weVCTXzdOxDWeW17IHdhN77TR
b0/vT+bDgy5fud56Ma5J/1lSE9RDTxvuI2UzDEyvMz4WcmGhpATrmdPZE8+QONvc
MaigklGrXSSxFTMsb6VUFIbsvwEvALrEEt2b3L16UtPwBC6cstw+lg+wdWqjBsg9
3dYVPAfKrSHcl/AJq2NSWZnpF9w+TR5aQcoH76bzS1teGTd+8YWfcqxzvRpNddj4
aXq3n5xgKmiwCuJvsbsRe0AMxZyenqRA9ytHLGJ1F28pi/XrZg64Fswkj6eHDfYD
KMoThehBScyV5iRWbE8Ry372fD0WkmE4zG1T9T9dO5MwS5CWDC8hSrbP1MEt+y8a
AW0wvlfbDSxtAj8O1H66iTDLrLYNEumghoAGTjCL3NVumyW7cTquOBv/+KHAvD6F
OSN9IRGDWpko6PiweZPHhrV6dg2lAh3EfF5bqM7bVMlMIoW7uttruFi5zsXNHHPK
X0j3IK2razPf5NRViLhSG7iYxp17WIhaFL4YstLZvMaMFA2aElfnbDLOOdjv168Q
HrxMOFMKCA7mfttwPcl8lfupPJr6EPIlfWh4pHurlXAvT4oqLycXeKB2ZceRqeoS
qOjK3cWw8aNMW+JE6UpKGrHk4YG9iOUNYPAVh6urehBhUiSD+ZQWoGBIbn1dmmq3
XKzANBt6PzWBVqf8c8bokwLXy70BTA8nGjuush/aIoiYus4bWZHIa3p2Lg+7pCQa
5pFSS3o05eZGLq/Yj02NQmzhIAdqyxGRE3ED6dPYSdWQlqTEtb+v2omeuY5lDy0u
kXEXnWfKUTmlBTMV3P9LLE8gkF2Oc/cLHIrFwNS7h3a2Ran2pwwZmGpatSnRuR66
Vf/dTnZvB6mzbFrjfS9on1Ak+Tnz1Rf3FT2GJ9Y0+ZL9zVH8dt/f4QqazRCvvfb9
92hlCTYeB8aK8hPJ4FmGBkpQ7jUNuVOFpAvZ71nudzai1+GEAHjyBh84XnzCAfg6
FIaKDj6EJgd4pV2TwaULODSZbMwGna9A0TNfyssIVxHbdGtcDDbIkLnZVkGCx/gA
g+FdSNvD+XGnhBmCPXTQyvDS7jpJ5O6zYk0ahAK9GoHGsTcOYHOL/wtCi4SXv1pX
/d0mWXVs2wQmB3XcCqJGZ3mxpF5ifuws8wrXyhZ74TA07LxLvE+rPlElgEQHGgkF
YMJVTWWu+0ByBnfQDbhxCr2b93BN+zQD0IHoVh0q/j5oyuPwHwiHB1aA3yr1hzNE
Xw+sU6t5rguAJcruurZOdGPGIWBLNjU1uUsiw/wDobu5lpK+N+0yUX0DcT3EkVDe
rR3i7WNfLnqfg6KthTRR6bsN004l9rhPK6u/Km5HQcm04o7423EMAbVWMffDCXIj
597ou1sjKx44bLBDkXGlPbWgmrjujrmeDGy9ibcM4e1QJlO+U0rZxHD5qsSAMN6h
0raKZXZ1NowWUs/8ejEGehpNGVMiD/FKjVvc82mPMGYNx16P7H1tDX0L/TBOaj3k
3lniKajvFQI2MnLHav9IgGAms8QCgQnSigjziYOAz52qSaSmDVD4ePITo+pUmUaA
hKhCR4BBa8mEZPPDGO5hYfV4Gvo0tKA0UXlSxEdHDeQtPPGufm4TetqVimBBorDW
nV6pw3c+fsEdVxXsbaVDxbHAc3J6MnikZAio83UTSNV8lgd7fLaiEylGT0tG6+tA
IRpRHBbEUGXb0ymhwbb8NOcoTjrVTWOXXDfLU4JTEtUF+1bXMKWuxMaYPiepN/IC
whe48SxJEPivVlhBJ6nTeMpJrId8lE6cLDBaWgICDpMajAuHs6Caw8/oY45gadLT
KaKxjHHmWya+nIPpEEFI99ovxm0+ePJS0utFPZdM/U5CErmYQL/r+Cp1eryEnqcW
kMYJx+HAufvOFElvOYd/Vn26FICQV98WYkepd1roMkwdaeDziJUybsC7rI/E8G7/
bhcYbbdt2nYz2bKVU+naQ4VMbdGdNM3scBkpTATkm/04+hhe5GzNhmON/w6V0tMI
wS0LqI/bkyDXub1Jqrv83iHG5avk1xfrZ1IEv8rIGnKENJ7yZDGolE2hx4wBWN9n
ONcwOHNDlBPxG4NViIuAMgrOdwfNB6ERQVGmfi8SKNsHaO3zmTHX/Wre10UhIVZV
KYj8q8ppPCcAX3w+sJIq643EjBq9b0KnYDuj6Mfmim3Yi0Woz+urmoIr+OjDU2rc
ZQCrCfPMubgYDJGkcfKIazsjHf3COMrDGL4T4LUwtcQaAJN0l1N4lSwVOEn8NbB9
+2J2ENp/UQAt/oN31DbBSHWQP11xPzvmfiCI35EmWiBP9S7pZZJH6QBzFVq7POyw
FqX4ZxnqHo20ldmSdrC7xESiRENnlso2tIY7Jkxz39ZwtvBd3ZJyoJ9qC22405HX
NPyI3VdcmFfLtWnuP+WG39OFwa2a52S+2HGcWPZqEQVLDir57VOAYzVlgHJ/OV0q
BwA2kb83CB0fnxcy7/tefnuc4v7n0J4a1hmw5QJNQjFyR4fKi6d6SW+mhS1IjaBR
v+m+he4ll/RsrFkVbDG1vqkda0r7C4aDQ2InN4axDC3fC2pXcr2ML49kJLtKns18
ukHbDEoxALvz/7BlS5LSbn1GFGMUkj4ivRzYS/yBQRZrKvpAffuwwGTGKm2LeEtB
OqHyjrnTsPmUdNTm7dAmlj4TuEx+fG+wFUZZoBY0/SBNBW8CiVj9QxDaznMcDDuL
/ShTKZoJAG7DDAn+QE5JbEEqMhF5AxknLhbn5IgwcikBm1UMlcMzA5V1O/5BnBTe
0fvpj6Uqaz4IxVA0uFPQsPBtBxuuMdncnEyIPhxvt7AE8rn/+xnmqfruydWJESaV
JuRksyCEZ8+GPmn8n1TeVz+EnYs0QGfOp29prFyXUStppy1v7/Erht9wdrNT8WQZ
fCkmst9S6bhiQsMNYmj6L1zL4hGjdrCOnjrEzOZj0WBme6SKxNJHKV07paNya1Ac
lS44RkOF7M1GQqG/pidnRbvhLSno87cpm8ucc5spxHZlq2+1Av+d+dr0mCysfoCP
avSSjk2s546U9hhjJ9gj5jFJb/eHXGCYtN13ldFOJJIrSUkQvghmwvCjK+DvEUEJ
H2YDO+7K7nY2jMTRTbVBhNPrwq6s6HRHpUABLCv3rBYLbkAY5D+u5cq5Sm4QiE42
1uovdvc6XmXtbpw2iWSu4hg8wOkBSpsi3g53qc2muR4MUPPIX4GCf9hUn56OGWtx
vKYZRHI5jnC8X8iJ8wbJ6rbwFsvsXIDCNgeMk6Nr6vE2+bTXbOoD21uITxMZMn/J
aTnxoLeAGUIRqT7GKmTE/RpH3y8uVFiOalpKPwA8AlLMsJSBBFLWsGXqUen23yQJ
0CFCuuH4PsY6jZmhK+kGhnmfW9VZ7JgGCpiAtD+RI/fDnXT1Rvs3jo4FQ/ugngti
n8bUmsPbi1oFGlHb6OQlsAtx8AVILvqI8m/x+EWo7Hi/nOP1Gtdfx6CGbgZxwqsX
DJoXLw5xIatE3TfSS1wHAuAPnEmn+a0rnO3g/LxjgigVrvN+884tDNEOGajydNzo
o5QGd6DAkJ+Nr1HAv/qg8P7NO286PnteyPSLxzTQsW3S3FY/t+eBxGz6xV+ZoNq9
6q0wpJSDtPHVpV+6xZ+ZC5cgs6F/LxnfSQLkon2z2cPwL1aVLyvsUOyXfQBoTcR3
F98KLO16qrfdQ6INiB3ZS114gqIyJSj9YLgjidkUuk0n6IeHT0RFQByrD0GXUMFe
+II2XUE3NGktUKMxXqaUAWijs7t8Oleq866cAvY8tVBWhnDUNYuoYj75trBQ339D
cWy2+rCgXBmI/1UQFSfp1Yde6M9saEjNdb1gpAqo3t5Q4jEphTVTCR9PQ9CYOzqE
V+4jqylqwnf6ia1XNQRnuIaQYiFeoxmAycQgeJWdKxoWM3z92xro9/FHZYMeglwl
wFuk+spOl9Le7XNsL/XYQwBgKp0K2QYBmABLRWPhphBycKDZC7Xf6pZIweNnt3VX
kK2XAJW5xaqUArtFrO9iH1NzyYxoIRVaommEmFl6K9f8TfMKE0amSDRzXCICfhSM
G8Dxa31Jg4s6p7eLWalVJTEb5lLG+qy9DNkrvcZEFTHLBtgjz6OiTdv+M5TbxAxX
DiK2zRTTCj14Kc0zyiLWZJl6b8+bRx5CbnGf1JANND6/K1RZsuvon2Cui31F9g/b
Rw6QM3ybrNYaxR835iqIxTKxij9Upag7oRo5Rre66wFzeQQe42zEPiK2vOOnJAV+
FORhHuRFf9k/e9amVWjrzAO6eAdcvIPOz19jL7EcWhm0+c2YS3DPgyTFpFkEYFtb
vs7yIpL+TVU1tKbeanM1OHfSi2AxaQ9ZcN1BwlHLRWIpHrqVS/hHpGV7xzhj9vYX
Nz4ut5rWxWX2tDhd3TW+72TO5fKj0bB242aaghkEqj/bGGsPnPBC5lF68DJIixwA
2pT0syy4edx+b+8ozcuiIpliG1d9jM+h0Glg9ce9VEzXBc8MwDc/RruMQmOpr9K/
ee6Fd3DqGvsZl0UG1T1VBZ6EcwmXtNs+lnzz2DomqDGQBRpBs7jq78rak1PulzrY
2I4k2q3Lt549LJRLlACEAAyNcm5TY8RtBpyPqQuOb8dtBjh252vEeEFabIsYKYUD
YVX74pxZ0YnMIAx0RYcGjNgWQMV01oPRLAo3Itm50tqhtYzfG+hkw1dnHUbW5GxI
jfEvImU+4CYGfEZhzVecuxso0uY/fLrIJZZXWEITPIEGlqPEKoMg5Xgbkw5uIhoj
6poKVrZ9QpaAIcTnvD0/C71xri2uPAUTm7Gk5IJKsxxcVup/hAey65ygY1W+97E4
qiusx5VIk+3DQdgji1SPRPDmhVU4wheFuHPTyuMD0Wxk93VeqeluMC28syXoasc7
MSwHzXyrgukSAXHHH/uIET30GAbS9QaNIxKT87LmMFI1GXvGpJBzLLeTSSEGcvIG
O3tYhUq0LSIXsFrWoSreTR6sffgioQs40aZkVj/MbAKUYzgZng41TkmTD2UOsKVD
+y7GA+08ZEStjMsbTpivEp2kPaw/y1emmPtpQ7wWN+XWKZ0XoGEu+qQ5UyqmpP0P
8dL77ldpq08tKelLdvKvS/UYdxdT4o1MGf+6urNKumvZTdV5zZXKx8Mgf730gnG3
WAFIqxd5DRHmuj7/7GMz3U9a2DPM1DjgWfX+DDXa85QBw0drJOFwg9FGFKRHMCqF
yjyHVTyiWqrjcvTzm1RzSnVWsy0gfquIzi64yyROIQT/xP4Tr1qFWyPJLTaTOFhv
Qv7wZf62TvQ3aDdvLycEJrhktALLrdLZd/ikY3KMGK2rSh1ewzkh0bSfuzF8sBiH
CnfDzjASZXfd44egArL4P4xO5zqi3Ia3T4XIEPR1MzetVVx23ewDBXtdJG4zBiU/
3IKUpGgIiTWkYCZd3lMvuY9kxwnUfgv47pthilQqqmv3y0irLgxs16l+2lpqoOpI
F7mpGN3vD0babxgnQk/vYGol0ioGGrtGy/9EsGYnFzq1Pzgq8bpfxSdVNHBZRO2A
w6b49xVSU1gx9cD2EXD8/uVXCssT6IfL2SEqx6B8A9YmTHrwXnVrTrNPMewh+7fO
/i1ydokTp993VuOjlN2QtC5SPbhi32kVEgAzMwurJjwCKu0cg0RbM8nJnujBVBz+
fbkI4nMXtUkGYZ91GayCC8SjOjwqTGfIbrkJhvrAafjBo+tAoNij/NWBqF1ZaebO
OqZa4yWLqli4OonXP2Tl0eEgz7lR/P3oThJ6r3myIH10WTs7Md9MrSFTdIH+xY0f
rhuCPXbwqEfIWGUh7RQK8KWrfHfRRnh71bi6BTp4Dp1dFUqv/hRHCivQbXrvbj8T
njAJRnGkGq4CTEcWHSr9aWGQhwmlK6+lHQIl9zgrqyOE6XNcAVaSvHd2pRvbsCRr
vj6Qx2R6iFoc24x3r6gsi6MYU8f8j9W33e2Fw4i1IxDUQLlc8j/+hp3sNePD5jMN
wdqDzrdkglUASrenPfbaBpzo+933YqqDwoJjR26gL3g8UOdJ4Sfv65dVrK5aLtev
k5ENKxmQ8TBynBINuZE5AhUUay4bgzoKQ00/Lyh/G96pNDUJn+grkQ//Tepbbaqt
SUMo2JcD303VaajIp/k3WS76Q5J58WLud//5EaCFeAjYSLA+SOs9HPI4yuEeU4iD
0OfefrCzVXMVVURtuGI2K+FdpahXOd266aAHKwC1Ol3Rx+p2AxGkqq8UXUV1Krln
MHKo0X8EQgCkaC5TP6n9f8sqLrjERI2sTfiGLPvOfQah5Qq+vZfto6+EMGEgGsBR
IivbUCadWz1dT+5DvtmNKvRcHDxoRyLjA035aovNXeddbcWCdXmrt5w10gz81JzM
8i80rKu7awmnqZUU87qsL7qW/W6Q+9nIA76knrgRFKvwrGjhXj8G/TszgXyZB0yt
+LVs703saUBaWHj/IsJEduCEIZHjV4PVSftHqOSJd860+lKlgGX2bmsKPghT2dPX
jbPxjMX8tgkvHIvFqjfaMlACaha61tiIs1ZNCPPuCPt42H2tVf5o7tLkezZxgzos
fgRkG0A0RK22HPtLBuo2x3n1E8C0IGcKqY3rA4jx8tLDn6MQXpeKChLm7PV6hQG4
/dnHu+ZPFm8HLWummY4mmx2nTXPsesXHJ1tqxWdIRxL4Cxko+BZ9UxeY/HAP5/3U
CCJY6tzyBnaphlykz9pRYH0061sr8nRQmpRru3Zu8qP0D4eg0NqeSnTbc57qX7W4
lx/wCEKNtYbOKLT/c3l0/cNA6Ml/CW80MiCPD4lY/hXhCyDlyr0M31FNQcvBox5l
ArdbhXXot3Z+NUQDfLJv3QoG1234CicUVLbSTW4COBD56lZP0fncBJGOqnczhfR+
+wfouD1bE/nBtBb/+oASZdZUB72ps3JIPdzLBzUNLqPq+h/EmBh5r2da2a9YT22d
3K2330Jsc6DZoUtKCnf3f2LlJL+S+UR7vQYdmLDBXZRAMNU9ZoLhjosVPg8G8LYm
ci3lcojyyfKDpEYJEBIQ4jHy7IkFjZ+OvsttjEOLUhTQJk554RTZc4BJh4QI6I2W
9JotrqeW2UdAK62rwJPc8jgTo9U+hqns72h5UjXQmCalW5bENm9G38MHoLsvgC+T
n4Sccq5jGuShf7jqC8+YY1vz5e0PI3ZfuBHFLEn/aw1RM/7dXTnqJUJKk306NbrI
AbM1JGSel9iqkH5op8NkUqhTjBLUm67vRHdSshsPzmDjGfr47TrrjfVmX0/A9lxH
rR4onUx//3eiz6Zyfpdto8G/897/6itAQy74NzHvH9PNKhXTvQ3q2kfrflJag+3Q
fmwOvlUjgBy+3VkUJo9rG9gVEGMheh35jReiz3ziXmKWXt6wFixA4OMzyAN1J2KF
BNwk+q8rvjXB03NF8VaCL1KP3AHVfBlA+kBsHqLhMBN3N0Giu9R0mKUiWHKDeiIP
l/YKAubYxUmxV+7mC71qLhv8KvVCpAYVD0xlxKju6XPf9JCOuZuBeMAZgBCFKtZr
qJXvxcDLQ8+/wR9ScT6mz1GGIWbP2GQKmQjgWHsZ4rk9JF6VXEflT87w8ZY2boA1
/6yNV8OwVPVWooYeAUjxLaEHoYFzGZI16uQv8YotNL7dGRj0k9HBxdOQsBiMnM2I
LLgeozqyD0dIT6pf+bx0Zd9Df59HPQKu7ZoFn1oxtd3wMB5Qztt3SnAq3jn6UDal
zUZgwp/q43cjG3j4pk8Je3B/TLw3aUOgFUbRzMBJNnmN9EXFySQacd/0Znu0U+HK
spkZt5cCAryHqS9RpcrwuIidYut+FxK7IWcwUDoT7c1HR8Jtqmi0x0TlSI/dg8aP
XRis6cbbpC3OUZD4QmcG4KAFUqgRtujJVdhImVWmCz7xHSqyNPJ0bmFYGOR+hgDP
25NhHO3DJBnoCKqmqn2TkTsOwRk1Ekv16zpcGXKORg5Kcrn++yCkSWjCyx8dg4j4
hTvTGHL/pzjm6f757cO5NtfZe5hB8ft31ff312d37pf1BE/Lmw9VnUqqTGE9LyC5
dh7M9CD7Efxzf0oPkfVzfDKj7mkhT9S/eIgnhTFwx22JcWAnNLE/fsDhwkJN/t8I
3F/g2RWFQF+VW6YU2k7DtM6MwpgALQPP1XDt9KAxUTxcNtnD2aqO2f1OuIGzb28r
o4rSzWZPEqku9z3LiX34DhX6efu4EWFNS9QpZtStne+q+oSPL1AP53Oq7VIFh5K2
7RLbsABmrxAE+moyRzPMB9ov9JZN0/bcbmjX2tYPp8AJTZd6ZmZXdrKV9BJBYraL
3QfrQciakZ5y/wyldoDq8ZzOiShp2BfruJbmbn3ykLnkmLgVj3YItWpm4MPQYD6J
KPQiHdeeVmX873D1ZeoQNAuZlWYbjn2RzgH9EJLV/+g1oF4Gs948MetllDeOZfTR
eqvtO21kPLoQHJ29oiFY0biDbQtS8op3ROe0FuOQclxDHDSQr/+v/AZfV1TVxyQw
i26HDr0KFnZc6bM/qXgLTPgcCS8KU/kCWmzidkYdDt5RQrmNsEVGi3K83QX77mSw
MI5xY2uVUlmzyvXi9a3IQmWI275r0znUuVJByjomV5orLpMwQhFpFWA2aSizdl7r
beCgd43emH23hStdIzaaqw3dpHO61UYwE277lTCK+KskzDjxn6gMAkzf56b1Rm3K
MGb/Cw8R2ni+O6Z546+n6I8ZEJ90dr6R7eeIVBDkAz24BUMA4aRmimxRNGLp0Azb
ffJgYruunfWpxXMM8Ia5bwz4FTe35Stzg4/qM8vpj2grCRRNkukDIFtruV4aoNu5
EaR7vbZLQZG9nEFQqyOSjKH9B3rOGzKQ0PZZh4eH50f+62hGOwgnKg7JQK1CV/19
f6iGSAUByjXk4A7sIYML8oDuQdPuysW7JVRFjGJ/X1F0Gp40W+OfKUHdqcGWbIDg
XpuU6NeBTIdviZ0knd5PX/1ENkwEe7ij1+/W/4nvZTw7Ggb9rDRSOtISfKmBNhbP
rNGwspJb6ypuj9MT62DXPK9+WmDgekxxn5KuPsZgkqSwEJPbDkubD6BydUUfI7ns
mGMKAv2amp7LRY2pvkFyXq4U9zVvNZTzUQL8p9Vq4t7qf4IXvV7bZ6RdAu9tRaNU
MIAs7pBqj/ovA3Fl1atsTjxYULuLBANduteRlTpe4tZex/2wnp8xwBJk0Onq3A5B
ZCHKzBecgD6jroMxQrF67B8oLx2AdLGMrQjBwwwQSYvqZ+3X/PqtL/37dDrJ3qEf
Vl3XNpococnVaqR73rbk2mHfoUfZj+1PoPwG7O9bwi2dl3mxsY29sCnfgLSnoOqv
/3FKrbZhYeWl9St+K33sK+bfaqrg6dYjDG+F3v9aiez5Yd7PM0UxAz7td15chb4k
T/mQp2OLX3H/42k1sQXhN6nb3l4rVqLpvT9ZzKNgCgh3JJm1RCePOpTiIVbAhTxx
0x67AKrLFWZ2r0dvTdBKnpZ2xIRwJJFNcMI3R70sszt9ntIbQnbepHapSnfA9Dsv
7sT2NdsJ6q6tS8EpePRexe+z4gkUs2y76pYCpN0nomwSoGOD1/s327alCyiO+OFj
5DS9fRqLoSE/c6c695vAe6x/0JNftOQHU6uWWtPxjjVkANU2NaAI+tdqtIhauD6w
HoCFy1Qw+kP0rdLyIdvyAiiC83HJmyIq4rUuZeRdE6/3BqVxKc1qnKBSR2XfhgjO
DH85bcWUXA1+HlPCIBAoPP6QS4tmOHhhk44mb6zLKNfRHslBZj3HjBTgpBbQdEUT
FcX/j16Xgu/v13MUzYIKV08UHLiLeY6usJbhdmmLt/7cE2DwpoRRJxS9SrIGqkYn
Ysx4TN6Ij7cQ4fAE9gIuH+HOERgMxraI17OECsG7ggS7DnUwaB8pAZvaYvrQciHw
zgiwcXwPj7+/FqZhGXKiTi2jQvIVCZYlcNjrh/9NwiIWKAB4lFXUdctT+CxRoTqK
xa4Q13WsGT5SyxML9Hu6p1XCe/5ubBBt2Xj6nkrrWcchCZjjvNPhes8vnNZRfven
zqh4Fl9hqCGWOYf+kRe23Ph9x44eAt4CTBl5ZV8ydUdStuFjtwAbD/k+weFFHP+x
SoXCNkuWxXTEHmrNPNHbdpbLpONBozBt1gkiJyzaNAyaPxj0NNW45VKDIa4Wc1TI
cl4zoPG5xKgcGNCs3Clgnmtpddo+BuSPS1Nhat6+XW3jU0HqAsRYM6YroX1MoUsf
GZqeExIgD/CxXakeMfUN5ZJTGUxzUxc+rM7YjBUIrt8B37oZac4KCgGJgqWowBZI
nyKJJNTQgvyA9hRwikY8L8KtLtpcw3AainJA/KfqvPIFK/qscJVj3e9/yShZkatq
HT/hCE7Ch1soCW+Hp/WkKFmzgJlxNXVoq0riJCty1JuR6CtUYfj44CCUBtAwEhVS
jZDp9E++YNENnB8LL7vyrnuQz5/Tsk4NpQ0+zSwRkNGNJF/ADsW3I70fuFhUA04v
P6lehm4LgNKaixVC0js12TwCXFTGfYP3X3tDQvp5qliESCek+pVvSVnmpigrN6KV
3WJRqI66Q7HJ/CuySOR79LEfeNrggV7Psj5DfHjGyKQmG3FISiNCw6RfGcDdXbyd
5hVctryAC8et8tfX9wiPAa//GcoQza5pOAfeBjE+oTHPsi4xxzJ684stWN6nsrE4
BOlbeXkYFCI+2i9EV/7JVU+lSKRVhLC4ystcW/XLQkhXC6FZOZJ8714DR6NQuPry
pppxjGHUUYBEetZ0WVi6zVT2FZtnRHuz3A0GhsDe/qm8FS5RtwR5Q5qyp0GedDBV
1IXCIbq3XcR5Tg+Q4zh7j4QAqoWAJEg8p3KIyX+Gkdi38d26wFQn148Qm1rgOK46
9vtUESG/znJ0H6AXt830RtHOIS5QoxMZFfcFpRBlGxNHdWs61yB27/VYmg7yUs6P
mWhSC2nTLRL2UMn27DeEVDCB1DqherUw8IWjcFqzTa4NLez5oUhiwgrilAr/GiGX
DcSgwZHCJfj8zqAXLBGVLUblTOd5eLxz5DRBY4CfeWGdJ2xdLBGv5onKEmUiJRK2
N+o9RYQxUPiYaD+l093lHJaWzzHTu3aRYpjE1RIbNeyJe66kJ8f0Lck0mpFtzt1y
THUbtyfuuWqaONGZSQA3CFRAIlufMtgwKyZ4bhrbD+0ll59jFge1ZlC+owgKj6TH
ZGGFKI/g0ySOAZHmCmAPfiKGpkob69NAApOzbpP9Y4RmgVKw5xUoEwDWNA8k0PWD
p8cI86mRvX7XGK1b1PSycOitqkFctxGf+PA1vE4Rz34WeAF3o/hc+hehLGM71Kam
nYTl2gJ7/DFvgPQliRyQ73zY7TVim4AoZPtmx9Gz7V1+JLfE/2nxsytUnyp4lgIa
w8dxRQyjYUTXploNBpupcDTY4XlFNmNX+T92V9CV3zqmY6RB5Ffjw7WKrMzJ10NM
MLs8oFHlQtugo0nzkXQso9IbyPiw9/EzN7x0VZuCB/FSuJGp0/yvgI+5r3R/HX2N

--pragma protect end_data_block
--pragma protect digest_block
R9zAUP3uY55YQdsZAcJsTZvAQoo=
--pragma protect end_digest_block
--pragma protect end_protected
