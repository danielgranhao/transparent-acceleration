-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
nkvMyvp/jrnfWxEGcGY+6oMxm4x5V4ya4mpzvdoYXyMbSHPWtJ4c5RUvcFDdz01R
mJKXGqigVZROvEPe4pAbmqqpFwJFB1mjDm8Zr2SygWzP+ORhJYdPazdqLtDV4GTm
0XA8QpnnrAw7qoa92QiZ0wKphOMyeS6+hZ/u3eFZPeM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 17121)

`protect DATA_BLOCK
DJvV8MpuM/IYmFdBtylNZJ+dc/4We7DCmeVe9RunyiDWJIdQa1j+kV1SmjFMUAzs
Skd23steH+SZuK7+JvtnobfSYfxug3Ei0BzvYANA7P/jQL/ZiwFumed7zlVV6HXR
Sn9tfVd6UVPgL36wtwcGcVnElJ0fAtOmGB90m9n/ehhkY4dNX69g0znC9YsY49XL
x3riqiak7Yg3270kxkKdAvpGlTWLpP4qGwhFwBMfh9AADW/NiwGkMbgqlqxIhF6k
b1dNJ3GmFiAXy61uLkxHKF/LNLYVUB5xjfwdaX16l3/+wyTLHbyuZMzFSv3DrKDg
bnDr+4chu0xjV1mX61YSpqAxkoVAyvRyl/q4GwPVm3tWlo8eaJC2RRUIUqkhNmax
+9tVc/vOZZuFYkwmtdKSbRQ0rOkeT7Vdujo7SFGUWgQ1XPLWKJpoDoNk00HpPYyZ
LU/jYJNvivdNlJJ6c5uIFHXEnH+6voILlndfAD9iSOX2/tjSWacw9vgaIidKtE/E
WVjC/DMlvOnjaPwf7ny34gpKqVC8xTrCydkO45ufuppv2L5omwlStnDEsBzFP2Pt
YBtuW1yQqCp5HcYicw8d//W2DCvwpfIhJ1jPZ6IA0SZ4pI2RJhrBUhO2l47707T8
awRM2eFOxRhwgqduDnjGT6d9VjtMGXcUQL399GtjyqFtsxxVVUVotp2f3KD+vJXq
IBYQWs0zQ32pZGvwT/lwFwRVhdK1fOQSE0elGr9qW1wpxfqQXWnUA2+P2nGnyLWq
GXHGvAp4sTtYQgs9pQ3v3TGz3rzE+asWQA9ZjuWUts5BCE4leMQwCcavxvgkuCxg
5WjBEP14rb71lPfgR6vx0z71tc6D34f0vUe1qTUT5SoqLs0z8K8ZU9im0dulr+MR
U1dVvi5VjCUYFDnP3FgL/4EyFUUt2c08cLD8EPKaoJw3v2+F6ZQyKCbFl5iAl6IW
DpjGY6U2AAYxAtt+gZLRm8jpuERWtQMBsXUeRSSJvPVca8ge5QHWZNu1eIw3/fPt
C5BpED8m8IyZoBHIAZQg+0FrNwpXhp6nS9omRt1fDZPO87fz47478HY300CtzpYG
hhIRotOOTMCRFi7RSXFG0oDzp5z6aYGBnsmoXqzwV0xdbuZoiGZJS3UAt+DeJrVa
r+x0ixxKIUY3H9IVdTqS+KrX8nCZ5dlhjXxHL4s/m8wQ2izih1hKJyYel+SFxJ2M
fb6YDSxXZ6EfLp5gvSZPQ8kjWywoeuBrLDQr0DjWOMC7zx/RCQSmO1Dg7LiT0r+p
AEfnhsQR4T4jCUqoOHRF/fPaVlwANdaq/tMIdLMvtay9dm0yLgRt6soS5pw6cByY
BsuirGQUEXvdQVyETabwqAFpOHexXwjZ89zLHoT7cq4oeQpvuHL5X1xFe+5Zagv5
aieDH8lMYH603w2JX18zIQ6QDB/8keES6vsvtGNGeAIIfOIe8d6mxS5vvbgIt5K8
2yVZ9MZLZvcEY758q7TDBtUApVn+8g1odnc+QJR8AmnyPnYadIV36r5QGAKZE5Ib
KqJi8VPjhZVv72jFVBAP6opDzyG/TJKq6zEpOkq6Sy6Uwe+hmTQvh/2+C7TXHHYE
7UpcUJhCtfbxSeegoKTTm0hEttPjrvw4xuB/h9PrSDg0yKIFb/gt0XFShBxtMbfA
f40pxo2RkF1jZaVTR+hnoHYB/dX6qxJQRsAupsCNyySRMmnMr0E4ymUccKxCYtql
dc4ICeCgBg46F444ba2cQweXRBaoqbhld6qcoUVDqndpE4NnxF/lFrq4wg+qJXk3
Mj/GZrROOAxihhw4fx1q8SIowjjvGWe41D5X9o0rvvgazX+Cjpflz1QEIWx1VPUQ
hy+7/zGRIgXz2mIUDT349dqJ26yNxEpb8DQzbIoX76yl5v3IPe1d6F1P45E5IZPO
ty+h+Lm+8AH1PBy81ZaqLGxsCmRmb491rVHuLYrfqJjdRpQxSqcpK2rbtYJrDxMj
+4GOuPcyX/UBPCZg5qV4KKqQaEtAViM34pxjQt1LJPHsHLNsxCnEgMTTzlzxVDhj
r41IYh685o0vVOjCL9A7cEab3C4YGXvgvCNIXNasFJXMaaKJvFF7vnaXQ9GyUNOa
5Zdbyx2I6XfSBsLxsfstQr0Iolvp+S5HMU1/e2kISCS/z0bBD3bGwwqwWHY0jnJH
tVQgywZ/BFDyuoOqZUWC+pZdO4I/rCmUZGoD/ZKweIk6T1/BeaOYdLWBfj97vfAU
WqDbR20AqJYto6JB+RZccl9lno1rCoyh8g9//ozAVZ/wY9GzWxf+76W0VJ75/2V+
BFrgOyERbKRHilbEcWy99A51PUarq7OWWs5N7+i4Ek2h/LFMOmRqU73OP9YpJ1/c
VoR4crZyfp1HHY131tiVAhK6d3tVj+QYIY8NgJ3MlubOolSEFN+DiJBPeYpIFc6B
z5MeIxXBqyjKw4wr48FzWTaEZ5/VbD3YrEsmVzR81XTjikqikbVEctsUzZMhdqU0
XXv9xQK6xflu1no+34CALbQ5ScgplWdbyjMjdPqBpzQLe5hIFBgxqw5WhJLQOlOA
VdpS5k6RUwpY4EYXbTi8jzHw3pkEztuK047rlEXeMybTRY/BNl+16jjw7dDWGzxB
z5UEsJOnZwUzVwMHxxTAZICQZlP45sfoNrYJzbniSFuLZtk0LHEF7Jh87EjMNv1R
3G05M8pwSbnN/oDvfcgA8W4NvwOC1mtvuVXLVWWs8qiuuVu7zsIy0/aZxnCAkxZI
MntAL264kFMyKUdLbSWSvKf7QC6+AyNphu+LHlsUywfc+20UIw35W6v7NiDaL5sg
cRdPo3ZOMwFVnY8ipNCSdkBAUMuPDfbNUoGEXrTvGzV8fJnBN3r0jFb4aIsyzGs+
XMonUFpZW9WrpRxRrQmXa3lcXas8FuhGn2lyiAXA3ip4QHW77Q+M6cNLcJfHn7+c
G23t+DXzX9sIRkt/h/2IEi20MIThemDncgRz2p/sK1jtxjOPWrduJb4sEhO7elna
S9KEgHwTjzSiJjTTpJb623upVE09XJULiUpOKTnYJv6vqyIneJg4nrAgkyxPgqv7
NMaBsMdx4jg1vwYPeJVK1Bdj8RvyYuYsIBXRzYbxXg6ucBkSc0wMu8WVkXZyCN2f
3zafqQ99fwK8dhMSWbO3KuqzZgkET/WYWWGhFIn6OtzrJLeoz9MvDcAnQzbZv98l
SOGdZhoyUJzQS+5eAlu8adS5kFJPMOv0YSmLbDYSVybK2Ooph7UC1p3KGLErH8Lz
ShbizspwR6TsOf5SMbWtfTjnO+M+uNZtvChwTwoM99a9IHrXFV6tEl19Qc3OspjD
tz/AeJphrg8EQt/V4FVihJH++yxU7dUikJO1+4BdfBXWBCbU+kM9QuJzkwOAgScn
A63O5wWc5it6iCjyXOIIENteGtzhVRo6T/SZxzH1uESu4Yue8dNreiY0JgfAQTiL
1r9XCcTmfud++xS4pSsUJP/xRhvmmMalZgZwhoc6fPkM1tJS01jbQMv8y5RKvtyd
tBaI/ySq75VdjlNbMsMIpL8QDNmmRU7hnllJyW+pqAR6CyppM7RJG0hmccTOuf2z
q31KYDmUm3SqAVIVNuQjPU2UiIb5sGwCtGOgpF24dqlo2O1/xjobY9Z0qYFuC5rG
xXIi8Ih7KY71BkfMgME7qVi8JUSGLRJWmImkZZFoKaiPSriZLm1s+jYaDA3U3o1j
QVPCiDKGO/tOaVAvXD+al41uKbxn/f0kgeEfHIFkSotwaFuu0ji8rTE9gCpqcn5g
DIyy+vWlLbmagFnsEpt0bQdMy6JCLL4M7mdGFtH8twMhcCGQE3e3z1dv4uY/V3P0
Jl9eW9eQfPQwLbrF+RbeNfKqJs33JtfestadACGyLl8q5crNAHLdiFzO4DVM+sm5
zgO1Vyaj3lV9FQcRmXrK9Wy8aphugg2AfcYGq4r7lXF/ksEYgq9p4UEfYShQqwHR
hsaAUvgBDGwjcRJ92i83HcTFFAMbQGFCsZS05tYuQf4UE1pxeQg+GA8Qi5xZosdb
LwIw28L0h4808TIJbUWW+WIcuuFY8Tic3j5ZlfYhPumiVI9UV5H2Afpu4WlaWhzG
oqv8/bkDnwGYrYE18INTJ5hMZd1XRVR6H6c7/2Mt4YdAOfyvvbb6kD09MSg2NGn8
REs413G6aufSeTN+9Yy8/LFmfJzdkmgtakrCTalIEN7Q5HmNzzryILFW8hmKeKg+
fYtdQQFU6DcS/7U1P17xifB5BBWTaf5ypUP1TkoyvwSa6Si+7Mu4zJrqG2dLX6Rh
tosLY9+BnuuJ48S25KQqmFg8LbE2UWSIXw+g/apyUk6FlHH3QjN66xuxW9IR4Z8h
UFQvghMNBIE1LMYCNZqufveUFj7UVtlZhVbm9eJ9Vc/k1soxCvkFVrxiyKaWVGZn
4JNe2j8q6SJdUuOpGLJQovIjGea9xPM4wf2EYdKeQLdXgEX8m8Tc17ed7I2mJhXt
eFKMISrPF9NE5XWBau5ePcStzBxVVEyjOUfmB7D5bdyK04Vc8Z6g8eih9LBX7yV0
lBxmXNNrY5//qQvIhCTW0/jwzMCbzzDCf7VREovJo9IsdTAXmodrgsLsMWMhiAuG
SCT6Kpp6To4DzMLnvwSmucE027NJ4INEUQo1iQt0cUUf3/ylV0lPaoVKHvS1gnzT
HKVMvYAiX/ZnWSQxqTfpIoT2IiDxYW98ZL97lGHbsPaPy9L+U/abE4WIm4qH8mbL
j34m8FNiXIN57govKtBPOentOCVMRkJEaHMvXcQvR32QyaMe/ruzznaIyzZlGaD4
v9sDHnGwChUZp93ii9WFp3oPuOOH3QHQivtz2rTMvEKoSn+vjWYabClAr+i+Tg9P
SjD4Bp3hcsu3dp4dEcumQ0Ga7x6kC12hONL41JR9CWgUpQ212RdozpHdNFOtFfK6
tuWPmGqHUNrU+XVNk4zEH7eo1/LXUMUSkR7Aj9X75n1lA0fqXuUF5eVzbO2WhXu8
yIMhPsvY7aPlcl9nhYakA4p9nF8EwqbQy4kRIAFJ8rkaCF59uo7yY9uv0FBTyBK8
XIpfw4AY3Be0qJ9w2MUFfHYEY1o89M3gPFRymvblaR3hJEwq7wO8BFbwvUYF+2AJ
AryzfkwBqv7OzNJDTWUx4SHFSBvGGcP61qr87X1mF5VjvtsDQxe9R9lqm0MoD20z
lz+fwUJi7gOpeNso+qrTH+Da8vCSW0zPfSgpxBYnNeSjaaUUr0hVuhY7+U2Grj4r
TjxXpsWpq74au37c6whviXfWMo+Mxbhndj0lXVQfnQHufGPp2oNpgCf15ZUcp3T7
Memtxfu2giYHJqZ1kCPLM8/+o89SmK5xGeF95VgHOqcojCda+mqwxzqRXtK+f75Z
RYOR3szfPXhsSGCpS5T6Ar4svQeAeyRtg7ecm6KHO7iNueXRwkgQtJ3yd6U3fyuR
Zhse8vN9RKRXu3uw0SEBJiYR9pQDnlckcPFYq0mwqinX7WvMXoQnfGOaa71Y6D07
S52+qkHdjZYSerAilt1RdAi8D+TDN0CD/eX089cqe9/t+gr+ab0y/tokm1gqrj4J
PJ2z8BMnJVd+iMMFjJ+OPbbNQWsVH9o5lk50U4cDy+ILxycmnXnQSqDaNYi0KLzn
O3jPekkCHqaCMiSUogEYw7IFiJfm0kKbr84Q5PTNIvwXFbxQgXVFhDUoGE09D1u0
TbizXZ0sM95d2/MHIkWIghxcHMDNKOLkje8HsRxhwF3whTDyX9UAhJl1q/xW6lMF
yhD3ctMVB5aE3adMlIxegNod62VkZ4Mb5PeU9jVbtH5bo4+1fCyWTovS2vqDIkSz
iDlLAEoqTlkmJKdCvaRdWTyP/PpZROv38h9hry0BXQln2sIcty0Da3zASa1/dSWS
mzO2xMV9RYa5K61hxO+cksQsN7qquY48v+Lc3oZmiWnvEMVnNhIf3Lm80/2BJ3zL
UfAJW5PTNrvhupO0kUKqw1v2oTggrOJKGaHznE6ut1X6bJzss2TfP00/d12GF57v
sxklm36U2Xn7zKlI5vJ9eEhlHFQESuwwm+dK6G7mtOjIlBA8o5sJ9K3SWw3V1J3Z
rKkrszr2GKBPXmEmNdmS+5APujdyRLcs7P5VbzKHj06hyFLh19TO2B6Qij6hUIM9
R3z/yxtsMsGNHn+5Y5jCO/r8reVPOQo3QPT3P85iwgvKMl3SpGEWhsOjgMux4hcs
XAGC2QfYpLwbAanTzTL8rw09IKkVYvu2jZncXY6iOQufF9i8KfY6vHTUhygkFhfT
+Qnmdt5w2oxZrcVE3Pm6+9PCk4CbvJhX2NVhYSuukRNuSn6pVI4uPQ2RpnGWmIos
xpl+fVrNeysxTpI208aKYVE0LqX7gBEoZA/R/XrXn4PhoAiIP8dwXVuZ4XhxuSOD
x5mICRU290SDO3m5Bi9k05nGUkIUC/4rbHNMOJTXSUC44kwYZ0x1x0gDCow3m+Gk
7m+p101+A4wH8QJsA2h7RLnsKRNuWZ1QDueRcqdDhBQNdqhYCc2Br9BiziBdJOtr
QNmBrdc2vZGUXpS//nmFQEBBkG48ZKnrnq3dK+SdJHPkmSpoeiagPneJz6oP9ZpF
M//CbQThaN63mHfLGTwscwoO+Upig9IYGfmnwSHwy2SmG9yO7RujGu9CGuH5/Wsa
fAFPNHVXTWb83OBwdyfqz9O2X4odNFJlf8YRrYYUKzXK6vfEHPCa5VHP+Cx+nDB4
21WFhnneLkLb3gpSUcUuzOy4GDtlfokuv5uWaJpc6F8ylxTsxDpudWvbcBcon/+H
dJG0soW5GjQRYBY/YEZlV0TOipAGNNio9M8D1TeE/B2gadIy13FsoUdRjfMV/vFr
BD5Joruasj1tmwvNmcBPeoBdQZn8rFZVFd6YS6VhaxaOWEHPojWsKfUM20S9GfPp
L/DLw1PQRA2SYlUmMT4LwGJKsCdcDjj9Jw0bsFImD5Bgzii1pMj+rXcgZYbo27jp
jayXwuYY0Cbp2b1CWTMJU+Ua7J1EGyvG/QoWyoF99Yg1RuZ/4tLDslu9hNu3iR6/
AsOgvPIIfm9hNhDx0B6GyVCwqaHLCH9ex9ud97NIoIPGQCMTxKsHp+/T9DHGGrIC
Y8aoUoBAABJQWvLFpQBGfYXANfU4wtbEgeuUNlfr2f2oUyI0AduLECyzt3W/PEI2
jOBjmpcq5Z8IIPhugu/2UoeG7soRY8ItW0fkmwCaLQqpVblLhM+alU+8vbTVi23M
u3xdyRnRMaVbXlxJKrB5/AJq/SfxnkeN5dm8LLO7UnXinP8AAEWlhR/N/V5WKSMZ
haohW1scPZVh0ApXZqRW4sttQRj0Wyng/XboKontpdnbE352yv1OcOVY9KymoACS
Ok/MKfyR+WtwiH12qaWNXkxqap9w7CCRsBBHjHYaizljPrPg8PdykxTPgsbRD4SA
WpE+/PxpbZZryv7ct0GuQkCzWgeK348r36tm1BREU8bZ9DnLdXFJ5FHJ4IHCICrB
i2GpQd+DOL3T2JBc0VA03cImMoAVV42xnoPi69lCniWGAu52TIdEVJu85XbSQfzD
uzpJ6q9+yoTztd9D30Dx0HK3YtKRuDrwQpsMfLzQl71yFkNQASQBsyzXnETzHDBi
62YO0uiHFuR37VI5DTKNUoTzIpXTIIllJJyUzK7QUGhpS2Oy/OBChGv7XJXEQeX4
H1rrvUoR4y4MQ7UPQyNHMPwP1CEwV7eGw8SRKnJzFXMAg74lSkwBTJPtf7KZ6nfB
kLxGkDzHFoYb01bbJmwDr7X1R+vXA6vqxZEptQSbMODS+CAVCUDYrLokYeYWrEmt
zeaiGl5JJKcOKovlcOgKS35t8z3nA7BJ4Pt1ZO342C1YJVcHdH9snaoDV5MGVk9e
L2XsAn3p+Adf7EJC/l9reApAC5vPIQHn07Pe1t3X/kciu4o6aIH5z+b1wxyAaWnN
B31gwbMGfjzIC4g92Q485yakGf1+XloKK05xXglOV0lq2cqdLcL8+Lgt9LG0EEc8
4HTAE3UT12f6ps/Oe2ekhjR/CWgF+AI2/nlmVo+NP5Maw4NYgb/NtPOPRV+kdEv+
toyEeKJIfR+XgO/4spxsqswxZM09xLGVefZMUB6b9vJobTveaJfGYOhIv17WvaNN
o9qoTPilYRrRfO2WsdqK8IvEjpFyZJEwFdqNaqBttcuZxChlYsi8QBo2YLZurscN
RXxOucT+eoCOshAN7/vsz+ul3MqXiMGxMO6SblsgC3+Y63AbLN079rHwOEAyDovg
wop94bG1FICBSJcWRKTXnpesCGqOCkuXlKj9o7ADxeSdramg3vFceWSvko4xLb4Z
nCNZFb3UVGKp2qB04GBFMGBn7tC/S2iO20vtN4+ph5jw+U4JS+B0/dOxd/LRCc8k
sL3CItXKKZ8liqXeZkY1aYLLFCMhMIZw+5QjVYorGlsyRU0FnYz4AG7eOiCfnMUS
MEb0fahYTpVA0RJYGGb9qijpFf2HsjkhfUZa7y5ZUup/6QryJYymGPWlpjE2uInO
mqqLUPIvuJmOwDrizSFQnIXQQ+p4ZhkzSW7GerGwU9ikTsVvWeGV7B3JO2lJzl9c
/0ssQihEWp6X1CRfsvqCnstMYHvHtLCBg9Pqe2xM7YlVU2dHk1vVe5OX3i2pckCz
PY50T7ICzh+5t5ekppuc3AmTEDTcSESRngVdeaejQvG++NawHFSL2/X/vih2M7lv
dVKBtkzzxH+iebCy4V0d86N76xsGcubPXeWUBru1YxmcFTNpKq39b+31txF7N+Oe
YSSWDN0pqKBwawUN7LVNxmI17mds/dYbzwYsxD4KIINkrkzbYqfoDlU5/4OAsjHe
LKCwGUnY2zqKHbHniE77AMfpR2Q21J8e3oVS7Yb/X5XmwaFMt5wUckG4b/1b4JeU
ezCo6Xkx9fEDYETWV4FRlkG+hmgbAjguR3OfrmJrO7YfIuUaxGENgGWHKk+lTKmb
ntbGrK+R/asyStBpkwkupv29phbYvZnEyhV4LdlsHsZeXu5A/wm8t96TQ44HTnG+
0LngVVNAVcEl69/Ql4a+vrBTbvaZJuYPL7w8inTZichf/dlcRuMycrrIw2BL+BY3
z6Vwa0I2i01761Rzz04XdZwUtn00DRVuSSWYEHI7WtWAcZUtl7gIh8QNyYmhzfyS
rsJ3n4v1r6O5TknqwiZFcA3qNoFEGsA5pnyOVG0kvpcm19X/JXzvTeMCTbgCIBj/
BLlMzcMt9hfKKjobycDjFVBg2bBju/usxepoQyddAEtp0nexXvVR5N1c0V37OGXE
78I7GThf7h4TJbqvt6DPgCtq5PcXjF80n+EqG/L95Eonehb0rUbOlo5DPXHt5Byp
ntDpLkghx6Obu1jV9hHZYbmiiRoamQJLIu7w+RYRzamE1JUDGqXnH0PlxubnrWF0
KErfrEk/hlFI3L/kF6woxgUMEiNrDM77zWjfgHVxp7T/ORKYMtA2lYdKaKTN+3NK
CuNcar1ScSPYkjL+POOUvW9GdFtbNYtRoUTFS87AS7YyPZblcwZF8UzotblJttaE
GE3PF4ZsrGlIyVmTcxVo/MzsDtmIu253pV0R9F49QuUKl+nGZUJVV1NPCGS66bAl
XtH+78TxJSg4dONocVOcdYcqqisqXGLsLmwOLfrSkywI3rgodHxtM2NpfyRslVVD
VDV87z/laObguial2mK2xQ4mYO9f1fyWMCN33r2Fv/wnUqIeobBgGP4E4GEPyOce
MfsGXpjPDmfo5j5CTPlpgDd+VJv/V11Tu+nYfH495yNe7aA+vYhUCKsPaoUjuskk
dnLxRFr+cyJkqPq9jU5bBC85utqn/33GMFrVpkk3xOecox7j++0i9eCi13LQJWDT
vHGmWC14s+6ktiQO3mELMWJ4NoOf992px6aNVVpLX7zfUosO82IXrou3T6rBQIw1
8Jxu1Jenbjpuu9ApsFaNX3R4uJjW/mo+7lYCYAFuCkOu+tQHbw6UKytSmk9tFUvF
5/xurDhUz81F97dsDSW6R9soDny2QbDduolfUlK3gSbANK0n+HXZccLGIpJK7qLb
115/UaiXwOE+8NaWDbIok0VGNX58iZeO7zVeuDv3S1wEwz2yCq74wjCZXEtNsLm8
Rcd+6Kt0t13cqejXWK1vdqDqsNRM4P0QVQrgFf9Lb+uWuWZKS4BKtkAbWu9kH2kG
TVs7Yc5Nb1yl0M/CUMrUjF67BrtbCqwFvGp2xMRqD1zEUYADgQfdXGx8/S9xZW+E
iEppUD9y5APev8GlBaWBJ72KJSElShCNeF/R+UT2VgxKlGstDmtVPp28qIOj9FeT
k1AZNkuyYCqqwf8vdmtBOSqw10vQdxArRfLajgf1hxG+U/e2uP7s95X4lxmsiNCh
3IUlnqxeAbbkyLJ/G1ImkfJHVbqpfdj4kepREZ6oLyCDqyS6N+keWTIgem5vZL34
XKfgQ51apJJDB2q/kUtUSfbamLNAXksHpjtd/WOO3F2h1rsIgf8ZSRtReOkTMuYs
qCPDAqXjJuIjscQbG05cN52Og9n/yvqvRSxduUHfr2xCvP0kEEC5BCD3flal0v/c
v4MEhhsZR6N3QIwIphmrsNZZdkW5vVoiLwlfI72WMxcFcsMVzdTenB8/fwEMBYPa
EqL9rprkViOvb9UOamdE47obGfwfesZhu1Ag5KeNDxEkyVOb8IkmT1jnEoQL9z1P
j0QkPMmFTfB/StD46THykengP8tLMDblKiQ70bvp1uSj1ir+Rkp0lY7npPqI812/
HGXWW5s7haLYdhuHVmCshM8QNYGl55F+Cm8RAEz1iG2wmCcmm42JY9GSzcTAuyO4
pRu/KfJOstmSsz56e5idXTWkXpO7tn7LIphR340XjvTduURuYgcsINaVBtCMocoW
REMVob13mcnB45AE2e81pV/A8du8Opc4eSLcMd0qFaV5pLHbQ0OM575sl/robltg
BfaMbNDX4xo0XeQDcRyeZQrg+49TKiWSf4ADyTsSk5nUOpeW6D6p36KY07dyCIZj
Ma3Y/gYoSfkiK+NTqJQs364rltu1BtNI3fobCJcBVidZTohbL1j9yn64md/98bSC
XbTNhtR9fyqwHR/I4h+g/ErDiIJvZBijiqFtL9ZnNQn1+bCknJyXJ6ZSDXkIkO6V
x4SbOMAiEU7kh84OR0VSelShvNd5Wt0Ijvvn5A2KiC9X43uhVSm48JoWrfmGtez0
KMMXfKl228xrkL7WJZ3vOFnu2XHBEH6UduppaOJf+Ol/i4NulUIBBJhCTuvpCuMD
u/vap0kgLy9326yaBnhK1XAL9iX848WFtS6JfmwgXXuC/seSEex/+hbFt/t6mFfE
Yn7ng9jf70prkmMO4oPRKvSuCXPA/QHljE/1g2GwyQACAGClcxARqtAnYWUYDypY
RIVnhu1t5F42awj1iZs/IBgVWLKPCZOjNQK7XD2E3igGGNJon0ATlwnCGJS7G9rE
Fa9751w/86bR4L1iMLwhcII6vck6OXH/+S2sg4NpuXIjUTb+keX8+j08XXQC3i8J
wQ6gJLkX9b1YBWNk/1uIrF+TyyQRFFShqmEfKjOrQMzBoVqhC7eWJA2kzdzMkBUd
9XQvzeE1oY3BfJK9olg5nAdZehg8e+yIxpThgVFkNErxYRwRcuZeqG05lByw3aJB
vY2b5hInue0wUjOpwrJFLxB+4MBGTTlGhJwKi0miEz8RE3fFvhRCynwYEeWM/CYP
QFZHu2SGo0/LeBAXHyDMQbasCWys/2mQQ0I+49LRz0Vu84RhhqlKhIkizSZAg/O3
kViEiQ5LXfNlzZRO30TDPdQ4WaCFqHG8IzQTxlDqvNr6TDdDM5/Yr2RezPrrLG27
AOfGEFkhih1sV+/JvC0DJTf7d9xNuzM0UtaMMGMwnqLkxpYwhsTnwMXnhbj9bLyR
2qPfJXU3TjcVIdpADLSRRh6a1H7Vt/deIquG96LC1f26jIdnYzYxf3QAByc+PHN6
Ws2LtpJC1e/azCq15mzL81GNwAREZ8s4fppKB7HS8xlghu1Lq+JaQ2IyhXxf9rJz
K8jESL49WGulc6glX/+y8ckTRHuoxe/yJgxT/mt9/Bq3Dnknq8DLza8xjih2nE+A
uEG85x8VLadYzFteoSSTtMx1KTruVmd202qiGuERr3wu0Pdm2fGZi+S2TefAkYZs
0IupX0q2cbAmkMmaTRJWW6c314v9WfPa3BelaLNW4KWw4wQln9gxEIMg+5SQ/nxQ
Fd8tzgMyGCz1hTjNroPA+EFsPHthjwJI27Cfo0retTLWZfYp887aU623Re4/eKjm
4ZD/IgiLfPFC/ysTqdmt8AZN1s4dijc7jNJKwk1dU4jjSXoHrUavaJZQ1+IJcGiu
OJNaBVoKTP/D88gFmAlqwpA32q3V3kb36pOIVLNp6WJPZrWCbuWjJlX4B7Nshh4j
gw3FNIGeft5T30q8iEWyMFB7uKQSrbEVsR7+NTrZeoN7s4qKIBIVJLJ7lo7Az8Te
UhEB9Tlf2qErUq8XxF4uRz+hO4xca/fSxieJVSLN4izwrPIr0UkZYfcSXLxBNOhj
EzrOXZA8jHyUBMpWqzD7qo0QnlWs9Y9N0sCNonz4VnT1FjpyQBTqKqqBR67lArBK
yN+RgFOwT9cnnY9f3NFchrl7X3jNLQMg1qNdagdPdshv9aQ0MOZ6JyYHGmxaFXQ5
n3i2Mw4k3mL2DaDbedSxzG969MM7VQOX422BW9i5EakKLrizAqY5DNb+Uk6nTsPg
bHoOhV2cyAMhO4rF0SI/c9zl3RzAXC1iXqb8aITLfuGosuOu3bH1Rdj5WBjnMRyb
gL4rxffqyX91t1FVo3aSzujRvYbz1PPery7DzkP+RXF1vuiSinik7Xau86OS+42x
kSf/o4GlrSB2+aPzynb9+mNzVTotqqbmrJhP+U0/xvoajDjWPW5qk+f661ScNGEh
HS9iwA53ptK26XTCAgXd9BgafjfOKrmhH4l0ZixTyfdYJelF3tpTmJqofMQY1kEG
fGf4vhpAKfnKfYx4NtIOnGaFk75/2v1JLbqOSKQPFkAilpEDXesmruCRJ+paWrsl
xXA+HXod5Ypba3t/ysPoja/lDeQ2X/fp+N1Pk2On+pDTrzefvxk0o8Hf0F99igWL
JHr8/QRHPbrLLTw6ecvXUH+swpWql7UfMbYF9Jr7QQAsrjfv6qNbz+U16FCAUybc
FeEK/K2fwOtALGw3EdgJfjECrfJooHoAWNd6KfZBSwROT56MadOZYvauycTXFOlW
A05a4kJ9wgZAT7sKb1wrEXwERs90WWrG4RBVDbqSxX/ChGKEVxlSs0sMmJUIv0oz
cdaDDt7139X2AP8swrVGJRVZx1ZprZF9UvsUXGZQo6Nomi0THNhfbWiGULBB7E1r
bbt9kYw62YL8DzESLiBGd43HQ8jqsiqMVI2mM50cStEmZRs9TJvGJTCwTHopSNA8
qXFsHoeF86BffKgwAreZIIZHmemMepJvrs7f5A/nWmKSO3TCiGLXLx6kiixADggs
mQALciWdOGGPQVEeAwPOKBqXkQlEa8DhzNhcURFw8QJI5ThdDeEsOp8yv4z2zx5m
u3AxH8oQ2lvgLT9BaKVS7NqbYwlk1fz0fkZI0obLL1qJmD8iOplel2q+vzhksQ6V
c8/lkgq8fouIFxt0EWi1oTiS5YIz7mRTOl0sM4HWwFO3h9aUYnRuTqfbUqdIeE5b
jfZfKr+2JB11G0SQXYOk+P0o2csBmnM0v75B4NHp5Q7c4Pe+/byyZCnakmNvTQ49
q1ymL4O0MPwyMjnSHg5gM7jy/boFlQM2aGj7nGoETeWh7wbLdpuF32Qs6DR8EkSe
hQ7MHgO4rHg4Uimf4UOQ8rxBaUjgSkVH0Kl15I8QvkGZoQJA/dTF9567StejsD22
/YYlveCnY1uTlojhFXtb89iZQ/Rxz5+jo+xI8pfZ6VID0iwQ7SOrCktpIZuGY5kA
n/81P3wA4AnSzYlSAgG5sJ/cJ2i6VwVGgJSCkA8h8HhW96/XsaQSVAebaRcdosqG
uI2BIzMfpYuUmGryD4TsLWTQ8boNt7I1s4lmRmLfPNtdV7TNUWTLuq/MhKUSr8Ho
49AXi4oWvlnylPvo37QqqEQrs2wkm+PgMdYVjDevC5ocSWXtAVXUoAR64zhr29Q7
FQxm2hKZHYItP98OEm9AZ1a58WDYAvsacfdgOi5i79y4Ge+FxtHi694KD865cpL3
Vcp7qO70RPTTnErxDVCbFj0BM5xgI1CNkQXtHfhtYTWWRMZZNSblNPI2NXZcO1eB
WSS2Iw898IT1RJDG1nc860ZsR5nLyCAJlncs3tODuUUmrC8RxN3UdQKy+ZQvgi/O
jpqLsfCHK6QfZA2RXXRBbpIbXvQ7QXDouxbDPOJTsNWBn0dFYrMb1atvaUDRXhdO
x+okXWT9/eiE7QR3OBg6HbwoyRzA3ply62RyTxKyZ2TgGtJPilPx6DcX0jsP7+N3
vnUJoZo34X0lzH5h3gPKojgAZ3lJ5GwBwArMS2mxu/tXHDCCAfnMWCXqDsb/UcG9
LBgWGAxpc7MV5Sn29n5NuWty6aHCo3+qZZVvkLwxlhMCiHDD7cgmHp70Ncf0bMU4
luNcDnjKHK+lyfcF8tzj6zd7nleSEWHows+ez0uuwmjzsSlYboJflFGdWHkfTRyv
KkblIpmR2+CZQuMtKIbLOTmuJG1oq985/C2jI/4KMrysXYb+dlWP0bM9JqNdCX9j
5yFXsCYnIZUymSHeIlyAUQFaBVc5xWUe/6xRWkBGQW3Zzdz2ojMJGAjgXOylHgJX
J9E4SU+lwXlKrPxhpe/xV2mLrd2hRGacNEdtC8/5212k8j+t8sEGZkMQ2VXyHFiG
x4EH/HT2noR4Gt8VaOHaCi0lsLS1lD6pEhJEOC4WLthbvbmtGohLvtNOSowpSA6O
ayH8EU+PdEbe+Q8UlvUcF8/6d60cmT9DREchMmKpgKMjR0pYL/zmXrT1CKJm1xto
SwesvWMoCNzqcfI1ThB5y+LI4Pab8HrXe9FhyENqwAWmE2p37h5gxSKrIge4JJDY
EnmnFuigUKGHReZSCdq6RExlQq3wtRdQn0KuIx2fKMb89c29c8DiySsFGcIMUeVE
yj6yQeGD94f04bTao3I74990Pq7oM9Zll6OF7ylafYhy70Khwa+kujfacWx/Obmx
Di/S2blsuPAalUpEiCBI/t2uQ0i5gHe3YKF9Ao91VNClwL9Qn+phSwPVDFSu6UFA
/prhlJTlLnPahO94JchF63m/Cmo4P35f0Rxe4YGG40DNJQMtltZE9Ge7VKRRTw4E
wGwUfKUPuIAspsIcSp7LggNTm9TXKm8TabH6j7MAFIONguQS5SeMqAX9pUC33YlZ
cWhyyAOU+iD8lH9udIahw5cIk5bcMG2FeYHInyMT7npU1KhpbkBRcEajiBQ9ebSS
UsNTKGGY9zi3XfdnG5IeNhFftgTTD2Kdu/cGIYV1ZBRz74frzYhQ9hBS7rW+72Do
/tt4W5aRaYfLRKP3snz4artj2X+jH+FVndaZA/k3yRlfZXvOqUiBg0oy0kinb2hI
dV2dETeUVlZ7UBHHse5wJsAWZFcZA7rd4TF3940r0qEALe1LX/XPuI6mA2hGcx9E
YRD1C/452FrAnOk0YqQliAY1tkvgk8A6mOq5+r0rclGYvFAykKcacU16gCdmluyU
9BTaS6Z52MwzwBr7eF+mZpteOdT3+EtOTHVSGkf2j6zd717pE6xtd8W3mo9oPPkn
WyE0qCVBw3dlGIIkRCpI5Q+nLsc23WOQi3VE6zJ6U50Bc8rptgq5idFPP8KtGKjs
bHX43RAGazlsGq/LKj9uZ/vvRvBWjU+VHavA9Qt4tgf/hkdEkH2ZCrP3hDQOX1Gj
/KYcAXi/7pidNzxuM2lmIE+rb0xBBN8nw9vDb8Ylhy5uDnRtURIagQH0IjpVrxI5
bwnCbIXOF215l8Wu+8Cat+gx3OgUaJim3l6Itz1inRH5zueIcvvxNFczU1mt2qzd
ZBSO+e1JyO3FZe9coLmgnbk9GQV4A/fmFpVt7GjLHeb2Ii0DnCcmRSXfFru7bZQr
bc+n7Jnb7u+9ifspFAZvVOMrFlDQEeUPTSnFn4NMMql+y8fA7TNSwbAMET1lMbw+
38wY2GfelPdpAwBJqoMbl4Vm+NAA8ZRq+8TEXaY1IEIXu3QF9So9IvavC+NhlO/m
tbl6EQ0oG6wA8Lt/r62wGUdwaaBolPPrt5qsmmsK1X7DV1QY07JOwOrZgWPfTEOZ
EisQ4MOCnnIgbnXZ7zHRun1DonFRn0V1CTv3NOzcnwz2QFMM3QofKrcGUS0tzCwu
R9vtEb8x+oOQlCPRikKx0vwrshfTsZsoHkkUB/2SWJ707sMd0v2LgiMILPMZKDYI
D/mFwetSrbzJUKvAp/uA+qv3XZG3Obr8QlPFuAWvKe/yXNGpGZCttrAIkDJO4iIy
p2umGoPMc2WuG9bCguUMlNJdfBPcdFV0S/sh3gfuMVTGwU9ORwo5vxVPcg9NPADU
3MGFGXdbCsFKnL0Ue2P5agZSjeQzuIp1zmigMiBbXv4u9qfVcGAmwN8oUhm6iqNW
opV2/ozqzPSdk2MqC6MtG2v5+nRZtl2NdVD01f5AhYJeLbTlie6NEDKuVjpPvhjb
Po6YQPav80Wjw9sWTWOhwfYl3AKh1MeIgLumxBTey6ZvoFcuDC+sognUPihP3gxG
65mE3DEZn9CeN3M39g3ZI9NMGUyOBq8M94+ZR5vU6MPJG4LCYrE9LJ6UJ7PfLMMn
pjyQfHVaQ22Ek9wjHklsVpWjyf6iiFnh7echeFAJchZkmfrand/Nkzd3yMGvjRvB
wCeDm+75eNtuAxxJoIH5vGUW8xvBa6M1yZnR5DBNSHWa4XOE/rzrP9A/T/4kRmr0
KVtLFK4OgC9hh5H003S3A9K1Mo1UZsXfdsg/4w/i9WDYtqWcwqMFuIJybWLVqj+Z
wVDDkPckXcw0qwOQedtmt1zWgBFf74eiEC/+QaXrm00SdTw16C0PwXjDY1nEHXb9
0alPoiH0z1vCC2CLx4lpuSLQkYqHJqQpEPP/IKb5DCs8CFHL6whdQx68E1AqMOf1
dNTDyRL7L8n4QK8qFh+nKu0ja1dEl2cNY744lwEx0Vxy433ykUgt1SSjPZ136YWG
CsXSDD4TnqI8Ek6WY9PfRWXAECnVajx9ZtphsZkFKwUA7PfGJzEQpTt05uyCICQq
lmbVaDYq/isDQI0K9nfVcH/germp4GutX8easJsJqp0B63Kw+rSJjF2US4cMwxEk
9zhBrcE+dzCpjw968+a6h8QHmzHAwV18PFXWHmHlY3veOJvoPAPler9zgUlvPCXa
sV9kfA3C96MV+ni/xxL/8sTGYmLZxhaFNgRPk+/sfSZgjnis+DER6c15xXmcFGtm
xbgNfkCSdMIKdwW/Susu3kTLUbxfXfz88OsvZK0BqptrJPbOjDhE8f0BPZrw2Y2E
1EqwVF5VaiHFE4TA8j2stioljETF76wIKSjOLWsvEDHhZvs9uhp5fpJI5YPKnCdu
mr4hjCfy94URv9v+TPCuXYborBYXAUXUAmW3Vpz/2kfjue8oYDSEuTtQKEmAQ3jN
9ACstoSfQ5RI7vPPI98/H2Sp/PMr7qN4zSte0TGD5/GaHBSQKhNOexx+qKrqvK/C
iduQzS+2E9LyF3iHpe0CXzISomLtbUXsEr7t6BxFimszoP0KsiHfX8eNp9ETvAfr
CM3cuhtQ1hXMvaehd03lU/aYWW4J8CM/UB4gmpt7l+Vq6ibkSJEHZ5z3l0gzOFY5
uu7UHy2YTbYF+ZPokzmKb9YHj6HLpB2tISW7gm6eFPjCfShZcQ3qRH3tmW86Itac
zPkfTisoQYLQ7jOHeyRWH98wQyeYsZvykpnGqNbCNezderfLf070A0vd/dwFo8Gd
QeBaUsQN5se7bHjRacdkXFyAj0ovs0oC9M3j2nht8dlehygJ4Rb8xqexLzYISovu
lPH/GjeQEYlz5chLR/81x9bqnQM3hvWYTlbAV+Pvg+w9Wtm7mCwto0oALYXG9ze9
KTcwtolopx2+iLhXQ5gfGotyNr+kmZg7or8wgCCfIE2nYxmSyNP7ZnFAdsAy3oDc
CvjyvtYDGOnfS31DqPMbaCqx+xTdS0iGv7Pl/3Y67+0QHLW8UBpEPDlzVwT1BSeM
GLJzlDswX+Gw0XQllp5AeeMKyxmPQyNPRF+XBhNQUHn7xljbivuQ/MrOA9FiwrOU
RPzGKxTJWlosfazIsaGPULsEWUCOMRO1k6gkqOZVcfWytGwrWnWGILDHCKX8oKJI
XRAjR5zC4FjycAdvDg2BMcxhU6QVCbCjMLlUBz9e6Ruejug4Oj96ve2BlZTlzYQc
bzq+zvVhHKFIiISJlGc+2L9MgZWyeX2QghI7D/Dp8SmTD1yir1cjIHPbMgl8vy0Z
ZNT6GWY3ToAw47+m/vm6SVTgef2rqlm/qA/oUeQl2lHlfxPeuiUFRcEel1UeYbcD
Dq2LLGfcrbKuAGVmxXjTXt12hyae9z/lM5CAvu16kdlGJWNrSEXKShTWLDUzmTBV
EhPyCR7XK6Swc2MP5IRzYd3OrWRQWj90HkYHoXjg0NYIeRfwOqsuoo8jnLruoEiT
7ZmWT7bsYbZXDtExG8Un4LIycFWLznBc9NMqIvmFHWc19jH9QMYYsVCqvBj7K9cq
s6OtZzrgjZe1Fe1TNz6gCOlmE4oogq0aekxlInsTA6jMAO7q5OKw7PinZyBrRHp4
Wv9i5A3VyYQCyzwaUXZadkIaB/ohfEQ1nXakJh+w1SrsKNL5JpFwZsu0JkD6ocQV
tFqc6MaCzUz3y3Hrcy4FB9GYTmwMnK0R5TLqzaidnpjvBgBkUB6+SRtOQcJjqgI3
SRnMDqMtqbNTJ/Oe4gtcIlpOicU4In9TJDYZFtxFv7jFRhGVk+/ju0uGTw6d8khl
t7rNgz643C8pcR68u3c7k9tIipbzeadCXnettlQWDOw6Qs+m5aOLPM7BMTOMc0jq
9AB9OI9dAM3N1AcQJJQrK2gN0EOBdhicaJNZ/+FQhApmupnc/A2A0vc2+8tru/7y
1uTU83pv5yQJyaXKqJRENLhkQNULVOhZ1zPLpTYQqx/QC6NGHu5+QJTCx1JJo0Pa
TPlQtr9lf/km4+bnp/60+GfH/5wuiKud9wKUs1SlSmbb3aY8xrTNHQpmH90vx4D1
uGprGUsqGzaSaFuSmrGCUczQC2h67hGyWskWruWOE10PYifllaFFs1NSnzsJEemr
L10YD9VHpOf9nj0jwp1SqOw2K0Wj8ZDgkrgK28a0zPcvtjMmvsf8FDf8rkHsptuy
jsj2b1dETC4dTuFEgPmfaNCnUxnJoa6bgIVjQdKBfx6JpOp2Iq8VG8sTfywEVPVH
YQ8hyc/2f0ry80zAQcD7BsUe1LgeQc++eluWsV3LPd3nZCEa/qc5zXL1acXzGwbX
pM7OwCAwq9pNMqAE4x/ShQsYZeQ8cA72MAbXxtwts1JIvPCU6yt482ZxiMoa8013
1wViuOGyaxxDR3R5COC+sHCmXy+LIdikThaDoYG2sU2yHhBtz2LtzztwKvTIaA5L
p/v427EXWXf06XdzNA76RdLlRIY3wORpTJE0tNTyXFIMMKJCfadaI40oJ9eWNrVB
M/N1qcSQbDXHPccYs+j/Nqu/3+r9O9yTS8Xp140JFADS62rHKukRE4jSwv+wXQ3V
jquPFwlDMpsOodB6O5aHJOJmUVV9rFr9ILOy8heDX1nC0QdFj19B+8DCZCK8F9BE
6XMmLw/W0MIqD0Kg8pTpHPgJC7sWBSPtlRnFGUuMYfw+tia1gqBXmEhIt8EtMnuW
dFlRjVqjhfyfhj/LlTVkAbC8p7D6B5KDJOiyUMMecneqooWcwj8DNNrKy0ftBDqW
RKrSBVTylEGN/uuCh+44/fIteAVXCqGXTx7nwussT9na75D0/UvlMLWneUIzivF0
b+mzBXLJ96Y/8zv40XQOYOWoVvwlYaLwI5xADkMi7mIHAAIJFpIyCvVbiyMSc0gV
APiZUtJS2BSslRESN/0Czsok2q8FyXTV6TWAC+Z+Lkf3Ee25VroSvzAnO27ysInj
xSpFz7Mg4uCe0iaVZVTBxxFwliE6Iy/3NDmA8qh7L22pmH4Q4vK+SnGbryGLokyD
PRykibQDGH/bT/71hHAmXdLmoTdzYRPgSCKTibAu1qVQtgWMAJvZYfDneV6sAMwf
O1M9TW3TpeG8l/ZlFE0kPOu5WVdxTBu2gPnX0q14OMydWVj0z2ByIhK16E1+4zew
RRqs54UZvqFcKM9QzycML1e4Z+AEmEna/HFC5GVP2lZFOWVOa/guVUr8y15T9lgj
/udjEpuU+lKLGxS0G1JoNJamc/Q1j0wbyKEgDrgdctx0FAMKVfGYGcxMWrumhh37
VWfg27KxEaFD+4MHrUKxz/EIQgskze6qUgpFRKNzwCKp6o6q32j6yVQCjj/pPZ3V
ALUw1BavBVCOrD+U/Dgq94DHMZWtimjEGDNnqENs+KCQs15uS6EZDua243FpeRQ9
iVFSwBcKgVUBk8Km2OscUW61VbyW+c8K5PEZ9bM0ry6tJLH2odxGga4sDaWtJ3gG
oTKaAWimSIYb+D0/DxzU3Egwpkem9OFtc4ivlndfMYz5AX7krjEzNECJrndyw6jt
V+j8K/wuQV2U7TVfvvN6OwNp8ohb2yt9GX5pDOyRYayO8syNZckTBLHaxbz3/9a9
TgwGQoPtRf/n/F4w9K02BTKwdSI5lAl/cQi4RfVrPl82x8euPLMlMu2WzWLiFtfZ
DtqKWvgnhFvVwu7B8zWjMaEgZDm855GBFKS1iL4nTWAlCJOBDzzmsOtWHh37Fk6j
C7QBD5QaZj/S2mm7j5cpL7+N9ChhcFA34nd2PxzaNUiZDSOfABz7YskYVbxVNUVs
3USJnbKDoIH7/sg7N2T2GDa40gY3mFWAYaEpTBLy5jGJTseePA4vFzf+A+kuwhqb
5XShliGn6ALLrmh+7HFMBNOyzCVFVY6Tfr2AkN68W5T3OHZ5lYcF/fuUfMRC8IYl
vkaQiLewy2Uhchd/KaXrSLuRxCALPU0gC6HWAnpRu7IwC5IuTIPOyvoe6+xDE1gT
bIdPHQbStDoNt3JzVEmAmAc0gD1+S77V/QbYieI4og8vGJlxp43RBwFph3pqybul
QpqyeKOKIVegBbNvqY4hw7S6AjaRkTO+FBGwFLxmC92Phk+Xvsi50Frngagx9CMI
gKetYcXyDNs00itCqWNIEUqZIHhC0u3s2G+dmS4DskQ7ELR2luFfI/wDozy3oMQd
OM8nr9Nh/cd76Wihgn3haKBlIcSP+Zm4GihAGJ1rDfN+iGPgNQ6lV5H8UX+SqOpW
1rLWdojvfNTYpQHfoSgaX7+PchIzBFU14SoFLFOZ0dT5eV6lUmAnbCBDpjY26ioY
Z/j+C8hpDOA7zK7NwIsqUR26Q1omgKXXAntCVBZpZpTL9rQDLODHYgkk2MpCwb0+
EOPIyqbsj+sdp9+7ny326EqMtZmFXBUwJd6o3c7npVUNHEJGDzG+pupnJFtNIV9V
h0EnW924RziTeShNrzzb8nJATYjXBAfT4Q/Hagztj11F7iRrHj1Z3NOqSZB9E+Jh
K6sokSFmyp3W8QDmP+PasHU/xHJDCX+cFO3EO11CS6x4ZHBhMLJvQPq/T+rIBKuB
2n+5B+QoQpAM5wEGGYrGwTNgS2legJPjV0vJTQTIw1vGgWr+0YjfTAneqKQJkO6Z
4mSyZI5v6e8+uYMKXVf52F6bPEl6epZygCbgyou338O8tmV/l3pIDtGSp8tuaFt5
W7Cik3CU5tab3kzA7KgctPe7bDryca8mqtcgee1onxM6g4D4ed/qjzdab4Z5LIbr
KrwpR4vRsvb7WZK7ERVR/cei/n4JkMaLUuqd8MR8hGp5+pqQ6XOsLDR/NNea7ddf
AMDAQHgqkrS4s1HlQbT4KsqpRMdLBlLn0NB3amuAANbd0UT2g+CZp4ZSA/aj8+nK
hwImyGaUrM2yuuwlJ1+HJMS2o0nqef3/hzXWilXiUQj56cos7m/2eYd/OhA957CG
eOKDQg9qVxiC4wj//an17zKtfsNld5bRJbC4vUlfiX40jHx8yippTCZOGjycKqN3
k1tLVQOSmv/jFx3RQRnS+J45MB+XWW1iPQoEfNuV4gOsfg3omaxbXw0GrJ48D2rL
TqRbBjwJraVIhXDo/tajQapYOGJgVHFGbpjbaHrcooj7Hx+LrvThMB/i9zz+qTN6
RQiQ6xbhBDBqtPgfOA+VHXB3H7QRA4iqLSCy++G3tfruRgoGVroTSZ7Y0I1q1RHJ
DgNOXhVV+c1fEZlbT3PyAf2080DTKb1FG4C6cbLl2Ogq58ZImMPx1lhN7PdvpYwJ
u49+ltGRNLJebPjZPu7zz1K7+/+BTQio645uD/IWPncZv8ScoP7KmhqJOhR+DgHx
sdz0u6fNf7vc0y9z2/XOlOxN6zL8kgahXl09GvKr4dcoxMuA2joIxQxchOpuyZYr
5sXUYiEFwjzgcP18aibl579aUNiaPIRL+LaWqXBIGxiXIFkDyqLjdBQoTmJI0CK/
ShraweuIFcsckiIq9/n8JidDhS+gl0yacaeWC42leMkpcVmOGQw/6nQZnH2ZD/Z6
IEGYJ43JahSUp0puIkesX87j7O+DP8Tms+9gfuWVWU2VKZ5Jx2yqC+Co4k9gFS69
x5BFSsdD2Ib9lx8kR9qeTUx4qQKFvU6E8jiLdT58aytEWaLlofwUSChL2pvaQ7mu
46Uwr+9NHbODuXKDgm632UALybawBbu3jAEL2ZOjusl/xeVbKNTRnG8kOJbk3iQF
jzggDGFc2YzW/UA1KP+yvQ==
`protect END_PROTECTED