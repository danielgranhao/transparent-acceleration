-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
yZcMAFm3PLwsHMBGlPE3L1DIeWZ60dOFqCAS2nwMXjfBGqfCFKWYKEBb+fsZduVtOIhyNI6Tkklu
5qLZlEkCLWzTj1khxelgUqtAmr1O/g24LAqDQ/Zu8Epspr2WblIi6a6+va063i0LwUMtkiwyGQzm
FdNUcYbNH19sJX/nIBLhwt2w23jI7EX9DLNXEsN01oCutV2iLU3B9WW7m3/qzfZN2l3RoQn/8fhZ
MNntLdbummzMORorx6AsBZWeOYRWEQy6L7QOLT6mKoXKdzoUTWtJXKYo5V4ghABdVGv+5o2EdbE5
TPCQB7GmsCcywdycrDndJYM8Fv9jnfwpO0NIfA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5488)
`protect data_block
vs84W8hGiKt6733rqWBMp2L/g+Ek2qvzkasVW7jO9cE1wDjtSms/bTsTGh9ln6GKfeSxvtkZ3u3b
VmYCXGrUvvFKbseGzsReNk3kE1jRcb2k3iPLxNKqbNjBiX06fdZhk9KgsE3fpgIfmni1GdVtiPNF
QFFsSp/lZchQLrCXGne/hTKmbD2d2K1n7wIFJAP6dme5jP8iva02rpmWZONfrc0fpuqFfxmqjhFZ
OszYdfO6MwGUnOdQSLUv3L5298IpviLwYfx4OHPomehYLzXCmZrh5nwgxRDHnAXKF9DfpKpl+L6c
QRN7kVtWSVlHAr5p0PWd5WHNkFxAf8AeDyI/QhfaHh8+DJm1eShHvEwvAyT4qmY5bHYoWLd4xeHL
GhCHgCm3r07OUBR+eKxCgWHo+B50iUZPRjOm/PQf7ZXrWWd9D7xGISVJnemjFACNdqrqHLmN0gaw
ukvrQ4WuiNmXk5vymwwb4mU/aRTRuT1W+FOEsLg8z45be3TIhuP9m98/CjEgSpzRhJVeoNYm/rcf
zYkZR86OTiEXnYsHyyX7pmN+x7df49EE0Top//R7MhN1QegGWQ7W8UdGGTBy/visN9QnVq1yTwon
D/HX3XAeWaEa58DwQjSCBVlduzy6/PmLdVByjO2g8x6dKfz5NaO7rinhfvrlzMTMrT+hVWh5LVhc
XCRucFQNWmDZzv3jh5OEQK8uIK+Llciw0BhOBmM3mFN5azfI/Eh9CXlkhU64M0UqTS9ec2OyvQv/
I13md4Wr8BwvY9EavL6jBDYPF6VUbNoT83ogGkIZYj3J5P882fXiEaFbH8fwT8bFIM36e/rAjbSX
q+s6DPljrQLfWSdGdezHKvhmI8NTEgPlH7vP2JNM8iVFs6MVAmiP2zq8xyoRqCid4f2y9UM2eZJV
iiX/xrdU5WzxFlNas/aIIJXpHmfQFHxnqug8Q4XVeGVHuwtS0d74eFxz40vo+5Uctk5bsAi92TJZ
XiJwQZbMcA5uzjEglQxYh/SkIuGLGg01DDi1uYVZRGOVCnqo6kWRG0ZhdqUUSC2H5/CTet5T8SM4
0LlOzKNwr5H3Z7umh84BLRoESeyI9qK71lzGNdQAZS1ye2SzOuo0bUb98rPhJo7UHkUmmQdDqETF
IHxhdELSg3sV+ssjQcSjnozwPxBUPNENngH5Bd4E2UXN1PYB7LyNN/pLieD4NZl7qvjKEIwH/z08
E2xHNc3REzCvy6VbhsMjLUnmSzvE+o4su6GmTZSR1iCvrh8Wagr5Ju9gbHdqUnOVY4ykyVzG9pnl
eaZ4IIpa9Ire8nt8hYLj+Ik30u4EeFWJC2uo2EjQ2PMVbyb5GUG44jPJugjH/9WSWgwG4iAq9U/s
+JKSG6TZ+Cr57oJzgXbD8SwqkIlSv1GaMBMYJuVE9jtz0MxRapm4xoyn3gV7xEurC8Qwm7UsXa7S
8Pku7d/+qkTDgFwvWXKqZlgxCde5OeolyO5CDT8JhEdIHlhgtY4HQLXjZ7YUfZY0T2H85N0vdORy
I+kDwkHJmSKeMOvTdB2Bn2kntfvh+DeKN/1e8COwDvP7ftTAzJUoSdZqkrlT93/0LvfuQCfzzrVL
Sid7DUvMvh4+bc6RdqnxZ3TFf8trfflntsaipUaQB2rizyu3elcLlCGoQZn+pkhnFkBd+e3NDjvL
q4xxn67brLMBWSOiYs6u8IADwPe9du4kwtYL49NaSMjiA9r8NhlOH+7OPIMNLgF9bFJFk7ZPX78E
ehoBQu8Cx9G81PomNx9SwkYpyTdfRkG1Crn0aF+eo09qndQ5w74ystad7D6lt8R7NhRAizZIYQLJ
6hb0VZjLkaga+5OSV2MOJqpASB6+V/pXyct0enb9iv3IC99TyvWHhL5UBb7lHNc7u7YEk7sOPfbI
Afn7xSG3PX3jV9rDSEdfxj5EJE0qBAGT5OFv1cnpEK3S5YsEgo2s4tA3HesUWlLIK6L7KSFh2ANT
3JU6Z1nrrNDVmyd+4KbkaESH6z4jdrcjv94iqTxV8Lz5DGTpslmhfaLyOkncQiMIadeZpeSysDeW
zRUrH1THC/DFQgMPO1H3g3eGXJtXKQxnAA6LjyvpcfbPqsKW2btJwL/EAiaARaFZGzvSIkio/C/N
DFJf+TzZG7DuAR79FSqeQo6qTw33HY0zzRqHpS/AkJbwNjmSKuo5Oz/ZPN9S3A+bMmQ6rBAWK/Qw
SJk+6+lb8wnY17tf9J6yUe8E7f3ME8vpp6kulEqs29pH8j4qcFkm7bVUyGvW8w3a+dDLG4A2PiBq
Rf4BA9ZtQnInCbWdA3UGRlUx/3snysoi4ZPZKUFVhJKHMa5q0FEjBUevRFwa9Vtv0fsYherFZMgt
nBNasyKHtYXMiwFRPSVSAtnwmUrWoZWlenfD2XLAXj2GfvGZ2f1p4v7qs6/0MfM5JHajQK9mcn1i
w5cGnnli6Vm+MNEcxXyWHrYecrdhcz9YFHce2EJVEyOBKbXpsiCJ/d/MuqS0R7UQgpSdFafqr0ha
ReZx1qn5/H2Jpa0oUo6NifNfIYcCxzlN3+YAjhDN5wc32RK3ZcUf2jLrJBqlwYNKyEKu/7IMzRll
Hijxj0SHb90wWk9E/IIVEwF0NYdlcgifUlFfzmgk9KSCF74M5x29IEG8fi2mxpCmVs3MNbFEBbh6
k4MURTCBYVBenTMM/PkiKrC2aGmngIgG2si7v9wpYbLEt/DolVdXyR0gpZiTj0ZgTJ3IwDOLRtfO
g6N8nHHQWZVUU1W9loqiXBuoREriq+cG5seWBPhvzzUYwzUDow4zn4hZZnHm0TO68hKw6XsDOhSU
Ku/8q3ix7Tvv9ohI9fv/RYkeRMJd0vAxyEomb7fvc367pnLTSE79OILhKQHtVErC0TERJDd/0dMb
3c3mtqzDA8wjRlYQsOjGu7zq6dHnk1nHxI8CHgiHSeal3rNPyxiQ208WWpmaiB7cFKo3igilKNJl
vxMkzlNVDyNV49XFuGBUUgM0Ap2YoKMITQ6IPtQ4MYFKb3Jnmbpa/4L/hEEyY6aFnLj6bkFkLxcJ
wYQYl1y9nYzEiu0KNb219WGRI2+XtrUKwar/3g1NE6tENnh+NRQPxpM++SaU3kvp3N8fwk2W3G5Q
Dqps2PXzYhIqTsP1McjVuxQUSjsgsb98qHuH3dQOxSdA8e9EPd78h4zE9Qj+hwmTLp0XJxjZpcfP
zJAroKU8oqyNUvMni5lk7GCTXfII1tCw7+/kheU83lXre1lOuhu86VwQXqdP0epaGFWoTmU2P2s4
S7GYqIbB0G2aalLxPf1hDprL9l8EwWwhgmakcXEJcjtX80ALJ2hcU0Pykkadd1zgRCsTpXd5kdJj
X1nVss25R3AvuDOG45SB3WE51tgSAJh78aYbtKJdc7GOWIRjPMIA8Jwcy4mg9GP9lBsT/jsQFBNE
uMGAf5IAj4VPiBMPjwYed7idbK+WDjj7rPeRpBPfpeuOeaeLbYYRuy4Em+EgVoi8cXA/SExpRTkj
gAsaSzuWACvuB0U2WGkGBbGJiFwb8RRqcThEhvuw3ukGnT1+Cw7eNb2lY1+zZ9igoXosPxSREljh
XkfCCMx8VcGY4jFwWTG9pInVSo0muzSoCWmTLy8vabQmMTf4LyMRogw6gKU9+bPmy9czQM7KAP+s
YYpsHMUyA3gkWG8UhkDvqDoovOQgIYMcG5ZsMxWhg+7x17U0E49lc8b/XwOz3bo3j0YMuO6WDzVg
voZaTvPiM+IL/TeBObsfWQIa/PwpqylwMm2kUNWA2fGyUOQbkQiqTH9aTHAQWlfyCWuelo6nQKAj
KGLLfi54HAib9pNHg94cien3rFonynVWYfooidg2Bwz84WQ4uKpOV6r/hnquE8Ns0x+MM1fNE7m8
ub3DlHtg6LDm4d9nTcsguFIqqq+UZjE9Upgy4vtqAZL3WnmgQSZxbBNMO0jz2sCB0wkrFhaIFZvN
z1NjGJ8ZMBSX3sL5gPXHkj0zHL/Lu1mdOLb1aHhUiikqeePkDfUiV+SBZw9B/WWvbPza+4YtvDE5
C5aO4LhxyeQij/lWJkA/BIDpcJdj1Al4GAUY7CQ1qs6U7d68WL8O3q2aves1ua1beWb/k3N3Rhog
s3VyTw1z82Cz/PEIJ/Qx9uclmXpq81UlneEl3vErdy1M/81iKop/LG0LvuaE/LLEL0Wkur4jp9t4
QKT0SVvNYDYGxETuoZrRqFjIkL/GFDqm0Pk053SeGWyv5K3W9Yg+bRqtE3m1dILwhuCmF8MHoALG
//WOsJPfw3Vmr6FD7EqaoxHBsN98ar2hAFI40ouVupce5Etv7itQd7o1FMnrMZcPIOg8Pm7h6srE
ADcjIBZGSpbXzbl//l0tUkBuqxenCudYhVu0j/3g84KHG6ghmbDPZIz7Tqe+ne9WQX6YrtCDfyEv
cOGRacwMay+M04sQZeoHXKLtyg9iIAVchdzGI1DLk3y3xauOZyrx+81wDmHiX+ydLC1+K3DeMA5x
2h3rzrVpIcuIRgxuwLNOjOI9Y+1vlTa0+P2QhGjvXpj1NtvsN8ZVX74Gmy3BMa93D6S8qVZGDs8Z
gPl7EG+5gRrYoTGaKCzX4ZpzNZWRnssxYbYe1LgoQwOV10SRza0DhBWWFsHr3ofAE/XBW46KlDXV
kd7zuJTHJI0Zzu5ZhlVPPMas3ZMWJu1gifWS5vdceF9MN3BAa9CtCFb2ITFYbBVm9m3E04k/Ta6x
3A6vcYC4Ra/CvdxWaHZZGrIITMInc8LhRF1FHp+bkpgXReleKJpCYQ60K7W2OHw232t2XhVF9odX
wJSc6XbOf9yeCy8fPk1/InsAGgzh/LklH341wDfYOzPW7OxjM6kB010VC0cOFCKcvwf1k0YjWnEL
+JzKioXVoWWNxXzlX134LbXWO8cIP9lBe25NW5U+30YX0f2YRAS5pGyOEm/ZkCuc9hETtHan7qTE
VGptGMTRTXV7ILDIjEJyyrn0IF/ut5KEqm2hlNhxPujnCPOlcBWD5cfHDJzkp3sMtp5mjiaiwWss
Qkb56i1T+H4+nOgjwBGbXy46imcmI5HGYR2/FSz3x57C+A8FmWVP03nPh1RhVU8q3hFohShloKtT
PoKsdTLVh6nT97Hju4lHnr5gC6AcZscwusnm2TH72Zq35/vOk+vO5e0lhSF5/8CRnpptqnrhWJr2
xFu5mMjOiEHHBDEKD11S+6fcuvh/H//Aiy7heAnlpAohHRXKSVFdGcojizrwTgKMSQhtABzOhfzH
wbuHI/hZQ/OuH4JmVtnv6GvMWHccP5RQtcsUnkPFLkEnylRJNm7/jwmsJB0b7TPNvpJMMq/4CCuk
o7WoW1X/EkGS9dOXjQa9ngxAKC2b5R23UZe9jaxQ4nCs13AsvxmMzHSIuzqJgANrJo2MU/dD2ZRB
XcEtVxd6aq9qptmCA+tckV3wMfwfUX1qU8HqYG+SLIQVxfEEkJDl34XmB9e2L1wj/NrfB1I+gu6o
7CWvai4VFSU+1PMJMBF5+OP4OSonSDjyinJluX7TJkzlczZzCJHFGxcPWMvT35tS2944sNFju7Lt
kUKQM2TMGtR1jSOCf1yVpuJeiWU/cjHcgm9r4Q0YbSu6GG/zHyZge6md5ZjIM1iiVVm4HGZx3s7y
tA+S2x/hr7v6Os0IEZN0mKTExJZpEb7TEANnZNqUTCYjlKmionB9vjJ7HpwNCdDYVsRqb/9IW06u
7Dl8eAChFlJpMWOA9JQWgLBGprs4WHp2wEqIQrQGR8BFE2hWozdq23ROb0t27R3IK09CoooyzO2F
PJd/ru0QfA9mPELuBWglaK5hSn++q3zp359XRQwy1bZW7COiLVqZwb6UuWR3B23IWaLWc2SSgU8G
AFJfSwh6cBSZOoXM/eRLighO1TuhkCext2QnM2W0mS7g5KDOTOr2cyaO4KVwGlzoS25e3UrFQcsd
I97zt+m00kf14wuz4zoUGHjzL26h2qHdOckG/h+/eSO2Xgp70rEtB74lQuy0x7NUBBqQbipkV7iL
rstgtuvQxlAoxjOXzYK7rb5JIgB5ZRxgBZe/ta3jDGXZDMclwwmWpHXxt0lBF6V1PuHMUaRhzWdx
F6VEQQjwn4gm33+JZZp0HtNbqkHL5AzW6743p3lCLEbTpDaJEzpS8AwFreSGCSkDf2onFre8mIGs
Sne5cB2LHgwccvXF+dCJF4b3tKRHVQW0gjldXNVYFReGePLjLXY+dqkav2xcYnR6CfO323YbfyVQ
CvstUHlLBlqydR/qh1yQveysx5mL+5qAoffXsgWZ+e6sUN4Mpcu4sAktHr2Nr2Xa/nMFfXCWG0MY
N6XjNq5ipCr3kcZVtqGkQ1nipb3uRE97W3m9WoSBmBOlv+5jN+O/nly6U7VxlreGFGF6agCbkUWx
VvC1MC3ggmNHQ/TxHyJ9gSnVj0Kzd9eQXp/pcHhPRfNm48W+4EDstbIi9TH39vlK105KTYmRUt7k
KLymTQKZJKqsH9c7R/kwIo3J+CEs2SCZT4RMhHya+R5roIbhN+IXdSkLGGqHepvrSgPSJvYRRFhO
idSnqJFw2D52sEI+glcHOlzlOv3wdjNAKfg7a0TBvErHAVNzd/jaRILdebzcst5ZblBRenHBTQEY
ePO50rnkf+X5YxMBnzjGiqPh6SGjOO8r69qG+OMxZ0YNTa6t0hNkIr30AqJzsZdPuCS9rHqnBsbu
VbWrIerqi/GO64vUq6luuPpdV0s7xNTzGE1rUOGUyiyshwKDe6vWAyo5Es9rnwb7YnjDYJdFBHUi
Z4BKE3Xppn15RdXtyyo/UDfwxDXi1CwTcBar1NorSxRhIZDODYPzLCzdGGbkh3rl2SVGvS8goIJ6
AzNWDpex/Zqi7wJTQ+f8U/kcgWgzrWIVct7MZ5Q/qNVorb1dx7frNMk3xdw1zygJml5NGsFcoW5g
Xi3ryWJ2S+0yg0v5hqp6mH4BHRFqGdgzXaYd2QSutI3+H1qiz9vgn89fStMg0KTF8LG7Kt5ei3DW
yA4NuDcDS1dxUO8R51e5tHFWlIzrrjqgAA8dErAk8+7++d4dRNkdB8TkNeXYSkNzhunq3PLVyaLK
syfRh5AV5T9WtupEzF4Ld0rzvfOQL5uABNNB47HvYpqkPvCvfefRQO23DGqub/NnEvP/jILG0aqq
pLeKggv/MS2gRsSJV3mOkzwfImH0PhsUXFWzWMjIGXNNi4qJadHIIgoAu8REAex9xeHNGeC+KIBc
565bqyPuxLbT1QkG2nRVypx4Nrshm+pLK7Mt21kDnjsukZbRdQsKngo6ycht98BSMvMr5pswodU3
uiEyLiR5nLpNm7setb27Kg==
`protect end_protected
