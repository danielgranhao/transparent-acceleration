-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
aeznLeeAKeSc/Zb5KgzfO6DyvYdIZFG2VShn1hEV+Hm4doKqeXrCleT0iybKsXWy
lhZ55TvnRXJV7rRJkUbBnrRMDqS/6OVU/VN4gd1J7l8D49rNqi02+GnqRe/Nrgp4
YwQYU5Bxo54pWp4YX9WTeQvkb1ZTr8ZkvaRtqjGeD5j/xqeYnEbMPg==
--pragma protect end_key_block
--pragma protect digest_block
eoF0NFCvSa+zqpDS+q6s8L151WY=
--pragma protect end_digest_block
--pragma protect data_block
pQf6Ma6+qyfp3Sn+RPmnUCYT47mX4+ZW13XKIHw1hSWCLVWghALpXzv0p/6f0VDu
88ZZ3IPB7gGySwWL10IoferC8+zacxH1Mn8OOuVH48QakVCYAalhdSAmfWy4KaLt
cvz2flKcI0u7KSbagSbwVifT1JvrwJ6iB/WNTl5ggbFBXPVRb1XOG7ZQL1ZQDKIg
SIb5Es1l6geQn+MKNEBCLVKAkWu2iNlFuHM2NXi1sQ7tOw54CsBXqxczIYnA5fmW
plcsj1LtEanuJJa/EWbrPXrLBXDkMMnvu20lwlkaJKVcXpV0CWvkQ1tr/5cdBu1o
7x8Qk3l8Z/5uTDfhV6WKlSXXg0QS1pIawqq8+ui6YcdjntTZ1iFErgezwS0pjE9g
2MRyJmlV7Q5yqj8Y2+LEZVZb8kldV/QgphWAQA8Bp1y/lTBxTN0TDdE1flv+8Xl9
+yqq+TJW68xCoPI7oGYrsvkKzDSvZ1dCUA7hWBxX2NVcljknqJqeU821B/XAHEAz
n0iG6zHtIUKwpIIzCqscHR7YMtrD+TQNs8TELZUpFUhbiPtZINIBsDmjcMmQ9rY6
BYlUMPNb7Bnwf1hFyP5BbwH+VV2kv7aIkKpfAzNCmY+tAXxPotuEberDatdzSkLe
FzK1FTQ2yjFupHsoGzcwF1CWBQQ30nRSWueXRtVGvtPwHZmS3ZAwniKpmrF7Koeq
Z/dSOKI226KmyUYDhQfm/ouvTVKlVDC23pFFDDgB0IPeXLDBRK74n62XP5aiVW0p
AfgojxcYlwvTnYwzXRK44rUqlJwkL8h49g8hZlTSyQzGy/qJTYY35gK4/QF2ZgJs
lC/geLKBjSFdvipaf4IPTW9HwONiTQlZycAg3B57AwQFWcQTlpIqv5ex3JTQjLzh
yyg5C5p84uMkWwCim9UkSPjpgUr0SZWJsLv/ykySJcSLXG1TGZO8gMqESck2qfc9
bJmtxTH/DsONbgtAS7Nle3KXdR4U0pWDDXZfv+Or+IrVc0XVtEyoawFoBt0c+0Xb
kAVE2v8xi4/U/fVOUBu+Gf50xDLwq/B6IYWrYsEL7c2btvnBGs1ycHa1RGJh42JK
1Xn+NNe/W4YHqIz3l7j8KvDu7fpsrGuoE0EFrZoRzJjfovcZ+c7U9JqZfhT921ET
o68FkjmCW0mOdxfTxZ+BlIebZYpeCb5Zrmf/+DADhuveGoQvh1+GV21a3JaGi02I
tcfqkrEfP8XeFSPrhR27atWp/bJsZ62FwmTvWgqiaAEiUrx+EX05emdX2jlEo1yy
lwSuZKjFMMYlbXeLKp8PD0qJHzI1PhEX3boSMgQSiDaJ2GniBHgvdzneAgzbwPJh
WrztHu7ZxTH6XCMKT8oV7j8g6P3ED4qaTaKBS3j30uoptxq+LeTQhV/+z2wKpX0p
yRDsq1tYy6xinosl+fGmkDRX5UBm4ks7NMzX/Jj3f9oMvBfm/S5P78FUMYY6/xnm
zfg3pbh3r6mcRUnO9n5Mk67BZXcmkiORktwDDtr+VqQYERseR9McPs+lrgAYlP/Q
QgvSj5GGxO7pQ7NP7LaJpV7uti5AV6H3aQKVcy9tXjaJCgBihA/CAfaNsHUVtUO0
m92g7JZjRSsHKMaP4zMiTghcBljOPowMAMWc3NutsyfuTp4qjBJ2Ia4nUXpXtXiT
PjPT9ouher+cUGcqA42LT1mezTbfjQjfmHncA0CS+M8uRgeFtpElAYA+iU/csiX0
z+hTJRu72ie/bEyeXHPU4+TNipsXgVNEaQdvFLWsXHArLJ1TFcrK67zBExS4furU
FuyuOunnU2FKe36KqLjIPw9KwIz/urTbvYyfQkjgoDEKB7aaXzSQqcIg9cTxzHLQ
LN5wc8fZBAEkSWVnC2pEfMoZEh2kwj6WqdJNfyYeNC580oDubN/n4EWyBz+rpzKt
l+X73SX664j6RrefHLeCRp2uHH8QH+z5uQbRdvgGewMydoM5ybmf+d0rOZbMD7B2
CQCviMf7yGGJmUVSKDvzKK6XnLFraEij1zejck5el9b80MERvyd0aGPxVAfCY9Xw
nGNhR8HT9oKR94Jh1G3N+z26XGavBlNRNlWFpTalEEQ+OrXI1ow/Y6cSc0Db8Q7k
17ZeUGlqFe+OXJPXo/GjVE1z0zjpTXiZkWB/lygzn7SkgMUQbesb9X0E5r2Dl6j6
gURxqp1t4WPUoHb/0Dl4EzyXbHj15ZSfTTodafTZgDSc5/O33TuLWxPlm07zvtnR
uNWksb8kGr6l7wvGMV7DTARZBpy6J8JRnk6U61EZBx1Uju6ZnDCmLCNOdZ10zA/0
YhFobhpYxFH9aQJXli1mgMR6xjXJgSE/I35sfDslboglIhk5mUsx1bc7owYEIsd4
pqvHYTPfRig6YXlWliKcm9F3I9L2YEWCsBdAK3OVZtrxFOMGs3cbPexMQcCaKXOY
D1jyoSBHm7+mEg/XROmzBucEiYzadYlukeJJ/z6gCjyDMRk3ofsj7ApayGr1GKU8
oj0eLirAeIWdnMv2XNr+eKNJvZhH5sqr/5I4sZFlFMWdc/umtQvk4FBdenGjCkCP
nhdL1/ODwZ0GnThZmY8Ehz07ARV++S94wwff1p1ouPakU0LgMobT4CmdO5oZRfEg
Jzj6y5oXwL6U1cQhVh8EdkSw8Kqf60YnD7bh3NNQ7H/xuQ7E8IcV8glP8BVgubP3
4t4Z71h9dypgQaWL3fgl+GAoMyxw+KN4LMR1iLQyJElKZHQ4g9ETxoSegFViCPjP
vLpMAhlFXWzmta6tOlcCQ37UVdK9WAmqFuIHhnJPkJGV9PbClA9czOyo1Na46DD5
oO27ur+5f3V3NPJ8nGif+ChVvAf1CWYmXuP4tE3nhLcZaWY03N2O3wkHekd2nHPK
3LCZ6PD+9oBD+bSE8V6PggHtTDaReol3VAobvwdHlcMEVtrgXwA9G0Se8DouRwC3
HKhMeFkH0seQ2nbUcO8htXNi/GCCJ0yc5UB4Pt6Ij03LgjaeV/X7PeKMY843F39Y
7q0jNQG7dUZEPk7P6+Udg/qebB835iFfiuhg1zQagxO6tCwio9tUG/d+bxl817Mf
ua95vu/sk+zpLCGon5S90E4rJQ4QxqC85owcxNBhSaWVqgaif8sxem9nFpI16DBS
Dv+bIkGb8zdlVIBiXN0TStAWW+OsX9iHKBJtKCnBpZQApikdTegomdc7OpLr5m16
3Wt+TJKL3Gww+fuQVnZUyzmN4x7gAMDEYS23juGo82OBc8mN4SiC4imLu3zAkeKd
hL2na7yeGXLlrX/KPxyyxrLX+Efv7wr2YAhFKpvX6AwJJ5uPhpR1drpZhtuQTqTO
0URlhHErN2FzZTJSRn+7pmCY6q3m+RV/Yh0GNdQBZCSMFwCccp8gDTHK0NHN9mvU
AoYZIWxqw4Jww4ui0wimLfrgOWt0Gez5HD5g0i6fkni99mVby605vlrEx7pAFTrE
f+ojIgwyh9tBgy+4NaqzXtOFY1xKp4Gk7Adc+fgl8G+LGM/qGbubumj1SY36MOi9
TqIZoFHskPUdz2JUN+fkr6lj21rI0Xv1nOEscUvRNh1SQi/XRELvEJggb8K6Vf9z
KYTG/8pNbqjqlQQXSz0fTBxpl2wmoZneWuBlf/mJvR6MOzH7GGk4XrVOQWV53AXw
jJrM3ThTJKb7YpjaL9hHfhhjvUf2J881m1+8JJvjZCdawT9GEzgzW7MtDLR0y4g2
AwsDZbgWTewVo2ZtmbekJckpnAXxZCrx25emOtWnxisgc4D/xQp/+VZKFeOF8jOR
mYIKMBlnklofcNy0qjfNaupKjuhxEeEnm9lb9Mn0Zw8kbOu6BOD3qHtuQ79yppze
pnJf1zBarw+oOEKHD5zk/hV7QRk4rlsRk/lIKPJ77LvUtJlBX78hfz3x4ejQT4BN
IvcoQFIvyKSwyS2CwXfUBJvIO7KncxV6RnhnEaGARL5+MMM5BMPMUJz+PnAxbhcs
z3bxeh+dKY2gNP5tcIcOYqFn55pGxCDHo0WcnDT5Ni5MCiMaq1etkuokuGJ0oZO2
Lyc3DcKoOieOjuEoafRcjT73S4sGPxxDm2NpY4cerp4dPQGMKDGWOJI/DT7oUh8l
cmJ/WrAHYGsiMtCoTdUFV5fsgl6cy3yNSCZBv8TiIJ2KBO1/mDoBcPTRDoAmhTAJ
qoJ/+XogmS7BrL3m54usSyxMlZyWcCGlNX85zaJ/OY3EKWLU+FigSaZrw68wqJZ2
SSFMDBy4uJEg4Ab+T18ckpt7GfX8obkLgrrUvCv0bWTm0RUwT4JLdBHC6yQOcbDn
EmqMiXK2bejygUmQuYcdbiGGBK0WAOu7WrqYwewCT8uTWSUJe7d2EvE3cxZUASeq
RVhaKzFHPBnG+wuoeNR0ISABVnBPLqKZafuDIHHtKxwLjQeQu/vo5skjXhddmFJb
CMkvanXSHFmhq9iumI/+KMGIK9z7JbR3XLKnojnkBa4El9M1RxqLTE6eIBFpliQq
wIAyVAxtXz+9IkaHoK2Ah26O7jRUHu6AA3oGohY5teWnXba2IThQIFNWrJ1Ql45Q
sX66m7WboOuYpBvPZYHcbMS9e9GlUhANqsk94S+VrmXPxtLZ+yn/m4rYvI5K5WUC
c7snzEqLZ0OAW1A2gjCMhMUHasxuH9gzT0VXWq7G+WzYIkeELeiXurBAou5qwZBB
WQkruq+dyTdmmXYKYBYcVziP0YQ19QqDYr+4+Y6iUSTtJ7M0hYLvVyaFh7iFqMVj
tFQamBgkgDCQkv1zPZI6FKwuEV2IoRX8b7wheyrX3RPQGvDFauMpQgPcb28CAsZ6
T74b+990Al+Y1874mO159U0g7dKipDrhgarmlixCvElFuIqC6rBUpRCfdjysGE3l
z/OzZfODgcqlrHVlWOso1oxK/x4PisPOeeNKP2v1IH2zqNkUE6nsllqNco+wGTKh
bmAOmPUVdQIHZiS76WhCJd7iGS4rlP2awvsWI59nxf+tF1zP1ao3APTjpTNa5Ucl
Tr46BV8PGaGsOWIiDtRO/BOXTilFsqH8faUEz969HfGBT4gX4Omwj2jT1J/z3WIv
WCbCxTpvEryPl1f6vU34EkCb1SzBF00tesTrGp4tjLrczAff7GiP4sjchwFaCeqv
VPvqfANWmfsqBQTjq/skVp+1ss/6jWDwxjKWvhccN0iwvNR7+cg4B19n9XUYrHjy
cg2xyZXXGDoj994ksOwzUzikciODEnNSe2TvosEC5EFNP/+jaKLZDVPWg4zq0+nB
jRIVzZQywkWvzdW/jikDgEntDlVK2EPIHic1AXyWZ9muH6drQvmAnGgCh4EtAELc
lK6TpDqIwzr7xfKTCb+AaeREnlPG/kOawyrSARJ82GDbnu9ZgptUK5jKifvmBxlU
fy8lvomBd/PcURl0yUHCQPALJht19HdI0AdvCd1b64R7aw8zopnvqB+2qcCd3hP/
9b+hnGeXZ7VjeG5MV1d4zjAPbQyfR1FR+JDG7ndL3CQEBoC94H9PhDAMn/oHqCql
Hst7dsSPVyOU2QG3T9nyFtTgPi7j8gOam7s5yTiOu1Upily3qeSVBf4t+qt91twz
ib05nYNsdgwHM/5pjIAy6zta/o6Eu+4XmOkzcwP2HXTJzbYuEHS43UyMgevPN52E
EoNzmy7Hf2T+0H1LdCcU+5bSR7uX9URDr6f2OerLELKrZDw8PXLNmRkcc46IgZuw
Qq5l8E+x+Z/6qYJFgZ6k4MlfVvVtHL2duN4U9GlTwB93NhIpDm9c3FNLNGsRuHQX
+LB6d5JC7ZvVHiv+BIX1vf/YUqDYsUAuNYGkq9mDph0Uv9ZODtocD9lEF9z10fDw
kYgOurnNm/dbu+iS0l7NE49OuYO9zUFtSPuLsdplI9kzw1TALHRz+r3GqVBNRuCX
+J+whOT1veTAUl1amiuJqdzbrtnUS7YF4m9rEMq+7HtA1bhlKcuC2gJWZoJOR93e
M7ELtiYO5fUqgdt2YQ3yR6jqAR4PQ7qpu2VluCQM+W4qmz5O6J3C5WXKaWtHTFuK
RZqHY6jpSZ1MSubPo+w2JmCIfzeINnnWuYq0OqYbQcPOtgrQw9xGJIRn77tBQjzW
blt5BVO8jCxQTLCm1lVu4CIdoFa9Pripf/ajio9XM0xGOoO/6pYEpBQ3zlg1ZfUQ
AqNGQTTtVShYXfxvN5ih3w0ej9baFTtmVjrgW6kzSpXP3C7OwKbX1Ez3Nkj30d3i
0rKbQ9b8rJrZJkek1LUBraR3FNksEwVYOUanG7Pc4UzNItQnZfZwYbLi8I1tqVob
7KS8CVbsO+Bxzce7cHjCj0CVPOus2gmi3SXCB0XsBcASog34yBtELWxebYo/X3XQ
ee1VaYwS8oPBvieO59r6BU6rdtaNSguaU2nQDqIqo3UmlJl32ncuF54AYe22ZfHh
Rmq9xEQFPRO8SKTchK++vMwOk5A36Xxv+R5R07ff2VcvgmXENkm8ptX7HJVYnkR7
3Brra14YOfOo1aZcoKe0/ncQQJYYeWFAcRNREfG1BZtHVrk151ONoZeNRqq6hCtn
l6dRuxA2V1yp69l56kux6fFq8uNZGiLDo3bNhmqwKXuhWOPzz3h/WSMFzTEibzJk
r4nlHD2wvI79terO9QctB8b5mGqQkPyUj4RQT4S5Oa1lWEzS2QGQU0yArJvc/Dg1
7OJFRCPe9KaC7UPULqW5LCa1zwBfE2UCre4LK2B6VWVp7P94d6ZIRjpgbTf//TEG
x8QqqJi0iIL7OKSynKxjqjYHsRSIZmqJnfgcQIWgBaZjEiTNW99BGCWGQKE5K6RV
4j3F48oZD7Yotx+yMCgj2LIxwUPjLAZQMLpUBxBgfCHNTAB0hL8tIcdgQJmDWrgv
6sVudsCW9WrFYdiuDM6d2F6QIOP52meiAf0LkgFgM8+A1t4wvfEVg98b0VZLxLxs
iX5bjFH2ubxofnDzjrehiR24V3g3Jf2880bpY0bjmLaR2GN3SUTOOHbw/EECEKdh
5nq2y9mALldRf+mf4ZOvxDUTi2lG/8SeJ49B1JwmApUPcvWVkxg9NpmhGtErzbvP
KvWqzybV84im17hqmcbVCvy6s0Cn6PlmqXySvY1B1nNRttju8y+gZmzH4Zt47LOT
8WEzY3NdvmKCiLdljaHeex46p9JJK/ElvhW4rDlCw+bAEJSD6ckS+3v7wUdH5Kzp
hdirIJbIyL7T8ynO0dSQONZ3NRDfkSqgJ5Aqjg0MzynCZgFsdF2gWpgCGmKI6cL1
GvMZmAJ5b4noggW6luw3uWaufud/JvxS3JYQi6t2Jsq4Ji+IBuN5dnaRkkNTxMqV
mdPz2ANrOGUaBTmrs77l7s7kJllZW09MYQcKiiEpA06DEVcipjKV8MuUITjkWuD/
LHlBDfeomHezpkjRJJkkbfVwkHEqHWb9DikEYdSEO8cXgV7MKdkIfrXxvSl/1uUg
RAb1RD8jUHmxFp+wRKkEypdURfDLOHsluH3+UlwX+Z3fUSvVlFmAL0grB5MKwgW9
jG85NSnKNKH5OFfOedaomteMMUNnAfQuy2TJioxQN0/jBL2clrLfeeGbsxX5NVte
+/DzGNF3cDkPFcR83LOexQtSRreK7XHbfOjPHEoIakeb69uvOTb2TnQFhMiZRgNA
cQN49ocXtEVkevV06bSrBQpCPcamC16iUbiYNuiZ6Nh1jdLPi3w3pZqF5xHfZqtQ
Vyhwhr/6wiORf8xubOFvpIsjBniVnQbpPeVd54GAxIhhgfWqObU0imwxfYIXfwVK
qmhADT5/38Tt7eiEYkj74lV5FByIvoaC0nUpQRFjPnjZ3bRk5+2f7Ih4MKbUS5vc
hX3+n2Lb3AbSEHCWih5nwrWad5y18DrX1UrUv5sB+cbwkGKNkJSplJIYxbiKe7XS
cGTYxNKaDLBIid5yGhDlDkSPnvTJct67oUMPoNCTfiQ8bLu7RZlRzl3aRX0ZwhCR
MdvWSHs9jiAivgPnmuYM591RLm2uZ6z4tiqqNof38nKvPHmtAIxT2x3XyRlFqRPy
9AgzQLvQnkbUG18ypryPQCj3BwgZHr/wOhdjEki0YmiBtaleER/kPFxf6zeSovaY
R2AaKvjq+mJ8GAmWNHC3UJaJmAR9JR9rSnx6ZDGJ2IYEjRyy3mSEF4ryIzLy3x37
P8A2YrcxD0VPEvx8e5jUZzfcc1L8k11uF64kQvLg80tjRdCvWAyBNx8EoeBdaOxb
UA8ay05e0CR4PX6iQgJ7gF1b/9y0l+DI6AD+8C5KS37vLu+kz0QYK7V9NYTcGQXe
WUI/DltcKV8SmonzQvZmg6HXE6ZHs7YY9U3uA4nEPG0mPtIiqjHpk/75NV9gKLL9
PQntu6Zh9CmfLK0YFnhI3ClCq/oFe0WLdxIPTjD4q7j4c3NujJt0owfJ/4jFsZTc
8m43AdusyuL7OCUA9z8pf3H2DRnExT45GAm2stMYxR08m++VYJwOcKVNsGAtKmNS
y8zaeev5QEYpAdgFcgpYrsIXjpTbssRw4iEldCwSSMlJRUPf/OJRPdQg91EPJs4r
00T6PJF1OGeln7ILzkKt4KapADG5S5Zyr4tpVZgm+9cuNbozMoQeH7mSYv1usvkb
j5IGpdgHyeb8W83FL5yv866/laTYb8BJzw7inGsX7jWx2kpwXCDUhSWSJbIVbRIK
6HoOUoEYqHhAG11wPvk9f5UplvPo0afkfldy5mZvVt14mOP2vApLXuOkkHMEm0Ke
GxCxB7S1QvmMa1Mi2Gev3aIy4ykN9v44ssj5hcSOdJi2vpGT6Y9cG2Cqrj/7uAMU
IlB/m3V5p/szFDopTeJ3GwWOZZhw+TPbxMilHHOcxG6q8d5BNZJ6Sb4HyzxCofow
wUPzLWeeds/MdGdjVwpgnCKYcXW7cQEUl2e/Za1wg6Op8rteBiiz/KB63EoH02al
gWASkeoEdLuVmyH44D0il223cUs+ubrGhrwT0S1VY8RfrWcozu52X5k0YhuPo5C4
q2gUdZiph+Z4rVnn3Pd4rNXc8sV8S8qe3/sUNcVu8QWzy19WnC4w1jWO7bezZHc5
swQONjAADxnvLVDLetav0XHOcsETeA7gi3jHFsVYiby8f4eWXeqqEQNCloen9gBC
XF+tNVZ1PDEt6MzPLMQxurHOuT3Qxdj0ZpCbc6Y/m9VSyR1/uVFHKx1lqP7CnGzH
1YiKRYekOobnWMy4Y1z1xweElLZImCFHuBjtBGB6VfwPt5lZcAB4ApRKhSKNw52f
BfVW6t8HHbnvMyM6QMIY6g7pAsWNmohEHSTH1QDsoYjqppTokVty8N35jBy8bgGj
uqnMPbFPy6knAzZhladwHTlP91Nsvhc7vbcUq6Ry67U1Kl/M7lT/zL1osIoudBNO
ZoAECS8k84kjv4zElfjA8MD9/rN8j5bec8cKTklxWNcno6a3s/DaOhPnKnJ7QpD6
gqjMym9A+pBjQh/PcRmROk/8f4JTkmhwEfVsl/4ZlYpGPWBtWVLimWzBa9ozmDwb
GI083X+osRMKXuqQ42XOv0driO4r2Whm1Y1TG9TStSepG6owEPQOdqxzDeNMP3rD
wkcYh4YLkgcnyyvD72kVAdqdlOCq0E851tlzUKcLsYW9JhdwZ+i5dNyr1GGeY9kn
FTHdOQC5q/LFBPwYQW929gA0GfRIuUpEQ6PFyJ9y5tyFvtfDL90joAuNClHncur1
NYbRA31TbGFN0+zWIZ00egxUSeJ/JjjiuMHKSvnLjIvk6YZNIzzinBrDqB1tOhxf
llXiFHQ3FNi/HdzTl+1brqaZ+36rz9CxeJVpaZeKxn2BVvXLnjHnNq+qXq2sU9yq
KSll6+Exlxp9h/On/iSAfRALbvwhA6k7meKj1xE6DLuJxEG3PzmKifyw1WFBihk6
2C++H/5ueb0rP9mBpt5M/0CZbD2jMR7acewiLHw9L9QiLlV11ZovOoR1eNzVqMJg
iDxza4HfsXsOb7BQzoCYKY0bYLXenFc2ZZ4WwXrkDSr6nnyaYiQmceq07gDbJBho
goRKoWv8YDzU5WsOmeBR+Rhgh2vHgPXwzuhmEjZPFbmxsoshfAwb1IN3DiZV1kM7
JyDDmnRer2Lou+d97G3F/IUGtAnbbjF3ijpg7qKOcMW0gagYRmE2t9umuMkKE80F
B+tl97ur2YRepN5lE/53E0670WlYZ4kJxSTFx5pmnUNh319ouFM9rRmviF6Axuz5
X//taLVm3xU1aD1pb9oa/cno2bUzl6Sij/K4i8pXI2C8g99UFLpPC46QPl5Tu5Kw
FMKY/sT7mJdo3CKVgFDZ+EbABDKuQVnrb/8lZPsSV6SbcF5qj+Jj6Rpq66gYVd92
ZuiG9OV1/xBt/2g3G37GQg3cySaRA+tZii6xvKhG8FNp6nPDin3DFo39y2E+B2lT
2UA1MTseRxcLbIsucIglHZqyLbZwztVWwyyg3ErijANlNeP7DHyH3LJbMu++2Urq
5Fsc5bXzk69EzhZyga0+77p6QzaNsJwyr3AjReebLdmvDeG6e+t7oUkMPJzOlDf/
NZMiMJVUVCsG9fxsb5+6ftyimMQIvmuZ+hcPGu9dlFPIg9hjB8NyAxDPEZd0dOSI
fZwlQkmDVLuOD8hvxTZawneG61i78znFFyZJC22VgXGktuWwzHihLWa2HuCyfhO7
wQMZuPN8wQVHkFQCPYXg7oE3nCzROI0XRPMkEw5jlLYhKIY/jH91FLhAoBMW5K3E
nnJv3XPVoWTuloggI1X4XXWtKgQa5uiluvHz9y0fz6fX67PGzMlPjIQhRyL3+FvO
Ql9/vs/Kg/f2h/9x04yiwhpX8aZ30UvDvRrlOaTVI5ja21no/WYC3m8r/6X/gfZF
XRCzLmzqw1SwC+kynu6ViIwXWw5BJYAl+W1RLvnYAMRSDENsdn8VDwJIXiNCGWfc
R4jGg+8ChCJc92zhZlL6YvfX3xRkkz6os7ysl9We7RWth0Sz0XVA+OA93Csb7AO6
wSLgDPc/W+rUE8/GFo6gaTeNtdezwx+WDmXfWrF9ehlE1Wsx7vnbsewNMDG2ur8M
HqyigoaFuyPlgqsQJJSh+YPyvGM1YPnuJNFJSuJEHpD88ETsLWHGY0nsUxZPpR9/
1HJK1hofS/AnvhWwiDLCou9lpLv7fn1T3jaK98A+eW+qoIr+8l0zFN3xCK0j8H+0
LTfhWzz2J0pmS5MTYPFSC/16iQzoHDVdXLkzTjbq1uZ8SkivVEQOWxIlOTL1tC4y
RgCE+mjsJTU7gmEve/Hc4ru++luvW3Ko9zz40glVN2ltEet28Sl9AJpa3ZhKt2mh
q1oEw0uOzfBdlwFfbEnsW8ZlfBXDqfOWEISAxlv/FLBSB55ijf+/4/YIMvD9T77t
k+Kxz/nwFXuaDrxdyhpFkP5GsHbFmXqXAj8XHwyznm7yfPj13A1ylSd+upLdUVho
54GDpSf2g9Gij/Y2C2cJLwh9bGoebDewYhSspjPJD9RP9qtjoUNbEkITjrEufmCi
F9He/uvN+Sr/nbSrbYa09xgQJCZzqEEAsA5+iJALnjwc3B2fEHDw8OS+4j59HFUn
YU6GZImeAxKotaBCEDh753YpJaSY5FlSy3vSE6d+qn/4tTYkYV8jiwbPZVLl36eN
QAlDFS4oBRxPTcK2jBJVAj8lcdvFnpAx9aXT8JdLQvvzX2r3fAoBLaZmjqLXIPDi
EfgPX+xgwOnyMKggQmDnOYKtAwXDsUQsnWK26S/cjPPlqXMSknRrqeduJI/3/Vkv
xeLvZUUov1/Y+BGsMACvTJDCkmaOfVuIm4EtZuBgWoAgt6VWFH18xelJqsa1Go23
MVdKaip2XFq6SoerkQFjt0Ar+5SjaTIwuJXhXbF+X/dJmKzh45edCgZORK/vKdwM
73FyxYZ4SVkBSm7lE/tKuf1v2xcWs/LRv4G/DBNv5IVFjvguFG6pnb5KJ4Gb88Xg
1n1atuVw/uvUV5nro55sg+72cUl0ENpqMkpTuzHuOvrP0x6IJBED+vl8Fst5HNMd
pDZL4+GK1brI/9d3WvhtkR0HVXOWkseM6NdfCcDMBRKHCPxPG1OQaNqL9Q1VZvps
Y2/bbrRCJuR9D4t9YBnPh1KduexCDWT3iMwNtF9JRYtr6/VRUFm8z5N6a/rZcmtN
97c73jVhxUyhtcM1CsotOAdyz7m2/JCbRK/bk8hqOXIpTZ8T5Ai5hYeHpaow8m9r
AbHxLfLwZ2nbHekZyHwrjQZ4xbdS7MbsN+OuUmSedNUV+ulaEKj+OcVF/KgAtVvk
sN5xC9hUZMX02Gj4AVR9aV4optn5SSGY1sWvw1nEM4KIFwe/CNGYiICtSNhXzsAy
RZJqvtUcKkJKKm80xgbpvFqMxOZmeoSVh9p2YTbbZAW5M1gwyaXtTGWk0TNQkmdx
lLFeXsvowL9n01bGcECsOG6o25x2ViqdvP3iiohFXtYraUr+EfpnGR9IcUbvusNn
Hh9uWY7RqcWVIUmiYSO+XX7RbzHXT3d59FOJIsIkBXCh/rAx13F3gGczyWHKmZ7V
5JtcXxb5t8oYCpQL6cOGf9EtXV/5YT5bw+m1RSALd4KtZFc6W2vlKmBW1E6mbvjq
Rv/Oaho38MFWGOZpByY0gv+kQK7hjCkm/OaD8zgKkpGc10q1SBml421yJhJmuGrH
LQnO6YbsWWxgIYSUTIoyKvetA3Et9uuWiWBOG7CBPb47Ttg7FrY+kJ4TVbtEwp8V
+jIlMiDxp5h9ehL9NZ+qkiyBoVqOqJQZadKQHAY2iBkSB7gaJJ2iOLTAmald4Jtj
XhMXTmeo7ur50klQZuM/mQk6Gf3DXXKQmhe7n8OjFE8v5Uz/vs1MBTZmC0SADfOu
u0vo82J/WIzM2cjGKduS6rERfX6oSbTGj0qgzDAsvGylaKCYsDIP8oKD2xceSHP1
ZGhLf4Z0RSSTJd6Msl6rvWb8lxIzZba+SRd739bG7gcQ/OaBnFOSkQ+/BHhB7QEm
+dWR0JhOMDdXRrVh1ZdxaJRz+ksDL4OZppLa04yYdjO5Xh8MwcOEboineruwBTqI
4GkTM208cao3hDh1706NX9Oh6IXSTcIJD88s05PybSue8/nCK0OCz1cvDuI6mX9d
umaPzgtrTLzOHVtyhg/UeJ4rozbGB4XkpPSx1Hd9rIKAV09rrPSRG9P4JA88Pz/l
dTiux05COS4FYh136LtWNAG1OXyBT5v8VVuDEzfSY66kAvfqYDMdA5m7fHKEn8kr
ExGSc08PsyaW22UWHgF0DCfQJ9F1hyVQM2odsZcTBkmE2d/6qHoEkAOQ4IsX1btn
gde60GqzoKOYO/xRT6wXthzVm+t18yX/qaPl0qZw2KVTMbjj/uiEBFLdBlyXrQG+
dBt4GGenoShW9BAOGcxk5vKD7so713fWM+igMPZKmaWGbawBGq69DYDvEEXykEKU
AODzCFWFn4p/IHZyD9dVOg3J1+dxyozzLE/Rka9eWmTF02aTKCJA+v/L2Z4c5b+h
OzlS/l4Fu3ioTqdeyES3KppKCdRuIGTL7YKJNSWvkQtLmL5ZfwqTTsHpWiSQpvZf
Qvvm9e81Op7fsgG31+3CbbaPW6mWPA7Z1obW4Cx2inguo1OHMz9UZgh3iq7T8grx
s0zp5DH4GY5AuY6w/aCMt69NCcDhnmnZ+XcaQCBg3Pnge4MbG09ULKyhZAxl+vNY
ccGqNcGTGVWuTUlwJ1Yui8NfklKN+FjavUvwNk7XR1jZ/2xUDuzK5raLsa4OQdPu
z1Ne0VzPxvA2UKbRth69wXb35zVF6GfOsX2ZoMV8AslwonITCvf+6CY8hd0S7rJ1
IXnVTPj7Zilpe5wMPtJH9WYz/N6r7GWjFZz2g9uQWT9nMu4Qs/GcFEkZbwoCxybe
sRF9/SLZUtsm//X2S4uEmfex9Wyqmp64QeGLuEoedO/Zp8DCcwiF23Cn8WWEDwkT
6iCu1oAZczZpSbhoD/z48Kg0QUS4fTCaUjcJBpEUAbwLG5WcR/COLwPZoLSbnYHa
QSqQyguGUEK3W07w9+Bf1Vivgi/hNUvFDzoK0Bn0kKIn3BDgEsyuS9rJLxar+g2r
odXo6y1nou9Zy9PFyOK8BPXR8XZxinACFwjmrnTeee+TbSPhukYnzJF2uDe1Sf6Y
VpGopHssQtxVzQkNKto6aI0YToqvHhbA+eRr/tLUFnI5+u7KApQNqmuH220UZTWp
BoKkUyyy+fDmiaQnhV3+Off+tPVVDmeTGGCUFUluzBDSF8eI7ZMrwKqL4FZMA3K4
o9fyzooRkpWjjUjZpe/yw47uCxDaWUoxoP3bDQbW9R1OPg5Eo6l7UhTxDsSi6RCZ
gLqzZg4S1stFzVzrRLm8A5tEDlJH0FrawG7NxtQu5V0MhVnN2Shp5KeGr2EL15VV
qKKGjVlbGBrEba0IVHwDD1qFm/jlePNDOqDlWgUu26jddjD78sItXpZjLj9rVwrC
lKGUXnUwk9XvZUZy/AAQYPC42xMnwwMyLgpyQQiC1VCMZ0bEDKvSHfRkHlfX2c+5
IGpqjMWzOAkkCRtixysLI2IEx0AHLPaOA8jGw7YIgE3LpEP08oUMA3El6y+AIvoM
b1e5/DZ+r7kKdE9yNy1s5+mNV1yL0j1iOsqmfWmQgMQ26pn7R37C7anKiy8fb/+X
6cXBMzzFvJEueLncPebReHBwQsTD7ANgHaOZ8vJOY9z1ecsKhTX1vMrE2X6viFeC
5pDzFtco4ZCruMnWMgd8+GmHAarXW/ywjncR7B1dFTt/TiwBCfXzC/Tf7+sNIxPi
+c+7EPCpMnDGCypJmJZcM4+Iiwp2qmbR8vvbkCZsZUm0c5NOXAKljNlwPowL8Eb0
PWzwc+g336RxdLNQ25aL1Cw6w0jkMS0+JIOBsd2p4LsZRfLvR6QatuWSVzNSYoT8
oKEy7WFOHTIhTCgMn6o52O+vMANP1y9wNXn3m9jE1aji3E7oTTDKpRWzcKhe0Xyo
NB/rK5d2gEmsMVsY7CcFNYU6JmVMdqyg0/Va6Q9X6Bmcc4eWAvmqiaTbC6zTh2o7
tenDMJONZiRYFhobl/D1o8qXkQTqeNAjrS0I3iI/2mm7BuPANjF9AJB3F/VOJNZx
I35l2U2mtJSmxGLaXtMomgmWimvNB/TjeEyaiy0hGCC7jyJ4W4xR5HdkB+YiSnPh
eMP90IBD2nbmLNtIzr7RdC9+Nt1iqY65VKxi/Rl2RWjspcd6CkMdHndvhTQ44I+q
yKmGoyel/XALNBED2gjUaOcUUXRAHx0gNDxkp1kjJ1XKnMxggapbB35v/fcPfHSV
/ttM4HDUxm0ToPEOoaURiBFbezNa52f1Kn2BmQkBH7kVoVRX/6eceio+8q8h13Il
zOiwCGEPaZITomKgPEKIVS/P6yEUnZ0AlIUO+Hp3K2bWizPa2drer3Hnw4B8WQLI
EUAQ3ZwccH9Sx8MOtAEy2MlHTrUEBYpOXl6FSiD9GoZksSkzuAewPPG2tog06A40
+CMWzZ1/sFd4fVZif44tDTsAerJ21fTucxPl3BiraMHLvDiiBiHGqkb1A/bIqjzh
WLGP6EDIbfCGUXRuQtfodWvYl69QzzBqQI9d/3XJavYgzTtSRF4nYzLj+LxYivZJ
dI0UpGyXfkOjVvRlisRVvlpSLGv89SyfG2RR/OfMj9BHtRH4ZN1ZxMYMvAvXa+K8
mijua9yUjgI9F0ckad3gNn+2yvolMh7KvsiCGp8uRyjQXOyTbjfX0DXtcH8YMtFy
H2RgXG8fm93mLZUKI+yNzN+iPuzBYkMtnlAjYHR5MUh3IESuSylsJpQaTciRLk7l
IZ2UM4m1yqAmIZGEz0evzIkcm2PgWo0RVL2mbQwMHDTDMyBXifm+gYW2jRY9MLcG
5pI9c+RwDShh/eO4axVSMTgBSQl3q4wfOikIyA0sXzZy6a/uWiSuDd/xf83yxq6B
f2S8fn4FqOB0DBT9LdkqKSd6keoQXhh/v5Xs+XnurrOHIcP4mWvb/RDzUbqSSLc6
B5SQU7bv8rx9V5FBcMFzvquFYuwFB1NoVjB3Y0W1tkaAXoPHKTCfRVTylMTfB3Pr
PV8fEg4RMGeCLJt9YnfkgZ12HgdP7QBC704ztYO225QOnJAZVVVEEf2ox1uXL8y/
UD1/euddBKIVKlgVucvCCUPxeFFiMcmWfi0ePI34Nh0TpvmebWqioCPzsWQNpxwL
TZk+PBWVbSmbfqozxJWk0twv+t9SH8SYpD4J4lxaYrFkAtgZ5UiC69IfUWZObDux
TRsbY6waf8L9X90j1mTpO+rVwtbKxzC4Hyu6ZY6v/gBdqKCUQndEok+hPueIo/au
mC/9JjVsm3yGL6fBQjgE4RdfL5BAM8HXRKN2ab2vMx77XgVRC72hiZsFg0ydbb+Q
+J00QxEZTRAKJ/xTWEittcJT+LuWom8EXg1+5PwEzcrEuDdPKxKOYv5viqayiidD
egtsHqELKWnUFnD4OFpSVrmdOsocPyrSMejKCzE3QKXXHmp9TjB0PjfNaLbnwCOm
MolGo4lS2ywLHd7JyFvDG83kD7hc4ylXZjl12K6MdrFoN/QcYBSDlJTEqhhEKHN4
9WMxGSIYpkW73XeHlxWm64Ec5AIkyOiwlu47PLJYCXt0W12VCCPgqc2w7bJt4xsV
UsDAzHEuXr75sfJbm/GanBtO+sJUX556Ys83WU7/YzTvNvqbfBf7u+aUQ1EHrrl/
/89z9vTTmgPKFpn3yU5XHuPUClmcpFQkqz/2Zh/I+vtUY0aMWCynsJiHfzN7/vN9
cvv7/QwP+sykZkQcCyX74ZsUi3X9HJuxnUP9d0PuOyLm6cfYQV9rD8sUBavFXy4y
rUpPtXYwVbz3VOwEQFDukJPVpfAnrRzYbXKay8D9K4B0ttILJJfeBBni7aVSGU8S
nV0QdCx6rg9eJE7BTDT9gGdeOG2M6D7IARbYIapMvLJ7XzmFFw90Zsi9HaIoU9OT
i4YcTjIFBwgDTT7J96G9wigjvC2X/6O/XsOx50qJE2rcEVh/MGRM6pvOI6yfhMSW
tEBXre9oDrJ719ZvW/2h4vkwZjN6HRmPXhvhv+tU/PFUDHnjdzp/49nBtYq0q/tc
26XCG5aVaVsaYU0sRBMMzvXcTfOXYrk/Ka+Ah2vONuTIg9rNqnrO9DKmhlorNAJv
e++qT88b15v2930PrnKK8e0LiHFpQHLXvnFsBSu+xRXL4OcyWWyKnrS7g0/9Ja45
1RRXgt7qZF3hOc219vPNjuN2DVWtGOD+bvHPSmGUpI1SEbFivgIhEm5dQBtlOzs1
zOmhH0JOvjoTUZgSvHw5PKLbYXHnPaoHFsBQUSDzAZ8eTaKCxwuFR++t5kBJph+d
7X0NUif5ONTPsPIKeaGku+aq+6zLLfgS5KMw4XNUc7CVH70hw/WCVhv6+sM/TCBN
/3OIBkT9XGJUz5T+FOFsH6/IOrm0UBoCwJIGgUhM5JSdU4/9gls0YPKH+KwGKrBE
MDH1y8zxATXGyGufT+UD7VdkOhjQ1hMaiBgAPdVwBlWI39Ns/qlAMWVFkwKjpACO
InPqnRKOXMA8UAbHDA3YbrlL5EKM5g0Xz+ZaQDDZuOJVTnZJULHFomTsX2jhocOe
4uBC0y+5TwX6p86EG+EAkXTPsASYLmgbx09nzj6wdlsNO2aIW8uhgak/XwhNyttx
xsESyn5zEMo+/ow6tC4Q5XOFAt1FcBGWiQXtYo8jI3lhmJ6S6Rvxdbj5xTJCIW4e
P1YjoKFwsThBXBbwqs8aC6QfqniAZUNObaxVPK6i5Hn5EUWFEPiTwByDJLwQOViZ
TDfPiBpuMn8wjLuGIW4rz23eaoorSorDv582hi15PNOKFOi8G/IDfsKydSEiO6Jz
9Etww3paCDg/IoDH0QK1cHVNSv6A6lV5Kbkzy4yV5EhV2OcayyESOQRbsKTgcXpM
aeRK+iRzSnNx+JND6S1iPxjMrYK3FGh8K0k72GSfp0/G17yyeuuZW8UTYRtFbUOG
fzZTnjL3aP1EwvWl2BMZdxgrkuLlePI+EtxglqzV2jVd1V+q6idEiDvpouWubXda
G6mdgXZW+/MYD+H8ubT78XlpgQCA3Abj6MA2/OZzAHFF4xMEE7vrxJLJKYMAmewk
tufwAdq2aItK4sFjvsv40Zf1o1Sj0eTflDQL3ZZ+FaL00vS9GhIu4mu9TqXmDB2r
Bs9hhwn5Oy9UqUuAJtLI2DwdAjUdnnoiWEIWuBLZvyYt0YjkBXXxQsEsWr9zYIPc
Dnee6WIpPMzpCcUjjBw2oU1Qe9/tY4W514gqRtVcGv1DSpfc6yjK+26vqdpS1InR
t6ZqWNsuVGS9R/DIm9+NIu4KxsO4cfh6KdYLwrWIDvbz062vnGNax/JH87qgR5x3
iPgzpGYKYVOlxPAj5tl+iYL3EZ/fEqqXmN+b3nzn+NoUgVj0yJm2LxRkM+FY7Pve
m9/K+BfOOiM3kka3K1LJqfYG2H/ej5O9VphKvcIpp9WL++3cJ3TmIBwQkqm3Lnan
DvfOxzViP8+bEi8Bji+N9Gw1hc+hFy6XezutBCHiLootO/QO41IGXkodFM94994V
n7kKA7uzPqW7o75tD2qEZjdMt41izAvlfcKwzTBSXYec2GWfN68hlwl+ojzt/Fiq
zphIXWRuMxJnoP31px/S08yt7U+vh0HWEIyHp53gOnLik2HismObIcNm7kYd1qAm
OP4jD7b8rx1V/siMvL4YUOWkN21WUzNfYG9ozrHCYhE28fy2QDy1wq4Ks3Z4f5dN
KxQ0hiPyllPfYNACTKq9OnHq+fuc1xOqQ5YSFxMpzQDbfN5AvQtiGIwle2YyMX2W
hjPQ55Ak1o3FXZLWCgWocesBMtcxmlHz0dKZ70JsuS+TteVQHpwsMBELHZc9DvMN
ExVJuOsbdYwjABtbuO2cuN1JrOQtEh4acbGe28TwNEWs9fFQ7v5JGP80xD9/qZLJ
hXs2PAmjAwB06+eASdYHN+mch5bYqavCvTZfvjembyT3n56wUSr70eCQHjZx8wOS
nk/PJ/DGTXEitOxX0lBz6dkeokZC4mM2SWVAZX8zI8z+TtvSUcxfFPJN/HdHr/UN
CaeZLVibSBvUBVi21TUotIoGxDnPdzUBUyrI6IOu7XGyYVeWf3eupgPfh/nqu73p
/FHCfLP0fZwRywo8O9Mrsymd47L5z9o3KFpLDSLueVVYJJNStMJOmPZkkhiCDJ4Q
B2rE0sdVsg8Pk+utNw/DvYONaSdXkhHHKn7/OY0i8P0CsqKylKryGj1nmN/og6XX
4COMn6Hcat63sHj1biUIKQxZynTY4U9PAXS4SN6jIt1Aw7UfiZ7t35Ef/faHjNpb
chX3yufVeAws+NwT77VlnYxxuOE276wfexxqLEFgMSbpxYHf1JDvSDPyEzJT6jTf
1GDlcYRzceSO0N/9ac1tOr+9wAqnrk37tStBIYePZ97gPKZXquYUmVOoDLnFhbV2
XDcsB97G0jw+AVe0Frkrm2bry70lPuQMtS2EReBxxo4f/sEi8B1go67ERRf0Jk9+
MLa/CB+gv1lOpda+UNSennUPzZRaUPQZ6SCFiRvVhKlXS2wA7h1RTjspo/d9EEYJ
BleIJ5eeAeRVLDPnZ69hpjv9uxY3gvhKBbnTuIDnTJBM5wKJJEdqg8VSIWMrc689
mpyDGtCrIUbiMvagWOwGlXsz9cfIRacYoiC8TC4FqltVwaBjMNeEgV8WA++a8mDF
pfbd9NlEnsntPpZHG2AuW+k1+3SZcUfPstG7Y/e9zHKNybPg78MA31Yy4bh9sYKo
84/KS+bjIN/f+gv40xG7Ywl4lqRQ5xL+LwIecn+vZ7L+VttpcmY74oub4ikclEVt
eo101R/8cazCX0SwI38DzyW3Fa4Tp34oV24FShTs9yd6zt2DCmm788e6mcEARHn7
9IzGIEgqMcNdv4bO/uVKzLgTGopk6BxpJQKUKolGr4YGHo7xeQvrQuDZjB32L2DR
rs8MedOwJSNFryh3+lwBM9MjZthfS4qi5XmWbzlGWIuddxQmS5lzm9jbgoGOyBY0
4JPIUhVVhNmkZEeyvFCKVx162YSDwbnL/sn3T65yj+62eTSBnQp00usRrUl8iJVT
/x8nBNJMjSypmfUPs0By/bVZ2tbnTjbFeP4SJjLMQAgTwV7D7qImTRa7XJNWiRY+
EEvf00dfBo03RAIw8No8S5lwZxq+l8YLh43eyUvvZC2bCxf/hNVdwBhksG7fNOsd
2KH7b0rz3YuZLgMKu5d25zwGxSiWDCHW8ByHvxivY/+18Xzk+Ew/L89q5kY5zT0z
n5bLMETRkgNL+NQa4SIKifgN+1j9xOgHq3AsijN9qxZbmTtewkBp7blPTW2K/7Rr
/EfZpFsGLo9FwsBeVdC9PMd4y7TrSOpAcxNclnT0vqNvVMCJ9OZmWHiQm6vh8El6
jLPXGqBAfaRmY0Uf76y1rzGM9krnQcmk4g9T4MrFig8LkPh5aNPxbT/MhOJEJM9A
JocBo/mTz9FbgHlq2OYxNfsFoWTEazFHAc4pl7ycR2WXjukN3C4Oxu6wJbZRPhD4
RnvBcJExMphsN2B/Q2+zpFTuqaL0zp0D80FeXOnNDM7LjaH5U6UOpvvmYzAAEXOd
ZSjVWUP2Hbdi3rFw7m0siEGqVxJ98afn12kkmmYLT9h1ex7SYrH/f1QzgmMwiYH+
vk/lj2W10iwDX6wEjEYiKteGWiIgNiOWviSPO0CMvuYPko6sV6T3SOPAAxJvQTaC
B/wGRsuG7sg7B8e2vYhUSYTarcZavM70uOA9afkqxChcLn/6Gui26lIX1HSzdGVV
bMneUoekYWvX015772OC2ZK3ZjssI8FsXkiE3PA7GT4IrmWiQzYHn2D7o3rHgXuv
gESK9loW6eMIa8ODxdFlY50L8YG7QodlwbysUMUiuIQfGEhp7qAFCkN2mNmG8DJA
MM4Qgo/8mBkTxgP3nvclNoi9y6PwqIxI+noyNW2cfcdV0kBI5gldw0Mn8OsU45rn
+w6ODtdOxqyfp06OtCcLQNEBSI5kpjdXSIi2ue6rQjlC0ZO7rFNvmuiuyW/z0L8+
toNDdnDlyh7z9L4IPdQUV+yBBVlLQyFcTIfdj3KOjB+PyLfGNe3M17nLnGibF4mb
HTkGXNpSgUorWqHt8+BiVbCD229lKgR11P8BVqg9m4A+5UBBCIzVEoG1bhy8sUN/
4AsV+ZtYAseT8T6+gD6DJJepqbZSn7PDyr9sDaffxXCsbsEo7PK3h4jPzXBxH/1z
DakyWpQEL7Q5EcEzqQmkIWCUZ8ZIoEQGn7tSg4yVsucKmplAMg5cAQVYngN62Pmq
4AIQSjtoN3fFMHykdfUz4rsXTIVuf7tUKzfhdEPJDpDO0LNBWC17Sn3X4tRzgTfB
6znt5+VGpyFi0Jg1w3LNyqeL7VBYtXNx9w9fg0Uk9g/XxwNJfrySTOyt3oIMZqIZ
uyaxd2Ofd2iqmU46V6qcBW6gjSU9kK14TpjBRohVNWzTC0ejQVwUELfWnipgddfO
wPI+vpff1BEW93QYyJX4AKtHwrZOqxtymnfgL3Zf5+QMQp2HPNV9Cr8ImoRjoRUZ
kitKqN3TGiavgvBixYR1m6fMqgefKYU3hSPYici7zkXWq38TmurRlnpzmHTE8R2C
S+mJlhBoJR8BadAFlIE2IALQcXLo1MKLC7y0as0UfvyF2M8DRTh8uV6aKHqaWWQY
0qXft2DPW7vNXqlYx8oSBobee614WfrjXyBffuWD6cQu2f33DRZN6YaQiCT60J3h
RF9zyFAtAdzueUmk+R9nYIQAIDICUEahDBgb6bJFiU1/x34cysaOK0nHKnOA0mBs
P8lN7m60F99Hc5DtSm/g9xQxMm6TUd+SR7p2ah5tdDmNw50qFJUV5XsqpGN38bOM
7wd/+Cuqw0w/L2q3PypzBOGsz5J3RZBBcvoFUVPcq4awQXqDN3podR2qefA7gigf
Rc22m1IAcOqQ5YKrDTmNhsgNj4XLb/kdVWn2z6Vg8ublmeYcxivj8z4Jwgm0xyss
TRc68qegBKvFTLnjiacDLJwH9aHHZOZZUxhpeTb64Tq5p9lQhBJqRFYW4pQIEMKe
f89Gmw885gkskj0A/cr5PszwK6z1Kn4c3dkfFgU9I0OhpaV0c+h5x5SQKXLg+oM4
oM3ePZcYmOKTVugl9NzFBFMSMOhBNShNciIsOJpE2WiIVBs5YHFhHANrhj+Dp+hw
49fcsBCSMzwJksYNQVc81h0WNyNovD7LjNHF677lthNEBiS8hEsiE+0IaNU1kD70
iOOJJ9zPrxQrKAAXnUPgYu/P4yfl5kT0GyscXGAY6zmTMSwZ8LuRdTtVWYvYF7b+
b+6yJPhe9kzgvYzvDWKl03mAN9zLcbouo3W5mydZcnYWE1lP4ilDg3OApex0vqE0
b51sT+qYo5F1/O8H89SPVMSNPyeJgCQXb7rq9reIvqIA/QkwXwng3y3fVGbm1D3X
0E116znQENO7KT9DdyLUTi9XxHDL56WsnRGD7qW8f4uy4X6iIghoqz9QuqVkDLTg
qlQoEEVzeyYvL7ve+CqhclFkoG5xnHbxks+0zw7clQsDYtm4PHVEZBV83rUnHjAA
0JzIr0ZRsCYA5ll+N1AQc3g9D8ayBETdwk/+ygKLH6UBS4l9WxTX9qQI8PPjlyc5
4DnuLOSmibTF4AjXC8M2NnsKC2MxWnhER5IxI1jv8sU4xwHfKECdwrBrWlMEllcv
vWEyfnOmzG+bVVqk9yXXgHR9Ax8u2UCnRMZBDx0ivV0WXnLEXFOyg8fHFJ6xRsY9
wjQOEgSbOILtnbCKyh22ALF96jRtlqJRpq//1WklIa8fLZHZJDvlFL1k4ysMylEQ
nxGXoenIuMS3YgPPomc/WYFnm0Eqhf/H1agHEfXTLvrYKd4EGVBB1T+KSh8Ggyax
IJOGXTcQ0Dx9A5bbcrZkuJVL/0PW+maozCrWC5KDd8/CffnTQ2cRjPCO7F/pP/TP
KAk5HwDYPurrIQpuX7z2bD2ACTdaSO9avfoT0T0r6LJ4orZSZK7zhC2RagaKgZQT
7MbpCFItpm7Zi9iL7iGX+1rr4Pmhcp797yQpiOIJx4NmwZPq+3jmOMtVFGUAsWJS
A81svZ0CJDKt210mrVecKxkv2++gDhRVbO/u/4z3eWec064r+/rPg3JHsN21Sd4R
bFONF7cX1a21+wFgkhKEGx9I5FBI7jkzILoeK2xuEhKvrunpXN29q/Z9bUC2zwbS
ASWll+WgDbxYrgm73N/eLBF5gH8bccnF65cK2kHJQAmwdHkB2m0Hqst/M9o4F62z
5Ms/no7jopunvI/NFfyXssxzSl2MnJOTVnK7x26xCMFhKL2jhuxWeg/sDzIYuG2O
XiWgZTG/kkiQKwo7WuEaQMeNQ/1BWK0RznE28/uowTguEq+GSkkyVk8PgPAJ3uG0
2JU2uCTGox4PPkcBuHloEj6wi+95JYhGRl7RyeIrfov2wDw4HbfYcdbrtZJ0qbYB
e9bUqOpZ6XvRS2laZEelYnHP6YeFlzNXZNz84ZMrL+eqjaBZ4/+ty2YZbJ6GYLQE
JHD9sOvjSjpKq/bXVIILJark7uNN+jca0mYq5gKrysB5YKmmWNCccTPo3ZDRr/lm
o6CdTknIWRLlNJi4BKnKFSPqPN6Q1+JVpU3rgMZj99OPDKOVDjdas0eE4MgUT9uh
l9BJU01rYqqcehPtYwR8HXA1BFJDE4Xfe6/xQ3X3XDZIBHNWp0nDOzafpprM9Jd3
hsen1rM6MGzctBhFdKAZG0byOK00O0lcN7H7dOnFvBWFs+bBvcUmtXBmPdPPSg3Z
SjNrjc3JCqznlC/MTUxjln8tztEvlfN/Z4p9Z7lbucoC62hjvOuRJZGOrARtXnhB
y3LuwP17j6CcTFASHw1J45+dNgyQNN9cBmnilMiazTLrhowaSnfav7oNRf2G21Lc
hvpS6ZrZ63PyPR2GUvgIprhYzGyCiutT1kygkKkx41j18Lw0gCbeMeSXSooVBmOv
P2yYrGUr8+w1Y38Z/G2H1JlEVlwbNjzgLGSwY3zBI4sB/q2pOCMnsbOjdPJcHhTe
Uprgc7V26jtOO/z7+ZJYF0Eg5SajlAdh3hoV5ty/54HBHtwQOxlYod4+Wbt+YzGI
KYy/xcJfIrmFkogw+YzBzThTikD9TadjyiA1xNJxSg2EOuszLYVoOKDhz8z25dOu
YAGlmLmYDirctQu7E8LlAMNxG6sLP/ngqce2avT5T7eHzJyFuVM9U89BjdT+LfjV
najtocIyt3HS5eov0Oz68YqJnlFoCdVD89g8UR/tOj067Z+nFnXkyBxyiwalRu9k
phbA8gHFma1kYlocPc1jqSV3xW5B7xgYyZR/91MxSrBeHz8/GQp890aSRCpTToe/
9GobaOIDlxjhdKwjVQYM4VU04u7nDHFLHtNA7hmQoJiMZtsRavE6mrghNSGLxnU1
w9F+ocPJMYcGyV22Sh9bVO6jogHg7CnblgtJwz5dHhItbn6tjdC4wigHfZexvw/D
NiezIlUiXKryY9YMTMz1ypcVBRsN20Up0I2hxig0avYtKZSd2OXIJxASvAu9PNpJ
2oQkkaf5cR/rN4tFtbt2HwBED431POkCX4Y3tIET6O/0FmL/aD8e3ZDhs0CkbfAv
WAnoPkSk72RDdfHRONjdqskgFY6xDGYkNDvt0bMH4xdbLoCILddBXNeURBWY41vl
871xQkNcgNkGe3igK89KFL9XVR88PtSMYaHNUbngs8Y50n0L951yAbwGN8jPr0WZ
RH92hRXqDNGFEb6yAmxlGnl4cFK6e4RxPJWR+igJmaHiwepKT5Po275jnvIfCVxg
n12UVrIdw5vrHDWHfFg+hyY+4GX+u3bEsPJ/hvQGx5QBZKddBSmJh4JonsPHzEq6
nqMtrqNaYH9aScdaHOJUdEa0NmazlcZf1DGHQtOoEGFKzmxA8lWpoRC1vWxxZK78
DtrEwplxN+159ZGOzt2lQFhKX/NyyvEmeD8Muuo+yY3SWgunUGRjrE2is2wkSBEQ
umTl1ke0vBZuqqY+KdQVUU2Z1QJhhuCxivZd6zriTY/CAEDWvnYqdvEUw9Kk8ui9
oR8P7SrpIt863Mlkuj5CuawPj+rRjZtiS1jBrQ6AxYePsp/w3XRuapfSGG7NXHU6
l35k79NDKc727ZY8g5n011INMD7Uv3R8ZeOfESeSVminAe3xD/HYSzwXVOsd2wha
u01FXk7yJYirb3YgMjuz60/0pgiaac+0qGb6RIynJF3hqUhD2+yjlTKGfcQQAgE9
o+CAZwiAl+PszAw3uwYl2VeQB9LztyGI/OdXYLHPVpl6YQfcArkOBaPuT1nCSFRV
y7mmDGdPn8riKpJjyvn+8VomMO268WAEo3nsjA4SB2+qELhe01g563wv3JTZdaWi
1uBpZgqT/PJ8MUwJF9d7JVYL1V0en7yW34NvTqXY2OOasv3pxd2LMmKLWXkq86QO
UPXoA2+eCXCyw3TlXMr5lRN3LsXDGfEui49Yn7oJxT/Xc5HOQQFLd0ocbkDAobLx
wlEohAm3APTG/lwp9y8JbxghhK/j6H+r7gTBMkycreRlV8RdsGD5d40wlRF9uCPY
x8Vdv6RaToZ3hrVN3+968FyxK2Yht7d+goJANB/3CQyk0CVZESUm2z9zpL8OT+Ct
eGNp23EAUS8aeNLPsbtmtiN52R7EYORIjwqu+QiAgaaC2f0qfIL66rbEUCTDAjeJ
LOswzW4u6fefG2Uxb8qZSEkrAeMC0DG6sC1QsV1/4Fspi9pfWaQ+q2hbnmW7G+2p
Kx8Vhb1lYO/NNgyBKuxDZUx3dIKgjof9084qOdCZvmiIwXJ2pSbxPKEK8EgcMvwD
nDWwKCi3inCQFa6vcx097T+GzcsaVSoDL+sT8j/AFrG0Iw9t8Cn1kbx8M6Jkrz0v
8VzsITB7+eY6VF4fQHu3yyHK8AQczo5Epjf/Ipe31N/s8zA9J+vjvU43ebGaT8yr
xHn8irk++AVnJkowYqg/i2gjwjt0GTRxPeLY0tOyh+PuPw5/TyUsruKdyh6O0NvZ
DEgjNVdn8tiKUxHXu0VY2v2KwUArY8M8MhKYHGnN92mS0uWv3CU+CuTxxMn1qcQw
Dig2wNp6/sdMVJlQIe4luUAx0vGUngiPyBvEtXUK4TN6bEkgWwM9l/oDxuOVTObK
nn2pU9WjVBM78I9BgV71KhlXycosSlO9j5IjMNF7LklGMElgrJWChJnmDUURHMdE
Si0+TLScbMiEEvpphFXyFxzuJQKydZ2gfvvwTT4qltoSMibJ0k6jxDU2fRdEw8IB
SHYOA/rbyy3+IWrv0RoL6cPHaJvzRkkTLDt4wtLYbCrCgaeDYrXbpWRliAJcGLNH
x4vblb9Zdz+UZaKaj0rZkGtPGmLjnhOPFifKdkDNNALY+ymUFsWE2iu4hpO7/kKW
oME5YvjTy5vuPK+6Fjym/Nf+79o0HHumun0Um2uh89+TY6IoCnCilgLjezGaET/Y
fFokB8IXGVPs/EX4PDs0pbJGDku+jjUOehtdoe+pvpiPJWrmHMsn6bNPb+D/pwi/
kOziUvt9x/Bn6WER5Gh8jjtYwOZhXR3gRiwHxJahLZ2Nx87uwG8bIccONBU1kSrA
NJ5GymVVIbx0ZHJE35LkKxlMS3zYcb9ZglcIf51Nhsca3Q+6uzsgryBYP1/ltgMu
zPnBfgIv7+e10qFBS3wAGdUdf4kdtRXTeQP9AE3lE2r8P9PGE3PAOlnxxXxip6wV
RbNxuVjphIHBQ8GJ0W7zQXsx5X1YS1UPOjJTs2M4hesipuI5iKEjcUil0IoWpJ/E
XEsLGlyt9hauoIclxQvuhrj6jDxwHFX5rBzbutEeVF5Jq1ww2Jgf5MPsF2yGMFYn
nDcJqGMVfCz17eVIij6NkarVwsDN4fFAi9cMBK2b5hl+1gYJ8dsZ6JIy/f8mXUJq
xJpdBqsME3+SxP5eRB/CnbODp5zDNzEzB2a8eIrtFUNwHHkwMdkRG6SwDxGiJDVB
kN9TGXXPQqJYiT00mevoIkkULMwo80T1Koa2mW7M3HTDZM2hKjzGp5AE4hlkG+8X
x+8c5YWLbkkc/G/bNCk4GMVSIH/brL6jbFX2v4mbhNtQT4Sph+3MmuWCjnOBPnjq
0pDwQJYAWHECA0TIzgT1lw==
--pragma protect end_data_block
--pragma protect digest_block
VqXWUYJEcQoymd2NwAe/Lrr5Yyw=
--pragma protect end_digest_block
--pragma protect end_protected
