-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Y2rOW7ZNEf3IUjbXFEHI8pftiMs4I+xlfob3A5ujxKR+hlASBK2boTffyfoDC5ogEcezgY+0kWtI
SmqI5w0/1HwzNRroUn0GwR7vQnAsMC29arXKMQ/B2Y4Hn0HQ6R1udwogc2rqDi/3kXbngIJyb8RQ
VTACdrzBOC04+aIDjd1bXNIKDp4m51A1MQK4Xu6QR4AVTHPwr1uPpLSAbu8WxeaWSqEBfGEehGIy
3NLDtQQBoHoYIiyE69fHaLwrg5PqhUwkK00VYeo5vZ8wVagOqzVMLnBAh/Du0lhg3O7xVlXh4Oun
Dttoj0upGDT/wNrqOBbMbtGA0fhrYBfJK4J4Nw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5712)
`protect data_block
QareY3qcROD5jTXjo1JzAVSVl5MrqizctDRsUdeJWNlJxU4VvYEkSRJorO4/rZcfu1aqzH3Jt9Z6
X7sTEcpLDOkwM+pDLlfeoNJMpsHdngKBnjva15zesg5yvcW+nVZoWXiwfZdnHeZqMjkVAbFVQv7p
o+QrwN0GEKyssPDGrcnnIQiawc9xAKmzsDPE/pv0ZXRVkNPPQEX7weplSgCtfkv6I+1n4a00Qk3q
jLjcQdCk9fBOvaHwO53h8Hc+M8i8o7djBDzqwjUgl6qiTKjfEfQCXQ6F8hiQM6CGLarX2nMR6kYp
Zj+NYfZih6gbYzMmWuA4Jl9rGraPKij2atkqaLSmAlVWXv/f1etugC+C3NqMqxTYytAbU6N4Ykbz
QgEKwmp9WcfyQlPSeGqBOCJb0rhfZJy7IiArjBHHPM7mVppSZK9jAzRwLIkdZbTCiLj1afv2B7u6
G0plrdlWRHSuEt+cXK9ym4Au0wyAvvTnIsvXZfpTdjgouNf2Gb8s+E9q2CdyZHRfPoxZ8sO6gpEs
WwomDMEoJVsKMup+8oJc+rY6j74hLgdpoSd7JPm5SZMOOaUGKKf/2Btfo8QA3ohh904b84Z8xL+8
yipQgJvLN+/bx7fIvE6b0Gh20aIhjjCrYDUK0/0pA2SmK9jrVLQCizNTw9pPmBzo+SxF/QsYf0tX
JGqwcnbL7Y3THKVgPRy5aE7x2L32DZTFgQbmjQ2GEHFBBjejikzGdbRofYP4NPSNkDufWIYz4kNH
r3DkmpXKVqPN8sqYNTojdrMoXlj71KY7fUk2NLNit/kwfI02D0d7zIz4hDRkFhuzqQpDUC2Q26Fg
Qdo9yTZimHM1tqZjkYtOkEpeA3FZc2sWrN1EoZq3GeLrBUfEbCdQZKRjGLOi3W6x0KvFw6nglbSD
1qfQOi6+jwFZG262Ndd0WEZzwDLnGQlhtYjqsB2Y2SIHf0ypVYuqZtD2hnvo3l0B3BUslAXJ3kss
QEbVmSk7miZSDYmlFZxNvZXhq0gJSx+dhuAKr3q6LroaE1cJ1VA10npDjTibfHNfcAuxREc3QZfE
KXNsp2F5rsrZ/Ry/KUb8jt8ld9doYq36Bleq8qOId8WQY+yZxQ8qwl9XgmQYBAhmcOKKWKCZRdBG
Xwi52kOdfwbPo5vawfV37fS64JpA22eMlhr7hixJ/54mQoXSC/kfrbg1Q8T216Zx/TTkhZBaQdRz
PP/wr1en5KLRAAqdsotTnRR+4cV8QdJSlnBi0gUDSVkppmDrcFxHHWFQ1voqDqu6ukp/EaDBQkMd
wYaWxZ0p737XVyYDm2wxU0E8Y3H9lKKaYy6Iu587P2YmOKDxcqB0HqnioOFvGkn/kNauvTnwgCzI
J720zBnXUqpQLTYv3EamfkihPerJHw81sF4Ypz2wnHkqSpo1CMQQYYVdRBBX77oOEij5ePYZJ18E
HXLnTCR/zovGlPJc+3cf81oxyGLf0N7Gjw8Cz0xr0CdpjLvYQPkkO/V1gvcgaa1+zonudEEUhps4
LFSUvnQoJeX9rZ37tMlPqv5F9Q3NGrZggc7ykSJJgKiAK7oKKbZR3igTg0HXPPRLpXguFZrm96rz
Poh7gfMxrkFNuR2pDspK8Z8/bfNijB+QyvvJ0qxnFYXtFfkNSPGbplNKnchhp/KkuEe6/RAccfmP
6qMG44sIPxQ4XOcnXwiqGd7NoZJdKGLU3j0hcVn8w58S4dEYwpMNEZvEOVXNAjRR9tlma2vA/chz
I6Bl/zKprzsacqpQH5hkq+DMh+8qT54KSlXYLgRZquG41jwXCYHLNiDNR7BqYRzL6L8+XVHeRjB7
4GZH2FDBs1KPhguv9K4UCwVj+hIanVSna/odmGHMK3ArfFu+KOO/FaUQ9SJU/q1g5j3q6pKY8/+o
dm7Fh0azPhl8vD314nVektvEePt/+GTrxVCbYaHG1QGFTD+XPkbLWu2fGwT/BNadCIomWa1R1vDl
kRzcDuJc5NCMB0zFTwI6A4IXu2q0L6KUIH5Uhiz1eLwcgo6tQsA+93dV5voRPtzq55KJIYnyNchs
1x/b9umYup+tympjRqKRY73D03aDn3jeRKLmq7eD8mA6uoFav3hmCWrktOrAnZ9p+T/uu8EPDTlD
Q3TYgx4JFenN2falkkCXWa+h77Ibo89PaVTz0r4f/p6cHuSSF/qzn0x46ZdwbrKidVf56/DTZdcx
GyzXkEl2eBblvEsRp9/OMxUm5nvRyqiiZPBsaL1ARkhMsTKKQ6hanYJUA88f7XbBKgTbwWsudj1R
gHeTfT5M+hpLcBvLmatbYqlNG7bMc9atb+MppTWbQcmR/33tMB/4m4CtO/53XMDBFWL4g03+cMHc
u2Ra9udIQmwh6xIWKqFKnaszHduI/Zy81DlJry0mP2D7aGKZNmFtQcxbwIXcQpUkVNSBWWMU+NZ8
lEKUqivj7T/rv35xh25RsTmfF6A3FBoWzfBRT8rRoFibC+CyKj+tWKLM2iK9SftNsCrmII7EI/CR
0uje8stPOwRYFyaPU/VIE1UkOwSATMm93C/DpKuyXEJW6zQFlfTHbrFwvLPt+6j6RCdUOuPRDRa1
dD1rNXfOQ9f6TDm4iwA7+BoKG65s8RR1gyoi7jKiL8ctQgdWZhRUOFJq4v2Pc2G+Js3+iubyCkVQ
zsc80lIJnGm2Y1/LDc+8Wy2UpLUE5QKsB75Xqo8L8fBRdAJkg5A1qcbNY2MZFN2zug54KMgCD9G5
1xJOM4Y87BZoER4kPRCVtZiKfTLFfbhhf9RFPZ3YPyiCwJVzOGF1cpvQ8+DCq1UmY5hzSkVphw2x
to37zj0jXvrutazJ6iKEoewsmVoSaxcm978kxN3O2TUvh+1nOF4Cc4m01tjvXxciFxA6kDTVMgWj
v9XrvZ7CWNIS3KX7w03sLjaKYISIfHFLJVCm4WdIugGh+y3VFqG/5d2fY8DDbPRZz3668EvCZhG8
/Xmp23mnvW8F1oglXwiBnGcbrp5fu63qomdmj7NbQ3599FxRZvlSwjmnm+9FKh7hy0s7bvc3eQK3
8tD/61BbFo92g2/tVh8BtMT7ddrKfjKIcT8v20Pd3ZWYp4Zzer/6nF10XvvulQPdCY07zu3qxv15
81nTZDHZwE0Tc11f3CYBh7aimH4oKAyfz52LdOy9jprqU2/xvMEtUwoN/t0Ms1UC2W1f4XB+ZvJ3
ipKmQ77GwqMGQ+kfjH8FMXNTxiOkEigcG3jRR/WXOjyzJ9sRbKlGCNyjy0+Grqw6admFqqW9op4E
myAnLZ2uE6q5u6qh29MPrG2YnQmA3i53fTQ4EbGfhdJlybewiHQTc2Y0tv8JSgkQHuMVIZDT3DEZ
TdPeNwGjnOd/6Qj0etDONNNUemAaxW+DLnslAktzOMUdRAFiM1zmCfLrLCzBAkwBbhXowGHHJuxd
2htYhFplKdHbvOhh4GC2o0yv5hpKnB0UIlxTxrXtPr0hRNC2f807ICqx//Kc7ZLiSbGZzXgqkhy7
II87qa37FSwWWe5HIf57bIftBo9yg+P+Y7iudS4yepf4Lj1tms6jHjwGudCgCfU4qohwUoC1mUie
VHaAjqdCjd03QszGaY0xIb8eoL9rlUmXiiHvTD19JHw7UbXkIyRynAqnxpSY9TRiAbTNDxkubVGL
GM0G5J0lSoFGT4+i5q7B2/0dOLxayPhQpWRdIBHoe3ehI5w7+7d3f1dhpa/xSZvVNeib7acBZD1Q
Z8d8hL8w7p1Jh/itgNeVBwRwq8A8iUsZsLVo/MmKzkB9G6T3IQ5ejml+mwj1nNQf/P2SvFbStKxT
4KZe1RGhxhvyimj2rDS0ljcOz5ThP6bhdqPgWsZ64XeBCv+BtZ3NsdkZ74nfYUzOsTGC69e+4lSH
JMnHuflOlVJmbZNIcAPD6ATTkff8aqOjd0sZlOw043aXdIOoQLN5WUk0/1mxzFi2LEYYKg3ijgYm
n9lQ94WgeSpkVu9I0rB3zrrMiwoxpaXIDzYdHOKx+DR9eO369w5IWszrK2asJq6m884THVu2VFXQ
pALNf2SxVlItpCT05OrZ+wlgRCcxYJN0mDZ24q9CJ+x50e5r2+qx0/+FUKNB+LXW5m5653fe4qjy
J2gaKVystkJQTpqOlqIfc4c+tdwn9x5TTnkzJmgDW4ei92WKKOqrw/TVUohff6O0Dk8JADqhnqzh
UN5a2RXxcbmthXk562A3pp20eRlZD/3yRz0CoLwyWCZPmeacmEdykkgQnv69BDoobM+cxOlIlJer
qsMneTWeCYiFA80sK3u2D+/g8xu9/HmtFgsIClj4KAGyjaQONTskIdzyMbHxNmg17QrEKR36ZqfR
F0UsUDtBrszk7ARocoqeiUh2pRWZU9bPcB925AGe1nniV/DygSGx1gEkPJ53QTrTAS3118XuKXa4
/ofaJoUfGCqsIoR5O9YjbBL2j1kqwnmCsL+atYw3smc1WO+V/yWst7uQW2kO0kU4bAj81d6X/ApY
ZgvS1BN5JLk7+e0+NntTHzFf5wRf55yA8w4xtVQprXIm0kl+KrjfJaIQBWEUjMmNfWRntljOq29F
lajIzxNPK0iC5TjLk1nD/c9eUjQ9B9H1G7uEVYuJYbwbl3Q6FK9Y4uiueTIfqdZVIKxlrdP2ZgTn
NvXFA4j8GR2qkUgarLj+bxmRB2Oq183qGUE3GqFnRavkG8a/NH/D9gUv/oPBeoGg0jzkA6eYJ39q
xaQkRx0yiUAVSB4irobiwORH7k4ufwXrHOMfhQ4GSOJrqrKvSxazk2X1Gju2cLacFqHbwoUtovSJ
/VU0EhczCVoh6lqDdBI+uWqBtkIRzumymRNfvALOs5qRlxAIRma/7AsjDciOZIHCwQlHnZHRDyAB
Drpa7E322uRbRw8HiVBrS6LWSaHZwGKu3qzxBTfhLb/qY+0FZEeVHtQwtK7VxpdBLuqp/+xiT/tv
Q6oo8UNZlOCFXrWVSCdz9S0+PoEHSFbLdRmInF608g9u5Pcr6PUpMRs3gHMtG6gARRFndqrFxjyJ
01trNRpoxpVmLG+3limpeFHm+TFyPTImf5Bh2uBf9KpLJOtC4XyaSM7jdhrirpWTMAE/9te1tt94
uBdd5oNiVLs8mYbnmxNMS3sFckaxwCmJeS2qkOXeFhA6G2CnV9mIOscYh64RRHP10ksWoHQgbfhZ
rkXGN0mOwDRGyWBNjv5OSHkt/+J9Fat2/Evfg3Uo0faFyUNfkzPlI/f3WBA9i+LT95ZlNr59Eez1
cYEMb8zGhgc91GZyT/fXBLHcU/I/g46Lt/B6NRtUg8WUFjptkZ2Y58PrR30pRd0WBQ70pjzpD+fN
CK9XO9dPHULcjdSerAuW7C3deurApdpbqSipMmtGbc78x9u0x5cLLP10EW1W9vuxSwWY0wCPcIeM
yAI55KzDb3BZPyQJf3oKr0yIwtTbAPGarwyTaezZPuLil6pp5HWqQPp46FzVyOqRhg9L6ezthKxP
LYIVYjQm4UX6gbcgOj0PwMPBKPzasIG9KhZhHqBwLeD3j6d8Upipe+xHlUH1xHxadVC/KTZBOV/J
z0xIbztVYG7g5lOXCbgRXrE6kqSEHRLh7t7zKBaVM/JPSIStk2WAS12LJjBcg8vYNnVPHbVhltHk
8I+jJmMenBUbLV4rRe0LrXniSlsm1JT3mcwkQgTrxAhCQCBnb2Gtj98HtEBsaA8wxeava7k1uA37
XVeQI5uZ0YvTKhMDO23ZuUvmwhiMR3kzmTFN7z58IpZIo8EM8FZiM8S2eHzUK7JHbjKmkUfYQHkH
S9fCzkkaLMogYiia7oi8shdpnTyW6Us30Izov3W3v6mLzYd5BSoTuvIsr8h6/QuYbUz0Hu9Rtbt+
R2l6z/bUto3o/1ijrDa+YIPygyRHmNL8WqB9AwK5c2GDwujZZenkAK/BZVqKKETwjp7KC+EkuaQ1
ED8vpB6F1TGKaPHNMRwqiF88XBGmr4Wc3MKP/XrSznyxHaKkyai4fgsJnQL7OLmYuilUIvbHxJE3
J24tWnumkVIeFzsSMtfOAc3+9gFztsgSlkYFNK0G+gHYp5DUIthx5HTMYEQOnCMlZtLJvmtraSW1
ea3GurrGE+eqpIX67wy/dooh+QZ/4nQlyZrx+z06HFVtqZ/kflQdmhS8AhAWS7C3FmGH6/nZOo1F
WKsZ0BNe9Lr+exGimQNfuMqeeB4YRPAxHpFH9xtAg4n5WMPmCAnQuIu8XyL1B+Pk1A3+xH5ERw06
ZhYhA7DAWRJODxkwPqIHmvCZfWZNGoK1EhHieGR8sRO5ksjrdj0olIrr8+HnAgqzDlY5dLCXhr7A
QIstZsfF+96xDI8nd1CDFHqmceyxKpRq9lPm6guWc84qWczQ97eghTrsTsIlZMkslFxtmDD00BhD
+fxPxVkBjGp/kbQt02fEqud3tfg9LDG7IJ4EEG/LUVNgPPY9xEKXBsD2mMX8j+edtaAFAvE7WKtp
Z9e++6+c8480KR3T+wZc/SURuHw+pt03gM5VhuZfbMJP2O2FAGAuWAdVzB+H+wEHNEKFJMFz/EOH
tdZ/t5IgGmgVwoaUgoHp+qrMn3N2gkkCOUzRYXzIWpeBmTP7K3edGq9qgrL8EVqEcIOPLIoWl+mr
5OETNLl4VRHGZPkpymZLH4QKqiAmfHEtexZIrXao0bWXmXz1otf85zZ+RXsxvgPkhC8D8w5WTY8D
wo4e6XKM9eyh2n3JJK8ovnNTdTHX2Ub1oX1/FbAbsUsvxGceuVQZzsZIsUTNAmJQqqqtA239jtvu
ndFRfWsxbfgfKiD0HkIMNobDXOd36smnMD+LLpd9Ld32W6us2tMVMrbclmIbDguu/ChMFjzgQFx1
C4F+k+A3wSxZPjZ7l5Z9zR9HUvuKR2EOb5J11Dpz2ZKLQhFNFhE6MZcTPzT6HblTmqwxSVEw4RzM
f27YSnmVzLeL4/sUFEU4okz4LlqilWO7394jdmYbIKfB660fqmCDJZFQ+DneRLapIRNsPi5B9mcV
hrLYj1Rl5493/9d4YlqI/OWoaiOZx4n5dHrK1c+fLCEz1eYy61wBFz3GG0f0Sw+85sc0pYf5DmNv
RE0GNrvsMxbDtGA18uYaOLuQoIfgnAYX4jWdf796i9YHTdFpzXTC1kSvkM5Ve41M1m1tvVErLQ6Q
p2ZvMHncehggzvmX15jiar2y3NrWs4anqrBjmlCxN+InJ/1uUu2t0oEZ6IdKVj/h5qS8KpBbbsKp
AXcFwidhzSbHzbWBdtfJQie+46yZwBAftlnx/Ogy+h9Zyt+F0XIMJfaD+N/djHA17xtW7GPKs1Lf
wyXjL7CBsLvY5Y68/l7SO/RGV/5syhBV3U7zvS4PFzfOdDpwAGZeJoVNiRmJN7vuem7Of/1yX46W
VzqHyvO6H7yScMkedslbigvijc2BHI7gqZ8F0NZf7/gMlL/1I70XKsJebzfxVbhmCyP/bOzgL925
EduSAqncf5Nnp+UZIqXVMufyzOC3V6aJnC1+qu6gzT3bTotkDudzzpHWL1VOemyOU9QRR/fxwW5D
lZbbwfU/Vqa+pSLzuaXtTZV567vXpFy5Ye8v4yXcKfUbzKwedf6vQjn6WfWJ5A5eAT89TYPovoa4
cYAoeUPpYTaG6bfE
`protect end_protected
