-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
sNvDpi7vE/aSA7sed1EbDzsJUBn8CNL1P3MowCDh9sQzV4IYpm+uGicAREv/mV9H
DRvmmOp8qIQc7l7Wfl5vovVkEPKz2YXVJFjXxCXV3IdBSW+V6ZA0glZbj3XNc4qZ
0dO+rEmy2Iqa5jak20BLar9dCk3bJbzADaMJMRbelJL4+zpMrJHCgg==
--pragma protect end_key_block
--pragma protect digest_block
9C0TKA/CVp/P8SQjkYyvCP3ZfnU=
--pragma protect end_digest_block
--pragma protect data_block
z4xr5wUO89OsArvUimZvD02oARkjtks5XkjXYrFFshJZJGp+K9noWmXPJBKyJM0n
FJ+YeJUD300+2uY0++Bo0nPedgKvNtWIaeV0em97lawRdY4J9MjHlEeaicH2jAAl
Aljtrnxn0c+nbZULjTTdEIT8KmGrTqO61KaZKiTRaTtQIAPN5WBoADloiS/YDUX/
kvSCjFtGpEc5jW/XYf61vafgH1rGTa9qE54XjtKhtjmA3+v+e+FJa+iAXDUQ4Rqj
luNDzrc9S6QlkY5qjQkLrCLJjCrWvWLZA57CT8o2StrkY3v3ft+tXkGv4Uw4QKuQ
fWD8XA2ew4uarlqJGRxZ5nhEd7LylGkfpE0DdUOhxezVkFmCG8dyi0tQk8jd/9DP
PSki5sdZFtH9RsCEd3Pv13MhMb4bYlW1GC0SguLd+ziJnBFRv2RQe742wk9fzlYA
z1H9uDpmZZtTiu9FQAr5un0IDOHSM0Mk4S4wHOorfyikLmlHX2JCQVGY0dmZQAtK
e3DOOFctEozrBw9rf43jLLXz+1faJdXBzv9qm51XP+iDFRLYBZqPBjOqGzE3rl6S
4BWeBnnTinTiijGkIQRg5SzSHkWHe8QQQJHIWFGiu1ts6BibwmjO3zOVZ6hSzvzt
0YTczr6t77J6Yut57NiHKLjEzXJl3g6FXFJX2+q2FK4Dz5z6qKi+HvkkAvVCF2Qf
9oUphVtmbtK+VLmA7IEN5RWeOoGcdX2eIkTq2xbD8i6X31yhf+eC5EnAHnaXL5Pm
u+cWJUGb3xdq1pqqRmTa34DB07DkYMoqdfVbkFScbELGxF5qH7GtOpbdgFZk86pG
LaBJ5dYA5N0wyD3P8hrG2ZUu4AYRyQU1V+CJ8SbtqIGseMAFQu1wMska3a36xjj0
nB6aS+U4E7EOce9GNRPa8BMu0NEvirgI4wYJI1ce0/XOZfy4I6g6LzHo5xao37QR
Kel3WgLyiOhitpPLO2ZpGeSH20EUyJkTgj5lH1GX32q9dkau5Fbbetkq0o5OtwmW
XoyGBYAhOHbCy1dPqo/Cs1bahR8QW3QbXL4zx1wISMPJHoFLfp7iTRbhKQN9EmRn
dCgeqTf6i+CtkS5xnLCP+JDwDQemjHKQvjgnLYKxlbSpPb4PHrXGupTOXiKKmPgD
OIdjMOELJxCQILV7eYswGvT19fNzOOmT6Q/4VIiS9AghKTa5nIBMwmT2HX4T0yCd
ju7vZZpa+acOmICI1UTP4qD9XyVz4ACclwrFq4C3u6vsxO79RDtTBXx+XTYcaDK/
9S35rW4aaNRAmZdp+MOrHG+M1kxVuJiS5juNTYeakmkBPNCjVDQVwdD5TLdjjSsc
UqrrklF2B82OB01sEoHHoXUDHiex551CqXpc9zZ085x4FtFUF0hhNDuOh9w0H52/
y9jgdzU/TOS9DTjh/Vt9wjf/t3NvgFOA5GxL7DK3M3JMPwNiVwEJove32PQNAD8g
yRNJRyhJwvCEJ0Q8BzGW72SO1Qmq7+ipyV5ettusBDBroZFShr3YJr3fs91VMDKR
CNFxe7WdPqxhne1A6Okad1nLKWx3PssKjUTUcEMeUQ0cN5bg8EzeCDU5b/AAmlyr
1r0M8s/oa2D+HD/XUqu80DxeWmFtVXfWNwYVobZendtUs/m4ptD+rLk1qeS32Gp6
t/ny/P5alpjRhDK8AX8UKTXa6oclkvBB6HIvbMLcJb8HhgRwPVu9w0vMMcIzvFBT
M7H/0LPxO0NbDgO6+TAG8nlwXbuH6kt2sFKCluWh/0Xl2KyecIcCptT08v/djt7p
RI6asThXl5BSSKYOwrA6AUPQBbB5IstbVYHdPQLEpVxNV9L/rtqTs1C9EvGLX2iT
t7s9pBGvFvGLCVuHbHIK3Njc8fmQ3FuDcvxcV+VUJaurcHguLM0AIrY8yvCMx2DB
Gof4/dWoXs0Omhb4pEyWDDrSDYnW78TnGfbVx6pZF0Ywt1VLo1sNKmHXo9aTjCjE
WnewdMQh5wIlvWq4CA03pH8uF/+5C5E3ZoYmGnmig3ZHC4eTwqXUldUiWApJfJlP
jwTLXrQsu8ctKPrvRrsYgYjNrsjLMD+Ovc/EHONJGmgnMWrt/iPtd9LAQvGaJByb
vq4r5yvnjTJ5vGI89eO1lI0/7uELIdTkhdJ3QimZpJtLRcIvT+RlOJlYbSwLvB3C
hHL0uNgQ0eeZTtzZDsEhNGfa13A/nrtyEggdqMrjuWgl4P28YQ5iRQKcr1Rz/7Nu
ziWs5NbKuClXWM++c99h7XFQsC5pZHSyoMe+9jxCG0+XgNd+5okZhr4U9vB9gFLd
t86oxbTRIluRGNw9OjBufUwz2EzBjcdaDbH6N+hkt9anNyeTr5qUmaJKp16V+K9t
uZ370V6YLcDshp7YjE+PEiy0eocLWD4C0A+vD+k3mf5wr+tWm2lE108gXIXLQk95
jgRYMaW0pGQk6b6YVFU+Ahyk0fcMrr0P/F95VZGsvztrciOY0wjugTD+FYyF9KlH
Qd9F8K7eEe46I2NqxzCBKK2znB3LFc/GZvfP9nSEXFggefsSZOkNRXGJr8RomTwk
ew/qyq/wsI84fNSrwdM4QcJGtgd4uPIyEVo9YWdd7sF8Dfz9ELV03Qf6w2WGZ0wq
BVOGP90nhmiEFc6IDeRxASJc1xmRzD3w6X6yqXMpeYOln/bGRoO/jlLA24/eaosf
Hypk9UYCPHjjOKbP8cPl2i6+4wpiXTk/KcizS6tcguzer+vMsgawNYST0Peo1BiI
S9PGqqjwus3IA0FbpclgCpaLT8S73vMYgCPmozZXAKZr/Lo2Ao3rZ8HjZ0cmmCCq
WQGWOW1gKWNREVsN29AtK4tN2ig9Wav3bumOfgfK4AGGd5O2SVlEAcevS23nU5/p
eXYSdOS/nifhg2YfWDuthptGIGrphacU3NKiPqKrsC8+YtJ40+Thxw7vWL3PvQpy
m5XkNbke9zG+RpPXDzbV/rilR5u+u3V9hxeWyLHIFuJ58brXUU7zcQiPUgeAau7O
twp+5ijBXgclu2obUaeyWtURfwjm/qxamTzJoC30MsAAn1BrFVKtegXpARy5TdMy
i81iDRcJYiFkXr/S3HKQ7vk4k+SGjBvkUXBhwOjV/dL1HYmkaIGIC/p/KV8BkYL8
c9U8LNC71/rPyT5rLgxXRQKMrxk7Lv3mhC40WMFT7TEFrrFWPhTLkNO83954zhzG
TtyyuP17PrBU/dbbeMOAGos31zJS8KFSGGvroGv9tFvajTJ5FUhZXGu7/5Du6ZFo
rcbehvyVoNYKuEz4J98JMARwR/tLEzqoDEc6Bkhk58adb3t8zFym4I9Z237CciQz
c/IW3++1dCXEttN56tFPH5VhIIwNbJsHszy5TbH2+Fw2pOsEsjmoSKhQ6UJ/9VIh
4Hbt3uNu9N+hzNDYISjeO2Vg8vtWmTB1aHi0nXB3bmdbrXqB2Nb0k+lV5nxUs5UV
G19zRSOOjHmViwIsflEyaOJbArwt9SgHFYnLhQKaq8vUJHhBOvGjyXKh17Hk0vLj
djN8W2hetokBe1tAchXiwspKEHs24+w9y0W47n1Axe7RmNLzRQ/RVUwjjScinWls
XdXspW2sV2ATojjMvbMd6tWPXxipru5LVKBZEb7lx8Qiw/k09MlZlGHc1SjHNbZR
OD1dWjJPc1nXvMLn0MdDMDsvHS2tJp5IW8mKvBOu4DP3bO6CYpjsLucwBVw5UnnD
gZ666/FVYoGyZXqn7p6gZsrkfPrt6q9Efx5KJ7Tnoan8ccFCWnGPcJ743N96/81o
f9wUN9bvkZ6vQlzo/sZRWdKsBd0qTe+DFHJelkTo9ryLbFdNV6KvfdzWwvw4r8G1
ZReXbmmb3vp/zU1sGOsxB7z5+mpU1L6HTwOxixbYOEq/zWbmZ6Nxc3DOkN/7rLcm
QpxHHqVIV9H+bY7HNyzmFQDLkR9i9lisVVYR4e7Y8aOGcaBL26fj2Zfa8rzZPplz
Vr++JejE4U1yOfI4JOfXl0UljX8dRj7u3qDlGJ2Cj1R/a4PJUJL39kYK6um+QN1b
kxK/zUF2wmlO279bY6CepkTmuMZ6KqLgg/B0icxc9CxOBRmGcFEsTgx6mrPgB4Hz
BMULNlKHqZAsbnxHZl6cJ/8gx2YjK2lrOIoXPkDGQregHU7J0nBl5/komWIJqlm8
zX7hQDEY6n0D3S9YA9WiSSQQM+QwqCGxb9aTcwaQzkFJmFLGJMwrQuggRtyPJxW6
4NHYpnnYOKV6esIqc+f3C2+ZQquBGDB19iZAscBz2ux+BL7MHVjgQDKv/ZNMogga
px+TkqWfvEVRMffXtdBv5SnEnxYRNIUmfFAxrCGWTSJ6L45LSIyBJKMzDGN9tY8H
vwWrsa4PzYx2E1rNIH0RZrpCshIru9okzGIn8kGbH6rNGKGcrTI6fUsaz1lJvMk6
0N6Lg7KvwcGFhHsAAuLdkz7aLOkL/Ghal8eCe+8yqTyKgeFgjx9usH0tiwCMhgGz
BM1VonamOM003MvET879CGrI/xbuH1pZrUiWntk22guwejrYdIwqc/YZ3aoOX/tk
j9c1MEzrHuLaFcLZTzKPFy6N+feAzhHCmDPqux7knaDkoAZInW7S6s+YoXbVYIRo
iYgz/zviLK38eZnqxuOfKnBnFwbKrzNWH0gxhtWkmB2VQmyYuzvKykSgIKNY5d+Y
nmpyeqEvpeLvQFa5yQe46o/3v19ahtWdqw3PE4iTq1D93P2KcxV2JvM1NxLqRFdi
q1VTrzBktQ+6T2XzYquLsCPS2qVNro8yqsQjdBUHZxvL0DxbyLOyiOr5UQGOrSs0
tTzj1bhIESgaM60CvJi6ON0sIOtPQFjYYLXm5a8e1wCxHHFMlUrWXsxLDs3B0PZE
iIkUhSbXWqKabixkSjBq45H4bRPiXB++xBp4ALr4h+K3+84PyzrDVeAGfVmAHGDz
baoFfP0gItcB2dllJ1Hf3NdFA+lBQg3BrrYvJRyWZb1rmOqVzp4u0D6x8+tXu6Yz
K94foVwUc/IKRLVnkjenGgnjQ+aq2nvAIhjZ1V+h7wbKyaB9J1MoCvMDkeus6dOe
7EN4tOPxT6gsSIdTPy3Yhjc5ESiG3hMSkhR0vgPwClnJyhN1WUVE8bcZ9JpuTYR3
5i8VPwpyuRR56GuqDea/4n+AHumV6FTV73DFg+zEzI230I16KNmLu7j0eAPpzyJE
VHzQ/0bEe2S5R5Mt7TKLBqaZSuMwG5DvyZ+9ci5H2lsKEyd5kI5aEJhCRqy/7N9v
VgSzU05+NdRSC2imLTRlmPATnYjelroTRrkyBU0eZBi5E1XAyLkO02SotNh36A62
eE5IsgbCtEOWNzhG7Xy/h9ip2yLPisyKyDiPvhjvwr9SsxFWbu4e3gKFWxEFyQjY
H9RFHO2eDcj8yYSZfhkDfryFdYAzVFK+2eN7CPyEAjRFFcY22PJy6vRag0uO5lOT
Pnd06+SBLdTVOuHLSySv7jKDxZtO22DLuE723X5/4ZDok3DPEgWwUCJ/T3hoXIsC
YxpELlZdvRF8s+Z2qiiiQgvudmtVmSz+CPCkTujeSU8IRI18nIeiiHRPVvuJD1DT
K8F0zrSnxYKVMUXiHrJcXsNZhX/Kaw5y2xSq80SupPm99LnzrVfEKX2usjaqts1n
ZYkZXtcBCZVZoSfd5OmV+95QmyrPb4pfPhNMPRvlmO7qmdgU8tChknCpN2t3HqkF
jNrT2g8K7yYizxCueoT1a36uxylyp4CJGwmGZsL8aYmhWFl3+Asl0PwZqOlWgfJJ
q+Q9oCQzrUb4oGlZn/5sgoiqts29+aS/m/qX2BdeXKoPzS3F6srfJK/XZk4Fgg66
JjEETGqojw4GtVy81Xkh0/6AQcelfEG3rzG87jrFUo4E6b4/mVr/KXY2nlL9k3l2
SY9QprlDdpO+e8fAfH+HLc+x0wMy/o0ZRRbvI20kmB0Oij6cEXCttFGyxsAHcqLn
GoICiKJzL/TNbjA0GQTMxeWhKR+otqP4TcqVGFv+wmbCIH1rE3eEEFtyrEvqrLyu
wnmYD+2IfgQI1N1271+ua+010vAVA/LLGnisBWhq3ddDmM2nIJGzHuFuI4HhCLui
/qmrBOZimNtkPoS0ucoA8lOnM3ruo9hHyS0YhQrdHxanh393EIx5vhPgaRNwU+XB
39BYCfuqbfFu8fCxsHWxxqliRZq30nWjpzjRZaIDwTO/ALYYLq1T+kZ36c+moQX3
qZMdJqx4U4+WpVdubKc5IBTjIXv4JLQtquFQ16u0LjM9SIvlu1bhexzw+wyw0S+h
HGIPTnguV/a1aggClBrUdKAECNO9c/kEGpOAmnwvHYUyPymj5lKq9QVq5k86Rdhs
eMYtsjbzOER/FBNiCLbCW1sd+qjUSppYiMxH+RqjIM/tXTjA+fOgS0OS+GpgaPio
+jO8J5Ir7zB3MxAviefGldH43NGZ5dPEDqOzdl1ru4yWht63q1r9TSjGDyAtr2jh
iFUD/d81UwPzJ5ABDD211iCIs9QdoacVg1lyuU+nK5Lg/AIy+bfJ6HWokfUQ9vpU
YT+sPJ0hur1JuwBrQywMGrnKD0TrV88Au2ndjNe7iVEf0ElYAIBH8NjycSOpUQd7
6f9IOrbFQKBJKM/1eY3ZVcOmQN2MtpUZOxsobihObvW9ApRUkqgjrYRDbnkizkQn
R2sW5GN1xfrHOhPnUdRFo3Gmac6pTYHm0v0Q5xuQx7XFo4lKfAskA6RL+V2HJsRS
2pq9cRhZjAmN41OLeYD6GvxtyURFk1Sml77t/FJosQNYYn7lnbeY+ggxQlLbS38N
lTgg8XyJJdj3LzKVwlUUOH5B+cd1i3L/zd7FQ1DPA4+KvAAMhwYGRhE97zatvh6l
iAbQDC2PzUDqoqtsOSXxTf0O2TXhvOxuPlUjByAISD1pvDL0hoEzNNWaWPFcO+DC
6px4wLxZ4p7u8/u5UclxJ5DaFTVgIQcJFMjr1SrAasd7fjNr9h+GOJUcbh7GBFSC
oDTI9nwJ+cIzPhw+oVH4oQyGBOqOsZd3wMpopF8nGMFDuPz+ZY1Y+Iam8YmaByW7
h2uAZVugjwgbKb9NTeLWHME4swdn62vkXB8S3qyuixm9PbllVPnFlHrfKxpsYf5D
x2wNYY9UnzUQD4QbuuAkcUCtX+I3KTmqpzgCrJSOCRz37EAwV+RHN7LYwmP/HmTq
WCzkoU68czqSHZ623ZhxHFnKINhEyRD4LOLpKpi3auT2xNf89H/jtAV87h+9avmG
uRh9G4rr/z4Efzb75zpCXALlIt8tZDXITGoX8UIar5KGawk3clPoxQK9jWEf+yEn
IuOKvsXeduJvuK2gJFdxOtWKcCVFdK31f6KJf+SGc56LND5lDaiNZfdfbWqpceC7
mPSJgAGZtIhnbDZyUmoqfCnGsTSAV6vjrDxvcCSWyyAdPxWjylZmNjL6GYZF3lSW
80QpO+VfCPrlKq/D5cEBVMqHvfiuk/b2g4ybdE4WBGCJVl5Nb/p7a3TM8bj+5RdT
ECklQgY17gONY4Euz6/DoJd99kfj68DSWev6j6K4sTuhZv5gFB2uiomiYpU+ZD0P
TN5syMtO1dORrHWOoqDwjFpw45TWYjZfTz7mDJlZJOJvULEgrOySIMclfC11ZoSe
KcwQVQDVUJbSV5wIUiv0yuqiLCHX1Rj0ONC8lMA7jaOgweXmbXXOMbIhOoZVB3jY
5L2at8Ke25UOOTwix7SrIVpLM5oHJr1Y9bVqweq1HL4M5wJKCx64/mK5Y4SLGEF/
k5vcilYbHim2WaEq9EB2xf06TdPDDhHYS03BF2MnwKIte09A4cWiK0Xx/viGMsNo
1/4ByEMwH4KCleqBIz1N+EdMEH6zaId26nmtiiwMC1HuFcv1BsrxTO2ZCJU26Yep
VbpssxiHezFP0IiV8zBtknY0eBXrc5RzdKJr6W5VIxbJ9XtlXYPlma8QGZWZDPG0
mWBONe3Vwse0QOeUGBxKEzGuK25jmS+k2QdnZLirkz+a6Qy1YbS9Lk3SNWDGlE0z
/izkcxv0a/kzQyygMqvvzApTgNCdlSNwBNC1WYQz7TOKzVKL026BnG142oSkW7Qa
lGozUZp/+ik7/UDfhlOsStDCu6CQbKumoQsxOHLHNMdpA/KuuVgkRmYi+PCUTR0t
cragSj0e2oZrTLtkLMJ0jwYC3d2oSTV9Ytb/mKSBu8+gzCT8XlzdltSqk0h1jymx
gzfLOPW2S6nPDmLamIAmWeIdyl3+UwnWpz0ADtYdfGZB17XjlyXtWYLS44EjXm8j
QS3036QxyWG4ZqGC2mjwQjdgrLYtbZbQrmvPviuGmRrVXvT+o7rBnY9+nKYIw8xB
EDyR2LYwduTOvaGiruu7KFTZJ/OEp/1STbBomXGIlFAo3TgOhAazCYWlQl90Aqtg
bXESOxwPqBCHuK9RCKvKMeBkUrbQwWFqsWZG2QGlOMObPlJ3IVMGgWc1ZRao/M84
XknL9gCBe2HtntgeYVyWizD+6orrubuGcGQE+peyEcmEeUhxDDbXaTSrINquFLoF
WZjhE39zc08W/l8rmk6X1QzIyCuho7T1PJ3GWPm1ACpIpyjeN44WfAEFaPuyh4j/
rnzhtjc4PtmkvEDCSkv0bZAV4RlvHRFLemt6P93EckQ0cMP4SPIDPyrH+P2SFLxt
axbMJRdzbx9cFl4ryudicztIwXnExikFpD8dZRDWrPC1gypmh0V6LFVPKAj6VU3J
6ihwxcoj/iomWrIlftofx8QSilsasipnX8EWdl6qiM51cfBgLY++YNbtVDzva1ER
EBTpsWLf2WAOgnWugX6glF9vrzNKc3BVHPZgE9xF9x/nYe0dxU2cFn2tgrRh8JZA
q7ZPL9jS/QiiGq2rTLEEWY2WGIYdlYB/UDBlP1TM4AFkyZqfBRXdiEAG/zhSVFKW
9LAWe6MJYwOoJB4HrAxRmcfZ5AWYdSQ/Kj8jxhKMElC5bLPLPgTOniBtkG8DYnKw
74jMNuyGtBJ3n9jWl+tXhEealmZ0Rg+6GyILcvEMKPRRgCQELGWx2IUK+GZmO9tc
/993j/NMqmNUcPzsYPPdR48BWUWYkAvZwmTtd8AqiXQI7hz0ETYuXSVTX3m1/x/m
/lOhYTxvoW9uEdzYoLWJ4wnxC3JybG9oyfNTFUf6dq3qt8RsShzXeTAFoqbTpqg4
UTb0gX07xZS5BfbQndNkpVZ2g8lzm1+o7DdHXlWClZs7XreCTLXwJmA9V6MZu0jv
ZuzMbjBkNOSRXOSGrGJGAzmjROBpHhCUPldKcup54KCwBNPWaGU5cXpwaxIlgVaY
BTertJCg37Tp4R1eO2/Vq8olnAeHxFBBWeY5adZIUgT2pjA0zQWF+q6IQcq7U0ry
iuVbpTCAq1P1pgJqiQM2QfqT6fxha4Zs05IJSse1UKXewi8qdYhk6r3RRC3WmRmf
IOkJly8kEBzhvSEeO4qPn2d5k7ypMdn1tv6/0XumcRGOK9gnz2Qg5cFEaHI80+NM
o2uld1c4TpDdOvU36a+ttEcYjH3tfjohk/m9ukq+eOt5NdyPF9XixxzOSXaD19lR
Tg4HC/gJdKh6okfQ6z2A5aLKzuHYFWMa9+IX8yoG1E8KZXJHr1I3/LN/PQCONr4H
u/RcsoWEtXWkU+hOo/A9Lw==
--pragma protect end_data_block
--pragma protect digest_block
2JzT60jBSatXa80qZFqOe1EktIY=
--pragma protect end_digest_block
--pragma protect end_protected
