-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
C99eoGaPkgJ5i0Ce2Ny7xqZ5JCSJe6TO9gCMS6m/5YDTkG2fyQ4Nn2IZHMxAgdUD
JF718GLwlDlXD9RrD55YvZhoO1sHAHwhnMd73Qn6VeETB5rnMle55ESQHMDlAuEJ
Vaz9TzucjAomhoXotoJtnarDt2oAtmgy0PoJxfCNW9Y=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 81712)
`protect data_block
iY9vmW9WFnMwm0fg+Yf8RBFsrS+/3kSAoigVWMuj+avbOXjwtDpQe++uv1JJZvD+
VrI56fXeFz9Rjrbs3moskTaZTYf8/VxWxxvTDuyBu9nA0RVUe8gSnmCvAP4ufMHz
ajuDuC9lFUJKzD8BeZ5i+gKpVQOCYmoNHZNgJOuA1yfiyFpC4EplgSQ25XFkwyYn
NelJH08cSnaKMzJLpBnYYMrifiQda205e80UKcM5g5CqAjCKwaZgyGr5ATBNYAOO
5Bzwp0shQrr5azY5qCCerrJBWl8RiH3xTTiIxCrC7+PaOhfSzNlSwT0BWsSq2/qN
kSRl8zno1Pj8+W9k4dKosZ5+/8r6CktaRw/wckFxbdmkFTyJ/KKIHpH6GwPH8vw9
18yk7sAHKIIKStv6dh0Z/jDihruLUvmPfXLkE7jLP+i4XHurfvxegE9QRzizS8go
ecMPOMlipmwRA3tzyJhbL4nk4MMlPPIL4dG0UjLECvrYkD0WpJeag5Miqioe4ddg
aIB9VJk1rrfhSoQdqBMyg3JYCEAQ3VzNNzr0Um3aaUT9MsrRnHVEJdHUbBe2uhJF
eRbEgFLwY1tOUhEUkRZpWUYRTf1NfFHwvbDS0KgIF53RahlRQO+adfBCBvbDDcBU
YGC1RC1rrBo7RA2fPC2yrYScjk4njGucPKT2edNSTIMXf0MuktRpCP6ONgjZ7Ecc
ftE3es4PjXp1LFZa4Zht3XpuONwjPu8ysUnmbEFxub2vCkkREU3307ncgOXh2xQo
x0YJuT3oGsapUUr9qQ8DL3uSgJPdJOUrDM5aDxFmp/n6NOvH7KA5sSw6jVJAl1bE
wwyPiZ6Q2llfwGxha1Wdt0OGAePH1Zo/U3SFN7RFwco9q5vuE8VfOyBnyGqVvRfg
0py97gAkdeimkgtIbUKCmpdAv+Rl0weJeqMuRwG/SRZTqMemGBYFgVjtNljQOs5w
CMj40tOSqDCTzEJqhqCX/84K1J5rIinsBu65TtQ0zDlLFUZ05549xDzWMGGVHyaU
lVQZk+L0ZRQykmTl8Ubky1L7298jy/S7OEIHHmXXiBfmvyJpF+zTNUrfj7irQYNP
uP8WSyJWAuIEgPyE7+byk4YPCQaR2hVyRvOWK/ORKonNNuY1fKBX7yL9nArPSiHW
ORz+mpx0XyvM9Yl0vWSwZ+BrPgYaGL2O+gEVLSW+Pb/dYLMD4PTWDOoy0n0qO584
0BAyd+SM2RzcGH7vhG2us91M8jriWdxNFjfd76e3PMhfcybgvz3GiJhfBEkQ9Cv2
7RYfVeg4wlQUb5QMynWPJrv3P+jDqz1ek1fdX7oQV/va12P2kj5plhEEYtAbRk/K
QsU53Pbb6I8Gw+ibOSiQ43vUoYwC3cxOs71vuHC2RXCTN7S1GyDoJSgk+ZjAkWLH
dcEc8ETPnrGzZzEyCDO//NpMhlElTFO1ModajLEW8OAWBk5VCH4f96qbHYgNlcCV
BQggSU/9LvJ54aiOtG0b6tadDLQdPGxX0UCH3CPoN5zw8LqYQ+I8uky0EdYFVA1R
Lh4nB6ateNvvmYCqvvtfthmpk+ZS6IsvGFvlZSjnZFTdUiFags8kcsm8JI0PgPLM
zPD2l2cKF4kxT7Kssw+YENPHSI1BFVtJS12k4r5UtogTXD+lOu6Z/9aI0YaV1+dT
0utXQHv7agHgVUE/nscQQ/+PNVjjiGkTZ0HlgikBzH+LjILuGPze6KX4wgaOVWEU
4qSBpEBx4a71hgpS64cNGzDa8QY0gJ4ZtmNl7m74K5eoLo3YDqE0ZpPmU4oTKgom
Tm02lLcpCzkPTOgHYG8akq8REqwq01hasZc9rRA0Vb2XoK9YEi9wRmDrt1dmVrWw
4uuiBJtmZrz2EcO0+qFsoGeyBW9eZf3QLCTD7aGIeLxrgg9vo1KEshEOFjf2ME+/
2NgVmYloq8BMRCbpi8hO5XjjMMuu+RDaBuNZhSOOOVPzZsJxm21yb6l/NEXkjAHB
4nzs+wmPLwabmvkb4OArqDGkGPxOn6AzZjLa0s1dcu2mwJd0J6XYHx2L2bqPBp7s
WoJZnunASREvBReAiVKfbqD9ebHQXdSrVz12V5ck2iW8PW92F3HoKOsWnrorHYa9
d2sVDK3jj7GEviJQBy0cCe5m+xpSTcNkkb9NGQUPAkfaA465FH3JWZbiqlhMLx/R
p4/QAhY4EwMuvcWIDSf38FAJbWJeK0JUr2xjgeL5lHCjmOFabdQ0YGpjjN2H0wWL
WIikZKsO3BI6h8IeviWuFR8jAlcpDe4veo0Jd7z2T7QU2XYEcoYpRaBUXkANuhI8
eisSBoMeX/eZGtCYVrPQpNGf03ZYc1YqXr36vXCrIhQ0ogzYCV2AA7Xf5kYKF9wJ
ES74zd5kNP7Xsy0gP7pHenPSZxB4Xb88M1NTpXA3wM70tdpj97k+63EhlIuWWAGD
AyF7C69y61G29Trj7VL6aqAXJijtzJdUODVUku/G5C1gHaislA7Oq3Vd9ESCWHcn
ledxhEu7NBjOf0aGZkDnCEm6M+DoaJV34/Ot63LoWxKJXkg+MBJJgBw7R3grX8t6
09iGQmxv/wUlatKi4lq8ftod/U1PD96/5Yq1FYUb88CZQuasVv8SBwZQXfpOo13I
Wyd5KUuroWGjmfzMzXEZFV91OacA3zVy7QTMRM4+HHivW6M6HHMEWBWf9aC4r9HD
qQUooYj1Cwl+8wfto8BDY6rsfhktZUkvO8oWmH34YbyTGCRHQUCEJbM2geVoIoR4
Aa1Ct14xQ+ACAqbP73Uu21vzrEKSAHXfKgCXeFybsYFJmlVVazv/ik09n7RldXiM
HzyuuHrZII5xIpOrCb6TJqcoGjo7YSw9YCi+ShthLfr+gP91S00pRrn7jxLs9YYL
9dtOa1RiQ6b1NIaLJPh7QaguS0D9Rs9m1VbpYP0Wx1FkUcvZe0Y9HEq9/ZXh7r/z
F1d5vCqT2Yr/TYGM8SP8soth/a11LjsUZHT+Oz+5Sn2JPCOKp8kIcNkGua5a4RDV
3MRWHFEvoq8zE5/LKgYOnoawaCeBAuSBE1pbvzlok3a+rGm+sehkhpMIL9oPIyJO
Qo14i0Jjqk7hSf3akJ4hCCJa4ltGCiSevRZ2axQel7TJ3CZ55/tH6YiHi8J+q2tP
WrK8SZTpNGUm29tSbj7hoypWVptplMKQL7T+vH465nayAnog3Z1u8WpNLNMnKy2e
MSjrIn4W5UsAVnUnKt/9oDk1N1ZuJQRafNvQ5Ezm7bj9qaj+4zglH8vLVFjzlxQB
1Wtg5vwjmDKbpWYYFz2n4aO6i6Y000bhpsedO0RDQebsJXUT+FrZ++37Aavk2vWj
1s/yPpqgot0bndlIp6thCuf5Y9nhBpO9Fdlh/h9ieNhRiq5U3HCA4CDxOA+yWFR8
eImnWy+ABwIZLXhO9u/kp7z7PDqpUOc71KSkD8he83MGJaOw2JSnpbsyjYtqLFkg
z9L77F++AmGR20DTP95nuhUEDF2C9YxnESV9gq2wsytomJwJdGZrPFX2QMnhdktv
vqts1oCR2NEKOTtqb0o9zKARbPAxpoV0QehezSGO1O5qBCKvAXQAjOB8TT8Cmmrz
mm0SrJnfl0Jh27vPMfInD5S1pF1aaSjv3tTWkST7QcjlZSRExJDSdDlcGjhCeQnb
b8FsTK0MUqyfexgf6C32DvfOFPdmxlwhSLSvy2rmObuYWEBWd6bM18tIDrCimjv4
OAhssAgOEWnrABZCnMqE5r3xFPMeaeMprT+y5/ufZb0CWeTrv3Rm/RgIBzzfhjIQ
ICfpejPS9rX8AC6mhnLdzte4v2ecKKrVQIdPP7QwFzkARH8nf870v7WhXhAUx9jJ
31p7fyj4NydpnmGL0bkn8gs01X5yszbFbp5Aaun0yZ48jOVo9Z0ck51wtbf125mX
jT4Ton7n/P3xYtAxhZ0n/ybfL84MKH2O+bAW8cV8LOdVzVpgDknONhIbU49OpZ2o
v7MMm2zEu2BUFgMIC598BLxQcvhh9o7LQP/L+daCt51acXhF7qQpjKFKFQogJf0b
LEdN5KeD6+42S2phdVqOw6ugAGRpibTRV+hIkpcSX5BY3wGrHx2JxCF7nqqsx04a
D7/WwqM0qlhoYA8yiwflMLj/iEsAdbwnj6lSv4KN9T7EHf5VkxVEQzj5+oHKv9XL
qDyn6XDI6juyGLBwfQm+0UD2QA7c4BZprC5VGgjojEDZEoHWKvJKr6CztaUE0RWs
4kYJD3aQx1YzQ/Cs4PZGiGa+6kQRgj3BqSRYpX2sKtg43YkMrjGN0GnZ4ejhf9Zy
9pT8rNS0L7PqHwj5Wx+nQKHV4BcswqN3dmm9W+HFNCShjrG+6nFk16lU5/6777hl
lFqvSSnkAchY+cWr3NswgI77h0irnf5Rs3vC6NYhcR+OjFv7b/NRunjW4yz/Bzrb
3cSH5cVhCfQ/D0/b7fS5AnM5jrN9gs5W4s+PK/wdp/Psvx4gwZ2c0EfvLbjxZAUj
SnJ2A8WVUbvgrNyhRCMyzEWIeFVO/jfMuq5qfZdFWgyJxz+3/HKvziIlElFCACbO
Xdu+uxDQHgw/S98zlSfcRhTJNEuu+xqQRCTaP8uCzrB+IaBxYn2FVDwEKK38dLWr
+NQep+lUsJbS3CD3Z/X+3Z332MWfHLOObGdVmDN6gNBm2iI7drjiDZOHQT0/u4fM
9+x4fh8aOoanwX5Zojvt1cHBLE2Mk86dUsMkseHSDyeYC1E2FJmjtKmlOiQ0bpJ9
mRi95RmQPpuNvRPqkWfjw8TJDGwl4s8HecqRzSPL9s7wUf6XCxyqA9W293OuHxQ+
HicaMTfukEdPjLJ80GrGLbGEEpSFiKAWmyHEcE5kIdCy0pZkvbxVfs1ZQPOIj8kM
Iy+xSogurGKC8J7quMAIql7oH7SmNeRyyo12KNcgCQBaLvoy3wBreiFhzcWNPvd+
H2RNnMHHsa5Jrxm1tR1FgJEWeuhzfAEDbrVVMx13zwRcvx8KvGZcLkSGdWKNHFek
W0L5scWT7reNeRsoR6OBJ8P7h00FDlhonaNCVvVDOxsrGti3cqNiPP+eE2slFbNB
Lu65e+dtNJyzqYBjHuv5lOyhaEYTx6aaRvK5rFPJ8W/T2/FoAD49qZbdnzU4a2q5
e3LiZpgzMNmnyG7CfbME9XTDww/CSt1/BuVTx+NrS5NR94P7eDj3cMMcfbohuxI9
fnR6phtNLMPZDNEpbeMiby5V3mxiBYWABswch/htILjOe6LvgvzRSawAB616jDYz
gdzaUEaw5DgziqYAZrKQeYQQsmcrUtWv+9jzk0NRvpR/f2fMSD27j1WI4jXCzT/Q
cj3RMhBebMQbG+gTfEg9slkQtGb2ISARDx/bMByZ2TAFmTC3uZUG1LV4abtYhLnM
ZQdZARZoZjPw+1gcO7OK3Q0WF1uU0OYJ2ZywTsx7Q3WqHYCI0cW+J7Q6tDNHdx2L
fE2Mbmu4obGePpyRu5hPL9DeDux8Br4Ujc86eMeCQVVREkKlSznkPgcHUnVKmVlB
jtbwVgmK/ELvpoDODE7m4iERNbIgK623js+nPhSdjWKRhKz+i2y0CdUXCAo3Ew30
tT+SIov5L7H8prckt3vJ0xVg0wm7McJ9b33g0fIkshd9KtzQBS1EWN33xGsvvx7B
9c2WTTVp94RGKXBTN01vB0GmrJzYKV/2Kv+4dLnq4pqm9iNjwOoR6X8bOP6mVMk2
CEaQXInNpMNZnKI3TjSOllxEs1BJWlqb0tZAnUvuVvWNws0ir8a/wo9feuQPg2+k
k01aIuNDrTi+AME/QdVeH9+MSb9oQRwVpzmVsE2SrN5h6pd3a5Zrv/wontJWfS8P
sG5A8t7UAXw+3zIUXafl8fcIn5NcPmae2RVTDPDT3ySXHEnxsuGKJ3Pe+bmS0kKo
EfeQi0Kb8z3TvckbLA79rrY3BYzSDQzoxvETzG58Xq/OLe8+eG9zaoxrrTRIEBsm
O/yCtPDNVwq/rMxGV/vrwO3XYukZcIUw2vwLuniUUlMXcXeJeXzF6oC2guGlvnUQ
iXeb5pDmB1zwHlaY/k78d2di0VLPbRN+dv4FIs0Avate/MZI87pBaAA58oExAtxy
WO/RevDlDkX+l4Qjlkc8al0wPO6DevXxGVwCsIUDMf7C6ESx68cCaX0CleBFkn+x
HLiAa9jG3n9Yn+jfr7QDiCekQZ9HSZXYspFxE3H7MQbRoAm3NI1cVAd1VKg7dYmG
1DZDjlm0nssANzorWNoxzkZoKmN3n3kCCXuUhFIVxzkm+OuiKLwDdyhHdf++9ZAY
Zfrm5bM+jkKRQGqspsLr/48iKDQutTNLZlpnCvhO8JPw+yT5ws1NB30lGoYz5yNZ
7QJTFoODyIsVeEks5f3MPN5wkIgR9GkQHjd+tSSnmlXaKOjmx0fR7RGwCRRoADWU
X03ve2/Mt9Qbjng52cW+zYpoljiUm9yPK8Tm58E+XdJEa9zZ6dvNiOc+NHKbKp3h
YLDkzBXH3Sw+2XpN4DS38tD8HfL/LeKhsyqYbhsqgDA1kK3oa77P05wY11CW/uT5
QpSeoBkdo+Gp7Cdoq7o8JBD5ZtP9ikLspPev2Mq4dM9Ig+e6GwErCK38+R/IDdWW
mpbyIpJL52PaGJ0aD8YY6I4r1ZloqCA0hcU/oTolF/E2xYlWOIuPkBklCmzw2uNC
cPgT/k7CWcErlEiPUOLbNaAl6UtpAXYykljNmpbCvOa22GqyBJywz/SoI6fkLFEK
2L9kU3mADJmACnbVwHt2Qx0ZgV3P9E0vGHNINRiL0n1tffRSlpNO7N9zVmhoQzlK
igIEgBXnlhmdPFkE/c25f+HTXL1RAaosH/FD/+yHqVRbihe0RFCAdBc24Y1kehKQ
2huQAFvR4ntq9GOkDYRs6IxsHf/LLuvcqYYZIHKwl6nTkqzDThXdXDWDw+4IP839
bfDNcUrOFA8mVM3jP2kc7tuKF24NL69nuvHmE7O3sasvUYKpseG6I/nyKW6X3geb
Jf4AdA/xfVvBgGwfb6HFEDYfNUNRPiAl3zEfAUcu39a8Sg5UZicejXdwjli80vGS
vPY+bvChVFO9nIY1AZ1uRmpEqiOonXGH5AEdehacEgSRlcJ6jN5IwqSPeTZQSn4U
5scnugRkZ0vz3GvDLOZ1BDBkVxZudPhbDBU/gzg5CO/ZOLnvDQCtRGOTbG9cnhHS
tZSveShjoPglwb5KULHoQDYtMSkw160BLU3G32CFExvjUcg5lbaf3NbV5GXpi1SM
B90vTAwQgzMV/lyvSulYmSiqan4en0moTdSRN8t7yuBLVBDtZxCq2Kz7B/8suvXN
Gapz1l48rb06uoCeiTEUPiOENPk9ZNRwzMumvn9GFjU2KqBN4mzNGJYAt6FX9q+h
mjrkA00Dbc4MxFQX/PiiwFvWftPnT2GpIjELEOsnpLzMsOMDN8WxNapbzAtXRj3i
bgmkbEdct/PyWbEYpxK4FCmXGOc9e0VfCCEd+K1aQ0apRXN6a/fjhgEhll+YcDoH
RfVCuiUc+r9PxzrYjf+M8pcrK096OFlFbbczU3ZAK2mLT4j8hvzOvUoRojdX/KQf
8K4gmEJB/ehV7FaV7kezJLvXKdESDTTlmps9TrPgVQ5Lx5hKnLWdx8zxqVSiS+t/
Z9c8ZMp90V7I0Ua2ahYjbc1+K6EF5NV7Gxfoq5XNl0qZ9WDxfXjP/ukF07tAgwVF
UyYLF0f0riW9nw8VcTtRnNtHrHEIcs6wWm5C2kxABWxQmQHW7IR2+rd2wW6zt38E
65y1tmN+1+7E2BAP1q7uhaFVqn53P10MaWvGT+/Lzq9jH7ZLSfIh/YSz71N1hZNS
gEusiQLW4zTDfXe8yEqPq/oRMDFMHqaJlctt2nV5cpRWutZ1xTO7c9UTJgRlIxhs
B5Lw9OpNluyvyOuFlgKnxbEe+SCulRxKE+8uUaUWFb4IF5qPqVKAviT8f/BbUp0g
KXQdvcoYDVP+ATD+ZsSxHONx1Yrs7VD67ZoS+L8t8lyb3/1W8MPTczcm6wDMrAOM
olKCBDGdnvUcdH3810BZDZt2E9eaRVlrwZG/W1I8yPxO1rYQuZoi6lomALPDuDEs
EO5Ko5WdErYMw2Rf0XXm2w6meUpAJjQDPM4AB5wV2Y/1m2l0mKPvvQ7qz67Pg7rH
r6liDq2OC+S/nY0j1fjCF0UXkX9zkaiS2ew6g8+WbF5CKew/oBJVCvv8/azr9TJd
x+SZgUW8G0YPj+sjEKCK4KD36Mr0wr5Klt+hDbax7sGREKakgHNO/as38KyJbImP
OiSOSwZDIzt5Dsd70TzLA87uqHsd8o4977T/4sGxoIrENx2+K6SoiUxOhiHZaHk1
w0tRd/+aqpktQiuz233hOPLCtZ4M1OGG4E+2xN6kA3Jla1nLxRCKcQHlttdbPKWP
G77Q4VDAl24kxPu1SLX0WnV+U0qeQG0CDH2wf4ElmUdZluDEUOO9K3b/Z8vDT5//
gyPceep11G7h2E7zXWAN3dzDLvnaJaLC+ifnweC3JLfjOBUiVskX33oensWhMlo4
J5i3wdPC33ssvP6lp9t8qHjVQQT8BnSNlqCH1cWbs2QAzdIer7Ll7G4Kd/L2eJ+a
yC1JT4fjhDlj6OoqO+XoPm2u8lmavED8xGzdrm4/gak9favB6uK7ZDKWbNOyc/e4
RGArN94vBnAtN/9bCS+A9lpMl6JwFmDHuSNdYilxrOw2qGoV/zKr0CQbCHss/EKT
1yoRqPxGM+p15s8wQcTWASFnSWYyOLWWsjo9G6024mSWTAx8HzII21eYkjQWHRyN
DBHdRPHTAeJEV6pvX2jALaiV8P84BEibmeeL/rOhDCZTk7N+NaSpBwB97Mr8BVNX
1ffW8uGVn8G+unCYZatH5Fjw7q1prJR+VhA1AcxNhI+JEZEhR9TNVphWIbvjElIm
j6/ykopWH8AMCCJ8N5OkAMG4zBuQ6HbPUYRYXGjpkLqjC4zA0Z6FnN0v9Ngu7e8H
SHc/L9IZzO9NeOWsJWsrTv143siZNDzR460CE3cR4Fx8xPIzU3719r3hWT5Tpmdn
lbvttJCmo/ePPY/PHyQgqhpCLsBd1GPJhRVYLpoxm0D04NRnFSJL43eeZfNSRy8J
TYrJtpixz4EIguEQpTEd5c3g0d+FvPyNsM95+8NP9mfrdJDUNRbXx20U/5cwCuSD
+pGQhF27rad8CRWdITMmjp9lb/+2DErV/SuMx5NaC6QqhOO84SBQSKZQP/FMp7j3
lYKSQ/nvgMiZYyy7yMuO7iFlJFNqWz63P5t1OqWIwiab2hmpRJ7jYpPRjpNFSc8A
6X6J1BiwLFVFZgNqUulh95HzJrHuiOhfDxzhRMYUvV+MCW0lHNuDtTvMsA+2755J
0XQpjbAYP+E8czFCX9Zx5ZbVd5g6m88GRE7xo8sgk5SJ+ZEfOrtEJcepvAVb7AaA
GqGj2e+vhEgppmEe7XoPlYpW4fxNxGaNuE0Zkq3V+2LZaGtiejn1/0hgiIPSpEVv
Wzc8G5/B+2Cz9Z0DEgsZblYIOQ0JiX7rJZibDBsHCvQ+hOdLY/Sm+1/7VIzkuBS0
pFSsmOxU1jwvydzqDtE9fLrDFmGq9jPzqqiQ3YGYXkcrdEjcjnwoqUVXh3piVwC6
55Tfd1DcP7dSH0iOKmx+UjVQvcRObcz0oHV8e1Gmx/Kiq+/Z2XbUD5gJFBYwg+Yg
nQ120C0/TEKt6idZQkPgmzVk92Y5WTVGJu+IJSgCcfO6t0e0ZOdu0/fTc0cB36VH
v0kT5Av7NZGdR4hrIP5n/ZbRiivk8dVLjTw0tDNLAq8wsRAOa/H9tQNkP1M2F+9B
cWupsyrksuAbneR5NRnf/Q1UZ+O6YHgy3cXVhPwlnO0ymv9OKHTEB2Fad9L6xi/C
wC6sNofCC8x4o4ZHoIvpudA4ZC+j9nqIuSIsunzK+naRjzo9o12zaUTncYE08XGn
nMpU60Ga3AkVbwVcvyWYrHOJHlyHe6AtmD19PcYVRbVKJyg6rbpTk5WTbtkcX5fU
0Ij6SKHCWng8wDnu2nBwXRUrxy8Su5dldJmsXMZkJlaNR9i6eglJVC3jQcbkoaoD
74w9g8sogyBsIMHrDYqEAWaJ9RJajDYj/hoAVLhJH3WffgZXI+vJO+96Uphqd5BS
YBVegTSDYN4aE9JRmVrEbihgOlNT5QQgLYyjyZyPiT9gluiYMCFIg2MQqghAEmQ0
0fCtaX5NQeFm+1rxSabbvdAixSIgexlAR3bAAUQ8i/MIpF4vZWlOHNsUr/+Yr6n7
I7XzDhvkp+Zk2CgNehvpvrpG6TzJcCCVU27saqoQefdSoLRkfRDiW7Y5EXQl4eWj
M6UX4nuejD73njAsiUxml+vEj18JWcuEVLjXBN+7CCLj5pthRkJkyma5p8IlIMmU
Zbz/Eh2dB3pZ8V9nclhxhswrr+QWDZ2IaQk5njaBWX0OyQEaOEPkbcTv5MIHcMOf
AESpWpjoACR6nxd7SOWp1DP6KVsez2aDORsyMzZ7+YF4pN1F7047EFwr98ch027d
ptkXF622tf3LyWpCfAJSJCZlsz17Rk3x4Sn6u2q8Fjwx1Lfj3FZ1qlec5ms9AdRd
EFZFN51ilJUZwZwht+J9OlJiVf41/Z09x9VcUdDqZUG/ZPelHYaJ4e21iuduQeaY
cGAbKOAZtMI0+YStWMScvZ6GfKPbRdbd1Ty2FQmZS59bV1vkCkS9Fb3Cck1lois1
O1MI+CndxeCHR2LPxpRH7HFDVpsOM1K1JCKEADYquMnPWgr9fA320cTK1/MSX+pU
o0EBpt7SCSlDi44rX9KOyiYGB+P4zdtdsscyjqB7IyMuTv3jJe1R2ggG1OfX3RLb
ja0UKsvUo+TWh//LbE3n0jrG1RGOrRUGRGSqVwfKJ/kOyVbpHFvLtVRisXxI8ih4
u9y9Vv/5ekoswZ2Z915/+ecdJJcXsipulJqhClrTGheGFvUFko/Ty/GtGnfJL4V6
YnefJ2E4PEXvXaD/pDiGod5zUwRFM2v7FsWsVG7GQg9Zx4P5454S+8e+J5OdBzHT
xhRCZ6ud7KodFZJh1Ya9TMTkea4BVl2mS5XsBgp0RIc135NHdRBzuJeFBTcObJWC
LDJ7B3um3HDzoaxEfp/QzwiwJ1KdtEuxGchStWMG8J4xG3Y4jHHwjK4q2aMSiTkw
iZVhLiz7nGxkn0ydxHNvjZsTfKJhEjXUA/PH63PfYLg/hB+aSTQJhosojeR7G61I
i530xyQOyg666b5yuI2w3Yt1KQQjqtb/ifQce9o0MC8bHZoh0NYfxZkOGUoU++qg
ctpOctCevCxcwZEoG4+kcMkuGW5Y2Q5ITJE+6EHgnIVEjVSLAco+fTvmrIMM9/K1
Gyo6goJmjUdffxEA6+4EVSXb4ZUlGgBnRg8J2XN7M5dyPtvQMM0dwIUHKHBDpR/P
HtgOOwY4Ga1Dh2zk8gcQi6SxM/tQuF9J3/Lh0Gb82tuqjmAEaavBF+8p52g5j0q5
pTdJKjicDUX+vfeKVRkXouo0tJaxR6wjT8mj0L2+p9tG2eMS4N0YCzO19tLFSAEV
/CLyLaHFxTZKoJZknqvy7/lYdocWGsz9qH1hXmU0gQo4tK2qALt8XDEBOZG0GFgd
Hu3gObDY8CwiI3qFqoDxCP1Kg+M23QJ4EAj2Gba9pA7x/5mZZ8aXhhaQgERGRASY
7VU8b4nmILdcKsExLm4YOVXhGLbLjREWQ/ZsUwFhkQxD3FB0spYr+xI4IyCMhbOr
IKyAA77cIhWw8R5iyyn6g3p3bIOG/qp8AEBZk/zU/QrvlXZRtAIKJ9Z31MtGYuKf
5QA/r1O5MWVo00GLear43x8SVEIzlQmMVwCbjPzMj2DTtfhKauM0VAizTjFbCYVm
H7v33o+4ADmLs9qa/liX8rUE8kZITA0ec3Ja+MToVLQuFcnNmxTidqarrtuoWX+E
R7hARuH+hZU0WAjxdVS/R2LruHp9KY2eUpfLbbg1CH7XgzFrIJlXU/xVMv9guqQo
F+PN/hYNfdkDG0MyhJe1CFErhg4SFk94dhh/jRKKSZVG5CqOxjn2Sv+fi/cNd7Xa
WDPrhsRvFCTLAQdWJWSjYxr/MeJcB0iA981c967MhYjXx92HrN0Lw44fGQzuj7TW
KO9LjuOIaTuBEavxZgREgmbytl57XQOav4WW8Ei0+WsPGTdUjulLsnxacpWo6ZF7
j6FKV4Tedn+ZztTREb3F1x7uJ+LXNZmlvgM6ebg0Vt4U2JHlkk7CM7y1l5xJG9K0
DrFxzsPtumBvssm9noK9mIES9LT02uNFl+nX92Cg7uKaMK6khyULjqHHRadZqtwq
OMgjL+fng8XyQe+EBYPAGXl9xeRwZn/Mi+pE51xxFmCTBOGLVYE/iB9Ae2bGSQ82
jyC4FAux7H0WU4xRs85kVnc432sAapj9zuThjYM7JaCQM8s5dx+WQfpzIA3LugBy
GrEtynCUKXZdqyLRRL3aqglnkdxEKr4bbHkiCg80nOpo9aI0WrBi05+IwgvtFId6
Li6jhI4JRObmrJHPVXmpe/vlmrY1MNzl8m5HC/H6AwXH3EatqiOyls9WaCIq9m7z
Hk0dtb6VjurSuuEYGs5vddqnNM6q/I3Dgo6Ue8cdHdNOmepnVVYEiD/LP6brS5ei
C9W+Oiz9k3GsJuS9pzM9IqSWUwIqw3y/MmFIsG/7EXPsetiDKT0yIug3yopwsE6s
jCptX6TxRwQCr/5GOmhnoRT4eQu3JP/neIBl102ZWzPlUggyTuZyMoHHtMpnigAT
pfeHo7p2m1ZRfxTjApT+rsqYilCitBQd3yzsFmXo35Vpg3xD6JKeV12d8cUFLOjN
ygtOv2jdTvFNSuCsw3gDDD6ONrTbsv6H5KeRxZp57SY1xhzr2jyIWOkyUWGbBbE3
JDfrBejZjk79qQrE6Mj1YVa4Z1Mi+1eOYmlaXzEwsKm3zIVJWQjdUc4WrrHhhu3c
N74vBpCk01gMtiOJ7RqEEsSZi6otkDZuyI2v/2T3bq7bjrkUbBAxHS6ZOtvPUOVM
JBW6sx9CuMDwQTQXqHcttkORw5WjVfB88F8mLa3nkGQ0LcvqGbRewRDQYEC4M9bm
grOQ4jp4GaaiXmv8uZZc7dMRqkm90RQF4mM/x4M7hQ4Rh7t4PdDTV/VZnDyaWnOd
qZ/Fz5Y537Q9ZJ7so0dRIPoR4/PTWq1pcT2P1cOdcbx4PSz+o73GeDfUXQepyrZL
J6wNEnK6daraHrxEBXZmtWBvHr+D/1cdO/VX0ClGokjSNJ2Uz5Q4t+/oQ31VQp4a
6kQ/8WCuzVDu+nIKjrfSatoXcphtCkeooHzAEGXjrSxj2vdkPYDdfMvdskUt4wl/
4Gg1Po3V4dykQQURfmBA+LN77oOKWsf+h/wvjvOADe86ZxzyQO51oJf6d0RL5zah
MtC3SDTHUEmIXl58D4rTI1wqbsn69vph4UidUEU0wI7hhxsUcQWURcMMHBDa/jCG
OS3MNEGoipDjDQtDV7j8MoqJ3QYrcpdutgNKlBAC0kgyZQoRfwlfTH4MrwRh74tx
xU6kVHkFKyemEF5PvIY3ijFRyRUOm985T/7h4S+4fUGrgM6/DRruX3/YvcfhscWy
VxUlpErqFFbbKjYoKfhjO41hxIPxGjVsqkfe4no3KEsXr7L1Hb95kfky4JsZDR6O
rsc87GOLqyyvsnQtV1Rj4TGORfR5A1JTN6n8Wzlo/3Q1dmoxntYTblKO94UsVe73
lWi6RsUuRJru/FHuuLdYSFXzJWljHIOHC0QWWJ5mFnemmM96Ue46XdFdsauXoZ9A
QoHrdlqaVXI8sWKQbQ7xkZEMYDnEitndeVw8jKbEWZl3y9a4o8joMuelAOcWV4lS
kQrhyyStua2dmcYAdaQo7hC7vNQdm0kngIJ4C2zF1AZ+Udy1eIy/l+6x8G+9ND6J
aU65CnCmxla5iJjbS2SIaR8q2uJ/1JAO+Lz/O+1HR8r0eE7havny/jgOSnTLejhs
sB9o34GWPry6bfXYkIql8Jg8j+Hqfl6ojg9PO6IUYsmK8qv+0huec7XZqOEDgYF5
okjXlByY5pWBLB+gnyO5zynFlZQSWn2n3K/gcKqTwb23ElNlQ63BhpOhLIghPpFx
v/tE9YHqCzOTD5lF7gHYfcJSjdI78x17SJM34q/TgqP1ZFg/8dmTcNKthyrUFt+U
KvVh8fsdMstJjVFVaLXm6IQ/k1L7Q71RUvas68vnQJ4Erue9M4Dkb5Nm0JO21HDN
fEzvLndWUZ0SkuM0nQEzApTqB1zMgY8Hq6B7u22Xu42QZHQo4655B3m+dWnnxnUI
sirMRNMsOfESMpW6HumalU4fpL67l/Y0+3UloefRJz10IdsUoCQCDcIytHC9q7Yj
68xvg3J0SfmkfHVxlFppp4yyDwEgC1HTb0bzN4NtONFKdzdlH6b6FELa958TxlBw
O3mvNG6K8EymnB80jDFCoN8RDXvGDwrkFwTAj8sdaEmwt7OnEBJOBk2N5Br350Lg
urBQ8NdrOo0vssubmxP6oO8JJurUljNKajIiNRbjrawKl70Wm9ZkO5/Q1Ry3d0j0
g3o7toCIEEzpiUx/CbnE1EgiwDk+5sTIbcVRpP25GlV7g/FzLsKlhqT7NP3qUGh9
oxnceY3Z5wM6uCcdpoYsv8RHMVbMIlhsUZSic1h7BHtH2mN5BacoL10VcfuTGDTQ
4GkvFLECAbWPvNAMb63G6jOZRc1xJPP6pz7ac1XvEZbGB6OE2EyoH+q4IJfDAcT9
rGuuUOLW/P2pKgilp7WTmnF1LcjPT+GTbS1Kxt7T7sa7XmNjSQUPw9dng3cTsNTj
8QXvHr6h1oY8BMOtOl0rbaIM77pBIjKHmi3yh3d/FHu6A54l7GbJq+ua4ucl0Oso
K4dZ5/ZgYb8frHOU6yX82mkgZMcfDxV0unVOLw36j6D68/r10C0OMNVIZvbSIar0
qVRr8mQrCb95Gokh3Lrs2Yl4QSdgxpS/z7j8i9eUXqr2eue7pdjLdo8G2hMZITfk
o5Zk5tQ18EwMYmDziA4x1cj41Z7vKKS0Q+EiVndwSO/r91ljGiv0VBlMM8VubRij
jwOidX0u6IUo1aLd5IF70rc30Esdu6DomxLETrx7nkXLFPJh9CgyVg5nQTc2fAod
ep1BF3ToAzGbjFrg85DnWY9/08UW4NJ/6xXNT/rNquTZSlEt/OQVT/u42wdZjG6c
8loiuP/rFcCzDhvcXDmw5FI5pFYZS6C8wCvO07Rn8l7uDesv8NGxJFUyfE90AtiK
zuawqpTYIlXcF/BZrLTFZmQTUDjbwcP+oAjWiTwu40dATxQ4bT1BCue4Q9qEy2i/
d4x6lqbB9/od7xltLNx8YTu0wva7gdoC8LaGc8iBR0pwnelhRjqg3EHkTfCwFLch
+zVIbHwwyX6/5yp6bAchFLCMj6NPGEGckekGPVIypLbA7eVyhvqOod8tRwK8j4io
fOjDFT9mKrFPPd5eHcx3BEcw6HRoMhYIn1EuHGYDgVU5Lrst4MPgNo+8od0LGBl9
ZjMmwKaVO7pWZr7XZTe2QP3Hms1LTpkAAYVLa9pac5VIyOnXvyXFZP7X3BmTSRS8
GbA4nSy80WJPNFmjuEo3pK1Pstj+n9+UwJhyV7BBjC8V00HbSmW95DRcELJEmHrj
Bqi1ko/SH8zYAoOpsgSUdayDgpQiOiUUPwyupH3aBLoaKo0ldFuIdZ+q7JCckFJa
1rQ2UUHx6a6tTrWLrZkOX7xnmjAhxlG7UcHgyD23rCg0o47t7DLjiW0Kpfey1ZDK
mKuDGyxwea6RjwrnJg10PhBnW2ai7f0tLZzM5cPsYJ+j/Eq8DJa4KbmROA/35y1V
bsQw9yXtt9BUAy4X9ES817GFzAmZpi/S020tucjmKnbv4tFSslgow4xa59kG/egs
kacyoK7ksY5BozDQjCb83uyzh0B9F869gnpOlI/9cSqSSpQE4QKomOIOB31XOxky
5TyUgfQrmxknNROBKI5HSA9aSJxA31Qg6nlTjWYxyiQwm7GWOgiRF1B/ozLCa8Tu
8tqALpgn9kK7jPp5mV8nd38Qn3EcZfGeIszT1o5xyRkINVmnqoM77mY8+42UnMQY
5HxipIb3Qnf6aOq9TU9mWtfX3Q6Ugxy/KSaaAHCHx65PFn8/wWPuwvWyvGAjWacu
rudlou1Jx3VHPu6BA4ThFfjsCGUW23j3WmjM00DAb6nRmxLPs+juFN/5C8wn4dRe
LVkIEhekiA8L2BSpeFade2D4prSO/1bOqpW6d7+sJuKFePwFiTV2NaP3bB8iWDdz
J2YMbLiVQGsm7Z9MLQG+TKumbgsWUJHgX7JgUW3MOXAMwr97625YbDs7QRud+8JH
51RuWxopKdlSxnzmZmggJTZ24bGq+6FLVPxG3A0yJM9j1eFKXo1qGt7PH8kSmSi6
khw+lbxVQsUvlWxcZKY0i/wqrpls0pyFpIxb2x70KkB7hd0/Jv+nCV0cQZd28jLY
UU/aehAT/QIJ6+RF8C91x7iw4yz6Yk9M+MNR0kZJYiqsWjj96R2WetWXVO0UQJOB
yOU7RkNYZNPxM0LdhhCv7dZ6OGbTX2wFTJElERQn4kxv0RF+tmNxwTVnmp3HXcfz
OxGM6CKCeEkyDX7DMqdpRZhLZwmQL4H2hce6Vs4VN4V02E/9UFoE7uA1pBw4dwke
XT0POqX6EbA9J14pSFsQ4N95EkjugYnp5bT9NU60y4tu9+Hs7tPnJk121T1vEgtr
AYGm8/avqb4YL03mVCjEcKkZLxZERhGe3iIQtszRwnsWkNG0oNU/etn3ft+pCrGD
69pinfrm9qiygSbb3ZV3QD+6F8L6+xXym99nZcp+ykqoyvqwryDwRB8s/Ac7xH6l
B/EgEjg8szkOdEgKzVfxK7udXK2Q49qtTWvZvPj8aA6WQ5TLjPF7xGxPbBg69ceg
xHSZq2/Otd1VSJG4iAUWQBY54Vk//26ksu1QdTbCIpfGWaVP5Lb1ErLjanClJe38
Zmappm7DRwjQBUoDyNE9t4q+c8bB9wJzE3PrM8mATF+S3Jk9Syp4j6DIB/xDl7/4
m6Nz87+EynQW3ZOLpHwFfXRw2DwqAuyw/8JVvo3C1sMlil3AlQ3eab+MAnDMKOcp
7i7axO7zBoraNBRw7kYmTwfK5zMZrXbHXIfIZCk3Qfv8/a3fS7KThu04SzzET5BO
Vy+berXpEDXd6cz7UBpGMJeClyl4FUNArxXM6hDmaSeoumB7SguVAuJaQMqC8ywv
oEYadj5aeaHU+yEybXjNV9ALFyGKiABXxcrL8Erzl9kERRZi95RrF/d0ft9xWISy
3YEyN56c8JcD3mE2XKNoUS4Z2W8LRE9CkP7ICgHIknrrr13/OWa6kQnsEfOUkVD4
jdq/Tx3J2FTdabbyaKKhDQrSonKi2zrE/48jHZEzmkQ5+PDS3SNNXsOcWMgwjYaG
y1huy3txkLxTnXVXxfqhk137u9tekqMw7oeR5t9KlMO3hqG80glkWtvArdQqB4Mm
QyeBn4QzeJ6W5TeWZffnPAaofLeQb1niFLnFOtoLzDnDjG8xJ5/Him7IZP1Elm5X
ECUaWIVFEO7njxNfzqKfR1p7evEK4+1J+WyrwUKo8qpbyrC639OVhysq+yliYDZs
1HEoU30LlYfdmxbREpAUPD8iNSyHmjE7bnHHGkTPXTBUFY3CzkYgwskfB1+OnOFP
JFdO8yDQVuK+ipMwrQAGJ86hXGubeLC5+33ffzLeFpQBe3VFHLsUnjWO5IWNDKKc
pp9Ttra8mgzFQJTC54OvWSJX4HGWucczuBbDC8ngeibcvZGb6H8x6avCGA/S6LLT
If9wRS8stn7fC30vneM0qHdxneYJStVU9WyX0r1KU2OVE+t9jXPMHVDq1adum/3e
dTWGCbkTMGmP9ER8hvMpFQI1qqtjB3XJIhnIMIzPmRxH179NCyhGDDV4ioRGkU+H
w+b1hMCCqCKcj9Onk3MY+vfWFHWombXjUX0Zvb/l/b7N6AOJWAGZvE4h4Gd2beJ4
BLLPV8pV3dMHwBp/e+RJ4i6u0ulDzM4WHRvxHwBkXjl6z3g6CkF6YmJCz4ELrmeI
8aeVULTnyiUCTuXzJ63dATPrdB9xqjz8qGmAsBhtoJXAiFqmWV5eYkRph8PyeOHg
eTnkNzoY5SCBDwZx05tCn0/wqRoMJBXNqNVAgB13hqaJUA0vGxoywMvM9OMSWGdW
3lX+osbDiOt8XPa8KSbeZMMy2hqtzowBs+Rxyzll9yUKmyY5ADJ9UDvEqIeVZUz1
ulXkAPLJ1RcKFV50hVpFPXqFov3P8cyp5Wl978345rXxdmDlsRcV7VBtfq3k4aPa
Zgvy3MOJXM8gCDl2MqgPdwhPoOjctLJYZv3ZewDgPdQq7LnWpxbY/HlmRDX3TDcO
igBBdjeFT4t1toPnqN65OlXhn+RnLeRvED9oFomqBIDJ5eM/2PjfDiw9VA3qTI/i
7/OtnsyrL7MowmN6sH2XwycGki4tQ33RmFfusAzVM3QG0Hcltl6X5BDXOCTg3BD2
iuw/BhZGGJV/1jSeKMTVJmA26pFRgIQ3RtwLjaoLmlpczfJyy7Qs+dyYu8Q5zFdH
hK1EvXgD1gCtZJxznQQruYmhR8M6hGtOK8yS3adFCHCr3QgI0Z3rt+4IcmkufCXk
nsXpRiLE1HiQ8v6DnABu6unQUuiOtnKeW3/sCk08UDGFTF10rweR8si0IeG2RJdb
9H+N0kLSoaJPNeTf4KBENkjlIyTFCtl6jbWhvi8DfOjVg5m8EMRvy0zQ1IZ3yFVc
QunaHDfccEoUD/wCHSyDsSb+9bbC7BBsVKgxsS/We7RmqUzcDzy0dlImgl1Lmzgv
mt0OZKbLSVutedpfcIZvB9ZrCdP1FfJhAFaHqdqzYfIdgLQPI0RgW8XpNVXroLoE
UsOJOjd7zAkH18DbEIJhpFaLSBaMvj0ndJQFcS0aifNTsObxzuSq9ifiZ0TF5z0e
RnM3kF6gumL61X7oy/WeMufQkZqYNk24YFxasls5ouUP4n6LcGN88sNcOsMJE4et
NFZyd1ExBefLEd0vtlqG4MNMKerilb3PLNA31/v5fgMKEEa76h6yCP/G7BZhG5ZM
Aha2MrmgeppjYhQMjiYFAQgjKtSzuErtImPoC6s6OfPu33ASLHC7D05GgekAemO0
PFz0BpdDll5Or8vZb5U07LLmb+agwrSYdPHebJl7HXLDyMePzubXuTTYs6iUn9wn
SKdigqgoJqJtC/Kkmk8o9q63MGm7t/d8noFgRe7ORNv1yjJG9Nu+ke0BUFcuL1wr
rxATbEe1U4+1qRN1RvnX3mH+Sv8v1PAD/xgkqWlfPLDUHxmNGiLJ19rI+1mxsoG/
Ra+MJXcU5gLWj4IF8MAaqSVzZt/rXl4kSqcHEHBYZn2caohq9vyPi+wp5P0cMn7R
X7YqlhyNBCcg3qgNvm/Jl08rBe9Clk6fZBZNlFywaIedQLqwdzSAGFnIFD6QHD9O
5JcUiMS16eG2408XtlW1mZLa9XnBkb8ZQhrmdrTQBSWiyNhJIPJSuaW/Uy+U52qX
9LDlo8QIO2BfWaPKUxqqW0zyGO0kBU6XiiJbutW6MEjWh3ks2OTyfm/Yj1UNsvd6
1XaaiZFY9kFC1tKwUxmuVscyVZc+l7JHdoP+UjmzesDaUHfA8aQmFibWdOD5XRzV
Gk0gYepZ+VZ7bmrFZWdp6ld7B0kbqkh/xg2BU+UN2rJ6q+RIcqIlRCrcpp3Q5z4V
jy0sQ1BcKQawDTcrAXynAzU+jelPuMlWRpZzPYZ74WclVx1VNQFDNsDKWoW0LsL2
uPT412f2FaNvDGlG9VL9v8y5TPHnL5iDpMzoobsK92A0vn9bekNoCH8p8Hh0fWL5
HWv1JzABFRBrZQ9lrL0svbvEELBEFaqh+mRpuePRBya1p+K9BSLJNf3wBRtwCogi
ibUg+LjpTyvvCI8ip654f2FgfoogViLXNgM1mfBfCMh/2AGfA9lkJl0Fb9VTlUmM
7ZNZ0unv5R74UZX/bhDhHcMUsYHT9NtspS6kQkRwUTOPbzdGaDDhOJvJac5kg71p
COnrntK+NbiXam8QAqXVu7iI3pyOzgYdqoLMe0EKyd3XtCtxzTu+yc87YhxoILse
p4PXaq5e3IvPr7JYfefME1D/DxsAWW2IywVYbxreFJIkZKcuJkUSZeJ/tUyHCQX9
/wyHCFy3pVdj1SnwIBeSoDFzlBaXjyqGsv5tawZIVrmWxIErP708C2F3Bhl4WHxS
PDOCDLKbwWIgP4nnPoEtb6A8IDNZpyTadhWtzRA3cIbX6o9VndaFl+9eJaKxDLgS
ah7ZIX9ehNeLe4ytMPpCazohJ1/v1l3DDlQdeztlsPuhNBDxRU/dUHSez2DGW8QZ
YVciXl9TqhAucL2+46NXV6bnrFYKwl/WjZhf6Bc3RVQBBjbqyPBriZubje+G94xI
66MQ3okKThTxWVM9u06ymkAo96cSW6Krz7I7vdJrBArM6ni7lAFF9u2Muvx9ax0J
hwIh7tMiavMrFqXF58FbOilf/X2CoVRlkBnbIylTdQ8OR8b2vBn0vAYGqbnpWAop
8sCOiC0RiwqXAUujqGUPlEwQ9RnLf+XVvDYk20XWqmFx3oT7f/ffQo2XjKp1r+fW
m/ReRS+94kbUgNAlLVICOK8sFV5I+GZxrjzItXpwc9V8hAFDti/OfR6T866QiS1z
5zx9g28hp3wUD+mOe+CkNaaUr2j/ndlkuYfO6I71hdvp7UoTVegUwigRfzM5lWuN
imiU1j+fowrY1IlCYYGC5VKkr6Q+FYQgN7rO4y+iiNM3QlNQ4J4SlHvhx1kpo7EA
DV+HtVZPqC0Vvldv8QCzGhoICbrV5LksaJ6NNNeNHJVzK4144bSB1BUCIngaxs0i
4N/lMoHKx0d6k7+Qa5b4HqeRV+gOY+0zBSBYAbXNNppzBI7P8SmWhIEXyuyR0UPK
dPvJ9wJ3vshwshPfxp+ykNawrAqaEuBINsxo8evOmpqE76dECH/xeeafmtYc8tkT
zACfaps1t5e5FAQ29bWaJvV8OhrsVR5bqSS8h2WJxR8l9EIQATS0/yaVwFx6n8Ef
iLtp74/2MFfuH/ewipo3KObmfVIzDE9B8AqRuMhDrd5AuZ0YYtLGM/UUenmeQ8BR
9xCXZbplf/CE6mT9XhSSD2Tyvf6gaxjs2eq5+xt61tPPpTYNX/2+2hXfP+0H+lGe
w4LRq/PXXGAtiOHBT3MLae5VuUeYlXmB9WL23QOrgzraSDqoF2hpq2dGfmaC4HhD
pAVIN5bZU+84SXnh1tKH0CjQ3fTlUUWHFNJmI9Fg3Wsuak+1GJVdTkz9zmQH6GMm
Fos2RyAd896WHKOltBMtiW6wm3hEtLcmCf/aFY/VOw4+KO5zvZKw1wv6KTe2tSG4
7I794SBXw4idj1fbCMxuAowkipIu/FaB8zPxsnLqbCmZu3tYz68bE7ip2SXVNdEj
RF9EatTZTsV0hXdVyGiFxC5LdZYRja/o3R5Fp+fORrhcFmm1K7GFJEwiRb03h58u
bfjpg8HkF8qIRZJv/R7Z7b92/idnskPRYYoPR8xQjc/N62jXoGdF9i0uvWP8yrvH
qBgHt9mvLyfBv1KRhtEHaBjYDzgPk08Cfl8nolieV8nDBUlXa8LQl5Qc/cU6hmZj
zsNpQD1J15AmQe7byQBFKbLdToOZqdtKwovvapXcfT6YsAXScXRhJlhMpilLMj7D
6t1oddF/ZEiDrTOFHA9/If4IAtE13h1movyTkqAuWhbHzLBQQeGxuud3/67Yi2Yu
05G5M11XDMh0OgQPJCX7IfQ4ry/7qOboDquVlCBDCkFVRRiEAqKHL2+1orDIuF8P
NVGpfXWKo59qi2gghfEky7f5drBZ/XnXER5Iiso93wNaZJlhUhVfmehhtE7YCGMz
9Vmf4jPr2eG1AhI0KhBJ587HEFdYOr9XLEL2ouJ3MtGSLLEhDfl8QbCC6EKf2bAq
wrZf8hZOz6+r7Co4vGesTiJGmWn5136b8NYqHQ4MUVkl+XWAmfqQHvGW7mPwy6Z1
scLBngBa51WdCfCmsEMncHGWXHsIqhwryuriGy0o0p8dou7nunH3yMlN1j5ZoHYb
pNhousmRdlQDrrUQQICSnDZl63DWZgscJ/zqpfsWdb4n1N/7WPP4TdIrS+M5vmT3
K5lRBrKccW2C5KH+qqULHwHONhUBMZidQhCXPIWfT14xeLRSiR3i4/JJepNjCL9D
Q91oL/WhVjgTWWSLdHhfcy+uoY1A5MCr0+0+VfS7vEdWqr+QhkcX/r4zaxiw23vZ
sgfI/oCRXNwlh6kqX30McKBIgLIaAtgzVhUUCm01KkhcIhiEkTOhlsewmk54Xtvs
K14ZxHEsJ3eHt+frAVg6/9+Ix0MfbakAaX2vjBXLRPltXoJylVgmGux1JpHNxj+k
zDOKyM8ehbOrwNdPvyWtPuVGPkqZwkeOWItF8/uJ5M932R4r8JOra3rfuDHbRYMD
nQZrsYr6GskXAfzAvbHWPss9CuM9m+vEdFKvZFgLEIBxL7BoFYyPGJcYGQIuJqf6
loVjmjYlcf9qdiQ5GCqf5CVKHUWreCo2zMQLszuK3phGyd+T8gHkEuya+SiJKvYO
oz5MLu13ZXxCpxNzyLhhXu1W0V2fgeXHPhY5NI/OH28c6DNQ1774+uJTfjzttoUS
IKzi9MrefI9hLVqjkGvkqW7rGcpV+1mzow80HvXJR2nbiHfQp+u20yyYGLh2HaLv
7p2nDIWDNNSjy03Yw6gNDVQYNV2U59doO/GXjrS9GNQp4Bd0s5mvimEAQ76Pm2b/
yn8dtNKKVaZhGVqT2+RmsdKaCJ++KT2AznrQaAj+tZ1acgixa9eSixC/pY3QA7XS
AuXhGoEqEUTb50z5DaZR9ApJoK3wjMUkhu5/8JKDzH7U350/Zw1sa+QE5yEbPNN7
XEWgkk2Of2+YbcTLvV4S4bUzNkYHQcpoF43xc0wiVx5M8J0KN3Pg4CLP3DmvGRZI
C6imDmDUnIPgxpAzgNhC8rE8mzC2og806KKxSsbw/ncl/eFBPNRgc9wbPbde3HP+
XJ2i6N4niFJzg8yg56AHu8ijs2N91NB4SiL0vjwH2ILAowCNwt5Qr7qsOQQVoZaH
R0fXg5WccNww4zDeaKrTBRf5D83StYjzI6FlU2GEZPHu2kl/MuhaTZlIKI8OJkJx
XO5caKh8lGliiL4bb9fp+Z2mt/mYw3v7kYeI91SBICsLAYwMTht5fDWfk0VXb7pD
b7T0X/Q+6dyqb6csRI49qbxQk3FJoV4MnqIkCdpUwqMn3Otv79ur8TmCy4Wsz59+
tu2wmL5qQHPjxnyZ7mQP6BhuQ/XHSzOkGbsAoB0zrnR2yWbV8O+cOGeQEIF4WacR
ibiLjIJZwRF4yg76ZbntqMpplx6rEdwr8boMneGeBa4j1PyhVx9Vei+DsObyI8PO
UKiAeXq+8ysJdKl2mOV4Mx8CgV82PCNM9BTQPBgQWsG6nE2g33F5B72PkR4R4ybv
d4ded1dMMAIhIeT7znRLqxku6HQOXGHCRaD4LSrmCCy/Ygh4N+pNyIvCpQTKW3+G
tVum+da78AicaKcMdzcIm0M/3nCaFpqTdQcr8Om88NJJiSFEXcM29qhA0/z4R4kb
0tB7EIzC2xn2iqbp4DR1YYaSfsFL4mh+NA3+YlJofysC7aQRKFevK1pHhq2cyILj
w0jgqwkPSctlmPj8p6DlqycVQ1cHoGP9SAGATgHtIu7IeFQhiJk8tWYT3CmVBYlr
aXo4+L/2IsI8g4wjrxcTIWNkkRvVNOBkcR4Mu+uS7WCmD5fk+EnGCrVNPvzdcegZ
bGs8C9GuPzNLzTAFnDfoBQf4wpSZiXajGJCmtp2UOSvSED75RnOruHErHB6uU7Rf
fydgenv3eVGyB63infPNM6m5hcDyN4XRnUjyzvQF8tdd3/Lc5/o+ov7YgPfk/OlA
LRLaO32gCf0bv2H+w8L85FLqKtZ1t4UriOGOXdk6eI1KR3ZA06P1PYJF35xEiv5v
a3Vdfxrd7t2fykX44OyYdiv6hipZ0XhjgrrYM0Ij+0TwCtsAoK8vAPZbBZAKP+Wy
5KaO6qrFyaaf3bDeMvf3BQbJ6doSWzcgCjRy7Fk90BYjqHmp388aK9Rxpl7xtGgd
KoHS33s+9CrnefAdzoJH/HkNqVtFnzF8aoNkMymaEk9NpqrIaFdj+ExYdBWrE3Rl
QQjFlqRtButZor2ibyDgG9YzQmxtH/OOCmF3dZAxUNABYQrgbz2m/i1VRAOTMndd
aDqHy3/ix6tKj0vyRb4DrI6x480s8j9MB6JbAaTTv4gaQoSEgbPzTik7apF1cYgf
IW0DaVcbVNi9QIXeb9JMW/eDsKnDP6TAuEcOjV0RmIVXFhvjkS3FiVgc6ID6E1PB
2SV3RBGEpMag3eih/SObEg5TP0HlzcFx16i1kGlQceiWWyIrqmSXjVsd7hr6FvOx
+bAZDdbAlW2OLLKpYiZR2EYgpYbbfF3q/ORD8HplBmEmB9NZBXHIpWf75nY85vsB
3GsQLYKEpWS6Pks7Guk2rF9BZJzcyjtsTSXg7iSdGYfQobuJeybJE4RbTMpOZIIh
wj+bE0ZMQwmyuoFM4t1dJrLFWsTYlXE7vEsW+hZvvewr6EkVQjWYDPTuQ5nA/0ES
mV1lPiVsESWdnPBVxcspknL2LlKMTkdJpukRAzH1Ken/QF8tPQHN3ehQCZd3P9Wk
EEffseEorI9px1OKo+2FW9Ed4zjNJonlglL6ML6UYhGcyFaIopXNR21UToc9mZ7h
gaOZcBor3Z7sevaO8vRPSNfTA5hCZwt6lCXdlpFf1vFMngOBlelzJdaW8xcETbvq
m3d9Cy80zcI15/2Nw/Gc45+6STysjEbQkZfBIUL4Zv/lVLdbSRYLp5jMuOwp9RIQ
N35ffcCbRvaTNSbhTp6SyBXNr8UZRXuc5eqoHmcBedptqxO7maKTgzEqRAJs3MnS
hPnqYF610uLa5vOVteszQuG0h9mpoxBs+JUm8rWE8HYKHyarkDPZfNdT1mZxZg3G
IHSFg8Li1hJI/hhg9PyWovYrBqPm+Yy990GTf9NjYnsYjrEI5xvgUngOqZGuu49E
jTTiY01VB6Qs402RYv5m7E/9To7KrCPf83IJFLdu011uHSN57Xhkk3cEh9DYKg4X
Mb/pI0wIN4Gn3yW7ca7EzCZSmwo8kVrG7Xo4wDaH2Fypmq/1+j0MaoiRt0kdny8f
V0ajq8+atjsrQygMkvtkEUhh3gXjNVNzGHNcalqL+g69SsdbWGQ9yCYdz5LDSf9c
/R3Bu3Ze2z4ZDshlYoCPe6NrRJYJUo6b73odogXD6AfigBZIXSdEZchTWCCR+MZf
RwO1kVwLEBOSMXyS2E/tiy1tvx7kLn5iUdY8L8LFtorgCTg/ClIvuKHzxOOdpemO
3cEBoPXx1ajQ9A9p6REQzqYuEYZeVE/5ArvVlvt0qlm+w61ETgLKwpwNcl7aJo03
hlpaJiksoyAto4+OMwco1sn2jhMYOAH5pDtXm3GWuYWYojqwPTGrhAz+xvzQzeSA
5MXCSZ5aY7DM2pTLHdRpCjTVk6OwwarNKE5HkBEH5rA1rAuWT497pHNrssYidQCv
88iG0UESUK5IRcF8Ca8ihz1s91M/wDVQXkxj1Zkh31M4XwEgFsB60nKLvrkfm4XZ
GS/xyZfl1GrGLhMpy0ahu37FMQu9BU4CO2j8SI5sLv+SChRdwxAJaQn5Bzafg30F
1RaGAbFXNyELD+l78P1FSSR8bFhk0qaVxaw10drL0JFRVtpkolNaaoY6wn/C9d8g
Up2wfc/e/uZxOF2ZuCBBvK5+sTyImipzvy5+NwIWEE98iuoC6l1Q3p4YdTGbX8ir
7n0L2ib71VsjnwsZmM0xsFkwGPwXkJvAXe4FDLQXyuhwNz2+ao8YVdaEqm32pAmW
a//uPQRVzCytDGO85IfvnpPAPI5Veyr/jmbdxKb5JUcVpUC3Sy0yRI/IszaF1cJX
e0y8+BLf8noMt5l9N7N3tY9iy93sEBmi9DlRofmGt3lHUs8UC45jpYMZJeC9dgFx
iySxgjUa5XzXxyDnkouPe9uC54mC9FMCU1SKCEqYPbS6AcpVki03F97h8YmFwHoZ
AG4zOdF8g1CNAX+4DXY6KCdLzcbv4uhltF7AgyZcaj3EnTmhAGQaSywOpBditPMb
ChI+MBHj54kQXs93vMxRKY9t/4EO3DiX4ZbawMfs4x6PkHc6RpWvC/pRrlmar1ky
IXLGnc3N7g9ozpSbTnpFrUROd9dFRFgNtJV4lYClqBc8uKuWjkDlQTg/qXkYpw37
pfzMbzTwzscB3s+atwfmaTT1/G8tjoOz3QbOBcTL1Y0JNbkzMyiWbfWfUuQtMyH0
LKKRe7WTV02VZG+yTT132jvRWzQLlAy6L+seDuI8Ih7nUIHePuvOdcCHoyCKYpOf
Pe0lYYVrB2uOEZ0bEJ72colBwiNNsxshCwkwSe++/w3x2PcZxghJcUrbOQtIiwLb
NPH9fWVnFGv7RMsDHogIgJht9zEKLhMmDZVCNR2VBiij71koTwQqvYFUdWVMwVyT
Xl6gZDuizJgqS0EMldUartIY3QatEqcz/mNCRHppsGY0trWxIf8m+I7vn+6zRw+X
mDWnc4F48jInwJB1dm0QAx7WRUt7bM781CFWoo/utKTVq+gKsazFOIfIjxOOoXZT
nGhW5LGR1N60HwVVlrVsEj3C0zrf8FSKJKjD5o6qOeZu5JPLrwvMrdB2OuJKz+99
oO+uXZFHkeQeySTZSiK+vrngG9EzRDr3K1/UnYH6c0xVT14KmqOvaA+boNIMAMqr
/4uzbk0/2lxhiSd3AdNr9ZyLZHLkRScniLuoN1c4Zbi6ma04YX3aMRLOvGpshEGH
tb2xzo/U9D0FEgkSIxLFyZVQHluen8Zowzzvyofvpi6ODKVYsqJB4ORAIFoc+BX4
jRKSISyNf5Vk+DbaRK/aDZJ9ICkJ/UxS19uUF6nBUdzKUXKMSaUwc2WDE3xZKcjQ
gjoV83ANPO44ln4SXvtH0V0mZGyU2yMqwoaQmhhkEJsEk4v9enFcfBQZTMwgXwQJ
ko0f2+yPcN54JFPTZzH1r/wFr9xCaoqx7tGTRgcqP5AzOp5Mgom8DLYfF9maorRl
WeZb2CHcaWlPurjFyYTbKeZ+4j+vEZO02vScDlrUdsiobUULpmNcOe0Akt1833ZE
MjR0ca7+i/y5R8PE7vmRB7q0Xju4E8buMeMKlDhZ6h9a61z655LQ7TVd/DU+kG1p
+NKRgtYx9gP9kFFNBZbxPwqHGvBoNdlvKC20/vibfaQGmw0QxM9O2X/Z86aRwjEf
Hw+Q3S09ocsISgs9Kyzt0WAkdlml6tos620pvGAlmJjtZvwLHRk1HKOJY+WnLN1m
Cfnb9uT/zMS3AEy6941pbaZJzonA8vN60aRXoNawfdcLhu/PU/50Mk/m4XDrssus
V5NfIwrwYBBAN5bpY2lE2bHrlBHYUSk6Zq9wIzn8rkaYf6tuDLFhebey1FPsWORf
/UMLrbLZCBcqoNVEzPXwbENYEfE4Pj3a42WRlL9l2iryyWAr9U0doSjoddCojOFN
7vsZ1SWU25VYumbkQwEnYdsZwsems7osn8pf1sBF+g4OQ5Ha2tJqMXUffWnJdHl8
t7y6cd3hsSs65fiW687Aev3eT8gCSUaxa8BbOEFeMEUFMedf/W1OvCDC49X88dVA
yMv5w2Sx97j+Hkt+hNIPkkwoUbn5NWFscMJwcaUHPncUMCZVv7WIFnnSOrrsHGvC
lB4KLZvSQfgF1bd6Lhx/Cq210UdQn9rSiKXOJGUEBCkNu9NgsS+5UPlibfHo86no
vuGILiA7pthQGk0BnDfwtcpStfgQnJ6lhNW/CW+Ft0JVIHYzy9biemCBt9tqtt80
7APfQaQ5GI1/SlfTxOwXotwcPoajrgU273l0En6uG48/yb0KI0clq/k8Y2eFCaJ3
CIP9WZdD7mG4tjTd49I8CjUovJKQv9THc2dQwGRHmbDeiVynANFBT7FZW1qYObpk
GH9gMwHBusjs7F+LqHvddlYYnu5rv971eJwRn72MgTK5dtjUktg07rZx28488j7P
KbL1coLDupWMjfE09907vlhGvER+7Cc+gQFDTF7JaL8sRHAhFvdY9/mPwn+Fj4jz
rdIMyrW6er1+g+EYGoY1B0A46qOeeCmjhxiPLxViWI0z9T89AuEPruBgPvO7HfbQ
ROWOyepazXIvXM1+TwIX5hKc2VlvtYmwbMjO8RIgtdYfDILGihJetmNkxHbeU9FF
Xg5kkkpiz7Yp3eqSz5V5favF+jsYNYHupC+jWX4RWae2caxs6l2M40gs5gaxRVVr
shZj40mvQmzFBG6mZ/UvnNfLfp7uOoco0Clo8AWOxR3LfKwFZCD5ywIBGqkIgqiP
YNB1T0FW9y2km2q3nnB+ToiZrfOyZEvUtS2Dqp9b1DjzmlUKq2AGk0TYpJMBFql2
TU8IFQu6568+viC5eIC+XWaJJuzavCctXxnZv7YlhBu4maC757x0WtVJrkGcn5zV
YbnQkGWA8Z1ZNI/m5sc9qqFnVhWv64WMiIHcdEddEDC+wKtK/Tz6f03nUD07+9sD
ioxteexBaZ+xTfsVh10XfAupxjeshAix1I1mXr2bjh9W3KCFhuLNy+08sofy5ZXD
svk+q93X3SyYqg3Kl4qByksOWoZbk36jtOa8jkhZaBQ95nfouEh24LqWMkh9DqnG
Zmo03RnCvTczRk4FL7q/V6de4OMhHwctEv6+/7zzJ7FCZJLZfAO1Im3AMmVp7wq4
o6qejfYYnDo2YeTEKKOG3prjuX4JHqkI6qjgUWW4vdtIjjwh3Xrj3lP1tUQDm1mv
bOw7pL9Bnha/2st5jrgIDThdTSosnRoIhNYtCi0Iu0jy/J0C1FEeE0XblFa6DZxS
n6FHhnsv6LpLxheRA0Hi81Ayq78K1PJM3wh+ROMdCkd/7owqcqvIk4hsXb/ToFXA
KYT6B0Y2go22R3iBAHOH2Npw3htKdlUHqJZgXYXqijbyR0EiWOt1Ie74p0kkN9Xi
FK0KqS7KTL5A1FEPB1b5QvVURr+j4x/jaIQcBeA11wGnfmS7bKl4hvvw3CCwLTpJ
EWd9oZuThqBuCrP5R+u/8npCkZXPLHuw907j6RABXEXGUISOx4nvbzYM3QbIymPF
thjF9XByFbPXw6ITlel3GkaQr97dq5v/zKmF88jM03aaRREs2VwSigYIRIlWNfjV
Cv7t9zC6BMsk5YApdNvwXUDFRAHy7UnYwF4JcVMOXNhcXwKcXY4rTJC1gE+MVkd6
loehxvQGSAFLKGZG56hiRSA9FtZpU3AP6WjauycWfjbENa9OhjddeoV+JkYUTfyv
aROXV0W4dkhMsGMNvbjaUJZnTCP859GucHPhMpjPGOr7EyM99wWspDbNqSfNg2iW
QI5HnlDDtzT2feWsEUOCn9etz6oxqFxvk8nvrJIppT/wu1MgbFpqPKGBSvKjf3XU
TbrbCOJgY0+t2vHupidDxSbu6UWpeHX+A10b8F6zgv1NT21uaApBbcK15Kj/NcHO
AxJO16aQtr+CGEcanpzIZjvoV9Wl0a+0WoborAE1k70KLrcE84obo87Xw54Ir+zM
CT3qOrvl1eGSL1HwQ3eoS1cX5G6pCOe29A1jmm2x2o5snp+/Jc95qeIkbfXLQVSQ
oBiC8ViRaKh6ay9ZxV4b51QzubK1kR/NbNognd4epqFDlkHdgyTMlN437TAORFTW
XnIhhMmhuvKY7pq1to8P+vm6TV/O7GT252wJ452tes2cSxDCQMHYB0OAH4ZTsjKB
b7S69Z+K1PwTNbPBw965TWbowyNwUr/pwPd+BX8GrBoHsq4VbkEvb/8BoQ9ZyFOz
JluMdOhJvftMeyrJfJhZ4/WOtcASrVgHqqOhsrHRMIHwVdlcuT7TiCx01HnxCkds
S9YD1HPuQSCMd/GoE/ud5I9JvwIchD8mQDbfnIjVX2oErYwQ17e9mDpVZheq/zEa
Wrekk/AAw4w7Agja69bzaoCV5QfTG1ODkDh5EEP3dhAgfiPnOiQMLyvZMfxW0PWp
C0jVXLnWelDnIuGrkIh6MqEz+n/D7rymqwvsFCJnKDcIa9I30LiEtzqlZU03nhwN
Oxdgfk3P4z6mXI3ATpgEwBijFebYFf1lOOsxkQUFUeFqp7pskseSTeGmfdGoc93p
4T2/3KuQgDY8w26jkg3/E91aOI5yz7DQtYRhyqCcU4nRnMrJy+PFPMn7oNPDML1y
MHYMBYS268tpUxDLR8q4n8jOqGAU2Y0rEbKsaHYHmVT1lXnLg6VgCAXZEZ2hJarS
BNpyIKSFc6aYUqxLX/EkpsCv1uTxnGizvOkyeyzvHG8VrAloajBoReVEIBxhBPj/
98pjHzp+WTLuWfItneHTpvnGdGLg6ofG5p1QgJ88UV0oYOqNkSJtjuQni4ZS8o8F
zHtBePCJu8NwIn0E8n2YhvshCaocBTMAyrsXuSg7z+FRpMVfzP0mnLVubYgdyhDn
xbtAtSqhySU0ExrGkh9sacD8MPQG3+JKb7yp0Qwh0YD6SRX8J9I3i3dvqFmVWsKi
gY27bLD1IYIosO/6h03cTZcU35AnaSVWF/3e3N95596DjLXD30l9dl55QPtICmuy
8azpWPdyI/91mz/GWybYj6/p9GIYWPmoJu8sp4/fEfh8jLNfOxeG1BCNuiUiCu0i
UEfEDMvZZeWAtZazGTltZHRk/44ABHeiiiaDCMGhUGbm4TsCxTiFPEVPgaewsDTs
epO53Aqvvp9CKK3AWbPaqzO5VlBcmP60nWn65ughiUz7JgxyvYaQhEiMjLClHtDG
2KxaBN2ajoRN1xRgBoAW71K/tAgvNd1OD5SA6x28uIotwwE+3LEMH+qmZzbvZTqh
vtv9s4qkbjqT4Yg85LGjeGAJBAyChKmv20k3vQ7TvoT5CdtDMkABxxtGVUvXnZLq
YmfIrTQM6Hy/QjJvSfFsVmoaCnMQrNb40CAAzhQoeJXZ7i+aORgpqrGRQ/WRX7BU
M/QL+JQnaJYHEbkfL/PMszyB+UlgXtApe62ap+s4WN2hvUsk98yHiBMgMUwULqDy
J2/SuqHZh5555VYOO8ivTy6cYI+VnZom1pIJYeJrVww/E7/PBpwBnT5R+yCGPPBB
yQ1ZtVt9de2vPb5sjBulfT6xdWOpKKipxwq+fJFfnaD2GvWa89si7VKIZYNgJYeA
lQH5iWGkc9DKUty+aSyPTd6zyjSn6EwkPNNozoS59tAkCuSZQrBeMPwJwTHM3hwH
76fMeOWVV7PIdbhqI++Vv/+o56CZHIiw71/gx4qFskyeSVPhysziJF8jEx3w9iwK
yu2xVUYgzZfVT/0ds7/rHxy3+k7ay45yWqut6yzPO9SzKdJP2k/ruH3jHsr6rry2
4KC9PMRGr1lsDwfCqGqMa6K6CMKDlZv/9Haj5zLsZK1WgZ5HeI3dGQuisdCY173R
JjgNstSJRFVoOIvJTlSyUc1OD7AwivROCrm46wingrDtUPzsLirZDACYc+VN1VeS
SJSz0VhdNN1GcGumCqNFFaa4AvW8Cd5Jl8xsvjMzfRdPdE/EJ6X4vEnGvE19oeh9
A/wnrCVPvNRhfKzrkzBPOGh9JYZ1ojLmv6rRrTlMQXSrNzbcGA/e3iHPnwYNmYJ4
lv8/fhcQ+dCNuBQi62nOiYinVBF252IvJ2fhAdowCAzV4YreDpO6s7lTFX4P+aaq
oGlIEcnggzPc0nYS5RKrR/TxI1gkJDpBEf89hXVUwFNHcUgzO9r1iutma9tl3cUJ
Garm+d/99QEnvdYUrlBTWZMIwwSD5lWQKL4GE/pv1CTqboGAB2LwaH+TBnz1pLAe
8xp1FaWJGNczeCmpJHgr1SMGbrKHhWrVj3c/uGFHp4chXv/BHPHPO6Xk9I/yeb/i
ygy5i7qCRFFq0KWNiqDNC3CAjemtBrGMIuONbVFWEHd5SbASIcWnS+COXS9V6T8R
cpJIgW19EWGwGjjAJ28t/5jXNCygsGLvNUmnM3lr/TMeZNnwWMiCuN4NTQX7wfr3
jkJfDKCLXAiZpj8RNZMeByrj4zy5lfZ2KxgWWHl7NzJnRlL115mb5Bq3E8R8FQ5f
xnk1xjmME0mwP5V8g5KTSJGP53DmUbzDFby9kBLY+WEs3KSuF7KbVuIETyO04wRb
pyX3lRTJ8dE+/eyVWsmuZnJCjG8RMEsR5Vh3xPhpF8qFd0Na3xt9+9ag6ea8YC67
25YJYkQcs/6FkQrahb6liY/Sqx42eKWZi+PDBIXBGn8Np8mmK+KILRuPYdKDH70+
bZNn+oWoJFHAPUz09dSGNXV2+Sa8zWj3JQt9Difi7+H8/06v49zKHf4obl8VrToM
eNXgzYahiOPMsRRJ0CTw0/Th7zeJ24WQ3gzfmvELZz29XJwOZru/c29mZA1Wrm5P
qYt4dPCUQ3rWOUGwpyVqdeEpeNlSD8rTPJI4RaEynP4KuXjDeYGIic5o1XQwn2ah
8eSp77QnLfxwcqJ2tMqFc56+t/TAr40XEVnrOA3n/NBoM/iYLApF9Tw1WORCkI+w
mPErWeX68/KF5grHhkAa2JWpV4Be1pobNi99duwMUxzU+h1dJ361aAPFNWqtl6/g
YjOAlyMVVUunHH8CDtH6IehWvO8aDZPaGIJQrNL5eKqXHApugZ/880aWHygHqZhX
tcHVrbctYZqecmfMQMb6//0HxlDohpuXzr+El+20iqId22zVjlFsoBvfqCZHHD6i
Mi1RSdC1PzhHQA6GOgG9lkvchK4AVQRsG+BXNNdkMw0pv7suveAS2LbWobkCDiGu
RNI/BsxTAF0fv3j+aynzm2UU7JnC4vAMq3neZAVfvIhncezhb6O5i++Y0mNVjV2u
W8Jm4qjQH2ZNLxFp7xJI9sMuuJ8LPO+gSS+vLB8sNpp68OcRSvRwdLNu0usKlld6
NAgu1lO/uj3DkOQQtXdgmyXEmC2lgecsZkHiqPYBJsxxJ6aSof9oHrpFEiJuZQJL
Kdr5tIbFuWyHozG0fZ8Fy6dhJmPeb5quZzQx1M6kYVYA98ASYQ1RlkspLRfZr2ZD
GVCPtg9C+ycwSsz4Ndmas8HsUl5dTI/Tz7FyTabMdqCz6QrMUoaehTiqo7jgKHcF
gUTJXiLpkWDJpUvaG5lOy52hkhClulMAZnlU+dYg3CNMwuFbFWGdewiuarwUjB6P
+NABiZzOhezaNA8c/epgaC55uEyFEQQud3pl0M8AEy1eRdeYcjAQCvKz6B+2WYSU
tJmAoZkBMrxlVg/OQz120emSv23/G+DXpQcPHbXI39TmrJ9qVyp2qESo0rhrWejd
viPZ6YTvmqqj/LqtTnCDaLzcC4V1sM76RU+/M07Rui4gtWyOEyNjhTbovRCv0rLR
B90TmCGAUBRiersGzuEZoyJCxL4ssaWt4GdkBcph12f0LNjLycaZCi2EhQ34NBhX
d1xdL/GknLe20y5OnxiZT9q59Zo6KXHci2Cg0sRujavaMPGl8i3IE4KqNAZ/ChQO
5a2uv8UXG6mdhCYt2Zpn199UEAvGq69V1D8KesG+xssNSyoR61uvq5bk9Iy6Y2Lb
dH07e/od7x9kIk4j8Vn3609b0JBzBqiPfO9pWnp9bnCFbVJtQnH/G5TvOqSSvu2e
Veo2rjnDO8XiF9k2/a85vUUCMy8iVlrfwIgS0uUbKjRDcYjuwIngESlGeXxIS93r
5FRH6QHKE9MHhaRAEipsjn2bJbhgxxmK4rl8vNvv418V10O/i1qnrIDap/PADwkU
AnCnawRtHkJvBxqTpNfkfPKQsNPoS9x/k14BGI0Hq7lZpCFl8vZtdj9EO1wjve92
d9lHvxG5bPe7UYdMzP9tCSz1zvZIQQc0GWTf5HYPlE8FIntV1mCbN032SqlN/pqI
CNpV1Jyaef42PJU4waUkyHOZJ63cYph18Qwis/jD2WEaExBNKzbfHhl2VCAAzyu/
q8vDaR4KdXeDbOJ3eqdZ+2zQkU3dS/kwv9yYB17qPSC8gwtnv3tMwPgLoEd9gUzG
2UZCaM0hu17cuT1qL890zmIo0TII3k5KVrblOCNrWg0YNSD8VvuL5o57dqlvEjWA
kv6CkXKHQtAMdEtwNFx8qXKEpSt+2Q17ACAEUxNwjqPN4YtogJ25jmXe6Cj2XPpW
0aQEh/YXlR/1Kf39NFZJl4RUYWgpalCwCGrqrEpG+1Eiz1NfI7TAWqnbpRcc81pE
e9byL/nqTTTwE0GRo4gqQ+lIauInYRhQaPQrZ4ffuFdfeIip1FYmaF4u40+xXg2E
96lw2HuHZf/87dUpA2b8mXbA1H84mu/fS6X61Pv2PsTbrsVLVPvjw+VJTvZqvwC+
7UxvuXb3utX1JmkWDma/zybvHU52G3S0DI9b/26Wd+MG4TL2u7FKLjROXIm12SOB
ZqE9rYjrcw4m3jswnimPa/jzH3ldHsLaB5yLNhrQVJkBQw8LoZ1PuHyE4L1sxqUc
fVGKmb9g3+pur3pVRlsr5y/hCISgG3rchA36vK9cxOKmJ4bfiRbPOm4x6fjZDcl4
6XIqcprxe5FVZ78rmBpoQbFZRGUaKygAdDir38G9rURKVhi0nhgmgmtd1g/pyg2M
YULz/Wbnjke0OjZDs7esNtbbFmX6pJOBMf3sTigdqELt/6gdug3wk1a2Jzy9gVGd
VJHkOe+4CN+2ORqowCuTtyhkhjyG5wI6WSa+LKJYy0piQ3qyjgBiO/lMnddK4KuL
xIFq0+o4S2U1NMjcqac2gfrbdTyVZtIROC7MtfgtjWOLWLFMElfDwKSln3rCdzGH
9AI6YdgGVxLGjxSjRvoK7nxuYHSzUDTjAFmjGlslwfCQQL3QAr1lac7yfd30egWR
tR6F+tflkTVL+jwkexSzjqtGfHE9fu6N/wEw2UNxSHUgdGifOPuB7mdpnP6eW758
OyHJxpg+E/jAFFNTuNaT9vlZkFYbhZ/1vMJ3JjGa1RVZYR7U4QFSkMDGnyRm0sVy
26yQzrKiKvsJc5SnIVA4Y8hT2iqWy+5Eqyr7kUpoePM5wmOcyjQzQTVhWNFfUXcq
9FxnhG0CAyP7Uyt8VH1treC1xOB0NNgeUba07dXzMTWS3rx/CLsPNDRTtb7bRDyu
0aWJKH+4jWhyKXqIxsUMK6nNZzDH4oJ82Nr9furzjL+V9CQU3Y5W6yLVRJgDzzhM
LDh/7lB5KFpk+mzusCEJdDLLdJEhiUiEcc0VCwbPTptlx/TLLqv3tAYqZO0fCchA
Hr7yr5R44VbffSqG7TBlpcl1p1yaSbVm7nTw+xt0dwoqutKd8hlosEPXe9Th83Nn
CNF+4P9EpXdFzTQnzaN04ZQLkWUW4oF2i3+fOM72AQ6ICG8V+mqy33tMLemsXIAU
ORLz959sfM07H9m/zvteTxr+f/hvUrRcjfooolXz7p+B7JD1bzX9QZtJcoYogPhf
WsfGOuOsaHG7m+YSORcCSwIe9aD8BEZr2GLqHKEEiCrKKQlV3DExa/Uo0bU11zAL
6fVVCgxArOreKvYohaibxWkspq2GjqnjDnmZeBH+Qb+/U99p+SeLEgrq8h8vdHGt
+E0/Mj7BqB8+EnsTfHsZPGZhmunLJaLJMH1IfZ2x3Oce3Ud1dI5P7kP9DIHGqlD8
X3TRxJmxOQvT3WJJQE6zTfDJnNyTqFRFtXDQ6xGkk5sMIww6dcM8YCeXwWUqvJUz
2QhgVZyVvLH0UpMnj8tPI06yR3szn0oWSyLHrlk3BvifC6SRO2fzKy+ukXvGCpcd
9qnPfFgFRq3eoxEkzvOtFglU51sATjUtqcLxIVAM/pXBJjcRSti37Ei8GuDprjD1
gznRfsUvNycHVcgsP/T3yikJGvwZcRta3LDk98j3pndYXVQv6jvpKXxxKq7i3yRS
qQk+2d+JmiUXPWpgKI3uyxSU/0p8577kne3Oo5Hp9RSOKWGXZf/3luu4cQiQd2It
W27SywPBOe4y2/ZjR0kNIKFz6RPGTSMsUAECudgpbBtsE5THFv4GtR81Em4DQFGH
APYnMQmv8WJ8Nq5s3XHbpj/83ykGRTwo/IJYE4a2Mo67gLXKJoyldBb2Fz9Us+ey
KRCtIOTiWMHpTZAZc1dlSps4xoUuVYNXoLfCkJid8q2Q4fLk/ASm8cmRonWwim3r
NS1sD67LeRx195yezIrQ1LMVa/e//QR21hf+dwJR9epLRPbWLazJ2rCCNc9IY+4E
R9ACyBR+i6rFdVR1ukMAsJZkI3bKHoW0wYBZSdgk/Dk19av2QUi3PZ4Eh+HSaXVb
WvyU0vJ6vt5xTka3fluKkLvRL6shjLwPymmvw9NblD9U9svGC3ceWOpeZ/NgQbXB
V3wdw1h8vACNj7maANCtWWqPNsvdscBK3DHgwN+a/cuXuePEscxYnZixCHAbDe6L
eqmEK9AEBHD58vjvdXKt055FS3MZDnfeZKm4hq48+kNSLQij4mzWaHZ6ow3NF/D8
k6GEcko/vN6DkIUxDvQY9vuqGbaqLvlLjxEsjigY0Vk0ZMZXKiPoYBZW/544e33A
45oj2AOO2XviCczFJubCrUk8+/ffS2wTnTMqZyuVQBHZo2/HQ4h88foxtqiOcbtK
2sLpckUNye0ALn32f0Gpub8XbB1lOHkw4KccxuL9kaL5FWWI7Bg/Y8TfPD9rGotE
AoHzBgpaiWG/kRAD+bbpadtw2QjGHLdDnKK2oedSYw9xlG6uMOI1mWicuRF0kpZb
PhYL0u0wP4RrWgXgssr9O7GOahx0QPD83BshSCvMMXNHDi1H69mA9+9Uenq9XxVT
FcZJsNVJXSxRnarlGthMJ1Z2sCF5tvgMG75v5Un/umA6ZpnIh/XbnRMRIrZ7JrIv
Q6pyzdmkI5xplvE/BF/Er3yw68014VqW2tzQ2j35Nvofc+O3Yekdir300FgwPIrt
EFnLZn95Fcv/yFw3U9tzy/StFsOe0BxyzRwbdyKxE3wYjhvWkT+MomqoW8TOLfOJ
Dfb15e/sO9NNJvoNbhYCd8YqJUZZYJgevVR8leQpMTzQ68NN5ODzd/CSy48wblc4
6CTcXFPbEsnJTjR1CUzFfOAHmUFocJ+UG+OyvbRaXoWLnxmfJFeoYp+ZIBb/+RdJ
P6EpClOrQTUaHOw9GLldS3YUYi8xBZw6JOHx6fzpkO2tbp5yaO0/ad5tQXzMfxw+
ynpmKOIpPbHBzeyvp/jkrQ+wrEpVPm/hzBBuGCoY4XNBKsvWvJinWAylyHE3K53+
7UQhQE7u2S2lDkWPv+gG2toqTNh0YSDubj3ASL7HOyZdFuLaZeDnZwLclMOqXAU9
s3WO9S2hfkrFAWTGn8kzAns50idSyZHFvM8A8aYkTHaapGMoneGMw0Epy3X8V1P6
clamW2bB4v6VHlgqRUnFnd7cjc8/NheHnG/5AJ0rw7MN/cE0I85Pbod4TCRcXJPy
am4dgziAWd/rvKpqpYv2ojuHYbvqn6byLeTrUvIZBSOzVWqHKT8I8e2XWW3XvdX/
PuAMbTogdeAj2qCjVxUVEAT0/QT1wsiQ4ik3r4kZu3w7Wb1jOjBFzzZOFdpVSP0u
vQJKHRIWq0GwARXFMAwrDQA34o8SYawXCF3jYbvkOHrnYPufRSGNIKJCCDh5B4IZ
aSR5PGSRgyk92t62eTyN4S8KMELg0FDXcr3I7LwzALhb8DOAs+VqVdM91oOaJDDk
TxqKnSaj1uqsSG7B+uvgwLXhM5jl1LLZigqE8PyLzfbyM85XkUaU8yUssNSuaKaB
wHFSWkhXuXVYlQ1LcEJjHcp87cvZmLXaIpwISqHie+I3jsdhS39cPGFekpzHr3fR
z2OKewYyIXL9VzV+bR1+etaeAudmB1/4kOr6o4M8UA1JBnnI7Q7apxA8XcTo5+v7
qqSv1cE8RYEIBuBBpgVKNZmjzgnkjD2odB420xVSyVfYD7OPJmf+4ayI1iREVIqJ
D3Ak3L4VtQ+bkQQ8Zp7SROdid+0pnU04r+XdSig/Qk6l6C+BsBeOQ63wRYqhQ/Hp
9UL3Ll8HwT1oHJ/9Q25YghVSRPA2hDohVemC5bEi0izQpxvfoZWFegcG5HxKCHAl
vh2v3ktWR6zWbhnlTX0gVVZG/7elnBrZHAIiR2U4EGb4ZhOT/NFymqk3SE6eghqw
Cvv39lWQphNz+AJfyS6UZvwJ38NbYszgKZN8QWZuaoh8ONDrrXjeyFDaFMwAauab
NFQKLshpAoOUpJLLMKk8sgsy9GqnXtQbgVp+KlnP5IES2IlweB+XJihvDDMJFswz
yupPg1pKpqEe1S3Xn/DqPNobawVnYmk8nfl+G3seOayibXzZiivkkcpfgQumDCFw
x3cAzG8rTjF0A6tZ37IfzyUGpPpjtA489grHE/zzE8GgJyfdEbvuCwtrSJLTcI7V
ehKMGvkH4vjzIZlLJeofjy4//owL6bP2f6Tzikkn0r9tidp4FHwgkIWjNn1eF5v+
sgAtDfL5CMAxR3cEDZA+mMVsqkuQzXTmlgzsbLhnRNaPDTJ+PlqRGvAlcERbsyHT
SxmjGNjOmORTdNUu3yzv+YLcr5KbiK6n4z8hoK7JRm9Ft6PpNoEqiD+Ht42rSg0g
D5ANvSjiezyCLG3alps9YtNjExn6c04OKUJ33zkHwE6dppbCX3JyrdMXc6ybNA2M
qVK2KVG2E4QgLWgUn8HO5mED8YXMuByDTCrA88IeJOqgNHExgYo482TYSPmJlKQX
1ei8V1v9Q6XSkyn5354eD6eHr8AR326VvIHCJOoBbW2Y6hj1VGrwj9Y9R9kmHQMU
Cb6Nc67xu2urdXJ1qAqoQBSjIowYj3dBD67sOVKT4FjIU3ju/dTtuo276cpeR22S
CijyVB0WB7Het9HtX1KyasGC91KHAYwXDesOSLSYrlUs8zpwyCOs4vebRhtygS20
lBC18LsenrLBY1Vwi25LDSnD4u1aHPhX1CribUuDJM8m/qK1dTs52klysVNSe3pK
eVY8W2U8PgSJYMfWZRoJUMLtoNCD+c6GdElAa0pmZVi6ws28XCYjv471gc65rL5f
IPRG+OH4JbhlJShJwm6C7GUMFBdxt2Og7OyLbTekxj/1R7w1AQKED51ztZ3grpvu
A1GzlI0fXIscAI1Dxz1hU6KGql6eReJ7Os5tJ4fI0FM6KaYL/QJkAj0LeXedTxQJ
5PWg+kRCI7XmtGBWZNXVlnIW+AzJ/nn+Y6DXqyEccKleDSxj2HAMwNTG+Boh9Xcw
3wYW/NZ7i02Wii298aA4ERKbc4yTkoj/IdhoTtDuBN4C0+hR+Sx1thXVKBbeHKdT
EkVTFkurwQiOMBRiM46Iyjx88hWR+eTyHoUQUEPkfsBIb0P1CewsPvuhpvWXAJNZ
IWOzgXPOU8hee2+vcQEeArnXFvJ7K8bsfEEckAHrjV3QTzgOoGtoE7r5NgB6Isra
SB8KpGT7QapM9L+z4qtVD8wPLdzOaqEWc4XpPYBXk9rop/PJ8UALkQnzeQy0hZbj
3gRmAY23ESTUm/uCJ3AoCCDLdqvQXU/zzJNzvA5/RlcW2fzPGQMMfDzrnHiJpr5b
DN8UBLBITIBmwGFeZAmYiw8iJDIsLIS8+Wk6fXk1lI3okcRYs21kaM3VYSTzite5
Wr91IbbUY24LXTOiRVnfMxncJZtksy1ZSxAkVTUSSpr+3m2kjvR4ozxYkyBqvV8+
zhMhuXqZ/E9mMiuma3QVmoGMlQzGfSqEcBT4BygeZsxlBROKZBI28LpTlq3p0OIz
TV2zHkFxqUMSUqnaHJiyNZQ/5GYF0kmVAGoth3gzAECAwxRTX9p7rW9tMAq72NUj
hm9fXTAAWZNyaSeDWNB6vo0190VMhzvGl+rdX89cJGZJhl3sIBBYVGz2U6Q7kqSk
CgJGGGNM7xxZdHYxn5uX+WI9eM7WlC7RRQABwveB4+TD3An2TIqAKx5thC2dWMcw
y2DJh/sq2LitukfQwvs7dOPdRB/GASQZ5eNX1c8SZLDi6lOc1mhPJHE5LmEa0juc
UWSJzx4Qzxrqv6/ny9Jwi8jqC227Q1jSCumwXaREh80XBgPzHoVF9ICAYUEwr5M+
A6xJi3RkmD/+MItLwYlZV6JjxRmtKzJjgw6h7kQ9sxFfczS1Ik8wDRTRHeP3x7IH
PSbY/BrJ6lPvV16gKv1eO226onRhh5xeRsJhudTE/n6j8MXRtOZUGm9Ne0hvvwwu
6nuI57z8+r6QO3+BTU/f9RNDMz3goWqMX2GmW3GvdIfSFT+Pq4uTiTZtcIpQE12N
ZsfrKeQiGiskGgflxPUfdM3NdJl+V7f3pULi9aToKJze3hiHFHZKCuscqoA7k4jO
vz2Niero9vwNRifpJm+c0xlZ5yBQzk6z7lCu7ZpMKcyMaVSzn84jnntf8tStNVhT
qZHEgM8Ib72ofn6y2yRoTdHk0AwCaS/yD+ktxbUkGNS8wkHBaA2R/tVkk4ijSaLR
onJ9Z0gpQYX3R+cdxrgrYHdRSfIjzooT0HBySPYTRInLD3RTtEzzH2T4V7s6Ss/L
4l5zr88BukEP5seNWwHdOfJJzj4J33UWrrPBgifUX6YhbYmZXKShxQG4ndPy6dHz
DiulKMYZZybp4RdW7wRtrLNmB27akEI0m6vcNSqbyqtpX7pYP8hpkpS0hXVqjw8W
eZ56G0s1gX0I/VDFOFinwe4+0rvQpUo0rcEhke7OTkoAqKSQS+nLbg/egm+GNIJp
9e/QUipWpRJrQHhe+wPVyPD0Dv+386WLR6Aj7I7+IXX+y49PQ7i0BnI960fY4gnD
owbHDuqs7kvVbgpS1WV4d6uIp+M/QZLwyITiPEJFUyzhFLa2n/OGgIR5Rq4th8Tm
B1pUawVRo95SJ4k18A6jiTDAg+pQlJQOKjymIroqFf1y0um6N6uYrL3s1MX4d4Qq
dIMAY8tAA5HMg+0qtP9LvNMbk/PU6EthcF1VrncypSdQ6rNzpDpxBP7HH8DbAarI
clrxAj/XeHH4NP5Dfo6Sf0/GWZAw0Ef7WLTTygMF8eAMUyFowX3KnnNX4MiHl9Z6
vXdsjpR4aIGViJ+jeJkwyei7tEf75pAmX2I8iNGdBf5pXcG4OH/Q9OKRgJCycOOo
05hgBN536JYHjCdyy0ZvO49dXdOQyh3jAIHN9yAuos5imjNeszKiyirs6ae10MqE
SmFvHmyhb6/LKKru8KVWv2EcuzojSGxN1KLSG9llcESl1zhnDlaexs/z5E50A3t6
t2EYWkzLriRYeyHx5p01KAB1PVL0RCHBd3yaeZ1o4qqZ/bqesOJ3zEeHCLwFd/6T
fdkVrVw+2mvYdwguYaJYtUy2SEUR9vA8upqDhczzQeU7A9Xtq3+5WqS8hWcfKqKL
BqSNRiCAYIuk/BUtwuGIpEpuhygJQPbhUgbWo2Sxub1ryW/NcT456WsfDK2PkpB6
ch4ehuc+Nnt/tKYPSbkZUqX1StzO8SweY/SxvypKErFXIBd4I/UlFXrx+DQAVJg4
gDVEV7RVCPGJ0m9J4EPVme3AVLVt98LlZP65F0+jmZL8scm2EUHQ7Hf7D0ladAA9
KCETrLk5TqSBgMw5Djr7AMwuDz8cYxPPxakxDC+6vhRjuLCbX/ySFgSyhR/bYtJH
g9N7R2XyaKr7d8yaDsFGcimr1STzSZiflPq/5oo1WioP30INULC6vQjKgFF7CU7q
Vzyxm+ZKHnbOT+U8BtvJgeo4ITIik13jUxwf1Pja6YlhDSgZPxDOMjsLkbJ9l5yC
8/dYG7k6GOp2wurZvadhX3lEzXFRG0LKSpJla8cJQG6uVaJ2jVh2cCOmHhzsVvjd
rBkYzSdolpzGzPMaTpF6Ho/gtm0PdX4kQR1BjBw9T86f96hoiHxt5Qkfy2L9wS1z
3+KlNzY5rZn5GAATYyd2pekC7nuCe9UXPkq79okcdKO4bc/SFcUP58bWvOb9E4OE
sj82eAbbx6mKbbWz3bUMrTHN2HJl5/7y7iPOC04p1e8KZH2Lu91YWB4gF4MAmXgm
iqPcqqFxmDdRXS8fsRVE9IiGvLHmkrCsLVmaCiN+Jk3V9kRs+t5Cev6NcRZ8iUlR
/+lca19uQkvrcmR8cHQMICJNzTWu5IjjVl/jvoAQDvBgu6ZSTcz/DEWZIpiwA7Dt
QULytamOXR10AaHXd6nMW+d4M79JZkd9d4KVfkY+W2wP/yDDi/xHySZtB6a93xoH
WixhDvh1cyNHb7XpVkDxked0pn4wj6VbSTP5Q627y+15HeaJ7d8uys6zzJdwjGQa
KZ7eb3Kg3E8lq7wJ3Mq3JGca5MlrjWbYuSQafRuKdR7yygq+lrcUWPY2gsZefSMU
Hv5PAnmMcmcN2p2WW+6jjx0PCZIo07xuTG7UmO2WZMsanwJ/Ydb3qcMsGp9Zv642
EDDp7D3wmedBQaGoyZZRb4RtjiQnQ7NllaPvTlBK6Nj5re6dFiA26UASdWmAPy8d
opwIyAmDUn0zBn8TpNfz0VaB/LW5FXNQkMC8mcqMlWPk/lJAsfbOvwbGzlfl/co6
MRtSXVOjJ3EBVY6m0yYR6j9boN1czoBRtx5lpzTRYcPF1uCGcePAEWouOkgJbYpp
PJ+raS5fFa2iBfHinCMvIM13467PHR95s0BTAxPVcnzfJwWoUh/1PK7HYczmBwqb
Eo9VeC3a8F1FdIK9Qozx6FAu5LHW2wHG/OZ6mheejd+PZZ3rgRsQgqflyCJdeSxF
ZaepSOMbA1TmZwfQfKHdMM2BppADdgaiZSOncaC9L0F/jJD4iyo63FC491KOxKzi
jXO2n8MHJgs8r5maEUhS8k6KX1DNjDbohlS+I8cJhWZe1zgvj+1ufCYOJSJGLr+h
M76O/e+IFbQoyTcn5PSvEYlwT6+TYHy+M+3jdavFsGDC9Jiyv2yRql2IXngU+jLP
vA1WX7Mfn/cVk6+d3xy+AGzhjNg2Vr+aLZwibfs5SW1qYDDnu2eko41/O2a9IdMw
GOQhJMGnJPUpu/hiNikAC5bRgyCbJqhoSCEnpw9egQ2Lvp94+KBS8XZKOcorM3CF
SlcMM6pe8VLLrfrde2pH6L5/PxZtwYm8XobSiCtXicpzcjOTIg2C9XQFt7QxREIY
tlJkdGcV6X8pPMFWqLq3meeAX01XCnGOoOo8gQ7TctuENcr1m2nr427GE3b8uGkY
oY+ayZq+BSLz6AelorSR3FBaioK8gcPwHqvrh9pSMFA6flD6NQt4qFoz8bkynhf6
wQgZCjG2bS3wxCoHSVF+zvj+zYkPxJ0MoNKHRe1g34/Xb5ls/5qaMDt6HOkoDOdB
LutNhNnI72lKvLNEsaGcNV2dKqPawf+gpmM0y/kmun396xPJUv064XgrnqHHLRZY
grbT+ou2dfOf1WybAkr7B4/dxjf0ZuqvaHSsi03MV0m14TAu9s7BQCiZezgHVePP
x1dqav84khwEBgh/Rcp9hN9huSh4PGnN3nZUgvY63I7XUF+8D/Qhzxqc2MhX9MMz
Of62nk+mE6fZx/HTTcMAZp+KWZsy4gdEFRsyD7M7IzL7ZhYWTZnDHsXEDdvTjHss
A7M6q9y+2TWa7GkyRlZp/VQXxsx0k5BznTZkCM/2G0o228Mn1Pwewc0YV4SxS1N+
jnaNAqGo61JRCo8Z8nTeUGGhD+r7PQxgoeC10PlXrz+yN6jfo0wpXMH4MeqRe3ss
ESHR17HT2lzHzq+wlCEdGWQ7BNSHr5wwv6Et6WQ9YHTCxBl0eLC+49PjkuDghqW4
eT6Dygu9oSlfp63n3fERZBCKqMM1Qfm8vOZqB0mLmuPFwQ6K868fNpTgzvZWSHdW
BVStDXF7gSlzk0SobRS126NFDAWEEcIWuoiELygM/dG+aOu1ei9DNYgDVlPQyhEz
nnlRKutSYxTpL3T9wkGXB/voiC8oE92GoAMUZMxcjHrY+S4T1J+HLugPdcd11+x5
bowcRf/oNq9UxJsC/ENycXuldivIfq4l1mbWxj2vV5sKsXR3ylw1YwNUcJCyPius
EVF3Wi+SZU8EXop+nduoFeSEQjabiOYnZJaOgWeXJZ61Jwhx2ec14ePh9aP899I4
s8DphOf4WZ8WmFzakm2YG3wItniex5LDxvLHkQxGV3zOnNtVVGf56R0g0smdoxDv
jQuGXoPlYMkgHAlRKp3xE9bp0hbLdnyY9vDJ9b/ZnASyQjW9DIDUwI6EYkGyl9ms
24/gj4JnZTmKWIIeLyYjMyRlT8bSWWZNO9GVf8PwIRTP8FdXzd33RI01XigQcB2V
+i1VoMfpRo6Sk7e4Wq8ElUlOVg7Z5gb8v0qOApdnvZpniWbmizr66PNFiEVcTTlJ
rhPCOZ3/tWIDpop/epsG5KYv01ZPRn08N7z3Zz5cs+a6xqEqTHX2wZpM2dAooq2H
6fMm4xaghhOk6X83Suy9GL4JO/nPobf40zGR7+HAwcOMdamH4zb1XxP35jwyfYqN
9AOS7ttxDwsC14YVpX8+a5oUFR0xcdjKb2rdZBdJPjb3rQq3Qm54G5mMkmjkAl0D
Lli8dxHo46L/VWf9A7E1yLcUWsslp65UKHJMkevCzThHBJH0lt/cSuiy0ZEnIDM+
uFgDe3IVqAzYg8me7O8nIPLHP6yiOXxmQYgD9CIBFAn1OAuBP1KpAmySp8ae4OKD
I4/J/aHRunJmnFvNuaTFjoN2FVDbhYThWunPVh2JwvpuUpXaJ0bPws1+dKBE9SZ0
sebgs6BDNmVUHSewDqAMvxHoB4vGyT7Rw6DikOwDQBJJ1V5MjKJihkd9zqvjQ7UW
wVuIuH5MzD3DAqNQGxMF9x5AtAOZTiXfA9Jf517VD99A0zfDIcRLDjHRO9mx7ZOV
HpPpgqppRfzkkQR34U3rCLQmj/hLJo9GPG91ThqTYSbEsGa/TS0zlQCHqY9f2z6D
LoNG+zTlxAFXRvKocCP/ZsTr9Hz/rXL6Hjd7D/EFFHi6IilsiI+a5v4uP8sDFWou
09B7UtB4yI+oPUI9VEf5xNjTIJ20XSgX3lyGf9e3IV67CBMOMGYlm8pitCbrOj0d
ZxKJzVAqlcR+XO3Rh7BhZdzj7Efo7PteJNttqnLVb8QCrgUC0l8wFIoWZJjOq8b/
8kSkMV3ep9Q7RuDTIz4YtLHZAA1EwPh9l3d7uVBl851ylxPBo1bp/SHneCPA4q+X
T9/UncrMb+UiFbrI5UEKDfRlYJuA3qeyOf5lSY+IKj8jQTBlvYuRoMh8a75ZGm5Y
20Udijs+fawX+kkDhiofOTS6aCvopWr7/4qzWxfuE9PRw+X3h1F8Wy38FDUqLuhJ
0uDNjhfBZw3FFBt0O/tMFn0Cl+mh/nxnlARfoBg4gLEuz5Zgg21c8+uUM+xklm4B
talG9MxxHzH3TBYbBJktwfBgJTgCBe70Arz3WzFocjrQwb2hLcVLrmha3MHTfgtW
1RehAHbpmCjgk6BNjdICvvo9txKMzAwioW7Tr75lhFK9063ovsi4Dni5IEhXZsbE
pyIbUVNvAF37edfc/kRGX/t/RNKO1qf2JgsekJTHYnTLT1xp5uyOhq8VezsZDo65
MHBiLbo8E7FTtH7OCI77HBwQinEbGrxkpVLPhLxBddGpgeZUu88t+YQwBSk/X16F
PYSJTdbe4Azv2PKPNwCBeYYTrmHRxF3udF2MX4g77BD8i8GLWjNTGwkBGfC5RYkg
gMMXtO010OuN1Kq718P1zzogetZ6MSQFccZ0tBR7laXyi2rEXpWF39JZz2GKCHyp
dHw5Y4N/hIVKWZGmaIm87Qjjt+O/uAEpO+gNTClN2FV8x75B96joGLKdn8ZgraY8
TVLS9G6LKELyOqeQEQQQS7NnLvzc4gKy2wyimcsQxxKahMm8EndSMzIMiIQ3WUeD
i8xJhl9avKdpNPVGhZDhy2reuo4e54qKOC1gLRPXhgXvuevGIJZslXeKwjM7KivQ
j9XYtj9nmHEypof8ykS77fTlGUiSVVvGVdfD8UUM7L17mWfDbFwY+fLjivGtLO8J
mn5Y6Tq0JLKUqEgLpALHUkKVuTxs7ASKaHm3YePn0KCCcqs2E0G1tizeH7AJN07p
sPt1XjONtdl0q9nni0uVtoXquYPwAP1Eu82YGd8hh6TjvoNQ0tFZcdng7VmQjIh7
Ecizuxhk94+KaVj1awbnf+gUEJcpELqlpGdCKpgOQmjxCMsl9Dupkh+pKOKmcTxv
dK7Xmn+ORxmgDU49DmIMCSiK/AJ01agPtqs+fIP63FP/zOCO+cvIPnXlPtWf730e
Ap14u5zs/KKN3gwR3iKKbWcGN+edp50BGUjLbNMy0KOHKrwnc/hM2g7s0cvDzh5O
Gxaip6TxgTME7bj3bilaO/Uc+6lODhhzwhmq9EFRYnHms13x9VQsPy7kfHjMUdcG
Bv+iBkbPbVrXKdLZJqOvecVXPE/MJGjXCEgBybOaq91ict9SM65R57ldfWuyiav6
gYYY24VfI9+aZfuvbrylC8tJAc3L4Lp7KJOE9qBZHIx1Wgvj92qDDG2dQfEQFKyE
x/OJt/kf6CEM77ghey3p8MLN35HTj/3nxSgBVtCNS4tTzYqSltbdEQ3h4g7rSa2D
4FIGOvb9+MzgqQr3Hh+nhHKrzmk5ygUpyshLwph6Vzrebc3wbqVB0cag/PA9BX4B
IeCTO0LOWSXNi/dmihS9QnvNgxK/DQs3rI+obl2kuNJkl0mc6+d+Orj6K55r2hui
saTntaLOooT4uwCVPQFpzZVCTMLuEb8ronW7PsMojSuvcmgkx0enhtSxVwx/haX1
GcMYx5VdGwcY81EvRc8jPlH/1gvkGbu4lGzC1oenPHt6+lAhjk6yuq89Uhz1e0Xn
3VOY2CcY9mL1GOt8sq4nXsc2kH0Decu6Z8tEAomRgA+p/jRKrg1LaTagfyVzIH2H
PwlmdwvJ9s6G8bq5P0/ZUBf91p2A7dlxJ+MymRfxUgx5uIMsU75oN6QE8xfDJijZ
qt3PvjknTtUwI/jUbXak/493XXa4dUJjPEpZ7RM181YTL7bE1Y0XssVIYOM5UpIO
gvVJVVH889+BxKxkSzdBU//v5RGxQ+GZGqrkr4Q+njq+csOx7/ttxFiXS23PoqNl
7AZk22JEZWfOI4bvdFF+7OiorrmZ/sSixuO1Ueol0yisxTu2J4+YY8pCMXAfqSRi
QZtahXuG3UB05k1juGYMaWFVVPIPdefshu7npa1t34JEGv3HyJqMDrArGGoPHTFU
tJs0pRpKngSsr9JXpe5/wh4pIuB6VNcWYPL78OQP4LJb2OAQ5Z+2SdFq8nnE1vlt
Grhz/3wXtJzzAbB033gkZgW/ymS6w4axmcwzuSmGVjqReaCyiHK/bgeTGRcTGCM0
rhBwf4pBl/CheFqNWhq/fESYmG5Kt7KX4EbFPwLnTkUNeOzFjbjHubzawJ3rK0p1
z1m1otKF1Cv78ufMQHs+qfgpqeZkfZASk36K4ADyNSRnFI2gElTY0SDubhLnOjMq
EGBMejoVRFRxxdV1blJZyZiMV+yvECvDD1Z9BCydpNvgrRoTIZl8f8VBi1LKAtM8
GWqTWPQHXRDvPzbKsiOqR1eyv1d7WHso06dlUHlsMC/AJhZxJJoQctO/inkSQi4S
j1WKHAiHDQRy6TXAj919iEQS760CcI6GxQS2fP6rlxDULRquw+jLC/kTWaNgfY2e
m7J9megzsNCHm7dmsmeSrd+OtgVT9Qawoam18uQ2whl90aa/UUJTpdNYrObIinS4
OFKvEU46jHFCowIslDnhkSsWSl6uU5HwVq4QViwE7QrZtfUX0ZiemwgtVE83XMeJ
LDhalYVu5NT+b1jmaxzWnrauV7DnYwWK2f9Pb48PRlcjyMSaYbQpTwR77ynGZhyR
bFDMjoci0SQHBs+u4lTtTO6x68B4Qw94VlyU+tx5Bwu+MntF8DSb9A3DrJgGCgCg
hGxP70yMuNAHPQ87tsSriO4aZkq81wR4iystXeB8Gel+YakUT/Egxzqq6R1OlLil
V6tojJCNMh13pmrs3LH+DHeqcOkYzKLHNyetc+vPn9S8nbJy0taYFKx0pw4O8rTO
MwvNG9USQLWu1PJ2oaCohcS5BgbzmAv9kLHoO9OwTI+EdF4UGIdbnOUbjQ738zwr
AxECOLQaEvzoD9uE1sXhdjYsIJJwVscmvbnYL2qI0Ln4fMmGLf9w3P3VjfjSoeBx
aSEa+aAO9XoQCEr2twMz8t3xCkYj2+SL5ZIBhhc/R+Iq6B9DpY/pcOCtEvaeGDIG
qMVMvbq/rjBiMu4vGxvQzg0ViHIjg4A6KSgguiEU6RCveCcBeT99MAVrjk7OeV+E
268sI1jB138QCNAxTay0CEW1nXYerTwlViGitLdpJku3x/Ap9vZx4BellaSTyixJ
gfh4QgngiYCSRkvu+NQCa1FVclFZQUqjOrwD2eSLZt2BRa18xsvgAepERt+m9a/Y
DCNnUs5unpKoFkzPxZbJEfTUdDLBAJH3ZSMPvHltu61GYIYk0uH/BEtQMAQPd/nn
4t8C1GMtwFaIMtY076EZeC4QHXiPyGEOMi/VSiDjRFY1YH+N1NOeRMckxA71rK7M
ZmkrCY+Q/NZe6AceK3NORbCnJhVUSIXvcsL3aqQ7F75yX3EgdrJdadmahdtYqYEC
udoYXBI1nas+R6D5zVYUKq6gFCSp/2+8IibtAnMthhg+lEV9yARPImZyjB1dbhxB
d53IIeh8Pcy5fC3cVnhbGBdd51y+y7tdbNadAO8VCSWm0fuuJOf07rjkSyLuYNou
Y4LIU7qLJicTxGHnKPGH3fpIM8jx+spPZy1oAXxmP8ro9uIi/OxvqPk7otU0d54d
SDkNKEN2crbvn0KmdaKGbBiOyb3IyIpc/JshuefjmfwIMxUm4y/3wHKOw9KpQ+zE
/naISvh/MjvUmHbNrcRlK9dpHEz65jSRAI/qAovQ1XHAyJLGXA+ZaUDRDHEVT0tF
IXGozIEZDUKn2uAVxXaUNC/Q2OcGaMFhp5bCgYQY2XEt5coI7tcvdvRtAr+pTYfT
VGyuHJYmwtq1qj06/eG9Qgdt5E5W3DS2J/Hn4PNl5E0XSPgqlPWwVy+nQTe2ctLl
p3B1+iD+ALYIYnzCa55QjlKyCDbhDwQ7vgmJX1w9dJbEbWlBsSldnAeUsEWq3DZH
VqA2NvWs2Hi2Yy85l2KMaUmyoSYP3lLdQ1YEw/rrZW/SCP+cbGyXhqgSGmgaAN3+
17/uFWWM/pwwQIirGnBFFjjmfRy1+BbesSHOZxHkDgWU4BYID7PkDh2tpwZyz6+w
5af2PCJ8lsPmTLhjLiozskJLtaTvXN4k1LiVNFv41vOVRfxzhdOrK/yye9XW1r9y
0fZL3qn6iHGMit78sCWuT4AYbmeCvLDD9S/QKeB3pNvurrSxKvEsJr5IdZfqO+0d
1qeBlpU3yZstCLFn7nTDPG4ZY5Uok3mWdHZ04jiGrHKxrcI8vanH4v5xhVO9fIge
0GqffzAUwbw9qe81COhZyWaUOPFBs4Pj5pjdK3f7kPqKBlQSjS0XJee2SmSi/fcb
tP9WQEwRWxhuf1QFAwpUGX1BS093wriQBMKWcFUd7erBaDgAxHmjvDmDb+KYK4P+
zw3nymdV4tXe798WjfE/H/grjPOUi8Tb1PB5wgL9igh/r+2cdzEOnO63zcluCi9S
8Qw7wMOJsF3bJPuv2M8ZkwVkwvFki10FFkKHIOD3lYrVEFaBTVrhO4OXH5l/cotr
OXW9FTGWBIGCpvnDrxo4lF5tmbUpEXo7aiwL0MtKde/PJtgNDAkn6SyoGrio9883
Myp8ReES4dvVQU/09/tAQ1Jemo+Zz8Xa63r1zLeeG4oWT3Q3NhOBZz3Kfx1OBXy9
azy486aYvEmtjT+/t0xkAvEK9UQSRqhMM614pTRV3e+MpDgQiPg/4WxFJtEjH87F
zibKjah/y5zm6vQrcjOTES6lNckefjd01t47S5YUOWAGAUiYam5WooBnJYa83I8D
4vWG1hcN2V/TrGn9pW22OJhN0dRf97UC80LjA11ThTEprHqmRA0z95jJPRQWyb0/
/No5yZkFsxMveesguVYidzZ+4sE34f1NCAiq44K7gF1zqnDRJUByR/+BwkcFo26O
071V3lho9tBOEqiPV5q6YpCfGw4dYo8v/G8ZUKXzkVVLkAVKx7aSsvtRwsZPD7Bw
ElIZNJLfKRpEKT5QwlC43IItvW06vTfJFRz8emYpsInW2AGHtjGTzMXd3EQsZ1nL
7JrUnhwBBWPv02X20oVsWYk7VHMWpQukj4e71xA6ciPKx6LNI5xp94VPsG8Iz7F9
lqLOPcPpi+bd0gxHbsakd8rt1l07igL4uBArv3trMjRUh9Eug/426YZsb9hhw8ny
m4AqmFhurNIpvTuE4Z7YCKBJzNeS+sVIpQWchagEMMWL0nRMNVj3AFUbBhg3ZEtv
Qe72e/QqcVKtHTVWKFI+1eoJVL5Q5TZoXtmQSQPlqIGBrCyfl/AkhVBA7mHFMIrd
yi/s1sdnRwmGjl9exR0xapa9OAPzR5cktEAISYSMgAFjSv3wv1SqVIXA80kc51NP
6H+RYpQmzcZOWQ64QXwM4DuKyVQDkRdwLor1ww0IOC4v0IRlxpueH3ZLijFlRPQ+
G1eREAKZxNI4FLQSa7AMvEaJ1I6NQvamtwEgP/hOyhijzpDKWzP0w7pV3uCHOlM5
KP9FtPMBgaPgOdwJ8LiX//q2V6EHrbelDAOtKjj2CfCskN0cPFYsHYHSzTOuk6Fr
GoKMoIwD8NA+vCtlK4KSwUQ8/MnyxZ6w75XluqZDQcytbBOHKwP5lh5cHPxtIBWD
1qH2159qmjpiuIH04o6Ed6po+HnN9W7/3/PKySwYp6Qp87c3A2xtOB1j0fefNp7Z
ySFg8iYAijvUW2/0iHRi/FNwf38VJPxafhY9AsQKQJs3jw+4FIF7tCOXAgZ1wZNL
AT7NAb71Qi+XXZJ3B1CLjWjjGPmEOX55XetMKy5eV7cOfGC0jHwquugvwcnZkeug
rpNcw6lZ6qahaM1npkhbWzgYnPFqB33giP+w1A1ftADlxT7t6WvnGrmJD9LpQXLS
AFd6zwjAcLGJxeR8ooPIYBw8erdY5kNpDRT/EhSWkc2NkgAd77rD5pKkluhtuiDf
hjTZg6HvMFOxUbyU3BIiWQ41jibCKCca9szMlSO8kfPXR+cv5czy7BdT0jljRqST
9/17/oqfGpMDFUWRkpWf+Kn5SPdRYrCa8LwDPx4Wm8Io4R89UGmmO2j34HLjC5Ot
lU0/MOUpm5EOgV6NMUF5HYnkZpDZbi/6nz2rNEQ92fmhL206bDqIiOSVPp4K1YFd
WjVsLJNS5vO3eTZSMqlIzaE1/HQ6D+gV75V9T9Mb1cAikXTBtIpYnZhz6oB3UW/W
aXvzT0vONw/gedcRtunu7scsNH8YcRw25c5/9unEsr8K9ppqUCszga94LtVnE1Gc
vKmjNze7e+nuVJ+kX/pqnV/pUR/xXU0DPkwIYRBVqq+aFJn0SjGFh2okKgrAOYNJ
RncOjYHOMLv1OZ3KGwKJVn/Ynb4bASorOtcsDbKCboCwKwkAXxZuSvKKyV2eMOBL
GNHKorUTy/roPzKDbYmxnMKp9sUqGcycfvFcynAH+G9cUk67iiO4kzs550CfMAjy
RuD9ktdzoJdlqIrElVdyZmXV2gy4ELGgErWO3iiK+nK/3jjgmqaseRasFvTi6zV3
0lRO5ggQ5Ia8JvznWkFptfyax7aCBj4+xQh94040UvAO/OVvsHaEvchhql3Tq71W
y58Cx+oZc/WSWFT4H5NVeDvJg0m3lRwDqNgXYKjwA09wi92jc9OLnZ923dhpLb91
zW5bpa0s7famX6G5GVWO2MQ7g3UlS6pcRXYKmiu5qdwjYbq8JRFYRqbyhEbFVQXQ
El+puoF8yif0p+VUOUCzzzYv3p6TZL45G00L2E9LztqHTZKYj5rHdTskU+yg3XIE
jiiQx3tupeX3kN2PqLBA7gFSutD0bP9jTQTEXVC5k3cIITBr4SgT6B7BcDmSBmax
2UE+TalgouxU4Z4QqAfqBSbo93z0CncW1GoRTTzFCv8VltKMaootJHh9Ii549yd3
wcl9tDILY8PQzpvYPZHWmNPeCq2F4CPzyonyg8OoUK1/VLU/za4u+BE5Ierl6T2f
QUdNaGrH8hWgJZXXzxbDm9oPFaXaoz5MgUkxXab/qpRTC+EgCkP4XGbNCXutg8OQ
N21FemhGzqv6SUnIy9bLAc1DtDsuEx1Hg94fd7UzgFT32uL2YkZeG1G7vXge9RI7
g5bF+YXJBYH4NJRYmIXZ2al56ZugJ8V+TEIugk8AgwIR08l0Fd5PGigpvhYwoNXE
USy0hio8bqDHuVbugsmDHWjzx4RuepIYfqqt617vA0tJIByhKDrkhqpjxyz8ptas
USZkmkwZ5DEe+jlArp4gqAafurp/b1BC16oJHOYDYyDlfdWn7LehAiTLT0CYiXbG
0zeFokJlZ5Ywfy3fSkwji8lxxGqLtO8JySl/25KKBChE3v4iyEo38Ewae7Vc6/T1
z/v4fr+l03zBSnhmO8DDvCi1JAQnHmX51l4CvLyPb1ZwHJAVQfXgAgJqQ9vPLYLw
L0zPfl6UraTLB4Wl9Fuhzg7mGd3hzJZuYrALUdIXypA8Vz+6lp3B6JQczLDudqPA
uNHDZafSQ4deF3qqvOCTuVEbrp+V7XsGwQIGijb/Fp83iP1KHTinlph8TD7IorST
zQXNksImmf+hpo4twXSuyguN/89eTen2Uh5q7UkRqqCuyBIHfipE1gVgxvo+6ew9
BL8+HAAWwUzauT3jE4DDwfvUazA7/2c8IVpGo/foEFaRsfqhoAW7t1m/cPG2HhQf
XuSWCN1SGMDiQhLBVCLbEgJu0fTEfiNAkCt7OhTYwGm6R/iJxRtvvjOhRdp+MPRi
BkKJ+l9BawJ1WDCiSaLmwYY5lsFSMQdVXRjtjGom/ImzgLzX6LOdFPf2JMsq2veo
gZQk6qI74qpsbbJelK8UXX59aIoxPtBjAIBxBvZcMLfv6q8jnE8BByscmK4N3+st
qQ+crxHPmpRBre7U1CgDmrZ7sC6kCbxyuRDshU0pIQMgvjXM1aY3dBbtzFdH+Spr
y/QX40VuMf6IWHCgYFyG3qPKzBN21PkimV6Hulb6WHd2WUgMYJ0TIXEUvcacJEyC
JTBPmDSGYnsEMTYxUUqLTQkGWLrfu9pXusISTn+if19+lYUuObeuMdoVxe+4kUO4
sjIJNr6wVq8xvRitV+TC0wrmIg76bzC88XY+hl2RICd7/4k0TlB8HqB7MTpz9Smz
EBnv/WWv4QchZPrKKILdyeAG2f9G+TPRSFmTvk4u+XyLTzwPdQRD0zLp+FbMSanl
sNQjcPSBFsIoHFYyDSIUjKxOwSvBlzd/HwiiR0388OfzsLdNRAo3us+nOYWpGVWr
Q2HNamkJrO9SJ0mXkMnV1xXAr33bLWJr9ZaybPAL5ujcUaHgDNvvx3F6e8KbOVTF
N9AefuIloHfN/0A8v4JmaSfl38sADaS/u3QLCeV96zFD7qjUk32MxR6v1Kt8va34
2MFzVV8kLg9HYo0ItqgyRCBKFrUEqZmsNyc6zvwL4f04OAi5ffOl/nbxf6VQiRE7
Y5RqzTOQ4Lw+zMI3XTx+zLkGmHs4Ou55fPM1lfjvuaDlxiEiVRviecx40ifGJkoq
eQLrjAg6YYnPoDB7x9Odo7G40SSp0ZO6LoOGNUa43d2ikkp8rOy9WRjjtMyRdYoz
MmRZKx6rKiMBRCyVKhlJQt7U+Jv4s/Dyp2tFXUMQvjrQz29OLc4tp421NLZS92V+
5T/4gxhlM5howvjwubLD0Q3WoqbCV9UajvhLN9tuvWSDDy9JTCf8v5CsOdqPMr5s
MssFivoPF5ZGD7gzcQYRXsxDHqdTQd7mbWpVVU1FfNcR88FlfZq0TK40/0H8rTbT
k/9YF17uNtcpkiLU/jLJ1pDv82iWQcONha4hUwHYIoljdUtqUd1wCaZ5qZyjTxVe
agpEaqUC2F3wxSVxQ4kT2zzdf2vpp6yBf1ynXjxYxQlNO/p/iq6iD+jM4ayynGa7
28j3BG6XWosJVNUYbiw4rUEjuN/QRrbEdLs7UArt1LfBCgPGrnVQBuR3P8ELec3+
fxt86bd2GxlTDRmwQ76d8c5bTc45/gMHZ2luZCDcG/ocj4bqQqlFF7/OTfM1NZla
KmxQoPJxOWqQ8u1W3l4WcUgAWf3pxlJXGqy3J2gjxk5457SNg+CqfqqcwU0JxQ4E
94iup8SN2/4SRniIZv18acC99XdifoaD9D6bz36ifN18jr3fl1bw9ZoaoNJqFohK
Hx0DdtiY11gDp1ISx6RmQz5osAkh0hgRNjUSi5juwHinnP8nYnKWFn2xyUYkM653
Fy9w+u58UUWVbYjuu3fxuWAciNpuV2IzP9Ws8mkhht+OKAk/AK654VnOOeT7tmjk
sYvCF3GLq2tH6/4eAfj2HLv8LtVr7xelSLBdGNGDk2t+/IVll2Gid6UfC4+8b495
TRmKiToKh2y0vlJLWAy2+6ha2469WYWSInCPRQ685uTOQ6BHwd41vl82rKfjjKDw
A2scgqVqsi5Xd52liWzhzs6pZhPxAZ7AwNc9lTWfqrAWnRcIMi6RHCpqtEuOnucR
Z67Sy1/OaFGZdmpjGU5KdreQGiUzzo6lFMRBP9q6AbeOF09VO5u0CsEXAtCkRCzp
Z1iCiztMQTDh1/9ghxlpTpuai1VZfGE9FjhK2htOVExiOYd7d4OM0ksgq9Ykym77
Cw99EsBrsw8OiHXbVJFP4Tcx9eE1UjVgJb5cNliRNNjqQsQQJ2920Fv4mpKXrfYL
si1bkNF6iCdYZyNmMIhlRUrEIvomW9egqz6I3XU54tSoD8FRgEsGUbSDDvFrarpI
YCp0jUXk6pZpR9oP4Jg71l8cLHY/oy02PzyPfYDW8kGiwjtyfWpzk77+slqsxv3d
6lbMQAvbL2uZ89aADPy32KXccxjFQG6/rymjuQapqcwjA2r5fi47yvo7ZNCdCTHw
xog88rXn6jzrMVvQe6+uFfoi/Ito6uK7IA4rPKV3rgzpITMEUHDX40ZIT3K79C/x
YIlS8Fw1QlmLcctRyIkhCHR+7P1fFvxLVghTe8F2EfaKe7qwYscBsPoz0z2G+iaY
t4BwI+rzMdHMrY8dBr9vgKvErq19iK7al5lCtIWurya/nMsUXAtZvFA+9RwxHAZM
yHhijoprUc15lafYkfhPejVFRcdzh3xKldhxJ4gAXDTWr2r4bVPd7ZssanBtlann
y9FS387sB+2+wZn4w+IVZxocwOBzoaw7mYZ1Mpf832Pxc1X9+A9dXjBj/JaoeA72
92BquAFZ32oPgLJkGBStduMtKA0qDgpZOFGOZeifS5ZiiSC0kBYNMpqxULNc5NvR
s3b1y15QT9a7LQOZSmYz/vh76IYWMz+ZssAJnpCdQ+VHrDRw9b9Fy86gR0j2a3tf
3FED3cyUNx7OqUjlU9NhE1UnNelz01qH0/AImV8du/VBFavHW8lftp3A2scj1BGW
nuj3gnUlcVvzA13JD+pluVMXBJ3fvs6HO1WEooeHNhlmWcAgljSvXgWmUnFKBmTF
/UzI9Bl91B2TtroUAlLgLXCT6KwwdjSf/ZpuUEXIi3HxibDxytiTPT3/QcPGlJQb
H6Wj+heJUzt7rogp6nJKxe2naL5Lym3mlTBP5572hQlMs/Y5ogqUBBrNygzOTjPD
7QKZgcxvKbH/s/QXRpGaGyq+C6vDbOAKWx4j/IQJ0WaFTNrgzvUOkE5ID5o3ZS5e
i/am0ExriaY60cUTCgu2gnjnL4P1AY2UcQSz1IKl7rr5jI13l2sWRBTpvQTYFDWW
kL8XLdM24e//o5KulhkTdPvTqMicBsOyC3dcl/tPVaT8Gsl5/vbz9+ryNha5pehj
hZF+ZsUH8ePkLYvPfgiS6NhCkY29t1UaKclRSpRgcxnJYvhTzwY9U5ucsoqbCf6W
b+yoW8cifEYmw9tgh+1vMHpZS74h0xXzsxk0U6Jdk2iiH60gjQuSkXPTbCsKnWDX
QHtNTh5jIKEMRzP7rD8U6EiJNmm0FykJggP6vJbCoqtEKAdiqVE1PHoJ6b28Rb+0
fjx9kLVImjN1U8qE5JsFNrjrFyN0lmCU4IFaHugqAqlr3+SPjBqoXdDrEyZkh5oL
knSWGKxFuCIYZlnRG6bStCjgR3LwrYLjljhNCQNmo4fD64oFJknFN1xDkZIHsVzK
l/WJA7lkGwvxSAIzN+/tsQgzr5sP6Mn1Jl59O8EonpPm63gvL8W/Scksd6AdrRtX
an0ncRFI19Knf1+cGGZ/vp/NxOu0rpk4fb15A5Ot7fU21GIG2zr56vQOLpLuPOPX
7yS+9aUNxEjlRUJYr6QHtJ9tD+eaUUu/D6ksvaE7WLMrbyUFfHIwr/fGymp7v07n
s8D0PyWI+W8Or8FkxMrt3H5VoOpWMfmEC8trFVyMJ4QH33g3BKU9mqlZ3UrCh9pF
0cVMOp6PMiFxdVU5gIctFnEue/mpUV3lkiGrLkdv5eIJJqTCPVgHB5IWSH63D+l4
FjVAfBkr6HGZELb3cePT6drsv6KBv1G+66oKbH1fLK+RxaIg12RCZawBMhRQRscV
n7MyQnOEKM4kIDGqtCLI2Egwxltp94rY+etSianRkngVOmcs6Ocq79u2l5bifqjW
/dlmbD8CN5ESg9P7AE1YUN8WVbkFyI3dYAjpdyta4/W0XqalWDOqCcMMv5LlkiZG
lBTgo13sfxrhO4aheSegWBUbu0Xp5ULp9bWpA1R7uEhLY7i7mEzX+zT4fWyaEZZB
3kTdiKmACfdkqOpW5DyHKmFy/uRebpxjljDfHYU+Yc53tcfhzbdW2e7hdTdvpWPB
orhtA3M+DUn6P+nGi3KatH/HFIrCKRlPo638qlluUfYSO5aitJOJTSAq4h9tJj0t
W79oZuVxLBhP5gBsPoKoCjOuYJdLOSmj7V3cCxvRIDBhNqDMVpCjfGHPuwRA4dOj
SpDkGdp72NfaeopPjLKaSbGnTTlG4YHXqKAZtYEzSGxMLEt5b97N9nn+eEHl8web
w4fXsx8Y+YMc21LVpEEzmXeJg2PKRR13Bn5Nt23wmjfW2OQt0VnnvsDY6HZ2sWrW
h9M9tf7nfyLEuuUTTXdAbFIuUsbzHjHe+29tReJ68/Mh+Vi5KE5VnSwEvhugO/y0
rx5/f5hPf+aKsWLlTMCQiVkTxuVps1z5LzqVoduD6ibCzFN8XNQAISUkXhRxSx1c
uab0bprVEsTZUv41x7FhAh0U3kQZlYSpvN4kFnwVIpgPsM2Cl0oFEHz5HLmObk5j
qs91hsk2UdXIA+Z6NsLfeVTkdRZyagHxTMLoHHCAv1tmXd89h0c1mcIpCJ/YxdJj
PMrC0Oa31Duqxdb1NIOzqnRS/Qbb5THgAJhzcd01yY2y8fYQ66irsk6deg7DdIiR
a10VOFH9rrV1++wlD4Vkq6ITGCjRiiGC1o5pBUwhFpg7C3a6GcpQaYINyWq9w7Zi
kLzMoUh/fHMH6ciSt5B5dkXM2rtM4XU3slRU4MJIpChx9nG3m28/Xb2kAgp2v5ub
lp9uiPXAr3Y9fOmk0kzSaY8fJ9FefTWoL/sxS6hGcCkI7932i69EnDG5LEK5uIiw
tH31KTkqXDVKWlaenpXMEfAYAAsg/wyyo4opZFq8iquHocvI7XKV6/jhIyepzvoX
n6ltUDegOLGQ4SQ4lW0SQxbS+PQuti/N3aO0bHtV6iDhEkBV4lKZ96C0OQG0TeVL
o6CQOWDu7FTvZYsXldLj1AnkPVx4Jx5zcjLyjUBuREGezpzSrBwZjbkMDHvjUJlH
Ig/TiPjV6G4OR2qZyRV8C8FqA+0RGOlktgerya9h7SOMCa8UMimh3KklPgJzduox
9qecI71jZzKWLiS4xHLcEEpLsaw1JnPCaT74XvVN5ZeCrVAJparn8Ge/mo/mOqBd
9HNRWIj3tuyKLFTxd7DA68N/lEDMtFc0ZvBsAMLXNL5PABj/t/3+kjavJ8FiGvYm
HAgU3KYOp6RPEbQAozo/oYzb2Dwm3KvH0U0oZPaHjh7rCanvenToTG3ivW9gZSXX
1BOJgkIEu4zUwVExVwnPJ5OQ+qPoZeZ9dPIpN/TQt/DnB/6zrHpeoh35XgAyjoxT
1E/7KSfYg7DByyr6ItbVmHZTZO+8HCHuC7ulVBus35Pu9kxgxf7OjOICF3rTgX+8
0XyX3xJW5soEuY7C3u7iuMrrNXXW4dUI8P4dKL+OiF/nbMY5Vrv1f5fuSmVCMNBA
YhBclSc1yxYdUEEKIhG3Fr+U7/wcZSVddHSbmovec5NAZsr12uvRNVQwI5GwcZkQ
6GLMelgav/KAK4TDFlfJq6ZuR2/wsOxf8D/v12xyQw/XTGKJLmiGikbbHfws5/CG
iENkADVvUVqn+3O7PcGIiwM3AaNpfyyXoDsBju5k5R3XJuXFAjczfPUK+6jwLqud
c3Xygq+y89lCfR6Qz8cNSvCcqBV8OpFtOJDVfoZhIRRbfBfEesMVibno+kx2fv1Y
hfR0PvQs/vuTcAeLgYS0HzADAKP6neuN7ykp3eMLib1l+QDbeqPg8qUx1IAC7r3Q
F85c79eA7qNwQC5hVlrrxk+o9CMKlUCAnSfvrqqoYxxohSTeUcFzOsA8dkvJf9Dt
CAlUpm81TTr9JH/FHjr4eBtc14Qp5kGefm9wk7e2ZEQgl8R2yVrn5ggfwZK9ym+q
ZpUlj1RAr4DbU7K05GFz7+SLTULeZ/poXU1ijXEoe94gsMtqdYB3QB2h2XkZE4zU
l7aeT6TTJLj5O8yZggkGbGi9tvpH3VMR7WULXTiQQ0j2ffx15bbYiYGQyWxfOp4k
fPbUR1J7WbHPKZ7OINrRisFZXMl7emdjQDjV8Oodbtt/zz82LcrK7iNn9M7aARmM
oezyrGzlCFJnZub1+tgClgFZDSuEgdHTs1y/vQgyp6QdqTFJF1JqDAIUsFMehuL9
jA3opr+3qTxnTsrEUFeddqc9qacSAK3lRq6JIpEzu5srvwBsEE+qnCdBXx8kaNTd
oYRzRqIbJohNlFUZ6EeOFMcdmXtGSfzqOp4NTs2b6BqZtEFtPIo7G+NfE99Pn5VI
fJay3CqUa2jBzMKZMB63GurxkeHWLG4mvO+NHvULyhAj1MF+UOeHo1xss4i3C+Zb
ryWSciVRhu6zyjpxaj+YGRh2FxvxfFxlvPTSu4QngfpwBW5tTjHqGHEciUI7BYZd
BIVksexHZCmRKYTWOQcCip2qIFjjOVL54Gr6dK596b2sWcj/QOTDLmtg8obWh6h2
doztvgIqletCjtwmKbUYNhZgNllRTPX2Uc+mC4cLCWWHytP69w7ECJKR0VauRw7b
TzB2/M5XbEWB9vARgPUj8Nj9AZQgKFysWaA7YEg5f/AsxrqtVzZrjxBqkAVpj69G
cyltLTdDWBNo+GZg6R4IM+MvusnXVfR1oY1ZmWp6167d1ewWEFCjQNfEOYLg6kTt
NqRXmsyGKijr1iupIl4cgDqnCqKlms2gbH0/TCcCGKzb71l6WUSaO6XR10H4WCLo
0BL26BRQfnRDcNiY5SU1YUYNVuRp6BaUP4zN40brEqObYeMF4aCebkGkqRMnFBe3
VMQOAzQa8AWT69d+Ii0/soU+og7iGDoBbbBNKeQ8p06UYSG+IZlDj9cwfPpFl2KI
sqLnIlB3KmKEWWIe6V02khfq5/Va7vGMz+WWanCtp2BAmwGQp92AjvD091FMxCVj
TdnbsYGk+x1Owufg5xayJ3b2JTbqGLN+rVQW28xvId4RN7nL7t1sGtt+rkfXQqQ1
s0BrKnkSObt6I/HYDQ9qYAFDexBOoA5UjoGzHUZ0hGPYAeDb2ko2UdxJs2vOYQTm
mXI555E2Ttr60DdVHgSUWf58qFCEwahQHsokMsnw6B2NXQX8UpbK2uQQLWGWmrwm
2G2n7bvnUEFYlBX/9jNz3z0K1ZEeNMG5AJv8k4ffNIS5acVgATQjF4DU+Mqgn4Ng
hs5MHnf7b3+Ab2+5VWmkO85jTUolxK2zyJYCvkJeRsYT7v4mnSBd/WK5Nj1ha8ez
BqF3myTMcQ+lhuY4V9SjUG7nhkt3fYMKAqgxwYNGmGU6F4o3xmn+C+XyW8TMd9YC
FdjFDlhfHccYEI9w6sngIXe5cXbcEXZUUdVq6NvcQtg9hMS88N3nZe9mYx0KVxh1
a6CBN1O/bDEsJWfaqG1FaPmdHgwrLNxDvjEM7ZhqR/TenQ+0Gs0Tld/SdvpRikSj
Ha40rE5gcjJDl9EykCwTReFXa4DUDCvf74w6m06gGA1s6IMJBGLHIl3kMhjhXWMx
5ezuY/SYxjGRTvyIwYoaCFeTNBxLUNdjV8DZVb/u5BCq9BkwqPIu5QgCIFlFmpjx
DyX2diVjInt/PPg18LJ9SGZp2/P+Juhpv+E1k9k3pA81IwRPLNmggQo9RKK1TlMm
QsiTQsfzjDXTu3zHtjNZ712uPZLdp9LTgqLAYuvubQmEGUp8jY4VmlryGJ8olWzN
X7fJcaK3YLLjtfivucZIm2gqAF9uzOboDm/mKr1Cb2yEHxv4PMWhNt7Mddi6U0Xa
9qX+swMcwO2pNzDelf++bIkvSvqdfBwtpUnGTJWJ/9vye19BGKeDyu89mb4oEVeC
Bu21FKyAm+33xYD6biW3vO9DGki1wmvIAuT1Ndl+KzGEHOlmaVrolYI4eCWBgkr8
bkDSdpa+EfqcpWonyh5Ax0PU0ICflGrz/9yzc55aah6KzBnaYLf9qabDkFAM0XDy
Ec0kzyxi2G+W2sSjuK4O6HZuejXFuohvhVG+L6SonjLlTVQrYcoFL9YFbNSSd6Zl
1WhynH0PiPkTKCSWusrWFdBs/tpXbpzC8IdYeCGdt+DGR2Pv9fo5gJt/pSMqI/Wb
8koesDoF1BrEok+BK2Tn7Od87uRzOQJ1m3EntrbuRHEXcIdmZiXyD1szKPZs5KtB
3vV9id8x8DB8IlgGSGCbbn0yxLbxMkCaL3u/gGLqtcsg/BJBXDLppYD4ZmOX0Cus
ySPvvC9PWRU5/lFldVKIjlwswsPX6AXbXmptQ1w2E/OwEx7c0YAzqrsbfednAEa2
Dkpsd+Begp1ZdOEiTcqkySvVYwsrI9d1PdNLnzYXqQ/vIYUnT5I186elCQNm3s5o
x41QKBp+FtdRAB1v1Y+mOMnOvexSs9gQDYIF/2kvaFUjkZG03kL2OgTSUYdIIovZ
A/PteJVCKA0fxLjSEAN07rKaVXv77+6WAT0TVSvKn+3SryTnEfOs9MUAV3Mvj34N
hYiDEIQmVeZBw9Xi44iEPHu/XNTPLJlSIFTJQixbWvYympcDVXdh1zbdr9jmKhHp
7a2K+7eu+qeGTjD3RXNi0ixJUPvMxM4Ml6gv0+1qM3+X+EgdaaY4Bh7Fm/yNZf95
MbOShPvmbQVBMeM/L4szHFRAITZVka9+wj7V3jbz66NXIIuzZTLwSPXPKbUvn9CY
nS/bt7eMhNCae3Rbv/DIIZrfsaSIyRkLzWWSuYvbbVob5SZDwEV0BEcnJO16AY67
C1SsEip7e2qROcv7748ID+UlrIBSHYDhd4hgYhNmgZntIQfuk5sfureNW44QV5jv
hheoZb64UkkZNX4wgje90jskX5OvzTFHcZtWZLtZYYGQ7LT6mMpvMFB+B39MxHTj
8lxgtzJV9mTO+SdN7fkZ6z4VHEXZx0a0YkArbOrEGkBJVigg16UBuraAlhBglW40
XS3ySJTVyUVInkzGE3bGf7BF2DXsba6vzx/Eb8wty3d5OK8Ok+fLNyrzBXpdbLeG
IQMA5ymKqeooDXSqiHHgqCGilmvcNgU54WhyQdPcxOu4f/0cB2V89xwq56SL8Yy3
rN9OVGPpyLJ/+2TL6/VIMNX2hwGiuMjdrzbSuJe8MRPLhxQ3oycKkxCYFifWUQxb
HqEQEEBwJKjiF0V1rUf2P8GjICNosPo/k/VUDnxh5bDvGUZEV3+Y2Znez17iMmXq
4jbjl/D5UCzmp5ibZkGYkvOU1bORQrYqpRiHaQWMAAHd7dfeGEJeXofLzH0tlpxO
v1hDxMW1N30Q6QXtoZ7QJJcAtHPRcpbETmMZGoh7tc8FVsbF6baWgmjJLbxm3YqS
ovwWNLNIXVzLJpjnLVVEy0bW+4HPtu7oG+W+mHLY40Q7r2yIDwFnqDiSw2dAEtGt
w3wVNkIKJ407G3KJq9BAbo2q7ullD9UvBR/kFW/WBiZF0sOqSfkhXYE+Ln9D1jqg
VMTHXsw3us7S6rWALYCWYkAfl8gFb3UBituHCH5bvM24XAhkU5RnK/KskoqUQq2b
OgJuIZ/1cMzgtLul6eWIdu+bvxDkk0viMk/7pKipSfjpWEDOqBeemx2nowTty7xY
dEGlZJ7yu8El5EjkDYwzILZAhUExnAwlgIts/j16HgU+Fg7dXfDH2H2S4RcqtICg
YhuvFySG9GXp5ummEgde/enGPGiVMsfxOyrgOwvUQ2uZOjwlEFwIUpQhFeo0l98E
wDUR55jL1VdEepArA55uc0ApCuxpEpzQU1bfosVElidwsD5ZNmcuUUMDIrja0IRo
S0yX/J38K37vZWWh/B5i8TfZcoo2iXcuaYTJ9WGGuwb0uIJyRfidfMKX0ylVJcQu
mXPTP55IDuzERWrONrwR8UkQNews1CxLme8WVFd8abeSTApZrhgDM4LkzUnljbuH
akGJAlEdcdYJpjrPI/e2zYHK4/iJGjV2rh6VJgJy73yQ2q16sDaYZY4jndDeiQ8M
O6CDFbXNsp4cRekPhGNaludWzOaKe00FyqqV8cOanIaVu/za7zKHTVlHRcg/ylZO
mo+ul7aiH1QhNa58C9zmzNoDDqx3VZetmyrCItzkhML2sL8aLX5Vgw+XEhp5hUCP
TpO7QVOHsePVm7+ZxzJAFn0ltPjAUyU1D7sUKTwS4Sfqzx7Devvb0mSrPmlylDlJ
tfdvSMs5uSZydHgoBM6/jzAEH3uKry3QLNc7ssZ9H4V1eYt4G+AKBckfzy5sTkla
9MYrf8ajYtv1bSwgvdNQmXOyldSM5hlPVVvXjs1zNiu8kvbXYh3C6ZzmRJQpQYKf
iYjXedaqeowWB34QvlyK9NEYrOr+tn24z9i8QG+73DT4EQbmUSaPo28ZglPf6SvG
20Wk4fxJ2QZ2/QeZNNO+gJIRVhBPqpPj5tGsBCDc56EloTvvubk2XEeEhbW+7tv8
8DT/3UeYJ5Lfspk+eJ3mWsk5JHWPnLZb1BuqRtUhFIj5kS5iz9N5/kOfTulTcvw+
bboCDX7vO4N9hWL4PQMUY5lajJwp04n7FuO2ZruoT7VBd9kTBoVoqwwmeF7Wbd5S
IlAOim+wuFHRoOwHVZt/Rvzi45D6JTF65WMvHAkNDfrFIEP2qHsHZfNNzvTQkTmF
OoC4lsN19OXPcPySN75IsvIoUdu1wzcmaO2183KP/wdjPGEThE6I1vdjM2IQFL80
nVnAynjO/OJ8sW3idZ+gacrtV03n5JvpihpJrvNBY+B08NHRER32wYLJexwIdHto
d6rCVi7aGNAbCXHK57ntwgQKLiRosxrsg0RY6eV4DN/dIAo2hpEhuN460UuoM2VY
wN7hP0ff3mYKAPhoLnvIAB8EgLgHZMTRak7aSJbV9a6KnsbWTt/JLVhAofWpG6q+
zWViMmorea1Hi5WkjFaS9yGRsp5+yAz7XG5N0Y4ysk9oAdrK1hrGcVcXSJcXcw1z
r2+PA1uH0VglkXOTLDxd6r7LSbaD54VGe/lyOUZXkIF55CC9KbqBzlxDyb/ZsKTy
b7qpXTkAlSLkpdr3nzbHqDkowIq87uENmVTH7OcOFWw+hczxD9GPQXLpQVMYd29W
R2dFZj1BY4ElQvRVT04aosGmkofyd+uLRraN2LT6PdTaNMRKagxUB9feILEk8zFA
zfLD8V+NxjOU5VvjE0DNl+Ov4Oy5U0LmDT85rcBS1E+fwTxhAGKmra5Gwu3B+jeN
fPrOSbCMq5e6w0iE0aHZ9FS/CsF5x/jZv1rozRikLLKhWp3m8kkjQu1b5Sbo3jMN
U5glcB7KPgazkCg6CNfc1W6Jc6L9D86OrDNjqAfm/jHa0/rjNI9A/0JeqQlZ+yHq
bQlfSuHFt9lcsyZRvJ5RpswdjAbQ/95S5qzMqsEICiYE1JL0srTXhJtmIah70x+c
0hdlM8/MHQUOlTf/tmIDl/QDgdpAL151ZI4MTxsOM2kTMCDHiDk5R7eXDskoOXel
4Ny03zrSqt10NPYenDpHd3Za04k4JYyOPDjQV5piveyNnNn0PSGZ6YeeWS8GQC8/
5Cc0UgKuzWTfyGC6cxnusIhKbvDDLFuWVoAMNlqHoXHUZtVYrr3fdMl0EF9EUnom
PXyTLJ9ZY+BqDwptxP4kfGsDHDpxcziZdREUmimaox8I4ah/DSQXlnrxOj5o841E
R0oOXM+kXHBIvCX1DiwuHaPnSXEj7xnL4p/mtkdN2A6wX9U6as/hHFBTFL2xXUXN
qWAoY2DpE4JkY8me+MwPK85XDjmYdfEP2o426ee4iCjPm7Fwsfg/k8qT9A12Oe6b
RBs4ho9glNHjHTMkzDyuKm4v7GqCgMduMHbBY+goSBoxoJouoDSFGXsx8dIA3P3m
DO3Z6t6QqrF7lOm0cVq8vtd18mLBv1w8+7unKFMbJuZnzJs7Lw89LmQ0eZsCK2sZ
p+E6wgOpFNtRjOdzNeTJVFjLB2A3h9JKt3yMVYWD6ILa0xmlfNl/6NuhQ3jOKsxW
krlNuzhcPBDE3AnR1gRPRKNWg0kK7XlMQcHqqjmN4J65b0U6m3wPXmef+ibPqnkm
lEe0QxdqhEAZLGeDOQDqYsuL1Tcdw9g+EADd0I31Wj/CsIUQehAuE6ZmO25OGyEe
973aS8+9p9Wbgz36sNiEoWS42Y+t3BKgIviS4cMF9XcI6P9XHiHtKgmM0iVtRTNp
OfGdn/AvOfJP1TDKo/RMyndHyqVy5j6Ab5ww0KgvZslGKfqHqfBX4rWSk8n3eK8Z
/LYrv6Hd3ZYcyL7fyn+zAY823QwWRbfcqeYUbwYjgrF6ceY7nBvXp466RhsVIs78
AXAH/EaVkJW8L7rMXQgcUYVaR6Vn9K4dKhZ4YFBvLN2+veJ2wKMj47MsqDeGNKaJ
vZ+za0HapEF2XMiA0NloBiUo76UFJRs8eZDp0piUMd12SWDjP+JCiNtvc+aSRoI4
KKywjLufwAio0naRotYcW4wSm+DVnDJYam6i4W1/oFcF12ymfCCBl4YVVWgp3vYn
5YSvJ0nHFKc4MfA1WRYicFViX3nQlk4fz3sNteRfwU8vg6VbvJ1bhWCSgXbQ0x0B
W+zlgWOq1WmaM3XeLD9wfucHXgV84a2NTv+YDpsibjUslwDG888OJWMzfr1IHvP3
CWzqfUJc1MwstFfeDz6FBMiiu1QPvseGjGvtsp4/T2TkJ7ft19q6k0h1po8oBm9v
MZHkFcThmFECBTvcmkxQmQSzdKlwRx+Aew/SSsqspCprU3taYxu13BF7uHSoAwMi
hmGD5F4GwfpzbAeePW8VXag5E64PhpWnBoqv0+Qnm0BRFbGWeRLWew3BAwn8M0XC
y2q4+4R9Px7HFokuDFPGKtgLlgNiPGF4cAJsFFfg4BbPRGQGHeKHOuWawOU++xwl
KK/gRKhx19uBBNLCdZ7JxHWDOX99uo9eaWKauT16v+UCnRj2jJdjShqS0SEWCSAE
JmhdX9CmSNw52lmzbR+ydSGtzVHiGFmxXOzNEZov3N3cGWaovYQhYtKNrX7UwGDU
YgZiDplSB8Oi82gmIcyJUIK0mDponxun8GgxdBSUyMwXp59REZzV9GXticQ0nq2l
hMSkwIA2RHPoD1FVYCKLkWc7SDPeaf/xKJBvpVwxWP+qLZz9L7vIfQKLlpgtL9Si
C/JvLrB+3z7Lf9PSDQsDBrkZ173cZiuzfzGbx+nlq5StFZ/eN+z7JmfSZHoO4UkX
1BmatYW9Ig6WmsKWcVNSpVoT3FqrYZM8sbr5IuQTOkjCiIDmCrodiPgbpp2UMebM
YsWQ0jV/MP0WgN3ka7nP1XsFEw5SnF7jWp1JfVwEl0HTVYfHPDX13UwW7nh7CSKJ
7xdNcjHOsrjNY1LeOIL7G0rDwCkbhU2UOejYcNKl5Fu6DP8kBDH/Wb6Yb6vqrtZG
K3pQhsozBm3ckZ1QeEkyWwRUfumPPdeeANn19ZovI39x4adEe+C8jdiOGojTrZ7o
v3jEz3mKAyck8hLdK3trcZjDs24P5D3bQuIKzeTw8EyDxKDXKJAQWF7PYfluOnfl
hC5YpEP3AO46poFt/1TwkZ51WO0L2IlFPGW3v7MSx9Y7qwqPRP9aQdW/TjMlyjzr
AZ5ZetKRM477r8ovtkzUcXtE47o/X6HhaeLHG5dzJbjrhg7yNmoc+3wy3fsL5IlP
p8ygZqYJcS5KCCqvNXKgwu/Pink9yjm4qS+7VC3Zho3msQRzftVN60FI1/Qd6sWz
ubh4i8j6ZSk7bGBkeXF2S8a3MNiRKGf38jz9upSVeW67Hpnw1jFJM6Hi1EB0FOQJ
Uj7EFAd6SINtGjWr9J2u1o3fpqrAHphOwcnOpYlkFyGiJIXtg/tgqtv8taZBNbhj
4uqzB++oSiMHuFRYtaP3VUbEZb2zm5nX/9+dKbhzJz9FDaAJZPQzFAMGS+qU/lpB
InzMh4xxxvZE/8GgaKaeW5ntRvA5uvovSXIUiPPi75PUKlz9YZf9lixxzE8v5LpU
E6JVr+YKwAI+RXc0Q9ryA9S7Cypk/S2CBOD48Vs9HkCA2j5zQZtHK23/cgZ979ie
uvxm2y6L/3o3fBZJdpcJtxM1XV/WBG3xJ8D7tfK4TbhFndlBsozsKMmIMFmdghgA
IFgIrl6vIPjf5QyybVNlNa3KiAhQGFCbFG5tXMoUFB+N/4QdMJhaiWfDWePy5OeX
Lz57Ot/EoFv07hgEFAQ9qUWdjfft4sYk+Myu0GzwRH6pBdvoCjfm8nbTzsX4KEtx
HIz/Q0ei3c/yb2r2LgQbmS7bFijyby1X8qO4krZyL5Q5/LiHxBLuTgbK3hmgRF2r
j1gfXcXSfRiKrxxOhWeqW0fYmz6jIIIxdQcjOnaQxz0bbQoOCrTB7y+zjcgAwIWJ
+o8yj5lfsX8Vq7+LnVKjvCUux0csYGNlQ/HPkPgCu+BcHcF0bot4BprKz4bL1b9h
Zcc56c+LXEYuRLcBND+V6aXu4gSY+LWAhvPmuRY7AHcIgkFG7GHrJxgb/FoMUM6r
eI6BXBHCZ+1piVTu2pGGqaf/m1e24nbe08E3AzPvhbiGpsYPPLLyxnkXivM6lx2B
Gup9N5qQxCTnLgTXDxN4TjKodC9PywcM69ymXiDcXK28COGp6BVthxgLf1uNJIhw
8ezboisK2Z1mppPOHZLCdJCsU0TXx6bU1bqtokm3ginOSMbYr8ZwoxpvEZJqqmLr
sN4yp6XMPsmu8GCm5mB1Oh/P9j428oX/WbO2z8u0fG2tr0TBqO6M92nmIbbH6zsw
s8aEeOKY+Z4jPIv8908bDbnnkB2H/HQPC+ckIC9UExPj3/z583PxbE7RcLGZ4gZZ
owTRttY/o0AK/1YgS978nicmGczRQ1N63mitoTPlM/xGFJuG5MlzgycT0IC+3+lS
DEDXh7JrBR6+jcIQne9gUQTo5k1H6qBMGE/2ddiBQIIQdU8Rdcl0XSI4U8467zU1
/2DjrJ7x7jUcwR/Tv5usPNH3+/XWiSUQ4p4NPrKYx+bBSLeX2u6hONp66ixHpn6w
L/A/wn7g5OrNuLYPvW5fow3li2aU6QfIMxA6F1ahc2Z3SvIRhkazTGpBXEHgRrmt
XK97CiNHdna7mkFZewz6LqYgvDxxQ03sgai7i9RdYYWQ7MFeLr/3qauicY/IlLBE
7yWljiJbCOPLxtdNsS9LapE13+nu2DwYnTWyY3gIeismhspCdD41nviNSKChI44I
BkFlocgMMbZsaLMjK6JGQLqZiwPJXfV/XLPLut+yVOoXHL7wtb60siS4JCwaOLYy
ihHzuMBiJe10XTn8wygqhEdu37BU5nSSFN5Ac7TS60KKByHGRKjKPKL2ZPLWkX6B
2H8YJgCN0JTC7NdiqaN6KX+ABF2JOpyjbdMTYiazMyW20ts6bE4bl3F4qutoO6zb
HwfgltQ2JM3UUkLBJ3L51JGbN5Pg+1k9Fip7tj1SkCSbT9hZsqg5IF9cL379vlj2
Ei/rMa2SWQi6Z6m/cJWyIV1nI87H5DsYnMdr420YoEKqffCZjl3IubfLZkAb9Dgy
92cVuPO9PN2Q5uofqOW6Sizy5y1DWFwAogWc41ad28b398kfHhdmm458iI/hATlV
gd7+nRAe4qG2CpoLZMQ6rhVTbAzPb95kZeFxBQZWNIiDskGpUZZ3aSnoEW43YFKQ
pDG1r1fh0gFvNZ3FpnA/B4msMQVUSokMqQOPEpW+R2MI03LGhAfy+29xHN0xHDGP
P/VUvd9P1UKVj1sAiFOkFLt9u2Q1Xi76MdtmrYySHGPBojYbzn9GgoE1mVx073s2
ci/SSl1dBwiGVfbbBXkoQ5jm9Sd4xNZYLV00jiVO9/RpwfySM5pb9XVelww9pb4X
LRV2tDGBmj70ImlsXFxs3lFS8k3hhdk3BT3Hy5+ApA4ScIfjG3xiTcL2KS5XZSTO
PyjH1xLh4JATc2tB3VBJUuCslOwvKbllp/l2bqd8o7Z8EdpWSweafB1rtyjtDqcA
4YLOfFai61+Msjn+c15MT5D8BRMgxs0s8c38yI//kcCK4ySy/ucNxUy1klkrRJqV
EwER/3APOQkDKqej3tg4HdWBH8cTv45Ac2tjf7E/nMz9nwQH4eRp9Y1GP2e5KCRT
hR4uNg17uTAHLnG+IeeVLgGwP9iukm+1gUjfyf1SN/Hp8NCq4Xk41SGsJhBFVJMU
Uabp7pfje5wToFu1x3MEyyGB4J2OymyIOvPT7UWFdafUGixvBbhd8YPBx6e1xoKk
gewK0qNG3H2036n9IqtoFYeDasu3gpwQDkZQU41OwUjnRn8kTOO40Owr97wMKbeI
J5j7VoU8Jers4Gw8KfE2YoxV4NnTSUSr211s7EzkWV6nt+AsUAGfCkUbQSH0zwGH
UqbREVNiD2RtSVc0OvWRTjCIUSd2CCme9kEQfINBFp+Ub26cl/NdQ/T1u+nzs5TI
D4eweeiHG5QpsxlHyBdlfGsx379oMdG4/GdkOonR34qZJ8zCPMg1aOEu3e5VMixl
zYHQduaj2M5bBbdHrNeT8LFajdyoI6U+X2cyiemDaVxmnTrYKpJDSUJI7DUDDQ3U
hPHN2joijezyF8bb7vU74xShhAVVM2BkVe1Oq+SLEMba4T0AAKhMAAsoa55wTjqI
wTnyIy8EyTn8Elnb8qcT59Oq7XYV7aynCtRbZp1LCgeR9ViaXi/XWh1AAYg48I+P
rD9EyBLe7Ekkje/WRepXu+fHmtKRQ5t+sqAb8qENEKYlUbCV4q614nnYj8T/l7VQ
lem4l9EdTYTfyW4vyB1bukRMzaQMlp5onCHmqTH9T72m1WiA15zxKC0X/n5LsDn5
fiYIyFNf4/zezIMmyPa1YEgY88S8ZnzQEh4CRk5L/Yfj3crGITXiOzDGI5Vdo6Pa
VinPRik14kMvQntMaGWfPjDTqs2MMOPZc3G+52jd4tXxj0PKtgtDk0+oUBdojIN9
l65AqgirAma0EwrwJnWHeM71php84wBINucYm2Z4fdu5ZTLHdj3DUBm01QeC4QyW
1g7B4BIr95mPdEkDiTEyatPZ5AH5Z1RO8yQ9PYNKu+PsllWGXc+qhrWcV3w6L5Dn
ltBL1qdR0vXVaRNyQiRw7UHjihpjoL11spgiYoKkJeqy+zFXlSgTiJTwMDzhYnoa
bBOBBzaRTiwR/iGpxvwZiLjSIKl1g61D/xDyzt9WBVJajgiF4jRg+PLpfuoYNYcr
koHd4Vt6GtIQTmQPpz39Tl4slcfmL9yoLsyUqnl0UBy31pCSl324LFQ8YIueB800
GSPHf1xT/ZGZplrCq8Z1Jci5D42xNlfKuTtxwQPHeVmnYnf9M5J/3dzO1eE6Qljg
uovnjQHNR6Vy+/NaNa6/w/iPhdChoe35zKmbMg0GW85C3WQfCylyqt99KxxbZ3Q/
v7lZ2edI4L3i2G3RrXBOYv5Jmx68Egv7H6GRiLP3M2RhpV6k/2FnScGkZKVBh6AG
MPknPZyvYo9VM2XHJK5AGEWSwX1yh4UUJUOrXqPjnpSRwLGXAnsZEB7eaeTFi4ps
WExBvObojIvrlsEuYksyktGi3zu98VknyIHlPqTcIWqDViE/yGT5ZckQrmhbRWxh
0JpDASDiVVOfUvHfet588emohz89BV2amaEFtwbvsyi9QAXF7tuARfhVF7ABJhQL
qJj6SGzm3cDE/l4fJQ9k61XAgfcPlfxylOSU8uQoicF2OevlaPJyQkvqwAhTzj1S
jlSPe6qhA4tEpyQLYkfdGLrD2LWNk1jG++gKsuc71KChV0ztF87DwJANGq41EKMj
t+vOtXOSyFBR1H/cLTYxRfZ+y4wUEzQ9WtMDXFUfD/6wlSys1o3SqqBV3jz2Defi
AiYoWdNBbfNRlnf7m4QLTyGEnX4fcN8XJorgA+ZcQTnI6HnCKCXMzKJ4Sn/SRaPq
o1az4q5V3+zKL1DtEpWHL8q3mHWc251tYUtqzwkMZ4Va+3Bwqz3dzGx1lDOFX7HV
snRJs/dwXCmTXVXpSFDhyvRwJVCFPXi088ITuvFI1Cq6W7UviFiyLU/vc7iU1jtl
7IJC8Ocr7iqG8kl+lDKQblhU8FuubvDYhoACXRlzOLqvJ4NXYnm20DCEGI6Rc+K8
zAAlbExGMsrYfDZyDLYSIMpoI0kxBnDyjRGS56wVs4HwslOw3XhwJTQXCO0tfbWa
Q0w2VhS2idyhSe6f+EO7fpQ69Hp0bpkMHW98QeRc64fJtcrtIDaJuEreHjOZhcFN
rxrct9S2yQrE+SgOP3z4yDMNCR9dFQshxEuMIjXzfHbPmTzHmqZMy6XWwGh2x+ER
7649j/afLEPadtP8/GZMLyCemoeAJtKiVcAr5OssZohuC9iYaaYF3xPBEr315+3v
kxEaZqg8v0uPY6R0/NtjqTPZOT44HIqpSyc3docTQTV4NtqC+DHp2dk6rpan7WGT
2MVhS2kgoUh19nGHDXYm/y1jG7XjDyOUtDDarY+py8yqbvFzqRllu3r1+zO7+1kk
pXETv28TSUTUJOm58HWG1zK9icldcb8dY63LXi+EtTdtMuE1TnWmPMTY8fNc9mkz
4a/4olayUXRQNWqmJZLte8MrzGYAmJYVuR1bk8XiJBNywEvBi/go+L/24S9W6o0C
IY+FqoPCVYvKVQngkxX4SGLxlbG3XAEssaNVRV24Vf2tQs1G6BGdByVY9TmBoZZc
TnPVdVg7SMQdM9dk+hlpB+hTJv2pOKW8RSphPJeLQtP+JlSj4HY8BVwuuwGajGcf
4RlVa3D42MQoDfQOLjJMenSkHtT5J1b6T+LPXS91F9+tqR0phM5G3yfR0i9VT+/8
r3jlc1qQPZsNNkWOPDosNnedRocIt0nvxUyQX5PavaV+tpvRUgDgtQMbefdj5xG9
0fCiHOvgWDiCMAEu3eabx2xMc1sv/v/p8RrE3JdDi0GY/o3e88wLVGggRRitQlrk
r7UNXLjVq3xNka7b5EsYNz79ooBotqygNQcXjT0AmiYTUvGJLTHWoHSitbPBEbKB
fePXev3NOjkRbqauMF8EBpxLdk1Ne/uwJTH7uZxlRFr1tZPb8K2a67h2oBKEPANW
lO9TRFIW5IaSjtLyerZjdIM0Gjp8W6vMViVGrSwoPvFbgp8hCF6xmDUlCRcPo5zN
jHuuLx8ydldJrgcGnpeECuZpzquk1FihYceotEzY0EwtB3Kc2c6ViyKlJqpc0wWT
/cl1fQ1q7wLXnDYAms+ZQXWcbdwPErXKgRR6o1gBRuNOJlNaob2RR608AZdwuVMa
NyX821D8T2oVEgfR0jJ2gipHuxBgoVXahg4sDf03x2h5GDb15ALaZuloBVR7ns8Z
6cXd+5x4AzjTYsqkmJLANB56giatS6HAKJDG/2GOvr0uu9J/2qvaDqjQQgHwz2Bm
sDrZxxeCZgnPMbryW0MHerJ43QknfDJEf+FbESZkRYXbno7/r36q5+fSeXxrW93k
A60XqId6n8oI15aXCT481wweHq21UH2t446pItRXnMV+B8nwNtxI5oYt3OOaBMFL
fgTxW0o1nUix7ff0e/AayZz6m7RsA6ZYeBHySTD6g1ZrtDGF7gAds2il+NH1jsa3
ISKtMwKiIDFru0uMQQrAMoX9CBUzwf5Wv6ivXTZZwEJvEW0goySituHtK5h9DHFm
z/maqoVvPfcUyYz/x25nJ4UKRo58W6af/eImvws8ah3nrAplhoGAwwAqadQ0ZpGC
irHQM2H0gA5mQuJd2wpKUXYRsK9gSc14ujUAwROxapbrCDZ7s2+4wTgdH2A4ceoy
DKuS97RDrsrWVCmXYUa+4y8GiQSfeRXjFy+JPU9UUYjAODNYM+mv2ZTLJdMck+aO
qVeUbfArvrtbTu7ySkyOBOTYhFU2asoDaY9GjMv0iZx4M/mLEBma0GdT3HkOcU0A
DVZnnDNC7W4O8c2X/SjeQgyplmW9mT2QrbdFmcdNykS2MgZQHzG7pKxls4HBZFBI
nJc32n8BYfEgSuz79MWFmQpJGgwGA1RyYfF9Y2t6aMiU7dECwsqf4idaphpviWap
a1nPWAk5fsAyHE259k1cst3SztfC8u1Pqh4kHNmeQTxs4f/Efcvpti2WPWuzA1Qd
pWnEuoCJem4Pi5mpR/AjSDR4u0Bs2uL+ALbSlbQSa/NmO96cTlhQJliIyxgMSWjo
yoNTaEGfUKCNt1uk9/acRPdcoSSTDjf28zj6U1yUhjj1wjPSfMlHiuV2TjQkVsV0
FzgaCpj1op2XLhIThwtYl6ffZRHRwNdj5phOw+1IJQUShCC398UV2XolSdtSGJTI
ms182ar4nc/iJBKvvjBN/UJynWq0aXR1ru3Puxa4oafGXWjptomBWOUVL2o5A/X6
JnWyQOyczAUfMN0H8b5EpNdtHXb8lT7hE9m0ZfbdhWafywD7VAOmVWoB1aUTYw9O
jTSSCmPE5vt05Oy91jPnwX0NAjXhp57gaXLCWsn4UgDCW08lkUkbfmEmPTIjR7Uf
4EX0wm/6OvsHI3vbMWmPEKmGpfjO1akmGGJ2V+MjQPTA6h+Kk8PXW27/pU2KacZo
WoglqywUGhKzigWTdNLFpCHzQOLOSxBIjwCi3PGpQVND4lGKa/tvkXV0kht+v7Jz
VT1+tuS519B7nsLcl/toWxV6nNiLdjq/1b79fbN1SCIZthudr4P694bglvObVPl9
BlGK4CSonaS8NJ0PTd0u0vsScUEm4KryJEeGkTdk4pEZPa8C0PaS/hbL36zdsAH4
UP7Z1l2fPCd35PF8PlgPam140Tabl0TVZ4QQeOahtjlA5DKdOl0wl3WX0Co5J8EC
8bw4nwyyVXTIM2jM2dx4oXude31fM0gw5lF7h58Qx8Zd/ucDxgOYRhAH0x3QwByR
yAiVlucBoDphmxFY8XVE8JjIL5/1cLSy9lt5mAYMF+avA06rGIeCVVTtvZWnBD/7
uB3bVnlWO9W0W/0k+Wn6oPrp+sZhcUHJQ6BCsqzOoiwtw4lEmYhLV5dD9PAwFFj2
9z1TQZt2hERE/6zeqLKF2ZuHw+7wwYIrR6yMSssX7cUOo33PKvHCITgk8riRa3/l
x/UgMrx2/nw5VE0KaD60Dv7kLZExa/unDcaISi8a/vf6rJTAAXMgSIgr8i08XICH
mF4M60iZhG0Ldt2/R1yvIzIG/ENP7ECK2kfAL2/pyCjy/CAFVsW8YcmCyOrvJzNV
42Qj4au9WSgpweMFSOc6tnPy1E1YnlD3tUVQS2PapAgrxTh9qfIHIn6cTgut9cay
wjo34WC4F0Z086472aCqGgZYH0oZC8wU44AfVWzEH3xdFfngrwDgogjPCFOVegqo
3iaeHAZFeURWs+5U9h9lOl00iWi8EB5q/DLajFtjAZ19xTlL36oKNDp0BTcXilYd
rLQPw2ldUcFJ2pXgpU1YesJqm3fNm2bDZTC26FkeayTDNW7N6skEwOMEjId/QYPk
EmAxvODaeHbjPwtpq0YT22an9k+2Q07BGjmLq4B/uLIqGmzSevE3WiznBru4y13n
jPn8OVDMACPCIRzgdARAPba6y7Vm9sPRo0CgYHlLEMb2Pb+yNalEADtWL4Db7hfD
pJpyAh+ykD14o8mMBXeI2xGhC+vsYECm0iN00h4gqIJVz9McG7M7Y6AW3ob/O72I
2jUrYw7vstY+Vf2zcObeBLYrtDMKq61fvbOE/n2AKBF8BunW5p1+bjSg572HKdex
v/PG2ercUuSmwa8MGypCuKJ3bnDCKDmnoYL5rnH4niM2JC/8zqRm6Aner+3MoQpu
pOSxIe8kUcIp2Ug1w5W6EwTUDr64gyPY13+K4RDAwImOm6qMP7f++T3LgmECb5O/
CGrkxOxc75ufZV+/I5m2xVmRUgnHGwUQYKGkeBBNJ/snpYgO7v5qQK2die1pkAhC
1FT5m3zaEfbOdT4+KVsz0UVnX0+FUB1HkUxoegP17yXxWGYXqSVzRaVLXRPWTIys
2PuiAvhqZhy2jJW2dGmXuOYC6kOf9+3NOytfkM1D4cioli7+laGjUyOUtVIRYRJn
6hZ5MHN3kXeBYRbuFNNWTqpNjQ9sT8PApRHHRIDh3eEABHMGbQO4F3yapHAjc9XH
ifRjRZbOEs+1T8tTO5GO7Cc4CgKW3Cf6DN1CDJNKK90uXEMmYTEIeq5o1A4bL1t2
RRVJjG51HeOojGCgAa6ThwDxYrMbbeYkkoYZdq1T9OYZ4qgnz0Qxk2Awl++I9W6g
szgn7waNxvg2S5FTQKDVmHy1WBbe/2a4FjXpom0HLfykoPDsTbBp6fScHMu864BD
DufrUypGYXXQ2AUTjXlNPV1JWjXwpC+q0JemdPDno77Vj2xYQF9kuTq0gUu1+U8A
h2CZ76yE+ekBn1TpIusZvlbEG2DW5+vzZk/oZ+p2mmNWkZVeKfoY1JCKcbqgQCzN
xJm2XSMFsAHpTZfu51RY5ihJJl2Wz/F10OZHpAcCjnIdYYEvOPdvWw8erx7G6iGC
qDTRYZMR2GFMu9sr5W7EF6ecQLszLKleoFrqmDKZEEt0JGdDHrkSHrmBnQu3jsrs
2Ytep+Blgz3/HVViV7ogsd5AshZuuSjGLWF9KFZG0fdM8i1wqgLAdUBq6h47iaiE
wdkuYCZnaOKpjPoOod7WTZzYbu4h9LcabyPssP/6gWTzyBqVEZZv4kNVV3gvkf8c
5g+yxHe4eAClzNGXJjlkPK4/SnW8A5Lda2dDGVm6pxGnrGb+uK/dvZZPkGFk3RDR
bBAw8NscZ4YiIoL3ajooYp8myNXt+7DvfzTd7V2XuhjVzAFGHY4V8dNYkRluLDj9
vhULKkeMGm9QLXttbG5b0UaIP4f+F7az/IwDxJNNizn24XRJ6Rj4BzvIcBBC/PNm
ba7LY9KcuXqHCLR1+PTi1v1bGR26BYC7cR5ICncrt0Lwx39bAmnRztX23uOUTGCm
UH4D0zhs7FP410OR0hYXCcZpHMzEFBONR2dfrSOLGpF4CxOta+RrD2k90BjNBF9q
55yZ7FmbCmXKM+hMnV8bDO/lpl3ky2x77/myM/zLLH6ZSqxwFoC+KmfoQE7mZQkQ
joirjVAKpL+HfhbfqZaaPSpZDKjTdP4au8KZe3MEG9XarPERXs74GtqAsoO3nONw
h2//J9S37h//T1KNxI8yc/QFRRyPWHZCKexWi4u7zeqlUAtariJiUkdZo17xDK0z
5Dx5Y3jaKzP29Ith8l3cebBHueOd3OIUGbM/nLeUfs7b3Rt5ClsO0Ot/1EPefxG3
7y7fOjvTKKn2cOl0m+yM0gX4FZVd0r/RN7duL/0rJFJPptNN5ZU/DkAHgmUZZJHk
RmRHARWNraFExCLr8E8ZZCfEoIkAF9O90NCxfrYA+PG/YBVdvQp9N8iPflHEFgKM
RgUYQdTYlAkBOlZVWfEwtyp1jesJPh14IKcx8CRr6ndpdDSV9Dxbqpmrau0vdNsP
by2OMniIXA57vAgEmAg2SufTWXGFOoKMFpqRBCKDaiobtJ38uLMCvzNZ6rhU5l3r
KNGoDwPZVJryU9tpLeWWgT3KTefnYsmY6LziZ3WRl+0KmyHZP9huoN/e6J8DMy3L
UsKV1D+1RjBsHbzGZB1efmxAZ5kKP2Q6pZDvTbK//LJp5vc8ejNpA9dvTalcA+Cc
AN3KfiQR+bXiHXzVTjZbVCuvcHSwGj4GiGp2B0pCjWYtCw+NUO72abkBz2SQ2wNW
D3Pls2Lmd93Fv4EcD/JNpNFHNT0jbmqkuQEJ777ECnRuzu+RaNSVSVFTbTcW48Ku
fUF2UTNkL6UiDRc2M5lqBfCEZH0Ax+MxIYErEF+DJ0a5vXvjZ5HSZkF/6agp60Ge
dvsYij6IgH4WtkP6kjpDuC/1pfzbbjlT3NDJC/C0BLhIpyKFhMINvp4L2s324C4q
9ByJbnF30ktA26QgLoWjmgL9lpZP21b3Y1KemmuMl+MutpV9BlDVOSsWnvbK45PA
lEhVBDGHKobhYckF8WvJNJUVrMYnvf9kg88/zbj06kWOrs+6/L7i9HZZ3KDoUH8h
WXv1lFdpZFrEJmSU+VAoRWDdDCQxmVNGbOO4ZHHpBVLBbdgxxaioDAaolvEk8knD
MBQi+VJYMBh+IppYN7xikJwHrGlAZoA3fdXtpUOErpbIwOUOpN8rAthhVJ9jTCcF
6icaQKv3jZNXhFs3cPLIUIK76dfeef8fJTkj5YBPCc5/NyzYvO6EHrKjHyM43JwK
y0X/F0mzbD1t8gY7vFVhO0LzhvLowqwa1u/QTSrjwPkvHdqp0JAE2gZmQhc8GwSl
huNrYsTJM2pZV6zRbrrhmfiYEQwh3C8bVPXcSo3r0jA6eZuxQ7FUcuOzrndyeJu6
3bBYGpHwi++i6i59RtozOdt9cCt+dUWEzx7puzADjvXBHuWJxisOFheZ2SeaqD5w
X9IN7axQlVxdlVSZLs89mJZMFvIZKXyacTY0OV3CFdqlxqgbWp0VF2zqXnYXPfxp
S0SEcuemGCzgpn2zE2zxwAJkceIRQLK+VbCe7j8nFjgiOw0Mj59zWO4Wn9qz75FH
TJpEYQjLH8Ogj8kbxSbAUsnPI4aYkb5KSOlPX9ig/ni7AMMYWgPrFKsaNiDq1AF3
G3v95R6zNU36z+YLV1YYeQ5+LIKU/oL4GN2ue3BEHiUaNEk380468W2eIT/miWXY
KxpC8x+KusyxEiC/sMK12DU+D02yei6dUdzZ1a1Y1wWVgD1pQp3I3knbrI4lvJy0
UIvrQmV4VNOoDA8vFbYKOL/QcckYGGNa6DuMYgW7FwYa6kqQtzGoSEE/JOfW/SXK
e5CLIJUsIvMbuS4DwgUMoqZ80cbutfEm0ZBmVepVtWcIyGCqEUWEch6JOEr890pv
ZP7dMm/2CFhmuldDuNcJ3ySdSvK6xWFjbhHPA5fYkbYrbhduVoSk7CClQlWXRxOc
4XIb3VXV5ASxCGNzzD07CzpoXXhdxbAjGyG2j5BfE647j0+w1RFjUKZH0gjSNbe1
M4tuVxBiP/q3xMbwBTFVYlJv4ocUylVpcEQM8xYz7XnCNuP4Xwq67wLp+thfiraa
JdxasS0DvCt/uKx47RiskES4RAOBDsS9YgL1C6f1ZY1zBWizxlPx4+p6EQfLEuj9
H0YJmhJqHIfIqwGxT9kYyvE/rSS+H+EXm7DgSfZHwt0BQF4cXjii4DQX+8GlxGx2
Me3v5I5Sx0g40lQyquvK8es9HK9WA/PyqM6vYBiYLNsmwY936ESTYwr9tybIC59Z
rB5lQCFw6eRtbHd3lmOUUrUKWQvkypcMfqmTMFms+rvZnNl5ec7AAfG6tlqCKrup
Grce7xvw6czUQLWI3vfbdEU6mGkx3j5C+iqNskibvOD5wSht2RS/uuqPa5tanX00
Sj8aTUGxZGvF3zBzzD6DCv/hJ+WAUqQMG3L0NZs4eWM8zL464OVAUgPC9rnmqUIe
QnqCdRpzYdTPYmiXDwzbV6d69lSMEosIEkflKuN9au2kbbgoBgC78/NhGX1Mw3CV
gEZQXKWSbbDsydqAs4Bdpu1KER2rvbKHGe8RvTU8+9Cd6oDK5ICLh7ILWrAfRyL8
BFwygV+xsitQmeGMpGYfjgDI3fRgiVwq1cut/11gbQQlDr1XPAiFvWJ9Y/XSRAuC
M7061hsGvbTEmwgg1D1xZqwzBjvWF/aMFo8hDl3A28MHJHFvHZ0i4T6LwS2B45vn
CCdDinYFB2GldGFa1gFMk/JBHhTBlpmDBF3qxHBW9U+PFyoJogmZNB/wdpsYD6kC
gfBhU2j9Jn8rr5hBhSFb2pWnY9vynTL8INWmMlKSGwOX+aP+rpJ3PRkRc6wPoIE8
qbQf6jlA8s5rdP2m+yec8S6ni7vRFiWug8yzkFQ+9crvcrw0Y/BQaY0P/in7ZFQX
ViMma8/4aN+SYrqzstCC2XKWE/r35fFc0yRKqEVRN9GXUKgcLphsTFsn+25nTIZZ
+sYuSmmGV1cpq7YK/zV75DpVocAg5hElvV3jCbrIcIcDW3d1MBa4yQardzrO4KNr
+xZtgiHuxFcLWJkl2Xk92P2KzjMkmZsHFY74EhZ1YGacU/pCh0SLyMtLpW4KOrde
0PQUkoORsbmepKfWlnnBio8qjHp90oo/DULSsd//1G+2I4IymXSv0iOdmiWQWjHW
8Mlv0/lO5c6zslYpI8OKu9mJNV1CNUfgT7i5JRr+4bWwKy9qmhaEKGufVaGIamF7
J/+YGUylPRnaTGAE2ZeN69KbdI9CpBBLDm/XdQcyMa9IyTWt0iCCVCN5M6vUQcpN
VCfoZLwCH0AbBOAP5mbMUMgJOv5+IRo3tSIPu2DohVeRSAA2CN7V2A2MZ2+mjVKc
ruzgqsgmVb6W8RWvCl+EzA0eXBBZk5DwVzMkgwmI6wQQV5MgpwlfCa2CNXnebxcg
QngKvSIbuSzsebrQrOC+hjddaYwv2NXh2d8pjaNlCn0z6fPASyZyGpgC4BwQqefw
Vijqtq3y8VAWXjL5K2GIuFB2Nsr789d2c0uDftMcJ5+Q/OpTX30IcBkRhlkPCpO5
zejuBifF+vx5J4uunOFCd1+zmxZc0TmWQ6Byd6sEpypGi/3HEPVhm/8LNqYb3uDY
2P4eRy+ETljVUUPCdv09Fw9sRuW/OqrDoU8pdeEF5LFA/ocPpiXT5cvaXtHK3qAX
nA3zIuLpTbjpIjsEcLKMGmwbyD1SzguR/4RG0nKKRMCJUcPH0RMCiDzmyVSUfJfL
hAmajiGlLM7bQTmxH943UkUpZ2eBenBtwsl1zR/rMKo6InsLhAXQlHVtG5sn2cWw
p9Ing4fJ2NjOQynGgisTEZ4iGiT4VP0gy6jvnliJm5p8puc7IqBqQ3JzU6d8W42G
BOBACVjwfLoh9NFgeHgIKfPCB+rRERA/fpV7PmUt46mrapIofwn8v6JGMiaeDjHi
yw4bJbfxGNBt80Dq97uNnTMMVYtptUt89Hgi+jwL6caEEtnt5B7PdCS39sJi07St
NMUMt9EMUlQUrFmJpXmnU+zbZFfjpbYZhzW73YyADUn8hq+/Eei/ilrajXOEjlLB
aQpp3LwxEKoBKwlG5J5g8wfOrcHAzaC7Ofr+UTUq+gfzAX1sccUHCQIg+fwbivKd
R7eieWacZnySY+rkAp+sq8d7HV7kQ8Vm71cBfOChKiJUozRsyZWdWGzSOOi6ejlV
deEyPUvWv6SEKy9lPv6z+t99CMzVFMICuKAeydzJZd/1+CZUutkXvjuZh/2SxybW
WRczDqGwHlq45xQ4FLLllmEwAc820ya+V3w9POotY5OyF5C+rCEVkN4Sz+t+zf/D
UmN7XViD7HxbnuyUwE5PnY1MCpdKI1EtBoXKKPHLDSSbjvIXFwJnTbmMMMHGJo9M
H8BRr0QjVlPjAvmLRCj6K6hFmMm8krhss27LaGbEmvSA6XaOAoE+EyUgjVA6I3vU
LkjZllBrO/Vvkvu/GIFL1JjU9g6KB4U1j7aO+cGYMGMlciQhWc+1A5iPyZZXFE5S
E55uAU2gh80OY6XS5papzg6l/TH0rViNfB8fnCI9fVGrAJS7Qbjde/mqIT979iiI
y/M+E+vuh0Stw8lLEJp/vd0HOIhb6BuJcJBPvK/wYw8+KbcenVgEVSqovRywnRFO
4Uuv4QIZnrAJUS4Cv2gPFDk+lgKBK0MCaNT6nWnruYlboxieP33ADCcZIUmej/kd
w0LgcN5H+6WuBI7DwKEKb4678popkzXhEgXNveq9Aa4T3vtQUazwjhaWOiHhMyNo
iqui23fj6YUBQq1wE7W0sF0XJuxuj8zYsnHOwt2IMNmgYtkaPWoW6aMhmg/RRbFk
ePOBRvrp04W+4kujXI3Vh3vAVuIhyuWesJHm+fcWnUX4AHvI2Z1/yZBpL6rlBCLk
eauso2oc3gAcxttkirH0Wbxo8kT8QXXjE4mWTkv3WBcI0LwSOVOa3Ecy7LAMGE+B
rkGS1jITcqm3GDFf+PRya1o0uSyuMFFwCHxUZq2F2pIGgAhHo/V7AECMwSOgK3kj
xialKX+GoU+st79gAg6Zv0sfywauTPLHM6EDL1KHKDpfbnbJ8oYukgbdeLOupDBy
QyFWQk4nV4lRIcuKBDf2iwWMswxlNmdEclaRxgyoY5iLx6OxcUCHXcP/4rtBUyyI
QrvEA+Y5VlCq1epi7Kz98S8O4ERqhsi1gsZDBiItmeQprI1KYiv0lshf64zCDlI/
pTfN4ry4dJUA5TU5xi63kfv5Bn+Uqt4J/lPveHSe1Ft6tklgVyXvzkhSTZzv41zP
HyOh1XTL93UEskwjIy6l4T4wvjjT1p9EVIDLjf6N5MsSH59aZV369E0Wi91yPC3m
hRYUTlLYxWjfu7Po/3HZci+iL5BBxe3bdfYLbjUYLrjuFPGvainemgaLuqd9gAg7
MT5UKQfZbRvgosip7mf2CeBpA0tRv1ZEu0MZSMqkmlTj+tqBCaa5kP9cqfqED7NF
MSAxrPcxm7epbxKjhcNwP/Nsxe7+vpNLNB5EZqk2Eqz2Zcpb3rcA11rgZjyx9Alw
ZXLc0ULkOLRxkDeWgcdIuibYaHNT79USTxv8LJpdvIZkY1mHsTaXFRHW7bD8E4X8
Q00lrL5U/Ewu4BLUcbhx8qkAJ16e32sN9jOG2zJnI27KOS1MpXfKcnFaTCcZqjUB
FGWb1gg4N29mQyjbXhzm2ejVdWDVduuIy9iTYpsEfZOW4JVoNf22ax6C6x9J/oXY
uZ3rLy4ZINFDHv6kYr9/vZGJeLWjUQpexIlmRiTflbgkl3904NmY8zOVDmZ+EJdg
o0CduFXWYdB0mSexBHMKPVeEZoqs1KXrvlkUvZ1oXU3l67JdToGbQDXWBNOQ8ukv
FZGtPJRUVfFgubVmk1YfZo9aJAFk+YOOrFP/rB6Lzar++2yHAJVzznHNkLzx9jwa
2mqXvITRwWXLMk5OPNl/4yp4dUmHjRh9q1c+ISmHZDWfnYKBPLx1WKPvGriHs2IS
zluY9PC/qyXipOqzoVhH8X19RWGs5yWyHe72fcMRwmH5QwM0DTfFQRhkikJTt979
bnkU/jdP+jtstr4GUCWw1aOmIFr/5DbuAss7pplfwFEd/d75h2LaTNvmJOCocNMB
34Nes5I6lde1iLyjT+/HeDqM8+CgT3JG+TNN18oEKvMa64dWoNzvNQy2k5R9sH9Q
CKHHZhMVmZr6h0poBX9Kb3TrKPU+dOOSvPgitAx6mb1R1MSJQrwLrjNbSfHkRV56
5LvDa5UrjijbbyemKmfeoCnZgueB1F6TqNDJh3Sx/LMHKoy5mECohcueGg7ou7xU
atxe/vm3lh1bl4Ty3pjuRyRHalDjSAL9ydUGMq84Utn0XW6RJ99CW9oUXGnDQ73J
xT/Nz7XXSMMJBvLN7lawU49WYu5ypxCrQISMpfzw0xEfda2CuACkITkgfsGAC82S
Xuusn9auQwWhct/kgIt1BkxO/R/Us6BfWBzg3pgFGE8XFxyBSRDZ/VzoiHqaAWhl
d55NMF0NySIdHJjN6fKgUvKvJidV6yq6UPtck0bp/5l0gzTl7kvNgLT3Ea/z7pBp
QIYhhbfMOc3ArP/94NueyD3iKifE+LL5g+YAShBwN0b8S/B6cAo1XSRa5+vUnx5U
Ld88T23rC5W7sgl/L6Qz44vVJDpzIYlutt4YfqCHrT2YztEn4EkrBtuAsK/zGoRs
Nk8KSlBdl569dY5vMaU1ImcQRvSV9Toky5POreioI9eqGVmHVsGrCxEpaW19sfyi
qyZSsYFUBigHlQ0HW4IzzPGKFsXKXz/kbbFEaDBhzz29Bt+GiblHjLzVSB5UPNzd
VKWFPYySCOaxvSSYUrNkeba8Rlz+TCRt0ITJHC8jBqy/baAUODH5fFeuiigvdPfB
ydGzBo+A6S9EuDcUjfGuJ0vPxLrd1b03IOAtLuk0plb3lBgDu0NNzOzqvTvCP5TB
kke7KtMvvL0Ie+xShpScqrjJRLXh0s/6+0UHuHvKy1JCATzCWah2uaOSLkJXCp6K
9jNqdKdhPzgB6HI7Ao0iYXa6eFzo3cjiqkB1xLP5QT3BG07UP+tXqn6byu2EG3LE
geeYdANEyklNAqnlecOeXnKPqUNvyIQ0h4PM8N3SRVtkrsE6ZK5sTSJv/922+JCt
NYzlPqYAx9SqRA+GzarHycfcrxG3KJebZoAyEF8wuLu8QEowvD86foQtVwiSjT6X
fLUdlUn2/6aLorteCCuvi2GlISdYadE09rye/6KNHkN08GxHzpAg9UGtnYNkY72d
Fr31Um6PhEpwbbtRFJCZYElAjA2aSQWW0HQDJnwyvYSEXmXK/QPDMee2TgpPenM1
VEss8/Ecn1jUzQ2/jb4m1R2eSVsDysWSFBMz82E+4l/r20gSPTmnQE4yKQEy66A5
XObYp5Gswxl4qX6TkAvXZedigl6VoFMzxi7iCHTB1DfciPCmGXO1FkCXzMJ3fFgG
FBdL91j2e1ccHSEiv7AEbsmoXFmgSE8A5qhQd3kb5A3fLsOc+UGGZExPO4JkSUZP
nx4rn8/kHhHcnvGhGh+n6bJbtl4ZIf2NkwIGpVOyrtdMUX14Q2xFFAZSNpIko9Ek
NMyC4jMaLXOrcNfd4MtMrEOVKWWGBF2KOClUNbUni3KqF3G7SOSCUJ0xsh++IejW
crPmD1q0kSnC8Gv4+wUtjMgoAznN3mYUXANneeMIwFdMWk0LDbgyeL78B69mF1Ky
DVofFsQx3U1EhxweJvG11VJCMOOZGEu5L8SQ0O/LUbcT+Lu52FWLT1FKLXAKdRwn
ZHDopYkRiDwPEKGvgtzgR7hvnaVmbslW/Q7aGDf1ZTpnoMCaZtCANn7Q6QSdzKuj
52AE3NVxm34yQ0PXmOHyfrPl5AR3sVnwHw1jEQqw46Bx4z0ldsSYLLKNReZ3vpU0
kfHVCmm/dMkztBIeffYEBa0oGBQXD905eq+LoQklLaerEk8jRgfrFXPwyzVbiPt4
X5ik/0YBf40jTOKizY1iIp2JetXcs2x+pMAC0NKuAqxbLbZ+m07nYe1gSvl4lG05
y7I4DR2Jb4FQAL8E3PYPxyNSLvwETl8/52vev2QngEwh3wWrqoKyFlcWLdXdnuNj
sGkh9XENA7X8Q6ryj2S6cmqSubinVy6FatmLinBqpaHywkGllYkRXia+n1lA2yPT
uOCdgYxzlApYNN9e0KFz4WIOc99SCZkG45jfSFnYnM8sZMooelcO710P+CaMMKNQ
DixyqFuqsJfefW7EpaxkBQhu5RsJk/rhHizSpB301ow4g8m8ClJviw/pPCBv/SMr
0+JqMV1Iaas4CJ2rXKVUPeN4te5X814flm8LmD6/HHaCw0BHni3B3MfyOmmOHJJ0
6E0COc48YGjE48dFf9Yn/Nj3RDrwN02dU682xiXEPKzZH5h8/saQV808neB8CtlA
XW91hcMeUGo+Wp40aVIu3rPi7Zck76i0xxW/pz+6UzKfzB+WWIUjytQ8KZuEZe19
N2e8kO5yHv+LVGzQuTWcCptyd0nItGxeZ7wNVylm4Fazo/kZrbpYk4VOHipnVgJ4
3xda2dDoYrrsLifDJ4gtT2jl4bIjq0Cdef6qVxo6FTgXZy0OYNNoUtpnGQo7XKnO
l2ZezLiXGQ4/aAJtzWePICxTh1rivxknbZkbRwBfYBcFtwI6zbgv2m2WwjtK+8g0
qGp2meYd6iaGg3N2nVO7mLSnzIlpYGKyEsiY8tTa9UOiVvwJkRcnIBsaE5ZYkKmg
lRzpe+4PXsfujWXi1mt4PUiEo0PTmXXq3JoVs2PMusSbPElgWamKxekxogZTo4Dw
TX5keh0f8SVtUIk39+6Y513Zr5sDbTfVi4ZfafjmFC1TNHvJtDxRm/xKusv5u+Ly
ZvkBD3sFHD31Gdo0dKKaCPua2A/8XMhJ/azhgO5Dw8+YCXZl1SFeVcraf6gPkNbc
phDsfmFLEFkp/5fcoJ6bTjk5TLRIWhKNG5AT1Xs9rZp4vJ0i2Fb2K91u62qWJJf8
wED3VqcaOpWceggKRJtlK1JofFQjx48HEKzfZpZrkTbPBpvkqss2m3jHiReZQxYK
rv4WfcuaXMWhpHG0yBSs5kvZfa18JzfLotFx9FJaXOJZHqzk77mjWSO3xv0gSwe8
CT8Wn5d2s5AaNQv4ldRhNiUN+LnaUx9nlqirmO49XmTDjUyrffXByefVTbXaKHOr
nv4wAHsSVkh5IOcXxqb4lFFZwe7iCr4BuzsV/zcpe5UaztgQVEoEfWBC8Og13tI6
eSn8CGX0FTd9L1ao4O93npPBuJNld20gAHuLS+Hcj+bTXvV6RyBO36pwjyx1Xjgv
Wo2f7kB/oPwYSSMCplfvB+V0bUsC4n/CxLonuc863rsw7MTAUSoSd07sCFaEYGL+
FTSy0yZ27S+12GS1Xvq+r6xajnytmMlXbeQ/tXZeofjiSVZPb1F8wur+x+kabb64
RmvKa8UYXbpjtiC8oD9A0ZlSpNXVI26cZiFR/QoKAjCyGDwr6sBol+SvhajSKnNS
zyScfS/j55VZWCbh2CMwINpEZFfSRBgYQcNJBPGqbERu8d6GsAp55Kmu3S1cXRJ7
iOEVMCKkTBGTsx/tCY1VCapv2xh6KtP6N3BUAQjhCt5uwaWn6uphyzhiZbxy9ndn
IwCzLZl9Dpr0LI0R2ZVSgfZNud1+CnTdlBWVQ/b2C5i6Ys/xq24qh4Lo0MBWeK69
eq6FV92lsO5U5YZjmQyIe+meA+bSp0uRaelnDEdsuF/b6e2MTjONAUcBGOOD7Z1y
YIWCC2CaFxgdRz2KY2S4qed5nNkuuZthSzdWGOc2CKPTwgvYgULN2tT4f/VSrPaQ
LQRkRJqEouh8mrKaujMfi6LQckouep3dgYC6JtUcBdETFuJT2KK/+ofSTyKU2FES
TCNrdul27aNlAsFefNVwgTtHZQbyqKDqBOC4kXvdeOLR76YkohjxPYX6YKb4byBk
0noZqEYLtODvJZwnE0HVUOkFIfw0PUxCvOvs+NvtzdsV2P4dBgL+6ZPSoktOkm7K
/Pbds7LDbcS1z0bKHx4HCWUTegzhn72HaRrIaulYhvQ6JcIaOJR8rcyu7lPh+p21
3W1W1NHyREtdbCgzXbLKcaP2JRlGhK3XJnQkk8s6nM44QfVM+stRClHvTIWpilWC
pXLl6oOfaGkZF/M06Yw0g0mGvjVQpAqUduHoXtdrAkjQ46QicRGPymcD3H09yIQy
cegF4ZLE/tYqd3FhAGEnl+g4GqD2MvvKUsFp+vgRjT3vUxDxjehjWPcrFz8HZe/X
8Lr6fuZf2EK0Rh3JOmMeXNDzf+FoEkJy9+WoEHcFAK1AF3HGp95lwX2W2EDQzsmS
xIIlzO42dkpW6n1xSTPCkaCB0XiGIockZd8VBTn3XF+d3JK919I+sfxMI1PtuDBY
Mga9/OV2n8mY2GqAqYL+7CTE6cXc7xjOKBQ9HmMiPsd0iKbuaKr+MIHj2mVKEnrb
8Qt6SaHmQ+Vj1T8BDzCIa9eZteinQzx16yRlKfs7HLALhmYm31GWoNup7rpEE5Ip
4OmPGD6er9oIxqgqg5hZT3PQ3lsSZv2NRDSWcuzl8PfaXE56DLGWVvcbDzcLn83H
VA3+Z4kNJN34pypaD+5+/A7FRgNVOvW6lpPk9P3UdkVWQYxq3163JU5gtkdQjdYW
Ae7c2QpNSyvhf+V2wnz6IIcCCdqBh5dp+YGFeCXZEdI5OcPe9VXOwtvPMPQ9OuFR
yN+E4Qq9mu40ffqkj8+1SVLGTfL0kgfre+mfpsBJ4qpgUWCJSKQiqEej77UB6ZMW
ex/mZo8ebcPNw18NRvQTx+PfsecPCqKss2MiuUvIF6dX89y+X5ht7phykMJQU203
W4FZ3OOgDNpKsNn8zFabjPnFzNXQ+S7dozCXncrjl6I+zzK+++EY5gA05mGSO1K0
At6AkPlDA1iuC8PsSLkav0NxwENAVeauBV531u0HL8FKvQNJYcVkEAmqaKVVeNUf
y2WhCseFjOKflDQ8IBPVXwCcu/ArwEre1sYK5f8lC9pMEO5TnOAlPrEGM/zsOhXr
rR5uLr0+f+/cCNtaT6hJdD5HNy+U01vI931V0AamKKJfIvQtgyCyeUSR8OhFCWhi
tPpvNOKerEazr0cDdCy16uTF5h4/xc2JzMbJyxn32lRL3DVdX8YNqqwfvB6YAdBI
xWORau7xJOmSAjXT2MnIZCb6OtPh8S3PPXTyCJd/FYc0tSsU5hUt3YlbIqmEeP/+
JHhpcoHid4G7VgyflrmP1gxoGpHfBv/VtGBi0+/wVP331mW1EfMATu9qwpUsyaPV
oi2rXCXEMU4uAAhkGwIPlVXGXIX/XE92U6Lxa0h6sEDDY37JN7cKMREqGWJa4zgV
I0tRndGsmAlPmImfhYQP1o33eVreH5MxCfBfdK1qn8ZxM+R3TJ/MviFDhSEgu4Q6
v3bGdId7Vn99Ycu4bc5HDPeJr4tFldiFr975lXN+BImLHCrrnRBqMjoG3Df1nM4s
QzWvBpn5Rxl2wDShX5UaRz2UJyFibuOZ8/rdSmCmOYRUg0ERR5/QRTWJQkkFLw5h
S1V5dCeEWNqGIr0YODIJkaJYdTEVZr6G4f5rsUHo2NNXsCU2Ei8Sn7eo+2wq4WC+
QENGvjx9l/7FYBgHicTUbekmHcB0EgEx/QJX2SizQ5ivH5O+vC3J0Ixz61bTs2xL
DqFAW//7HVEIAYHep1wvkV9YzjiYGPe58LxrxAln5VMhxiQaO9GTByBXNDAeMHrH
TmOXhQ2tlvNytnP6jf2PzS5Iwj4pB3F0r/XpGJA+Wb5qAr/J9SEQK7T6Qzz1OCcF
GuBJU7EgdTwgsNlkORXc89oNCeRvVGLCe4RynnFLa6+77y6TGNY0h/9ANyhBEuun
bpjtI1wNfcYbRJk/72TFIPwqIn7l0Izh6XENPRMvtXRPN1acothDJUaoiAcKEiFc
evULpVACTjqvMFGh8QMSsuUVE9T2vMYuSwxS0NQ9hsclv/fAMYzKf40qeJZ88pfE
nEp6aZ1+ygydjoJ5nioeyjQHGPkyr0Vt56ES8u8s1hVemXymYK4BaRrknmuDhlrT
uImPUwcVlJkKX9lKIAg3IfdTj36AfmpUJmTSy/hqTy8vmOAJJs7cxYB4L476QrTX
LCHFTI1LAHXrWRfih3Mt5/uWyCtJdJWMBzBxN5H+k6DnndWPtrBHQHFUWs4c2cpf
/IBi87T935dxc9iDvIwNaGKldiiBLhJ5aOdvgCDpF5h3pMx+G9FSLOhV9VSAKA8S
ZdmEMmVk9P+GkOGJTJvg2Zjw97jTVEiwlct60cTOdThPZwtXQg93yYgPW8vR22W0
se73dim5g8KQFbRMxAOeNvQ/2pSvBlvTUHMA8n14ZP7+Elfotw+BeIL0bAems12L
GLtvpjCUw6eLtD574DIyG9i8kw6wB7yo9PlX8SjoUesUICM1E8LDpvUo8+DWFK28
92N7KGutR5tCdXzqwYBBDAyDcLvF25ms8XvT2Y3F0l/itKaa6VIPgfO16tDzl+pb
IigWV6sQRvqvmQJ7uxmUVcRkngJ5MQ7weeWbM0oRxdrc1AdKOHM345ZSAIjgIHwY
GwjS1RIIECLZhn0xZ8oBbfQG0e0kdKa2K2hOOHdTeAniSBl36NbPg4z2RwPzcsXF
b88+YeSzIykz/HkuuJec6RjqgbiCYXVKbJNxVMrsEu8PmxgZ3vQKDdtHuRsU9Vt2
/JYjLXuwoUG+RzRjXECDGAgl5vDk68Ejdfq/75iqE49y7AWE1sqVfwlkr5bEwTTG
jOxd0c0pI2tE6/cgaIyFL+HzXRKut5NxLeqJycT2ahwy0eeAsWtH36Xd9OOHjhje
+pqNyXFq7mxbyxLHquwfr3uM2smsVWIZ8NqwPZeQXJCoEqL/MDMRPzl192qZ+Uch
lu+ssOKKNIzryuajiMqc1y/+zanT7jXIRVhdjeQTJCAYmKYH+QYF9j/KoeHrQbMe
A0VJMrcpYD5mneVf5WIDzw8joZpjj3wYJYAjTOCbOez60/sd1gjz6OcyXaDJujdT
MitxIk1ykDz88NR2SXf6f4o6iauThQiPIyjW8Om7nDcWhnh/9XoZVtEsafFdSNZo
uFfBzdTfsGsxxz8/WEqt4Gyzb6B27PIjkyxLU0kQalRB3XyEUiH8HEbLm2Tmb64L
zebXjks5QCmwTuG7/NewJv6Pkd3miPmLIyq7FopeswYAiWxIwd09E3Rd1Z5+eNW6
8GEtdRgCaJtbta/3w29WWGWzcQEpNSjjGyfsJasuEE4KGm4HNg8X87x7w/u+KEt6
h5EhNHg74332gYSPPRWyWIuTIceNySlm+8+x/r0gu5Rn2j3x1b4tqlZy4rJQeCJ9
zLEbgNK4hjNd4Ej+1eacyoP92WRapqMFHvOWaXliy2g+lVVFEBMxJIwWvLGCzsvP
I7PMD+QcqhF31c09AEgVKPvWCUX4+4iEjoQu5mzcYR9+BAotxWV4GWYSezLuxa7z
5SzV3hc8/Qp45Tj4KFsm/C5dmsIRNAHB5ElWwQD2++vynOV2XdMoJ7RsbJ+4mfPh
T2qFPfO1WCMHn1i4Z/g1YlHCloqmcK1ztRMqqwiBIMTcT+hlL2ECmWOdDSgiZHZC
y4gYQG1T6AlKDCYluXXhaKCdKT2DJFjXZvIsZIvUeyAuaj1qho7J8XJ8a7I94osp
ussZQtGWB2hAjswEQeYlZ6sYlPxoI0rpva6KHi0nuiVzZRRJ4YUdq2SIjK0MtUzW
JfrN/k1yn/YBKy6QqKQ9x0dJ6GGoSxCNoXscRYKtoFOUc8xiPF1AJSHNDrufGo2J
sZ4Oeh7cPyZh6VJhJ12yW4cUEvQN2EB7ZsYsvv6k1TT7PNMqsVyOpo9q8Zegstkq
1fJOFT8LH9Cfag83s8HP67aUA+X0JBQdNodTQFjDz4MTM6EdRlNOMdbKYZkPbykx
PB/KNs6xSg3BVR5IRF6lcYHqU75jqwROHBfEvm+/9SQnjugVvPFrN+njqdlXnX/T
AQbF9Ky7fBU1OYIqr5Z++T5op8H+8KGYL+Lfb23BLBk6RZ+dIwVIJWH0JOrmAhxV
AspFaXz90IK0qLWDJEGdV45n30W2k0FkWz0+e9VMSwST8ZvMOVnarOA1cI2oakYm
TB/G8Vi2F4euoreCjyMmxPl8gcquub93vSiFCCSzTwmuEzAp9L2LYwq0Pj87Tg1Z
IAMEm0gIP2bsKEdv0uWctI+he6S3OVLPWF7M4bdCDEg9NAk7T88cNqtDDm5dJwqd
2VzbNRWyY0kBG/2IQ22L96/u8VfpbCq7CvkfPCYiLlzGxfzzkcbAl0oGT8H0MyN0
XNf+52/VzG5QZR5Kl812tNu+53ji20B6dsLfmTtO0/gqW6AwbBg2NH+NaPa7P4cp
FZdRj5Fh8YQ97HYia+FYWV3hmdBagZbv6KmWNUCGB9f0mCh0KnZce9S9JRtHM3En
SosezCg7c33EdGUDNpija6Qcx6Vq8rojUzkXbfSNprvBgvI0GtFYLRr9Nwa6fUEn
NB+abTa1vYJd5OrAR0U72DQZjsW1Bzl1Hne5lHJl1wUTbyy2KgZMbpz4C6EYsTVe
Zh6utJY4ISCePPoLyRVtyynOAKEQZQryrGYK837CghNiYITKhEeD/rbOqG0UimGP
LOGBum6ITwt5Gk/1MxMnm0xL9AxT1/tlt7EzbIYNhyIBDxAoQcnllj+hAZiNDBdw
lYwrFRrjn1i/q3/MoO2q74WdN3CagcQ+lSeAAyuwHsMWZ3eDrIvkxE/bg0d/SIEE
3jY9Wif16Qjk19k/NQkpHLOsQSxCpg6VP4rcnjyCfEN5PSF16YIr9X68B1GC+hB1
CqPPXoC/C9a6vdM2Q3YcWq3wYnhWBmmOklPorRWi0zGYhSz+jvEgl9gCNpo//oNM
hd03LSwLBLQR/HLaZD3vXFzqe3+yaQyNilNV1crrdYQ8iJscc1pCmgMW7Hyrl1Ig
rA4ilgHCd7mxAwzCjeIRZQW35RrundVuj0wC+6+/I/MzuNwC/KHtd0KGA9f4jL5O
hngYWk64dZ1uC6ki4HSKb5LKKAFe7PPyo9172MNPVqcvAfP3qYEiB/RYp5o9Endr
yugD6TtFYEfqq55GITjI1l6xjynyKILrBb3aLpoFB0YF6hV25LjxCxclElC1I55N
NJmvchdb7udni6fZB7acxSWzJ2laREp1kK+2XxzN9GFf5lq8Jmns0hikVCmhj/iv
CvIBGu93IjnjpZ47lC0+W0ULDzC0QlbAfeUYCg6JpV8IXr3hFUSc5k84OHJQvKfk
Zqw3W1LX6KS9PpNa4qG9IDjj56rZW9Ot2f8uAAeOah61RlMJM1ivYkfMdU+Q9n8/
c1JYYvJfh65BAFuyLxybzJRv/IB7yPOGdvG1YOvhVrCKS4cp7mw83yM9Ckki9pZd
OuP1li1iQHWbIQyS5TmSVGMn4Xy/srtMLmIHG7Dm42taXgD8x9DAtypULBBKZpvX
6OEszoHTA0g6ngmeBRz0hxh4EdzlZTa85eSIsSDibxFY1Awm7f/TO1G14a79zbkO
y/wBkU+c4KpiGNn2hFRwNvRuaR0MQt3kT/gEq96gBbvnhIhgT7h9spPyWasCf5p1
XXAjYlfBKr0BSwfLSb+vLe7Ga6nmH3IGdVnAwkqMyuBUofuHn9Zxv1Q2hzNvums0
4zFI3r7Ctvx79sP5nnpdhI24bBdPsZUgFwhh+NCcb23SGRKVnwcaGBpD1riLRLs0
5uGI5fJIY1skzi+bUsvHRhOXlJYgRSe+63u6pX7DPev4boxKtJ4+zvI4oJydRAS0
x2hshTIXfxpmPeh8+FJm7zA6IncNM9bbMkIhgNwTJ+jGHlq4o1Q63hym+6ZdhVWk
/+ctqy/PpjeSQX/a5cky4QctKTaJHCwmHLQ7EK8KLzcscmtmQhk/J6jBYzzpp18E
E5Bk0QGXh2q6llV4S/zTBzM6Stf/aekGg3Y5r5qKns1AaH2RkjHvUJS+wstRLNQo
5nTV4mmr6ZqRmVqMyFWP5tc9iqmGTOorjnsZ9Fa7QN3Vqwa3rJrD3lrZNQy5uFTd
h3V3ur/KCsCnH/Vo8ehKaCujkwKa2Z6PG3DSJNAz56CmiKQDrH8koAisIPDcc5yr
ZeEryXsdtLUdj+nMYzb4Pyl28fl07dtwUsQT/aWm2R4zYF1FZjbD4+nxbznHaL0m
sbSRoLc9GzDuhnh2T0VkqHy1eGVD9M7EqB0PIGtgZFw1jOv8Mi705I2WC+/2Jnz3
XeEGLmXJyXjn5oUnZcK7FJPfiZY6FZ0Zvf2+/qKMoq1LXz49OnQHGPuqNAHHdm3M
/VO8MHUu6SqRl8IDyu2X4Ym+jzNIO4KmuQDS0JJfjX+Q2/hH/1La10P7xpLTtine
52nz1lqGxkOaQiepY1vc2wI1+7VqaIJ+IWMRq1pMJu/nhJPW3Pt5N+nku5vTReVK
e6nd3NO7BgJcbQKG1R4YbFpsTe0ThsBUTYpRrlXlrV1/rdmLZAyifF8CuIgADvUU
+J/Q0LKtIDanNXKD3DN1uQqfCujM5CGDgaIH4sEVrdqte2GqJa0SRDvfAreo7zd9
4qFANWnLNCwXZI1NuOAXwQUV1/PZ2MSF5rGIdMC8Tr0FhnVa57dZ92i6/bfglTXW
Gpxc9hQEjXMI4IWhd65WCBsNYNqUWP30qeRHYuFNoL3gQTxueI2i++TGTvuiH1Ul
7dEJndJwiHJTWenqRsDILZq35Yo3y0sA9DeZCogf0b4Qg/Tdn7bH6npygdXoqVaY
JaxaWgh4QFGrDov5NwbURDEBy7tKsQ7M13wDvREGjQ5gZGt06qXnM+Y/tHE4JT3C
1kl8N6ugVC5r/ZMVXNOFal1XavMAGnqAPDLFPhRiVumyPnl8BGUyHIonsf4rqYxg
EmCcR6OCthfsgOhyqzz8TeVl1lj111SBwJeWr2UHAb61HoIq8KZkNaCEw7wgs0Ok
nymDe2pN6ltC/otAc0s/a1MI//NyV/mbuH4IGh7jNNeCNnk82D5DysmZ/RhhWusT
ezEs2PeTVXBUKlJU7esXn8RPN5yw2XKlZO9yhv35aUw/mnW8yZa13R5jpTT7pt4N
bpmDSHdLQXNLmI1a0zD8Oka+5e91t4G6p1r7vttFuiE7F+j3eylD5rQUuGgb8IW3
p+rOW116ku3oOxaBTBes6V/64GoeHbU6p+KWEZhMz67B5KEBDufpqVGedjk54mWe
rMenhqaS5oENSXxZCs6/A8LnqlxNj7SHpZoKnxZ03h0hKaOX4SD+9QpnhMndYK65
WPQweZ5ty0Ti2ZYlyeBGhBFQwfu8M0iLii+Nz5zLzBHq9jvIn2e3eJcQ92NwtCQi
Rtlai8a6S9yh1gWzoGFYB8cL5kLs1K5jm6/n1j0TMUYSEHG9gfMasPNZktt7UQhe
a5LzGPJ/nPraUyjXjKtDJVhC8GJfwQD8xcbLNVZptZwpkAhzwPeExmJyXaIjpBs0
kqF/33bi9BziC9E76f5x84wFzLna96oia1RYjINOQcVBQPUpdKNv3UXseE1Jz8D/
b3vij+QT1qdmkIblSDuRK4NI7H0HZ8nyVpOXQed7JoCI3AfpMikI6W+aeO89XYtv
0GkC5ThURrZCetgmKZQXFaVnaFwUZYToxTZYMV5nT7xJBwWEzZlfLbmhfwTcUv+/
1ngLvhQB/lp2ecjL7Gxe2aDd9KHODfJ13DD3EprrBF7Fi2iyUTP6jJN036WqyfvP
1sdIczEPd/fQsS1mUsDgpSa6rstpbmnm+pseis7VFotxV0HIsxvyzmk2DgNhBPHR
pzrvABaskp/xHsFjPVT4zMo86Pg9s4uwKYjPXhwksAqk+rZsgUEkWbQlGz5h/2qu
RtJCW4YiOaLd3pwGb+J1gAMWqN7EC5KeW9uLrH6SrdZC0RAU+5NxAE47Ek2HfZTn
+EkySTkSN/m8piRUSM9SahGyLBqJToop/XzPx4crTod+e+gB7iQnNTMNlfp9AfLf
q39E4MbFYHsaA1IN8CIWvsU16+F3TzPDdp7LOodnaKu8OX4RKgxn7YQ6t5BqdPXO
s7c1mCXWkiF4kJRhr+jJzrUddpsRb1OIx+kt1o75s8tbT4C+xDwjOsyMTkWPmEsu
dDfS5Dc9QdEcaC4AQvNHqyaj6bm4adGq/K5HdISAysEnLHzAjktXbElit/szMS+e
Y+ygrWH1b/GYJhlyCeIV0pIHxx41SpiOUiWstNMVz4gZWKX3QSpRPPCB6gHcOpqK
eNj2skcbT0dkiXNn/NXP41z/HP+wvrVFzfxTc7ijcu4mvi0Np8tEB6naFor1qqbQ
L2Uj+p9IXs5y2GkjsAkiyRzsRe5wa3c9IEg0xn+KePqsfh4w7HKNzNQ/QqId+Bge
BKQhft/IT3zQOfGUvb2jn03AeMC4+GKLtwzL+l146vmIP+5GfL4IZ7/l066uR421
2JA8nsKFBUbjkaFi5fe8YKWjUJ6I14Um6TOT/0kKJmW7BrA5iW9LRW6kSzYmoECR
0GOxpkaQDbddTq4wYqPyz8Jn18MB6hbhXot3FAb3x0B1X3nlHXzfuhsolPT+VhnM
K+T8Gy/oLK0MgYrtqEqDiegSvDqqUzEgUb4da46VjJHD8l58WP3QB93ztStm0C3N
jL3EBuk3Q5Iikvdcmj7B/O/60gczEvPR8NMJBqwxuYoeVbYXY6QVw/7SHitR7iEW
3rUURHuu7jQPy+j8qZxunqM6eaclKI1y6H9gCZ7x2iKnZnKWrt6PLoADnYefSM2e
KjjcHRqqyPNrl738l7VOxPBM84F0JcGjuTLtpfje2CcTROFUPT2jqexH6ryfjaIc
3KBFu7+lBRyLeMZXV93zdN3jsXbqDuyJ599lT7wMd74oktH9zn5s05xwIRyjMldA
DK6YSAV3qP9vGF6M2PuXN2Ffxq5nQODZvQqcQCnfTmli53Sg4vrXAwvieZJoeajm
Wr9L8hytWBQDGTz6SzzWUsXPo5Cf+6Y1zlF6DG7Tq/Yd1jld3x7x7xF4oSp5tftM
otGuipB7uM21QRrZCCzYbY3cXwNbx6mkXvxx+piPQEnCXYGWM9ZGvTnoYeA5XhvY
2l8wkr/OIlXPUegEpjMxKjevuUpwOjF8fCLlD5Yjf625ty2307XBR3i4tOLzs+jR
WztSrefZ7dkqkB+Zr068q8BT1MPCtiZn3kVC25gsnCDZ3Iv0PRx/lzCJmwKJKZXZ
N790GVNtgSbmveJ9WD+Fi/xlRmCFNeDsd8e2rQc3i1iL2/IOxGUdCCx63uq2m2nO
YOmd56SK7UEElsA6SXj6b3xnrsG2VGFYkotVeB5vb2kIxZgdLBnzjJohuroAPCme
wtgYdMZcPfPoRMa2M9VvphalimIsECNyKZC6Wx5lNIjzwNrm2ZCjgVKLwH9fPk/c
/J6eRFziXseU5wBa6TkgEd1/dJpZSheerhza+jwwDlK3GnPdlhz7SLf0PvcRoR7l
SAPm/dxhEir4reHISYqUG8HVaiAeh92TWoF0UsVCXjiIVx+m1BYkk4C3RkgNJiye
0RkejP7t4tFbI5q/3/3MkjF3rGOAHA1N5OtGgyzxh3GlEsIfV4RSOYUFdcvgyvE0
swTo2/mP3XiSn5yL0lC4Q1s6ev7kM2rIpK7ucbkV2d4iMOXgCMth6t+p4tdtY/JP
qybf3M5rhUyzWDeRgsYPNYO0sT09mkFVKOrMDFyaHmOp0v++E6OvRAqe2YKBI0lY
12X4rebWHP+BbbTXjY2hgYXepy5UfKqQ4XZBX5Ak6dJ5k1yOdFB8EgAgcQTrhsC1
Sakskis88mehwuQZVMEoRxTqREPP8nddYa4L0mKO99rkTZ+Iyp2A2RXt5H8bA70U
B+8o4RAh5X8Bmsq0rFRVGso4Cf7HIrfwsMUJb2k+35P5tLLMMdm+0ZVb7z+ovTLu
83jw3hkwCvghYJb4pZOQputzLK71fyphG0v+QXsbH/KT5LISHUuNNzed0IC2QjYM
VfihWF6s2zQLE/6wYZTUiCYQYL0RANEcxRecoWd40sw9PFPglenEuhEJNHeG18zF
Np86YbxPcN6GN4T8KLAeEpnicbDGH1z1MNGTa5vZi0WnQ2in5lBWT8upf4dXhnOG
oIq0VcdQe1u5gucuJVvscCbBOhmcl0R8kAynRSMjqNRt0yPdTvCPm/5Qag1hr3rF
dICe/zYnrOYImhYmayD9dkSzJGalwLkckRXF4JSqXseY+wTadps8bldmjEBk/10U
HiDXYbn9gHzTwVNu4sIka9ZD2an7zE6nrwgM58RHvY76dkoVb2gvqVKAdhEmmZX+
XNrhHqrxeo93qZGR99GYxF/da2p+vDRlIKJ/dudVOmjgXx1f8NKeAbJK7wC1Oxkd
4GwFGSx6VZV18X+H4Kk3WoxkeYHRqlyoliSMjb93qmoP5e+YsT/JworRWAIJnxfw
46NrZ/dak7bgVdDuqiEFXCDfFuNYEHfP0txHXNg35l0SFqlxdg1qh40laYglbY1w
niXwS8/W3Sk3WYzMEbSNOeS8EdrRM+yyJ9ChAq03R+p6hKYljaTX9MgrPR1hKIQO
PEFMYgvB6uHmAWRDZdXyYVBxkBrRmgSZWpqp7jS/5bQMMBF3JkDIpcVBOUjPEAvY
uf0A2XQRv4nnQ5w5NCgWZ9jI6YwzekPxkNOXibSnbJ/LUhRCYdZv+b2HOtE8xooN
w7MWr0snXn3FFK/BtuMt1O6pullNTlnSL+x0V5yxg9hYdbjc2xDdIqaMLSfpQUK1
+b/miC2AfVyKOlIx2ON2pCFPkVzXg8Qxpps4lqegtRFATzgt8hchzEvS0KX3/zTF
sE6Q8BW+rCNV4XkQeWTG/57oqh32ADKBn/3Q0LzWyxYO6WVs8WPxgKYgb7Mr2kFq
BE24R8YElzORhFWvQseZdIHCVeom48pCRulmmzEpSlB9akUv89ZntdqmEDXb4kt6
3Y2jkU2cq81ayL8gPXtMQriKSOwvIUWLHAT0/ECR255zexe6pMcG3uLSHtVjIVpU
zfc5K1T/3v5ukNNM/x0VeVQ/l0MRcWDI2NMz2SLWBWArs5e+RLCmFv1mlGMMMr3h
un+VKBUUF+N+5ztScOuPuusvmkZlIegwLC+iroIcclbAwg0S80vlmRVY76neJZTj
MF90OskAmTPQTI68vaS/K7m7jc587aUSCCNLQ+BxEr9c0cZx9CKOrAKzRc2j4DpZ
jj6wzBvnghmjoLeQs57vOU+koxo9sMliS9QOYSqU77UxEYmfKMwXwY8+bDqU5yJr
s5mjMuYGXhCZtNLx29nGEA1ec+dwpVLm0RCli2Ij9GY9A2R2/NsvZTiJitfTsNf9
sMHwPs8Z4Y19aAAsFSmw2zTfmLFFK8vaFrnoevOqTACAmErveZ0FiZxJFR/dLFV3
LSIpmySVb/622Z9fy5ak+uZo1RfDuTJIpJOz0zn6uNnHjlCTGserHDUUIk6q/J/k
NY3EeSFFBArnud6Axb2EoM08p2J3uAXO7q0ip3+kMqw66yzSTAvUYPWwMSf7sxJ0
5peyCKcCrYcEB+Sf8ZPi+xLOrzTjcy+h13YO64ZiP1jiAw4CkgU2kVu9Zrnn5xeL
Aj4hQ9A97YgmsvbrlGPV/DLeIhD5VpzICPZaTA5/8va43sVnOixoIy2iQm2yaKAX
OXGBAi9FsZBhyDRy/LLcqsWxqauQ0J0XTOxXb6cde6ry9PEEO/vqmy7JQV6pO02i
c2M3ZvwF5vGjcWIXlv0X6XO9pcOgnpENVQsnaeXLahezEvn5PxmZe/QX/WhnF3uR
xJTSWsWpLINNNumRFDQ30EAYUIp/tKTq3IE4BdmhrYucMym3jHkJMaY+TT9Xu05I
h6EcsVgz36tH94cr5xn5TT0WlPQx/fi9k25uyaEVs8IpMppau5n/O3c9lMsy0d3c
AL+uMU+Q+u0WpgZHU9z3ehzVuhIYwV+UwRbZcRqPk1leX8gvUUZZaZ/qd/AFTlOG
YBgT4RA6u7NXCpHqtCMKnThNBP3j8xKSyzXY/e9vIkF3UzMB/niPF+q1OjjZ+X54
QWWP1WBDiF54v3KFh9PF4RPRawolNwGu4o/JzIs1Iy3s55FTo7zf58Z7fZsqVLFF
Ad5otetiSpOUBxQgfQfSX7E2i4gdyK64U8Lr4hswkSrMbNlFuZgUzTJSB2qjoMta
z8ML/T2O/hv3uwKYzQP4NgkiCGEnIEpHaXLxuI53x3JoBMEJReHIkPd2bkKoIJWN
ih1CWxvt1QfUcq7MqXVrWk+v4sWF3J1tzoz00gjje3Erriiv7ciD8ofQ4uRldeXD
0NzcIc9y5gIjCrPWA1WdZIyWHhsy8GzxSdtD0ZGgqwTSsa7XJ4h/KTgkLgjM7vq7
ekfNkW5Hi+moyLjidGVbJRVuReCteVloAZH8S2D23FeZoA11cu4Ixs0tO0FEbNM/
dg5yvdj/FJJo/drCWIAYo3KEvt6j/ao1tVnJywPwwcjJspYt7VeoJ/lD34WL20T7
0mxbyEzAlgdctA5K7tNe3izpEdcTzDLRGJe0TIUNT2FDZWwTbjhYswUHHhRvtcEk
SV/MNTCd6XpkOcaKq9azHKIWmfQPhn2opCpCHJryS9N/7nLvNMOnMJP3nqovgKip
ew90qNGfP1vl1siUtjbyaCjUjEBjlPcgnL/69nydXTEy6NHbK8YDcxAHPambOLRP
4ieYJM5irIkg+XSkbn/1HYVtKcJZFVGegraXC9vNei6I6NAbRCPgmKzScpS1bKlc
ZzTsL5brJgWfMway93ByBGp38QD0X1q53PhViL00T81ycg6nqzUDHjvnv7AG2+zb
utWFOLG4980lt3cndHBfcp8ZWbkqeOLblnAJgLoQa+CD1Rxmo/Srs7NuQQMeF4bL
VSmLlF2ednM+Q4yF9wEkv9InaFNgNxhpjZ80dTTlRMjwf6VyscUE1037xcxJ0P+C
HcM/gfDlVXYYHtnNBu5Vde4xMSUkEru49XfEAGxUaMk8ZKHdpZQpgIxYepX0Yb2O
VUUFRFGjGOkA4azdDhwp0vc19mwLhtG5cRSpSWFXCEJKPndV1jltqfVgdVvF47lt
RspTTbPMVCYWkrkTgtCPwBMEWaN0/1uH1IaSWQRf8p3DjQvNqO8mtkuRzXFvy64Q
MMExEzAb+0RjtxF+/kUGtQbA5ie/THTW7uDrPreOgobKC+ySCj2dyp9Hd5TfoOaw
HpqegezYTCcqcQRiQ8vSY5cd9701u0x17ixzn0pmzCkd0zgCX9nsj7Jfh1x/5Zh8
hv/gBl/fqncyX14YZBrszo639TDD1V6Dvg0FwmhtbPX3XTJVELhCWjzofqxdLwLp
RvPED5ehtyjEN21S+osUqBNFAlGmPyIZBxXDEbE0suLYQEz0cKV67jlNa01HKHgb
kVquGbaNFukVlQbttmUCql+t8U4jjuj7Qtb6lsj9cVdtCXmhDq6ttTGYMXVw+wzr
eOIWRySjB76NDDoIXBO0s+Kmm3tQGycbS+ap+/LvnGyQTv+4HkpIQBNEnTa0l6Ow
HL9l3YL3/dGrO2v4DAAGNQ6TaBC13yvwQCuNukT+lli7mLwkGdwOe8fzeEdnYFhv
v/9GMlQOHEqms89lfY2Oe7dBCHElpk9ehywWMKnqru5xMAHzw6RiU9g2dzmb6khI
T/6zSY+RlCQrc8yhYyYwW/wHEWKU1KceB4ndR41kIrvgeAlCbajraQ6HYdbpugHv
Ke+h5d5x15eq6SgL8InKhie7uXJ57HpGp0AHFxJyaosDXhazFl5wyiMD5GFuNuXL
VfERt0krFC7TdwCPZBAaRnyKEJVYJapcNGunBk6yZYe7XViKUZ3D1zsKmqp6YH2a
Z6jJLw9oR0noGMlE4FUwzs2VvJAnTLoXpVSLNuOm96H6lwlM+fCrCoHyfde8ChZ2
zRwE8+f4NJUv5dCc++sp1rC57Kdjtv3ZNnfsIgelu41yDS0PxScEs2YgaVZT3jt0
fRIrBCNaNXI2+Utg8NSkjRjTpIKWPHxJ8boJ2L/OqHbUbcapMjOhNJAm0ig1l7L7
+wdqSqs7Wkn8xx4JoZu4NIFI02oeiXol36U1AKVtvF7zwmceXAFi5SV9MHSXpdmQ
B3zuYHjIijbapkHKva3Dl5IChLCqQ8ISL3H87y2jJaJsyZjjh8zH/U/cXOndWVjl
+hi5QnJnG/6GgY0eKaqZ6Mz88HcoQVyetiu8WGURxYFqmRrNohb7S6J0LQJQ4Gaf
5Po9oASi/IlMmZTPATlQUP5M2x5kdlR0EZKc5N6Iod8QpyFFfzRdz+CalO7pLGYm
mzhTjPWrty1Q8UcNYXkvuzz+3U0seplSYnssowGb9QUPDh+3jp5PoMtbTWF7cR6U
vgWND2DTBADCogecE0JsmHX1DfOc15EYR0XxvUQn/hYMpDjQnmhUWbZhehs7mTGF
6OOnSVtaf5EY8jWBjrQ6dC1IrEbCaMHSMGDADYVKj2g74sV4Aryid5By1jgUAKMD
qHzCucqOc8Ts3H1x+2qZJIUtGguxgGr7jsklV7GJvQ7JI1yzRMjbkxPXLM1am5fh
DqhmcDSUiRBdRkRZ9UxjQP7hGS3z/ZA+AbQH7LkBQDYgcnm1xPlOr1tHXfoedzdQ
M/YtKA5mczWi3juJ0y7FTN3uKcIKlGbjZfDg55qSztK06la52ne2w0keZ55PB6IB
vTh3laiQ+Pxpr/awrNfVXf1P3udcGf/cLCaU7+HyWWINP4gRaPMZURson2bH1c5i
jzpNn63hPFN1hRI/rOiWzJnSHnWJprglLmX/ehVuanOXkVlrBA/QoTc4t2xAnzf+
LVT0CzgR6hJ7ZrzYqAik+stVwKh1A20Hxf2D6Bvx5Um6pCdTsXVbcqB9x9VN63m8
bFGvPrMTNQyItoa+oZ9Gx7cDvWNPt4i2ovexiaGRoKAhy+xbuWXJ8PoTCft/q64Y
rMJCg3bhBjn4SlhgEEpD5Cp6FE+BnBwm/AiQQiXRhAlYOfRRF2Vx2VDC68SHZPTl
T4DgSpwaSLxc1KPnK+88cQumMKWB++EiIiNHM/Muvlg97pm6LTJlrsTP8eSq4m+7
Vq+PG47AcqHtV0Kcdngc7hgk4xCtKwK4IUGbc1hLcvoBR5u5F5/GQYjeBF4oTdZp
8jajJLS6UIvmkIra2F9jmxHso1+dHGRArJQNx7pWwpVjseqj0AVp/K7+tRiutprg
n/Or0L6I7BGJzvRr8BxweIqE154/GC8UnOJv4sv4Hhz6vLzcfzXTRlDjHiv0YJjJ
09TvqAgHKyeyW6rmCRw2atXJIssOuqg/p90KQmOv2ONN6n3TVkxcg1xOqyPSt3aB
sbODjJlUKGtBSi8H5u0KhK7ExbdYZRvqedXkS5n2S5HgR5qrD+hsReRotoJrBcVl
XcRPWtfrTCc2PKd9i+iKDH/xh/g4MJzWbb4dkSA8oReKhHZoGaDRgbVJeRs+Asf7
l4CsvkWun9qHae6zfG+9TxodYT4Z7imtqEWyOIs1PC8JDulMxzvnODUF8weHoh99
6YG1TTyDM/UTnrBU3Cvnyk2RIobJvOZmkDB46Pla1QDBztKGng1og9SelBtAK9hN
enePMasthwNkhOfUgIJmiY/XbCNH/dT3dwm0fL1bGVItKHX8we4vWonvceWMJieL
ni74c12lD+yQdKWpPbsZm2GRe54XnfH23g7U83r5wzdUBWcuiYlTVek27dvRx2aM
Tui/s2zCz78fGXbVihabKhDxvs3H9Uq/Ke12Jk5y6l9DmtDZQLQU9BCeAKTgFcXE
Z4VSrsk6bahYMYVMKivcO2jb6SorvP0GnWBlTJu0nOh7O2XlN0Aa5rpyyClRDbU7
QAPRoQvdGlOmrbjP+k53AV6OnFQK0UTGPdbBBHFdwQL6pmeiUE1oHCiaWvUdsE8c
AC0ntRdOGKWksAn1ICI33xP6RgR+lKdG27++B4IDZ4IO9a4IkG/0dKOJoVWXfZBk
9vF7BLEMR9dEYtR9IFmRQjLL2SXMoO0z8sinFvOKD4Vb2FA8jmqksErF/EJpl+h6
+ZIM78PkrIHyyceandZ2x6bS1NejeJA0X487y8UQhCzVgOJzCPAYaTrbdxI1mjQd
ovBGqqGiIXKWhXAzEskF0ULSM+qhaP9SW/EHspVdyk0T/r+ZZu8wSVgJafnP++WW
QAm8qE8aNUYK6EPiYu2Ng03/6gT3oTMG/16iQd1g2oqZoKWbhZ8xhRzJH3Y8v0e6
4N8eq97G+OF5YAi/ja3IYkULtyyy4g9qecdyOEnd4o1dLIkCl476eoDldWQiL4nA
LFps/JMJtu5w4frR571Ch7slnimOq1wAXMwMk2OKKyJw4Jq393tu/Ag0lUbWco6E
C5kS2nYzkSUqD4vgoAvsUp4cAHGadJ1g7meOK1sy2lOmtm6JNwfzFfAyxD9wYaxs
su3Uor7yvIHF+ShALVgL4X1mqWHNPO8QpDJXKgmcNibdD2Fr+curbcrxSbMOCnKG
K4jJZyVF9/bKbIqp1pjh+4Ut7/zPX/gwSPbCVQgnZQQlrj08tlMtttBdlHXrhb15
/Esqej5YfB7sxlS6NSZslLZ4bzV81UyQV51OOaz77sU8r2czCVivo+gGb9AFhOtw
INJ83ZqphucKcrTY/J0c9N5+Hthj+25zxcYKiFabthFqWnQIZAhVGSBJjCRUFXX1
/2/z9OrZWjGW+eE2hL4hi7pDuNipB42HnKwPVY6aGPubesNNyRYee2Nhrxh1CLo1
8WlwJbUh2bKr/qK6cEHsx7stkTuhbOW2h0S0lJbVvsNr7VEyz3qYcivaPfTUWOzB
DNLms7gAeGEqPRG6htdtE2ylKFNyOyPMve3ukEnLxh/NNCV/Zv89kwtBO19LvTLJ
tmc2XUoGxBXeoIdstrDJg56j9vd1Kf1ko3l0/d8+pp4JyVClhE2d9CBv91KPcw36
YNcM6U+z1y/a8kdq073lPvbmHqNf6UiRsL5Bt0JsLHjU5RzyWZuHBCuCG+syCttW
DG32OYXINXLVr21ZVdFhvJnFO7OZjT8iqY6KRyVPitb4U8gkyTshjQjsWT8XB9Ry
Eiyz2qW2fBEqEBaocT+YJm8JKLXOBTyig7y7QpBGS8NNmhSlkaoG3saWY4TVtpn8
zJWbjWGRV4F0Qe2QaG3Ep0kcLQ8mqwNek9VrpASrLXvMkM7eIsGD6QG8xbSUesh7
nYx5PyohqlijTPUnMRvpUQQkd2g+dTOoCs5fXnDn508Fb4baua3RE7cdwI2LmBB7
CFmzCkJZRKYJ30ope00G1LcFKcud4DtIWsa0hTMVZNrh5aqtiqRlrpQUH8MoUXfR
p4Jc68nx7Oly/sPe8dMq2IqfiRh5JNMxgdgB/7LOqGauflEBMF8cg45/IYjVxH5d
KTTrwTM1RbR0eRvO8DS7+VU8okMliSzhwxu9JBikIzuqAm0uEc/AT65NDNLTTpro
nJqeYfM6Id0eQPJdguSia8bmVQ1wSvSLSrGD/gxycexMJqqIAX/N5vfj78pstlYn
VoKxto0GDC/eTP6biXGr6/zYN1cxi/BjtacYF78ckpje8zoJAz/OHFPDG7p+ukDl
WHfdzlWwAteGtabOpiNLmkr+siG6mgMJIba3r2E3VXMEVdosjFwBPVNmXxPYpZVn
TZO5XZGvuFQpfJ2ODWRLOokqkvcuV0bObm1lotP2A8p/Hv3qSR4ZmxY6DUnbWrla
IrfEAb2D5D25glXx4vBupLOhXDdBEUEhva1sooMx2fjVLREPtk63mmoEOFHmQ/P+
LiqMUs3+Y8bH6x1yTYHeZIwSGM9XSExPz9+UwPgBDfNtoAxTCfUc7UatS1iw7/+P
J0K+YN71Ar2wvat3xoYpL7y44tlIhwO3hzYh/XxZSmGR0E9w3f5Vo1KZMEPEk1RE
ondaRs9uKOCf10m3VVCi0hW+znYv5FOkkX9aBVJfpSs9su71Ebu6UyMfouYR5oMd
mNX3B6NN4BBCeFtjShvB7AKOeAg570pMNYBz6i4R7E04UaAZPLWaMG4Pf5iOr15M
QHUrs3N1Ir4/8LHEkLPtX8n6cwNeUeQxNbU7zwTJPjcHWiEMzhpfM61cTOtau/Ld
ZCw+hy73k0K5VJTz1ddrtjTKxEBYKMztGFmxMfw7SE8BBFzRsUGbQHOyVcGiBBt7
a2W+vOGyhskkYGHYKMjtxWk3ey6qOVoZaIaimBLhwPOhgkCTszaS6EeINUZHCbJy
4YKRvPhxKV2Vmf+F02O4cUbgaAdaULCE9BG6FqowMq6/kQTAba96ekeKcBslWkQr
3nSl9FSswiVYPLoY3QCglzwkl3owJWcQ04yNE9R65iYv0A0yZjx3ySNc1sWwyIrP
D77zCVbtPG6F53tPwtxWl2OdjdS2Fw48XZonAdRg0lE2GKwFkV93onkrYpQ5tn4Q
lK0lf1mX9t1W/iUfXaez84msaXRBhzJv05C666SYouYtDqne3/Wc4SWgb+M4qQCT
Qyf93RUrWQIMLeiQU+1bjdAlmOvs42BzxAPGhzNy78Nq2f2OLxX/JXlHlL/3gUu/
xaKDdo++9cYTKBGezKBub9vPHTfHTQ1TmcFB2jI/XZqRCMeh1TCyPyjWKlTMxi7Y
EEMK42b0Gklp3kNEZubnXAqiuZe8f7jBCXLtJX5sAWOY0WkOaOv6Jn/rzg+RtwtG
Ij5DUcw5fLBz9BJ+7w0juP2udeZ4cXlEQfWHoKcKxLgDhP7FRzqNYUmXUDo0mrMF
MsI9ozDe7QUeldETqMTizvr7yhOOQBHF2Tf6Q6uIxteBh5zpvNCE83Rnk6eSslh8
9dysbJjtaG1BoRxr768WLXF7/NeX8a0s8Ecx1PSKBykLwvktrHsfWiSdeoFSG6tp
6MLFZ/wZVdpl3kLM34MjueiWpnwTH3ulNOmV/qTLJ4onmtHP0T03+xa0vBdgH3em
Y+UJb3JnOe9xK1KH83TMrS5rzEj5U07d/oUaOx5ToPiUeNEg64rCIZRCUTakwxEQ
YxpK7GO1Mh5lPpaMVep+TregofBpaY2CFT7ZqynTbJ5PdW6tdn2m8hNirK3SnJ3O
bGpmuaqWLhmUoWiqisoTpH1Yc3osQItCAvnQq9EfORaszt/DRfZ9Kb+DOcH20y/I
3N7z2p7LnewMLqHPpoYhawsFk/Fslr2s+LszZrnSgZxkhrHn8PGZ7t5HjNIxPVyC
zjIDzGCylxjUPL36/HLh0ZFIBWa+fejr2FToeRdBFzWmUnibjplLbgEVk+Y26wLm
WoVid1g/MDINQ16sPQDsj0QQhbIOLYKqzG5zZnTFPX7bCG7ie8naHVNzhViG6EeD
yhHbv8YnKgowZKgpBgNWkwCl17QNAoNeJwllwas3H7+VyxaGz+cecQVgWj2AL3oh
X3aLZc03HkA1BRTCfP5fU4Eha6Ol0pt8XCVlFQ15D/sYo+rMu5CutqZBRpHB0UTj
s4UDsMlxcUuwfJBY97k8gSG+OayvvFMR4T7TIv3fJBhl9Wd4srn+Gy3fZ855BWcu
OqleUHcdOXOHcc9B9q9DFKx7Ccds2WUWEQNrXtd1G3ilrgk485A04Uq+R4G/T5VB
h773bZ2sIzdL8DRyN9casREdS8EL96u0QOi+UKKoyS+7ONtRGPWoHkfzQoEovDK9
Gv0Fsjhd4/NkgFw+eMLpfwOUjQlmgszqpIfX/6IFQpBjT6xirMUdTeEkeNJUIr4T
V6LKGdhj+8HzQN/DB1GhWZ5iiTkCMZK61EcwlBmS1/t4WfeyFzefPbkfsgJ9mecF
r2/dlJNsLR3xM+fnTZmCMOSLOwvfxn3sHei3DQdTFKk56VC3uBjehSNQMYXhlz1c
PSCEqrx5hvqUkgiUJPxkkz9kR9Zq1I6LiU9H0RCJYMi03ukDcjByLGiNEhNheJbg
aaLoqvazzUdI+d3hVP18BfN7bhMvVyc685JjnlC9LCYaueMMkp/aiO/brKYcE8gD
MKzjPq6FHlwTVEyAqkpO+fLTMjNzqUdr5QBoSXNFHf7V18osr/7+PS8TxAA7mvj+
/FxbivxmoNngizC3gKTbi5GBqns8WIg/ocLFZZ8RDMZnPuKodIUSQPAaCMdRza1/
gGMPOUr8myDAfxFEhzzeoBMuS/r3tfQi99M6XJkb6KnwYt+M4bF6KHVRMrBWtLNw
A6jr6eDaKLrP7o1jmWQlSMtSc5Rt5hzYm/C1omSa4XBNszJc9xZR3Qcxp8ora3YX
4kHh4Zo708lZFfzF/A5STa97C0+l071VSIzVHRs8Tw60IvwbSQ+xM/8QzbqQBQdF
kbWy17BbMbjQdibxV8aqmBon5yrgQj17A4s13UuuedIh18rXHtgJ2GcaWbdzaQxS
Qa5d2uByKxAw+22/vaKHwxjsopTPa1v+/qHSZHj4PgnQTOL9OO3NsQj4H8NdWvbv
nLAHJq3VMkIgaM2DB8tUKLruGx7GIu8Rh/Pbbl2xrVxPdNUjI7HXezsJjK9MzJNp
3ozZAB93ckKk+76ZlYhXDXWYWBSSzbhNtPW2JgLCLoKcnIaS/OQ0PkbVyytHywtd
3pJHsUsJAr/vhq/3sWVRHtBWVy+2E02p4Tk/rSgk7fRNpIIhsqbY9NmNinzOI5l+
CIOkahZzI76Rp9vnjC5bz4+5gq2A1dzQSZ/LEW+v4aD+82JlfKDQntq2I43pjIQ7
Syc4X0rExP1Be6DMnbNQ/t2501I0Ow6KYih2LmrZhl0MD2xdvKgTBAPqnfsOv4bM
gx/MfAs54u5VS2hQCZg91JYo03eysbaJksbaBgEkOFu4yGHeLtowbX8wGa2epled
lT4+rdkbD4ExySXOjiNTVCgVO6EtlmCP7xlpp51oOMrOp9Tr9umlNV5VNbw5SC+S
xrDiOzPQhPgTIeXoovFvFI8FePn8q+4YCTfQZlsu+rKTslxqjUyCnh4Fj2a4UJr7
f4I3tDQNvXksU90rzfpvyc+Kb1xGEShl9mJvlBbK1VLOBcG8PKRa/3fKJIdo9N+c
I4H9vsMR9xSZZEJhsDHtCnvM2ZkIICHkI8HagfEwksr4n70H4U72hV/cufZ6jRe7
vA0KSYZwhsPILP17xJX/Yppn0lUyg3o4qBOk4nqiv4wldI9ZL/Z9yqMVSvNfCKu8
RZKdY0wICnXxNka2z12q7cB8/2IvRp3ebu5qEPgtUg33u6UejJIy9Fh3PEwihZsB
wKY7jIN6my6JLSK00hL7Bbgko5+2QtmzudhvdlyfoPjNeE2GzAOImOCeApGapDI0
mrkoagh7LuK/ptV8gvKXFb8o60i3XLASkeKXCvNKKOl11oyoJrfcD0ncr2nQO6ja
KlPB3MX5arHdFM1UDFYmjIq6mLAYtmNo5TUrpTapJgztCngEPfjGQe7aBhymx7/N
YY6CZlHHX2b3WNXFKLGbGs1g1D2ckc1uQOdnWoR1NOgbsgaq2D04kfezlyOP7GPn
5TTUIe4vPmPAEyA1CTWqb/3c53gLYpdIySEiT0kEISEc0u6nZK3Zra3btoJVjOrC
Vos87ySpjXvsknrEqMEsQnhKxxhnEicaX4Jf06AC2UdPjO4qwU4tSESSo+Bdi4Gl
J0M2WzVOBiqMoyO3Kcx24FQwE4QIpTuACnn4M+9ak1VW0EpZHsbDE1gfxsb5hMzo
fQ49YhYrshsrj2GruoYgnfRVKmL8oX/6tFlFUNqW/IJsHVNskzFEAZliRklgzl4O
Xqckn9QRdb77HCe/YTAd5VEUmwwB+Kg+UCrHO8F/5VCKdrUTtc4raWArYpK8gbVZ
J0zdGfsemVtXDCZ2rljzPykzC59iyL2vCrRmPAIgieAOGvdulR9onBK0HjKqaybO
YXlMKI8tWfzey0f+vWK5lVgV6ianpVUrnIAuAQK1xefW/SKdtlg1X7zPlytiJSn5
hsd778ta+YWk5wus0irNdut2GVMN4SZC5rw4eRGxUUTG7k2fN/VyxDusg0uuzDrg
Ovk7OiVMhfm/KV/FMuEMqKzocq03tOH1ceeX/u51PqE1sJCuu3Am4jkxmzecz/AK
FLyt6t8zbGIETvFvEfFtTroTXl4CBVDcKRgMquK5i3ZZwC1+JJTZ7auTb+aevW5V
LmXxV3moT3XxhMEsQOKflQtXe+DbhzLTZTvAr0TwJOa2BMRkC5ByoMimbTkpTAWf
dXvI3xeV22YeBp3Fel7ZP/t5xyu5CI3V3tpKcUyHlHFH497/WiZZAagXK7zEeKXj
pDQ/0/XnZvdYIS3hkvWZrJG9H9jds7Qef2KmWL2eg1gXWKDWz3qFpXt/h+jNB3MU
z652vTWig0AqG3lay2dqCTeezVmGiVqxyIgeIKJvLl1/su791SyZ5lh7NcXxeaec
/YQQRX2NJHo1rB9H9zEzA7ZlExLJbpNT8ueltrHuXeePLCoPkAfl35KErC3P0uTd
IkHDZSNebwmXhJGqWVQV+14M1g1sssM+nk+vfDkM+pX7WEogOINtrjJEU2R3Hqwq
ZBXAhqeCaIeSyGmSXNIwUPEJ3lVQD3Va/JUAFkDPcE0XcBjkiA7gyuhuBhXq9v/D
4jkai6DQ1EOfJ2UGV6oS3MQjP6hazl3Kj8kp4XZcUXM0+FENcpWonUv5pjD9Zp/9
yYGL4kHTVmSW8BQo9j4bbo6bNsDfCDuTKk5QAs0IrJ9Ntc1BbbEbKCFTc5ajcdpb
S4OKRU3WhGg5/qWJh/U+UVPhnodLlXzaL2Q6Ff2modeLodmyH6AdmL/VxPV5nuDm
nmPns+qOJh5KCYPy2sHXw6ZPZyH+g+SRlMzA8+ue/anUKbxxhRB7J684r5RYmNEZ
nWTNeoHK19jJzNyPXVlbZU6ZP48Ec7nyPzOQ7L6a3W1BhdalsdxEGxhCSV85i5Xx
HAE4qHLMm58FsdQKOPz4ecQ7/NzIFGKQdakpG7xDlz5nJRSA64TRpjySX3AHC7DM
nhgPuu1+72KGjq4DpLW5X+W8NX0cVc248HfHT78Pq+7LVt1k313Jnf8rCSI66D3j
eNTaxvQHtIrbbEBva/fxGA4SnVm5aMDq0l4lvaUvIfNSkq+BcsKLwTknWdbLTnVF
cGAWWDF8DV0VqdAVditHF6k5lGHsJH9tztQ4eMRjgvxQ652AHyfuUAkTBMFDdP9c
my/xKYiK7YFcHrj/AHGGcI8o4eVKa/0zzMJnm9KxiRH6Hry7sPmv999IvUNXg6O4
WDhab9XvPkLpAT1t53i25f+D6OXA37jG0KID27zgv4grfhgdTwS8IRWccoMpkn1U
gfRuIowSFkPpdbeevY6DQvmb2mtgEHUV5YoyPYAOUG/SvNAfjGx32kb8sq0cBUhi
x5dVw4kLZClAk7xUVbVn+0d0vQxVyGgJXBzLNRHFXjbD2WOd/1f0DO0QEnBRcjVa
JJ+A44UnVVOQnxp6QNgYM68RmMqGjq1jDm8t73/TusbK6HmsQ0MjBxb/xC1pwvev
DngNT1YSiepcL0YrA/wgGQ==
`protect end_protected
