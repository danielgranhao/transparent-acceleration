-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
sJDnnmXP4gj8kxqTW8ISjjfcLsVd6l9hgpjbJYvGkYtSTsuj0sqNv3crtFv6Ck59
hqDOU9HABZIrITvSNrwbgsDhcfM0eM8KIh/Vpszlv+JxHt7B0H3idnaOxD/7+hGV
ZcEIVwLBKEDi/ukbN40Xag3VoKE9Nj0eNr0a3npsj0w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 11552)
`protect data_block
iQzlhdHxwnPoC8ZNxuyCbQ9OcE00xyfedgAuU886L3HGc0YXTVFXi5UJUG7Sk1/W
t8OoYBRfEN1zrck9byHuvusi9cAyxUHHljrni+ccgZF4QIZn/acEGFT3iGVwzOrq
yk4SPhO+2TC+u7UHjxYfmHjtTj9+LazoZQl2nYDF5YST02alD6R2d5c2pPklcJ3j
6NLVRk9wbTjxynNXZ3i/2TSGQp1f4HcerNRqwXGA4jjhnsJIQC1DVfEV5cC2dHAm
vKGso70EQ7jbFHcscKan/6wKuDvOo0rpZw70cqk4hNEsfXkX7vUs3knxRmLyEVbO
pLF/hG/bPK1WUuuqGcoI162alI6SyDTteMwXlekRUTRB9RwWuH6m5aqC4xbrTOq/
hsrhNeR85lCm+jAmUQKt7seWK1MW7XkkUJhCPKsRSiVQ0Wt1aWr+oxeR8eZI3HqX
I9aq/VZbYkegfslq1ojCsnbtZhVYF94uCFkAE4DwKWEC6lTaLSYsl7i0doZjdTFU
tT64HWWWoPqiNAc2c11svMDL1qEOAZ5Pn23eniiBxC9RX2tZfnQnPV+8M2joDfpV
JVMRifl5Xz0SIFgteGX8EYadaFRlsJ8XdW47qHX1SMsy/hzEmCUSvT3LV16Hzcg5
z8rrZlTqS8iUGLXcNO9wP0njHuBoBvNGm0+8M2osbanLBeNJbMFWW+SHjmy1u1nL
T0y5u6hTyFRo9ZY1VHl0eFYkq3KlSShS/8LQ8l41/YPk3899pSF51qsiGSPGfgZJ
LOSrHhLjCsehDZFu1HtFrPAPYO73go2z1nfGZ7CuTYs30DX8mkKp61bbvsnzsAvE
XPpPSWgNKgUXl7epu17EvL74DhSOe3HY5xa/MN3Qq6KcTlsL6eMnChVttgbmU9qe
BTIx9GvfR4MrFTxfbHVfICheuLBLjUtYUq1zSg6Xe2ngEb0KpYuxHYgn9Bq/xI3i
oucx+qDWpGxYhTQlFxuxwV1u47of55nz/LjbbVS+zMt7d+8pykyEZ8qu5YYiFOc9
BhUilOn3f8sGeO0uMqeopAOJCqNk3gb0lIMrJsnOLvBAGATZjQoBMibJwso2WIri
+vKetRbKtUcGb5LCOmq2d/467D+GPEnTy4yl5YUpwuRq7fP6uje9Y3B9xRun/gi2
7Vc5TFgLI03RSlziE0PeDEM4dWL99GdVhqxvLezVlxLq+fzF8xU1hv/aa7Lymk9V
0ZX6zu51mtDc/K5b7Gwqn8PPOy0jJ8qShucLzgu28M83lzS0u1oY0JaY3bz33Rhr
YQll8JlbIrzp2u+2r4yBycBqXPrTOw2+VtgvKJ2oPvKMJP4Zx2geDe4uN2sOrvkR
xnNHUGevVfFWU6GRHOu5nKwrXK4oTdx3U+8BcumnRJ0JnqP0+O53t52UBoqEbi/h
s2z0EM95DGta0dvJB+wEFamWTc53LJzlhH5rLzoSGaEdTcn+fPeXcXbgib4fE7FZ
bVWOUfV9Cju+Z+w1TDSAI6taiWh9bLnZBMenM3cCzLqnf7Yms1ciQr2U9cbj+e+/
yxf7oENvZKOF89g2WVwAlux+T0/UmDN/tfJR38ca8uscxNqDz3xigz9wkweNDNRp
CyUFNPiBr9AY/WnAH7jVmVVvc88Ob8MLltHRxdT/pAKnchBol3LPCTm56xHx7Z9x
3ECHD3PKqs53dPfEwEoa+6kgtd5QHQiw98g8jJIK0jaha67VM6xwmM4I4O7+Zbez
4QkoBQCEJ9PqTBMn8TQH+tuQIZXqhjRwEglCMKjmP6DDc8ecMh0QWoUlJuKdUh7n
z1jorXQzi5ggakkbjOuxi/URIyGoe46sMDqWnuhpRqgNyvkP00Bw1qv2Rx80ds+3
YGLOzQCcVj6RktqQqaL8XZblJJxRqNrZzJV6qBzBN4OWrdGRLlTDpdOgU7ivGF1Z
aWfSB23yWhSXP8tYK5qLdgYKEJA0FLvDR4UUwEXZ7Pn4ilq1BLbdajMfui9Ko4pP
g471dVbLyolgig0dD0R03UuaGm+VaMHQCELZJgHEe30yhQ0DDMLdyEt70vXb6gzm
MdR5rAeVve9NNzHX+VKem1OpKa5d1o8mFk9tcqpg/llxSmig+D4sDn3JLCeQ129m
kkaOk0dcmjUdDpafasq1ySU5bjIEZnc828tAo3yCjpnuRJNXMLHp0WffbS+0bkvZ
DoE3m7A4/V9qSJjz96lF5BeyLJAjaxOSP9yzZaJHUNe7gwDNxD1MAsJu9kuyeew7
3DQNtYAUpMeewWbXtSmoIJjHnZ0+ZmQJiflk5Tc5hTyy91w3+olwHEQBk8SnlWl6
DJDylux0h5fZ1iD6h6l2tUkKqr1PwUP0cmnKNGLVXUYn2ZmWoHZxq9sn+bZmGtXo
Xw76p5h6LQsL3zxmDeR1Efk5d1yes3f0kulCL98OYM6m/5XAcQM2wHnJao51Uvfd
4jnIaqCQ9X+WTQ26PWdsMZYEACoeWVWRf1RPoSvqrKR9tFZEaciGehN0saYWnrxn
L/Hv8R9OExQ91NwSIHfhspO5XY2HncpYhXlu1DCddpepkDr3K+nvYmj/r3LiP+0E
EyoUFnNksY69xHhP7lC/yJ2k06Y5FaX3veRWr2hJjDTEUquU8JoQ7bSwSETQ4OUH
T/TzYwLBWfopfLCGSUKivCqHxGY7TulqKgD8aGHJ7AaapDd7Xm6lk0wL3opnOBky
mZxM0lhXncc49gOqvaO5nLE0QXnkbPLcE/3TcxhE5CwQALNl2x6FPYdqSbY0jjrP
KgPa16rstQbYBeu60fMXXtvFF49VtNji1FLiC/qbmbJrSctdV8r0c2AguJtMlL5+
HRnqc1e4YcKjSnBH7LEWDDzHj0jucBTanwUQnm2hZL5WlbMMbArVjq7caZvABBxN
8jyfv9FdYYMjbGrg1ehIuAmXh/xv1+/xgJ/puwpUBavcIzVqeuoubZWVMXmhPXw9
Z8mofYqkN7WtBFcVUxVVsjvdiftGQuzhblkDIwjP+CwAmWddGT+PEOQbyseTIejr
3R15XYjDYAywPSGs5cNh8PcHY2RYNM3aTDNm+VGVDuSdXYqamW5x4qq8Msod7ODe
ytTURPmdLXVeTMW7yYOyYro70/JajPrNk/szks6JkSpFk3izxIth5NU8GD/0YDrS
Mw++lHxHK61vVVuFP+qQxoFlnlh9/CqTrPjyWrlJNZT3CgX5jOTBKiJzl8rN8typ
pRtF8PGuVZP39od8u6kabd8lDGV2M17zpTgxG/q9gNlb7tIMowb9lgVJWOd6AqI4
Arfc2AxD/rTNG9NomEpjze3aSYVZtFsBsSpsEbKpO5R1j2I/OaiQe9LA99enDrsb
yJBrUP+BbzucJFpB8ByjTf8WXYmcRznbohFOHeOamk8y5TSZSuEuSq+nGZPBV0AE
p331860aiy79otmvV3YHrxCNJPnwXWpYWZAM7iEKNaZAWdfdrI2vDjpbU+PfUlAK
72xWHvhcY3q9zDHL4cUlafCWPb3BbX9+lrNtAsI6f8jD46lkX1K+/0mBPaNNXhzQ
+3zqYAR451GB09iEvVWgYRR0nuWvL17iIQGTwWRu/Rq3QW9Y0u44qoLKkYtx4r3V
a06viFazy3bhbTKJZuN7p5HRTzT9DlGwbthVKN3i1Sq0JhWXyaiF2IsETR/QM5uW
EzeBLTQHslLYzikevjj/d0YSKDyNRilHQ8F+FThQhGf5uWMxAjapGgGUkv7hIuvg
fvU+t0/pUAzBfYYB3ykL+PhcHH6Ql3ZYG5WR0mlDPscM4xN6wDNjasg0Dmcxcdn2
WX8ULZUc0wMDl3a7ZQ90PV/iCWvuqFDZ0vYJmATQYtIXEazXUt5N2Z4t9XxB5nxM
+fvX7Roc1p7yjhddk6w/iW7LoKplwc4rbIs7EusN1eXxKDNlSmGi1aO+NvQ4iC2N
RCwX0UD8fLh7qDoXFDv+uj2RG26AykAnjbvl0Dl5PLGvQ/fWEPyGv2dQ9UAbbcKl
LDkMNnUubC/Ou6Goevx8lWCbkGv5C2lW6Lliacjww0SjpwO9l3l4WBiUy+nOlj13
idMHur4vdSKSfblYUwD6OygurGkdIN69ZVO5eKLnhTp9ePQVtlXzp4ipG5S/EdY+
Nk8svqVlTSTgVaGplm5qUf/C7GMvHGFuW9eaJnIEgI+4UqHgXPpGYi5805WOwmv9
CzPgICvl7PKmiZqNXoXI9YzyfHrudb2LD4ngsRKr41ovAbNJDK6S5qoQ0AB5Lq/r
kotDK9r9UBSid+4U/bfMyPVwWCy0aHKH7CEgmTixn+fLHLuOu4E+XBUBhekc4HyR
ogZznKN6gYvTD6OpPkE/tS51x+KZflmcoF4frSqf6BDn8pxnaEXnwJarj7/RQPHo
SeoV+4dQ4ZK8P89l4qI/rsDU/SG8il49jlv3xGbtECgURG5tNuOFpSFOqOktQZAT
ldRCjNPMpnIbtbDKYg5+MPceE/MxouF9cDZoU36gglStgdZFG1IoXA0odFDysw6a
34v0A4EMObdcn61u4j5Ht7C2bGYbIuQ2YtlfVP3YpOADEtqkWVDkFwWFAQdhrycX
rfcs3Yd8u5g1ApNhTPsJ3G3QjOmojIYxaniwzCX2v9apaFsfKJHTNOxI8p59RvYy
Q7qw5Ww/FcPlRTxx39BJ/sMrLN56IN5TIBdjE0MQz7+dnwDxf2CszsuchLxakpKD
A3/X75Czfyyhvr7lc8PibQgo9vghq1pH7Y9ot+tbmWfYbQOSvNOyVUWx1zte/z8y
vdgkSsGfbkY7wHJrNtdsMhf/CBLLZiduWugaZKzX+NvU4w/wBCHkMo3hUeOeoC/6
ilaImRdll0eATRgu70fy1O7wAdgpk5WGt5RZD9Zj8J8a2tAMLmrgKuPip/qo3Poy
McMnU4FJgIxYWC8/1QSYzHUbgDCcKX1O9BZln30+j9RywIjP4Rv5Zcyw2FYz+bLQ
jwlvF48J4tx3ywv9E3HI7ykpyCd7jeN2ET3Hfq+khUOmgeIkn0WW9sbnlTeUtZYh
b9qoSTSyFeSRDrS5MVf96UHLlvy0gCQtXD8hIMTUEJ2pXukEMLGqtOBixSiecvFg
iS6L4w0De0GqiG2QebaSIH8FThZlpv+1ftT/INe8sQX5EObUQn8JRTYmVduM9Bp9
nUXGnaJtKpxHy30xo92CfXr9XEWLUsL1oHIJvHDvnT85EY7aoCkucMtS/66V872J
Eq8zPJqaleMkspBjrRKBlwx7Fo6d0ymkIZ3cVFjpctet9DzwD3C4LTDvGBp53tmP
t3Zb9tfQwqQy7rRsKaxQ7IRDl/zK3OWu2/qiNg2yxL82Sxtbjn3BO54CFz5YASyx
e3/0fsnYrnc9ynEZfWICbdCfWEaSS83gn+m6bkXwsQVot1rjpwoV9jXAJOvmIASm
BO2f+H+nUkJkctOL3nz1zD/ezt+zwOMH5KTE1hFhf6BfgUjxsW3/7g6ahOdCEqq0
r9x1cvHS0onDERy4pvIItFgRGafbOgFRg+MmV4UyGuCNDhJFbzzdhV8ggWz6RFXl
gISNdeJ2iEIGvss3j57XgD4pDK+QV3BrDEtDDiA2XbynpQTBac/wq7RaxmEPzySO
zS4fnbXEHQ0DspK2EdHYdpAhH8Ih4WDd7BhRfgzPPRQwR8AA0FI1eRIuQLftCsAs
RieUiT4XqjQhOSYuLUmn59Iz6O0wwKyqGAHpnw7ZuEz4ajVTPwFBRYDx+1/1MNOc
nYYhC5DXuFBPRuoZfkGMCAXc+wO5nVo47sSeWD+ABBvoTDwk8tWcwhMGPmcJQtGN
vA3GxSlopHqSp8DL89wDiCj6cfZPoMxLPslsYj6NuI59+gmWsh494rAFodfKkQgt
xapXWmxAB4xVoGKYQgQFJUpNQxa1UQ6gbfUoF9FvyVT7OQ0XYIe8J6kKycJ558Ea
mUyxGGC13AhDjJofz0uGVXMTieKcLsLfYxQHXhOgUS05DgwCE1xvqj8Uuh8YYlQX
llJbtic4xCbRd7ie8NYFnGhGFf6qoexDlbqars96BT33eQZqDKPu0mYx+HD/f2Ma
WAmXNfjGmUmMmnuG++jjXkWcuNY5obQA2DinVRNsYdRt5/B0PEXwc3czoa9CIMjp
zWRLwu5AnuoQlIRVgbaD1gfPFitDLiJB4GuTFyo9RrfpuYBpY3aW7y4a/hm4UIze
YJkEmEvfbTjcyFJ0/A+ByFXXrGrXayKJtAAvg55O8w7YP3Bu6R0cA09SgBIKEBBa
M44J6+X9iQV47xcn8ogcf+aISfL8BsMxf6o0t95UZYKrfImQPT/gZeztVK/O799/
0epJCUh5Aqog1G2/lLxt2OUzAwlmIPz/ch+5Lz8pVlio59Hj/Ko+MX+ZWfSNqlf4
SzMYOqgMtjUKeP+lLmxDYLcDsvS4BBk/DO20rAFOQLhhAeU/NVa8u3oB5wqaLJSR
2fbeu2XVE6QQlgxg0gWNsj627w0m0f6GIi8Y977QFhUN8lZSwynooaIZkkF4uWoY
4X6GGNXr1SVI7iE59pMiJy9itrCtUnHmKVyWBv1qCpBdiCzFATfV4K5uAf45+njY
uPsm7ANVjG0PTcdVKCqbA0RzPoBwsivLAdPBAnzY42f8Q0IGcS5YZvJoyGcoIFIX
imqi7WoLMlvwxxfViURieRTOs094D6fKkKHxLzpGTAu2gUKdlYYGrzdbFUYB+rBH
6LHu1lOnvdC7cXECJV7PS6El5O38F3hKAWPiZytXWWoB73N3xOnosN4lpCN5qgHa
DKvrqZxqO8mqQTMTlc0U30eLI3nNy1VWbypSNqHMs/sqAmDGpv6CRFBdxmFe44iE
6HYfnqlRwGJ9T5aplqPd4fl0pF1XUdzC7bAfVgHh3WbjFnQT0I04fUj8/cL4LTo/
7oXDrNDW2SkRZDMOQD2r7EKFwh0aR6Yn/iMz/BM3SRzVrwd52UNjHQ0I7eADSwXQ
cOy5/bnTPcFcaCU8iIN80DfOe08YHmicbl96zKp2lPW+Dalv+bFY26tjNcZnNGVm
5u9LZiXCK5Syks0diFniAxjmoBrgMVOmiYMvGBze6AUf4BOMjCifVTgWk/gKu0mX
FdxrMkhd+eqt3/ICEMrICJ6IhdDD8CC2oN7kU7Kz66PZsrjNqiHVamfwMnhnNQUO
r1nC/SkJoUVhbumy6acP18YLUz0QpAtbWmJpBof+clod0nk6g4O92zZ6xkitiUZR
hTWP+Ap8+ec242HIWT6GEvXe2Xf9u3k73uU4unuxwW6BxKU2SnK6L7zpt0syoY3L
HYyOkIOxy9r0Hd7nvLcAoWG4sgCuqUBu4s3jRWmrI3iKzG/7xiPzAlXElHcKvxtR
hbuQYvVKf+FTEXIDELD2KrNLxxS6wQ5F/tqoioZLsEIGe7Daht4Mom0GZzCL1cUR
v7cMRIm1qY/W8llvG0Bl/7k889LgYRK6PfTurNFVWdY6+hBPNn0p6bVyWfuAG3gZ
+Iku86Tk4Zm5AWIly4a9ISJvR0kXorzP8Szx23U2bTbLSu2NMzUL3jwQgVbscTjc
TvKn4AIAri9Lzz2canQuvzcURVbO1lunNRAAtZyRQMhi/4hzOJN4n+JRpGz5EvFg
0STh0B2zN3pVPgZas8Uc0Gmb2JjK0Ni2GsFCg9d3ebZ/e2aV6gkDA0au5PoSFrAf
fySPk1MB7INi6+A46KMzsQOjfT47owgbd5fJdnFFrhu9qcIsK+L/HOEoK4KJUtHx
nRtD2upcDyUEdlGBN2SOfzbj13WnMyRQ58lP74z3+bp5thp5Sbk5DeCKpVLfnRGo
o27YsFa+pTPIrnCEwFVvEC6jULn49CniuYYT2Y2xtxm0K+txRuLX/Nk919JiefTW
+3iFSQod89VblqKGWUIl1PUNyGAISaUjUNkGmaJPa8zyrk/4nrZpagIV4H9dF375
N7RLENWSA/3S8pPjTbgHMlxmzx/4+/MFZIYfCnf7td/Wk1s3MOOKBCvmNUW5mtyt
ozs41eWoavSiSfKST+rXwouCTd9gKRO+MqY3Foks9EKMRLqOA9dVgk1R/hFsyx42
wvs+ZEdp3Slt+MuXNsl3agjKpb/jDz20XG1LxG8SfWKWGnTGOnZbrSExHuCUf0xH
00v8pgcLzjMmUM3vaaxxwp3T6nX0h6em7/HwKRGWkbYhwjLtrvrPwW7kBxOtRrki
W+rUDkA2TQrJLrSiHEsqYyKveQAFm7jtboeBhpLIGiTeqXmcRpAQJfQ0oTEuIcAj
QDPTb/JjdtA0qfS/dBjwmnp6Q8xKVU7GM7dG28y+TZchtQsLDptc9XsSu6I8Ftae
UtxThFC138a+oIONM3AIODQNrDIzbyh/fsOBjlEKMscQKaIkZ9+J9700SiJKDT5Y
BbTegiAi0rQlMuotHE2cFzlxsTX+mvTpT9NE6mzWpG3cAk+u+LmuuunExsp9S+68
1h5a4j2CLyHjHcuQRJJleFoDKz4yqFFsJlpce3+k2KH9D2KhFrPo7PE6o4ERgtVt
ZXWZoi7eb9uJ9C3SrHGjQqZoXNNGqTOkRcugCQ1kDuk2Peu7g53Z7hbG/REi9tkv
FZq6sCxkx+3Z/UMbJl932I+hdkbAB3ml9hXNod4nHVAoJyIL8DRfbDSLtZLd2C28
TeH1S1S0U2ujh2cF3FO5aeqOjDhgWTymBw0vFehgat6SSa7jInnAKwjug5bxIlee
PjrchMYhrzIMlBLEXEWlwl8xnujmT9n+9pUdI1LvN2TIm0fZQRWpRdSYOWDxHUuy
t5XiF7K3gqUQvNF2yOK6z2c0s1tGt6rlNNrueTgsXNLBwFINl1nF1yyWFFsUcURI
mb3e+WM/oOlWgFjFcOmJr8CP+mRFUmLf5sB4fdPFqK8ZX0L+lCWwTAbkItGZUZB/
OHGLqrXE7bLY65c5RAEpmT0rZ0IOURnJ8EHGjNCN7xPRnFRloS1fb/YmLtK80Cx+
cZsoO+lptWqa4m/87cGrRifbWqHd+YeT1YzrcFJff5b1UgJyPjUTYbdJSDwBespx
xP21LszhtAvehFJpflVojfaLv6a6evAwF4HNqCk4a6rFG9DI5ApQ4lb5eTG+FsWB
OsP2o8Ogj6gZEoxqSsFI+1NDJeo8AstN4PX0B7bhJcPtsKujEYF/OAlBAZVpMm1H
obvqKOjztYqJWkNgkA9yLDOu8e+RzOugolOgPq3SUbUd4xF1E3Dl09QLrQyUX+hb
+X5L22VUQxW/JAdgEJMuYRFxdKF6pHqI4RvBNv8R8rR31dWi0njGNYN01LbbXgVz
lrNchdeNg2F/prFFHTK76sZHHjnkiDjT6EBSe1BQ9T0NL4FvYznf3uKu+hQkpABj
AAc5n6wnR6IMwhY7v/nNBMVmNyev+VRRKr8+he0pbEGRXGLb4BPAp7KZcdL33mWx
0p+nXY6mWDYqym1t7mRlYyKf5mCkK+V4BQNRKDzRY0U4raMjf5FJ9xyF8xt6MMpY
Vl0+x1vuZ4m/AZs+Gmq8P1QiKf7TVOqBi0fF5Jtd1Vt3I2WVlVvAGzFiRIH25Hl7
gn9dFWvcGw3oF+Yr/zn0H/IdLUPMNO5RU3Z4CfVJ0UZsn7+48ZbxlgEzVYR/1gkU
/SKGLUDFWQnT5UgVbXJ55OHD0Wx/NRABQdLm5+tEzuXpBXXdyhr9OYZ8Ee4aYKl2
2WPi79X3pntzd4d1OFIrEG624qCMYDRFTK+Kb41m3wShhbC9S/dxlp5zvvu7LA/T
UNLjMV370VdUIVjnFvw5GlbazAe8rlAWkymeFgOtppRDax9+yKaZF+SRCFv/qDh2
cd4ZQwVD4PeN1CVMhym9u7uGDEhL/WuzkaaPeu9Jln8wJjG4maQF9RDYsrxBPIWz
dy/CFltmzaEbCmcyhPa8uiza9njVDOHDiIKVKCGrvMmdQOecmHq74ijTdeqx/a9+
8j2ylsHV39PmHP3TUCHzbi+8hRT26ObbkHz1eBch1M7pagTyAHFKrxh/Y+GTSnyZ
MuQ0x94XK7j06eZF5wJhoqF2AWLhTvk/v6gHA8xmz93oJqqYbK3248O84uRcYqUq
g9A8abUR70eiXwjySVgJZV19f76oFEMQ4SD3axJsPkvmrp/+Ik8nr/rNbxkzsXt9
sO0w3fWyCd1PN1qZQn/wRkWkir1uH9YJssURRwXVy5fTwwqj3TzHTfjvWEwq5YhT
E+u+4xxUPDf84ZERCP/C1mzm3WIy6Na10pB1Vs1+r0/0Fv2j4Eq/OzNLam5wYbah
Yb1Ys7phF8ahLbl40oPinmV4K+4YSndIRyfBy9gKa46CHzwOTel8NiVMHTOJVieV
aJ9/F+3RNYwYFXTyLDN2MRtbpT0UerUlu+mSZEo7988FYUj/uRgQLif0VFSqo9MF
gQcBe/65HDUsyt/MqTbqSAHtDHb3EBEyMGtKn5NORCMVQ/9D8l344A/7wL756OLJ
DazPDhiDE8y8gKAoVX+f8BX5DyGkWdcHSiWLAQtSMwXacPE0Ke9JFJqbRP1qsLzo
yS5JepeF0FePPfVDFOIBZ3/jOBqMh/nw6zIybkwSTL8T6w8XAwocHa5XZuaOuRJ5
aPFeQWQYF64disRPYzimvufpoIgeZ3dDZZcUZ8O2T9EW5eE9yJw7+LQLo1S+98w0
9IIYFFv9uhI8HBgYOiqI2729U5/koa4kUHJSPswoikCX5PmQ431hldiEG9wF6Zyh
MLbQII3w3NIHiZLGA+LgecZMu/zDq4JzcqHbB7tJGl5dZZCoGFUKfCAV55O/pdNX
u4kiQgIs1zfj/rNapbyeOR5rhU3CzIf3KVdSctkDQSrBewgdD72rJPZ8ZQxxgUBR
p199lZG5Hlo9DsSe1KfaKQCefs2zX8+zf17wwM587hs6QcFMwUtUTsmEkZ/b6wvY
3XxIygX9cEKfesUypz0TlN99a+888AO/qfJC/WFKMqHaIGGm1J/VR2IQXoKaWijE
OATwZ61cMCYI6VtsN77drnyPLm6MCt5OzpTyjhkQW7tOogjTcKOTn4rKGNrCuRuc
ZILuRwXAF/9PYrIB34E7L4iPjKBhnBFZrQSBtljaAyNcBf4B/PsXLFuGG1+g/Cmk
GjnWckUvlA+cRQfbD6BvMOuKf5m3tLF7n/mNC3kDnWen+8e36/GD++q6r/mbCrjC
2Axs/m0dDFlP8KMGLZx8FdcAj3TOunWhwJeOVJnEW7uT2LhDH7EehZUYHE0X/NrQ
ArlDqjL3bgDBxxEsDynA5nvqRbmWN3HD/WudXhmlGKPhLXg5s26t2wEcFdRbmmXP
MLGcpXlsdfyhQPpshSuP+TjY0joijD+YElyHYpyqT0hQ1YFtoHTrZZw/JoMuTKFb
hxVcrrPPshyjdOMSLUceVNX0h4S1GlEaZapijfgIbG0UpGBDWB/MI2CAm1G8MRHn
8rwgukbnB8sFPavYAqa6oo/bVLTZQJyv9NFJ6R9P+W9pZWdphBh0sb7xsZnY47BN
jDgMxZil2PeLabvpJQNqH8Ypb5J9/G0bzUZtGWG/s+1pmCwYb0cNMjJOPB2cfX3g
KgWq6PmIoOsb9JgGsHdedVxnou1t/CHcmVJUjy/nJb4h7QLayoBQazoyiUsRc25s
03zmtYfGokM+EUEotFETbjSDfESvg7vYz+sews77jrETzh+IUCqBA/cMW/53IjYP
Q+QeWaab3QlCDYniIRhN73m/hT9SJJXYG/IwuakT3rY3gerVDFMo0jymtJAb4PMZ
Ejy6INiaRm6VGcj87lKbbU3676DBTNHCxOZfBuNoWDkyjUxDRx6Jhf7MjH7dcEUx
v6UMD+KOU9Uma+7Zx0h5z1FQMRAitGvBJF50D0aUUHiLbXLpcR3YAW70QKoov287
lW5v9mqRA3T9jEA+LWXywvvFpcIsk5uBKl9tMlb7pjvPtsIaaXqMIeaiPpypuaOC
JVFUyAerUsV+M2oamFgQ2OdVSu9DEScem66afgvLkKpLcDpzBr+hBP+CmpasmUfu
1LNpOgFrSlRgH8QWR/+mmq/2Die0mcAHNBHWGshTjULLHPGj78dJTqcuof/CsI5L
QUWt8i8ofWxBO/S+FI7nVpQak51WHC+MpwhInmP/j6HVIfsBElSEC9AONH87k9Ni
OjMlfZoKAs216UYm5/6lVl0fRByOzvs6tVo/syYgdn/hiQ22Bv4IFgCV0OC8G14I
QHeVnGjBH8w2Ju39nwLpDKc4GZ1SVZTM6uK9KIrl0lkSx7BadCsg1dEXRGQAP7G7
hgMrxEi3xc4wtPUnnXIuyLnNlDr4DFn8BaenZ4Qez7e/O/leOcLGhE3n5e6+GG2Z
DqWBikt3n+njv2QkqP0UbAyaoLTZA1JmJJE/nZaLannIdmQoCtS+vs6ov+3s9mp4
0+tQFEI1bAdO85d0UjKyIzVYL4YVHLeEJICOtXH9Q0yuppoNXQc65CRyV7nMo5CE
PT9NE3h9LNMANVeJR6xSNQTr06WVafIUL/9I90fGscF7V/Hbeo0ubxcWQEwrZycI
K4tecm8rnb7eeXJOpvl3y5P5EpRaJjE2BpcnRe6aBobyt5lrNc2aCEihPB+ezIZH
ypRB4C5UV+Awom5E+feLZiQ3CFCfVBxObzZbhCNZUTPm+cREh+aPImW9LewPz26E
PlHQNpsvRMmDrQYqz+5RWWPZ3SgGbfC4AVUN7t0Zbd2y3lI7p1cCMZudwPvLZVuQ
ztVWB8EJve7butMfvEyUsdw995qLw/IuOJGOW/5zG9mVTEy0tIkRFR6QAYV1MXBd
v5pDHMMRKs855i/q8H4bG9KS95P+XsMRGFvcznTkcigXdLQkn0fx+VSgVLqoG6tX
iHr5wkpXDdjofBPtx+nV4wfra9MIIDZ438CBEEBnq3acZfe1g8lmq3QZaH2s3XFS
JaW98m0jTXgfqD6w2bLU1h1/K9Df1ZzXExCRynVtb+jBu+LCArzn7k3wCAxc1CNs
lIkCUwrU9ZzOqzKtyETTkSffwYj/ewmGhmJUUHmjczqB/UUqMt5c4NAZ2lFOeI3Z
QqaZYt08oyRmdZv6ABTupCPXAUDrxNx7iPQQOAWDF74CkbDY/PpHvGS4E9LMGRG7
loo+kXDeI5xMNS+6iQms+pX8gYyqCDTcGtONu4gAuDim7mDhNdO9czYVfYg1csK8
Pq+G6MXoqOZrC5LPY9WKUpnXO7MTeNFcOpsjZ+W3qJdBoJF68agcy0z+VvyBcPOl
PJ6ulE67nROw0CiCz+35HS1Nkx1kghjm703XS9fxhMuPDhht1PLmEQlrN+bXgbg6
Ew4LA0Ks0j0bXuXQdaJr5CMb2hEPUGd5c+9WdnjUNtM+P8+mN68u8ILDH6XmwYD3
IcudFamEJpENQp6v5MeMnUzChiTqKLirdz5C+AKM1Mb7EQNGtmJ+dVr44lp6A/RK
EypwFcFY6MnAWVy8Vfq3yrU6Ak0be/vg0HzMf9jxzuo/Q7QGe+W+FqZOlJXRYlcI
xwS1IX7T6jX0z+hawJTngvtrbeJBVbu0FnxuL2ZggqyCoJksWt/JlOqBf/W1shiM
URxXSZYuHKdX/R1o4HjyeLqcCKzQnqxz2r7fR2ZpZZDkOffO3BbqAEPdEmI/G8TR
TDf/nZS2+rCc9zYWykAvwKSwvIQvATO4Nu313HXhnA6cEZhfhyaws5Qb2wJf76yu
yM1KP+F/BHb6YdgcxPCjUoZufBRMLtWxIeSIbxg4JdaLLZ3jCtqoHXy+PLPOzfHR
DP8Z467c56OyAc1oAmtTDsDu9JUbxcOAJbaanpBgNKwwGTLLGy+QEKPbOLj74B3H
sld8dxVAd4cyeFqOdZUbrp1U9gdV2k/U1nYHfyLJE3xSoynpmm8faxERCY1N8ngX
Nhbce20HmbLwf5HykpgpqM4/pVXsE7eitCl46LJO/uJckQdOYFJFtlmZy1aljgKm
5FKmCWe/VFAECbOjV7G3hF3AcS2YlJX/r7UdqlbT201aJDEiR2dlFi4ahcLdOeIw
uXvjmBJxoK0OBpdXsHK4BSE6OyuLmND35P6wdqUA91JYr6CcY35m9gwdMviXx7bg
kwYMmwrOUc7w+gkWFFf8umg1bGVZN+f5p7mtuEvUlt0H8f8Krvb4uyvfmYhyespP
3GtReRJKLS/YeAdGONtStkarLGrH5Ws7Hjf8+1+32N127GCFkIG0pJeWYXuwjEDv
nJ65c15uz8LHeMhk2HP6Y/X9OEPq9QaX6bx4mC+NzOvAHC69Q3ELDH7v9wwiIylQ
/3LIv8aUUKIq25QOc+1u8NH7gS4R/x/JGFJOAl7S0WLHkAM+8G8S89b1+HAhAIQj
VpwRi83+rmzHUJCrSrbxZYvMSCY1SR5BXGj9b/jYno3DWfq7/akSrxWAXEYoeMDO
oyxYZNvARYF8YZSw7qjVIqHiEu44KpbkQ438L3qIoFJox3OZHj78MiTz7fM+M57r
fI/f+3DcwkYsWpSQORNeab67pFvziF9BYccuARmjQcwPX0lR7Wze0l94BmUWGj7A
ieoZuDVS8Qo8ASAqnzgLHCgBFgCiy6WG6Tj+5KvSAd1nkNTTJGNU9WesA3zj85oe
1WQU7ySpgzyVT1PSYn82GuAYvAKpVzrYPCe54Wqtu032/2oub3Y7RChNiBmrT1Mm
JVeE8hPy01Ub1SZItDHD+zJ1f0bv902ZDX+30qiJeuoMgDAloh/aGOYFA47bmANd
mF3+P7DPUGlzJ6FENYHe6ADtj1wiZc17OhnX6OiIkXle0nw17JzBgZdbU1o1U9NH
AnLMjZ9xpnUw+t3SoskYOXDc2rJ7HvWrQZpV+m+8Ae/aMFozu8FHpB0Xfqjo6QkW
vTJb6M1NuxqHsFWi6vfjDVA1TEAk8e1/95jPpYaIO4PCbGifEbYdYHYqMyOBcBuO
xd+tBxWkX2T8XMU8vW/A/t6qMhufQQc+z1/YOtYzppFettifeCViL/XdEv5mKSjF
anTXxIGGvg4I9l/zKRUSblfCzbr0Mx4214Hb8z3A0psFYx+pgXN8ehI7/V15V7Oh
KAL5ltCmnMfgOyCbEiWd22DhDgD/7XkRgcWZRxonEOxAydlEy8M0hn/9eNh/Nc32
2Xrb6XQeWof+d9WJqzzUUMbSmgmysrJMnNePhMbPMC8Cau4r08PGXUyfWY3Qz9s/
84RKOlM7H1Kso3j1hemQyjeMUN3i0MWuCnAyE8+fRqOpnQ30DNhYA7UjnB6nXd9F
fpEbbyjLQkxsA3RbHIGs9gLBMwPVdCM9EMNJx1WNs7BB8v8pD3l2cgKxHNsTC2jK
U9OjFiaTIfg1ZPj5G2LTjfL+RhysAbJWc4zzX2QiQ8Zx7dV6+3LLlFmCSfMoHXMi
/sUlf/hXeEWC+spMOa4p8kVFKAX0v130/ZynIU4CDV+fjWY49cKOtEwraYwrZ7MZ
b1GA+HWI7LmWXBKjN0mu32Fc2X/g1kCMSAjEQkKxc5mRmQgx/xHLPmLK5jTrZVWw
AGduodYt4+ZoT3DBFXMTgvmr9wr5Aro/QvJRi2XYT40=
`protect end_protected
