-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
XmQtfsOHnZJdVkAgnevje1NWorSnF2BGIP7cAlteehFufLqNtePzSdAftUbcA4xc
uQksXqT0gFt/t0nbtSAMkUyB4j9GTghG95SvjB4at17k8rlF6VaJmK4wfMtExyiL
oh0v36BmSGdW7qZI+AF7mDUJTKECMLfq52uchxLey3w=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6432)
`protect data_block
Z7EKJhVZWa68vUkNERcVZBLHgyIx8HKoODr/cR6tvroc26YCUSUYYtFWML28MLx4
CN9xcb/1eqyfTiQ/uxueFjzvQgdMJGprRLKnH5LYP7QCZdbL7mB/J750nrwh5Xla
HrwvA54WtNl/VFW4fJ8jMmFDtQURasgj8oY9p59boQ407aqj5bDs4B1MuFGu/IvQ
ADReesFXAJWwP943N/1uKRpzjjS9ht5zThufiuErsmbwr7lIpsIQjYTudfoExLu9
T6qUz2CtUrHLHybIjGELKjpgOjIHycZV7BIR887Jw+fcevHYvoNcsrSRefjEnlkq
IwpW3UGjs2BiAQChGxFVZCGCnngSYZWEzHUsr9BZiCiZ4V1BkcsX2bCH9bjIwGNe
275z+xPHxIpArDoS3Ig3xSzC5N4QlWLjcLHjEumRgPIXkYzsuOKNG6VPizQBgqPY
FCVIsIHaOliIYzoWmUZtQ2dfSxZFuAFbD2LU90r4zMu62wTrnTU/aQe6Oksf5Ubh
V57ZK0XF/J83NfGyINAxNxz01f6wgHAN1ygaKnmDNK+u1zPG9VB0LPQvct5/zZ/k
eTFNI8e3y1ao2uQDtb/ZZk8OyFZ4CHwzZVqFCL6INpqD32SLG/kacV76L7Pb+Vxw
VA7rY1vLOV5XztXieUePx1IT8LvUY2Oh3QulL7stzJtdZhpT5SO176JEpF8vZuq6
79VuGeVSYRxBf/pIn8Z9nBh+PO0hqIDlf5Kr7zULvJ53eTy0t3PVmF5EzW6EEPnu
26M0KLmQQvdfmHXK5Vkdgizpzh+mrGpvJDv34fj4AmTbRZiL62kKk9qItw9h63B3
8yNewAZIC1d6JuOpKouSjiX2E5fHwJ0x4AzqtCazI+vdScbT6M8OS+vB8RUPnImc
T6+k+LYY6x8/mixY2KsSz4sTxNxZvgMW6CRh4UgCgT2TVrfx+bnvlbS39+3Cl0g4
WENq/nDZ2LdoGPWtcvGJ5xaOki+1FCB+odxuhxTXXY+eNj6x4DyplqllOrVkwtmD
Zu9FbilEBf16D5V68vRtrTpdKznm70aaXyu7W0GosDHtzzCFlzSEwH/V3+B3as20
4BnvMuHFcP1duDGge21CsTW2U08RpfQsd8HMmzyLrF/0NOrA7We1PFVrmuIpPEle
PCd4KfeLftlWjfuorSkIDdEnCzFCttaCKLo28NMmS3StKHeyPak9iTlZUWcC6Kfm
IkeJ4I2hw/EO6IYwBEwaByrfzKaP9NDEFzCaLNChI0533cDmkxvYmwkmZCdRWCST
qP8o9Cj0TP3PQYPwRNA+KofzJT8XHtoSaC5ZA/Zk883CUY+VoGNsZoDk0a438iP0
aPn/8oEjbtLyWeHCg0u2z5Livjq3z36PsK5x/kzYet/r+kd6T9vXFFo9SE7Zl0el
6g9ZsdsMSAnvbM1JjTigGWrJS9241D/+wAvsqFWHRTpJM5RtwHAOdUZFzcMTXu0Z
FiZzqW5KlhD9M7q6ie0aww+25f9F9qsgsTYm1Kojo7GTK5ZlfggPAvGcDnUDtLlz
yVFXbMKTYJQbpYhnowQ4gzG99WpPRwRoFZKReqEQUd6SnLxYoeALE2mrlyfEkQRY
YcJUPd5qo+1m2cxUwpjgS8tno7yhJR5OAs6fb0GJjccJXOot77Bo+lzorwAAkjzr
SKC/VDSwKTp/2hOjVobtffzjZrrX2JY0hgwyeYUsFyFEEErmCEvIqayZ07zsvkiN
W0vcEzVfNcRl++uFlXZkP+B9oFWt/+0sUQtELtCA25M+H5/A9kjsa6DJzbk0ByQB
SHdNAmcQmDd/7kOjmW9uhW34P+m08gISwSXVAtRapeuObjjmV5/QK/WZPolfZlKL
IOLnmoMv1igNTq7BlKME7DoFCsRJTdx1BN28oLLb/1GZbF8cIHsrT8cuaKSSUAUn
TxabFX3xXXkRv995CgvSlX8CyKHUQRYsLmX10zEVIuG8IUX/YGysi6jqpE0kar/q
DrNtFNDASD55LkcK2XIm28nX0HpxLm2kKVFqTUJU2Q2jSmSrswuzTAeu5ODNqm3X
40ntvE2xLDvF/fmR0qL6jT36j9JUeCWNIEDG6MMSV+PgBszwXFDvc5341ewCAWQU
Y5wrT7A3OgpXuJg5O5C7Xa2dWIehSn40bv4BBIALmhTLi2jvdT+WE8v3r2kJbhzW
DNcFtx0Kk+AUU9madUdCYmsX0quCP6AmEI7CjH5+zRSIbZq83A5xLn8h1jnJSQXn
Ve0U3pYRHYOHLjouiCclUgE5gyDvBbVok7Q2WwNGU51AemmW4t/VGcTKtGkOLSRe
aBpcSgZUJ/AbGHUFitI+UWNJ5f3gpy7nwNzJJkhLsLSIltvQAw+3VKur3QWhx+WV
eBICHqE4CVXaCc9UESX+gy9ndBzxiiouexBW0jIbE52FW/GvkTErSLoVO587+6uM
+sSVzU08S4dIpZbYq2Ps8kBz8CvD89Ukpsrz8NgzncMGbLg+m3fn8deocnDtuZXE
i9h0FVwLt2EnAeskLW5CC5RgC0PNRRhB8CwNiaHRNgVoc3ULScAUnQ7jx985Vscz
Jwd1FT5Kc/d0TMtM1fZGASlaAoLnjCPU6OyvDvLz3/CgmtY5LBCC28kCnkQWkAXP
clQ7Onq9aehJANF0FcOdbZo8uPvxLTVEIRn4b5hHbsMajcpkyuKa9qb2nUG0bvbP
/JHqjPs3nvlkXeUAQEcN6CugyuPyVVd/8XXqokxBdsJNezvssc5XBuz1X8B2OChW
GhBUWngxWomDXrpOZWbnclkwMjTPf34wUS4AiiEfSCId97bm/siAedx/QQn2VPcW
YLAYOPROJu7XN6WaIoF0d/KAyuXp5BaPU2gWHp57zNloRtBNES51xTqcP5iiF++y
NI5vv0k78YO/6gI7I0XPDGdUzEShgE8CCcjk8vhqvcUbh+g25gCfBzQiRod8J9hj
PopY0rjqm3QUxLkRZRuR4noSMOHCPD0PwdEZ0Jtk4wkyJG3FwW1LELZUXWHtcgOX
gOZyDWiwZ0MjJ7Ns2+QaSV7KDqSziS1cD0KsOj5zXeQZgYSyc1WIUq7ypo8eEtiR
nClOVFD6TZrHbJ77XmXxIcEt6sEoyn65OSPIvj/KmSzPPpUkt6plaKzw9sPQKZGt
ggV/1Xtbk0K2BBnlyuxmkOZrRXmjUteROj8Hco8b1Oeh6OpHVLRzba3xJm34QrzZ
05hrm65DZEVpLMWFVoTCKGhCE6+YPodJBBxE5KfeIBqkO7eu2XZCCeYLADs0iLE2
5uO7cCKAYbv4223cuQUYt2llzezGucvlbHkZ7Ru/9XGsCa5Mt//hjXKAkqNT6Z1o
JfTDqqUVC+WSqbcLUMfMEAStFngPXlwdCTjHL7GDVb8S+/2pQ8TgzU4Wp+PkdWP9
MCHrJz8gdo48HmdFWrU9NKUPaSxdBBkwGAzz3eMOijjoiCd2ak3Em4dUpDTUNiJ1
3BHcbDMF6wpQN+pnFLUG7m/yG5eUCoI8P92DtqWBysERIaqqNftHKHNWzgKEVa5I
W+nD4JVJBHd59cQUdO4ToGYyvjU3yBJXcSWefHT0QbsNDPDkCnI65Sg5S8+Hk4QY
3bpbfK1dPmwdzO1VyOVgLk+et1AdNIt4l3VeO5t+bs1oA787Qk+EGDW51M2nUPrc
ATn1XSsx9Fwj2fYZF0+TUbTp+pSLeEPf2J9mRCuNLhcvsNV/ckHyCSUa2cCR4S/y
S6ZTGGZObTjtW6H25HjI0R68EfuxVdgZSRe1U0jh7iuS+pMXxf1xH7D035JUovgK
oTKT0vaaMHyAsdH99MXyIyPU1D5k+vjcdGRW75c/KTI0wu1euTh2L3GdcCJtxHSF
jjgp8d42BhuoiivcGLe19/YbplmgNfaKrUQrvTWWG/QKsfHrdX5mxfHU3WTJ+Wcp
1O6r05dGHqttLt2BaxOB3YRXIJ2GB8NGI1+M5RmQqnWRPRRPkAoVM9NRAFyxGw/p
FrEnG+YrhXkq7lPPhL8ZR3oFQG/bHcrXfm5WXkfdhUpYIx0XfjtqYyU4gmpWLwVW
iBb1PIdhxlKMf4WAAqtonoQlrr/xUK+8TV10/Hx0Tjgl9ichTpiBlie0ZG/Zq3nU
lGAqzkdzYmlqL8p/aqkHt9dbhUAvYnnI98k+gYUTdr0OfUVVciGyHnkRE8fNak+M
RpXnd2Kps85FQnEHm9UY3u4JUnvkWJvskiW8+BDFHwqolfhuCEaTPQKCIWNRP7t5
EIiXV+krwBx03fgDWXCWTY+E9YMsr8uwsYWalRaigd9nHJZPXMvwGm6yApf1jBi7
1pPAgj3kN8olSxQc8NT/X6aOSp2hqiNVRE3MFmHFGQUjb1gCPRQvnwzRAXlI+sPU
aqWStQ+SIs4qNgLAJ6xNUtKYeKcFKl20XriQfR3vwGr4M/5zYHveIcWkJic6q9BI
P6bccCDVNRv4lvB4TVmn28rGWmZ+vfZzlZsUFRGQsrg+Ke8jogUNnLMUPAxzFGlP
LeDuGMJpI4C4Tpb/st4OccOIHX78DYZMaN/tp9qsTbAWSd3CMGJOIXJUNX3qXVRV
FXMr2IqGKsnHRlr7wW0Q/HTvUKk4Dmuyo/dYmz2oPiI7hXYWKuA07If8zJWLwitc
+sNhwPEEVqfLqCVhLdIDNBy+R8Jl2CYtcK10jEFzukgACdO4Iv3h6r+px1yoNN6G
pyyXjXSkOKmOBHfYBLpXHCS8A6Ek4Ag4oM3Yll2Girxh+85Gbd6MS+M9OjYpU/3d
jFGArQ7oHvob28IIuG7rMtaXSDBVasDNKVFV1RUV+8rrZzJRKKuGLXSYJ8RNPi+K
mlKDaLkoOYQp0ju+W3AJze1VzbLf/NIRJghcRtXRhMNOAbqWk0lDNKn/QkpSaYM9
UZC3pboXrXzpioVYnkIMOWCqUFIrHF2sCWMg1+DzlI8PVTolJEKEb7t35VAeX6my
U5G30UmHi9uxaG9MRSUrPoUuAHEll0O5H65jLww8v0JmhgezdULVbPtmzwIy7jSt
kSWKEtAzBvjJR2ObOTt/yAvSIKbdc6AAKEeUZ+tsiCwA/nerLIdLWNSlX96wDKMM
RAqtLCX+knbMwPawsjVZSrgOY6Y+SdhHn8NFpHdlxDKlhQc0tffh1ku5u1kCoQdB
TZ4LEyhTMSO+xZL8i0kcUx0VbWSiGBjFdeFCK/O15r9tt8osZ0zWzbSLkD8L//GX
gVjpOJgA2MM7owcpMu5JuTteDqZmJT2RTmELtFCKAP6h5eaiGKTmh0+bKekGnwCI
XBL7ASBJXcf8aC97hCb5NqI+iANM5w96KxMqo9UeVmRLjmlFv7TItlBcKV3Dn7f9
JvtaHbjRIotIykv19weWragUYCTwOn+BCXYo9P34dRlcuhPnSK96qsSMp1yumExy
YjpagfaqGGYyImG+WQtOCa6Va9Hg6RxH3Qw3HlKyaY+PpMyBWFGpMWilCjcvCvN/
O5KpAlRNbhRdFtrz/bTAaCZpJET2HKvA0HchKJG16QM3ZZDizTuNbs9xcM48+Bin
EIUSs1mUuN7HzgTCcv7zcRlnK7Z5C8MY2GUGOQwYFUJzpiyR9YUXeInQEPh86Gct
YUXWRulku4uZNGqQ4y8+UsJZ50uDVKtcr6SNsBDbVG0o8atpV6tfVC2crKu16Qr0
/ARA1ZFBBR46XRd12uUpwLghoHfwlK8rXnRCkUwntTSXScta6Y6ymJDl7VYEfagI
5CnnrlOEOQcwChqTvJMVLHInz9czdTuwN9J+m2NezHw3p9qbtRP5Xuimyixueq0b
Zx9zzzxUOiDix4PnSx7dfibApvSOKfQtEfGOfGDpbNmGzQ+cXoD6bmsjm9G9IL1V
aLLnJ1QPA94wYx37wGUt2QVVLFLOG0WIvtjs6v0dXKg4w1Dh6P9M0qd48ythG92X
7FX7x7JLqQt4oxOyFLojh0T0w4Dc1MEvc0bWxc58Pvt08QQPkIhvMcJwlzHYjOcZ
13HDATkQ6B1hlYMaVaZDSgjagXsDaF7N5x1H5hNLUGRDmzik4UHSRKov8v9981dN
xmkYSvpxAOZYW/fUJI1I8JwW+jfsRHpCA7MR5IPLmgC+kMBC9mLB81f0+gpE5ldD
MqIniDcIndEtWQmswvOUOaUQ4Hp7kxeyGmWTEgOE+5bqx/X4aZzXnaHfuBWM8No1
9E8/WxRXAip5OSLF3XByRsIxKM/q5QLAcnQ+dpfOgpGQmrKG8dOFQAJofB9kAxB0
4jxD9QA+4QZg9tQ6xGlMH4JHyOjrHobGhR5z9n4PwUnOxgsKnfIBTYCVkivdXDld
7YJRE1FCwG108QGL8fd3kxlf/wd2cJSoaVbsW8EK6iFGO+luz4IGXA2zMf85yZZq
4CXmqYjOGl7BwpejP2Q8iIQ+bO5OOSCx/NxsMrJ5+BXK/DCETJLYqRjZRKTEja2b
LDShh5BaVkl7EBcBtJDYta5XtNDm6LniAP+qL+/ppFgw3Y4Xw188yIWXicw4raRn
qgJ8pTm4YrCikzIQG/+RKqNQUWcMoGRle3g0SEUhoR2Rj9owHa1kMHa+mqp7CG3B
eZcVbYBKujkYlM4AY1c2mxh8p0/NJ2nlyD0RAfwXF4HzdhbamK/n+swMkK/VLZ17
ajfvGh58n+ZyWCFjGVok9NI43NpzD58UWXgelNEiDaAHsrWVhm8+XUiVGUg+eyeY
a9UleMb0xze+SRXl6Apbs6iox6zvkS+7DxJNqIWSMCfhVT8fTG55l7wDv9548jqV
BjOMBfKoLcXHcPYhtBTXoeOEc2ODtE5GljBM3xXW2QLfrT7aZbfWHMr5q4ptXRSg
8q155odYW4WBMwTeqH2Y8vDO2z4knbhbwoWeIvogQZOFAIh0M8mmKO/B56WahlTw
HPEonNTTZuVi6b0GAHOntYkrKDUQhCEPHaihTJ+R5XUK4T7+1jKKGI4dfzRgYkbD
7hsMAdlWG7IGf3kGSRcEk91CX4ox47cgNnjstn2Q7O2QEKPSqVorTHBP+XifUkd1
Hcx5evUf4JRVAeXvoGkA47rV1cjyHz0Ld7i+5LTXVCkodTYdhrBGnWsAKpxyBfFo
Q2ZzKZgWv8JCldu28tgHBPJkW7aDYhqvRsCxn4ecMah55p1SQ6cNQ7hYHWuivD79
XDZQvG6WDjhB3vTKvc6El4L4BPTanXVjL2feiCpcK92QPsLQOTvTFX2Wq79BhlCl
Go9FaKY1N0NgfNA8N0k9G2Z0l8tTVqGnKzmfZP4ozDIXnMVDRtbQySB805iUG8uS
RSPAa37+l3trdHixd5ZLMycANiGBq6iieE9g+G+D2MzgpBAgB3glMllyln0ViMDt
jjJhRCPzF/P4lkUZU6L1cCgqrAq+G16UbyKkVVYFIqNcmnmZh/2kDMFZ1EZuooI0
WfB+jeC6Wfb/isj2djROIPpeZlPBLliDhyyu2SUuuRWxWXBspzQgE0TBq1wbR2e4
NO7cmME65Flq7VFfk2K9VrqqwhCpZyB7OQ3QACQx0UEPeqRjAA25Yk5hfo33faRk
vN5sOtIncVsHlhay7nD98uXuYziPDN+iJTQm3mrNPadtj6Sg132kp/2kxXzMxt0A
mvX68ijWQFN/9SNth0Rt83KFvQNtfYNNo5uk8aO0K/5HLg7z1NagoX610QFSZecO
hax/tT417PQz1zIsGtfmzSBcOTZvrhY1dbj2i/Q9qdAmfmtCw3BTlZSmaCxOJxCV
HytWNaBGgfbGSSr44wX5IvP9k5FDi03Bm61DP/EjVJpd72DuohJNw1N5BGXQ5op3
khnC5vXjadurj4ei3POmA/SNuFh+VOYDxGsu5MHOUQ/6no68iHT94Lcft6yKmQB/
IiZB1mxhYjvEe2+khPDuJfoF36IdL9lYFr+rlijNSsoIaK0dg5x3+RaD18NQIMdo
vZw6DKGoV7x9htEq8FqhiPbTZ0Xk5jVI4IrgusM1Ve/1X3ZMjRzSC0XpEIkaIWEk
2tZ7aU9kDy+SVRe7hXRP/e++tPqLXu2QkYooUwsIbMNKsg8/hLRK2mYAODi0+bIE
bMk/M0eiDq3rsTTKYVow2l9cB78Rz7Xqdwqlu9+VCg+UtRHzg1RFbzZP7INI8x9y
YMJkg/BwsZoJf7716YGNATjUCSLka1KLmp6jFJIAUYoaFPVsk2lG9J1qGQRRf380
fpGf9RShSrgEiPbYAIWHGkf6HlXfMeLnyZYD+mP31CRJ1qNYHMr8XyLYbOVsSZ25
8gt+cKefjXpr6DhIC9SUwZW0ziuxgeTu9oWJPlQz4ugOWexKn7fp9esSojoi6rVO
FgpfbSH+fp1GfmRuKjsJ47wYtOa8hnnJu6ilOFahm7MZqq7PHcWLAowke1FZ/QLZ
ohaeaqN13sXsfiGTxgpo+8bg8C4QD1LM0xCdnKQ+nfjR3A0zgXtAFPlT/oAoHZ5d
k2HMNoe7dktgtfwZBRgHwEu5F+326e4ndkab3H19jbKE04YNiL8zXd7vNDNdAF4v
wS8vJD5H5w5OjuTYKGV63yMpODv8IQhCH29qM1S4wIu5ccXuqVLlzTY1kpJwlV7P
VU7i7cS+NRncCDUvjWfwdpttsnkV6v5pZrzDMaE/LygH6eBO0U5JkBPA/Y5MLNqY
`protect end_protected
