-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
g/lqbRn30lngb0PxA0TeW3cimSH/ca19Y8PAs8DFhuINK8xNBSi2Fm30f/zC6dYH
WH7J0+4CDh3R1KwSQGIaQ7H1oPXel/Un91XfHGl/Q/ldhTD8N5wQArKK9bjv0TSc
OmiHA5SCiF38hU4uJbF4A/1gNnq9Jdzgi4KZiaeHpWHyox6qeJoESw==
--pragma protect end_key_block
--pragma protect digest_block
s6/noNA1x6DU/J/XyLtms/LvKxk=
--pragma protect end_digest_block
--pragma protect data_block
m10Gda8Ouck1yXuSVaUNzvcbYlwMx+080PJjQ3u2kJ4hGsbF/rJEz67wBGntFrUS
45BH0xDoiqY3qdW1FAUQqgalCjbjnJIwEBahtdJsbpOFT5wUavKP1bP8tVm5U50p
LnzD7+fethl9KVmr13W31AoTI1GCix0pzl1AFGhJE0sKfoyqFz3zkBd3tj9v416l
f8QgKxEOIGXB+YEsWBAc3z2KPYcjeL9MxGlCOFZ6hWADFpGPaWygr9wtp3yQ9ZGk
63dKzxmhrelvsXS+vweesKE3KoPtPza2huQ6TzcbtkbG6e6aNXN21OQfL2tn3h06
Md4PR9bSkwEvvcnvlDsrNJcndWxJVVmLhj1PyS5VS5dF+6gknN7icgPZS9eudl24
in+G8z6mADRXG87a0GWAo/0Pr/Z7vmTRSM/4OVUCqckvx1JoPIxrMZMm7m2pWrtI
IbzSBHEQXFd/1f1obqUbD7YCsoiI0dtnquiwhAjxXPj1QFaOZ05o/LoI52C3xI4X
m1MHtH7i19VQFUO6CrkHLfcv5mU0tUraV0Iy+GRiJQ0PYFkOcHc18KO9VAb8Nk2G
7//xP6zqgeK9E+fYVYUM0kvIutB1mwX3sJsxa3t+JQt2n+m2Ethz4i7V7ra631GJ
4ii1wnkeKWVuIywGPfAesFQ8pzVCTcnohrVMdT6UIF22r5N1yBS/ugN9/AP43C8Y
DMKNdu3OS7A6H7WuKCkkc0lpjxBsX3LyvfsBVYJvkK+Gzhjm1+ffj+DUw7k6VSwB
nAdQHb2aDpG6mx5rAx9B/8BdWCCZFJzik9baPWT0DnwiZGwCv7R7g+dSnnQZ/zMg
ZywRR6tvfawfwv8fRXwS2K29WrHrtRC3PGFZEZ1ZTZG31vs++9go/GpogJ6S4ynp
ajUVqW5pYmJFQv76av58g3la+s2xSVBLsRCb+n+9TGSrDTybjy0i4pC+DHt9PNAo
JOZF275Sq7pq5cX8w0HHnxmTq/dGIVTzu4jwxwpSLZd0mdIG+Bp3R5r2+um3Wg0P
njn1d3xOR5KHA6KJAJRd3LyVyiSunlDbvkOEfe4rKsLCgn+Z3vsYhzj5I1UUUH07
5Kw+BAkE7I84blk8UxV5yaMVuc5v0KSAUiorpLpVrgRKpLTN69k4xGhe3+cQZtm4
ZqkLF+w+8z7bsDMMbXSj0rhQLktbfIz/ihMK/WzvPqhjfWzzrdn9yxzrwSQZCDvC
ZxxaAfBZq25dqs9TQZESrVXDKUvkiaZ5NoFEoBQNmbfaz5DhUp3bsS5fADjDhxSN
Wr8WXKUU7QxzAfmJk7B7HGYMFfnjzWjnnBc6PWwspp4QF20AsLzpg0zAmVxmuRxE
k70Awm0dNVc0UpWx7UI5e3sxxhuNW7ojPm2QFNLWfHyN2trRcC4IBoLrPWKjAxdW
JCH6MCI79cPg4sOqmppvYJzOiYUkk+gzGZZsgUeH/vhBbJb4a8/F2zG0w46CkJ5L
wUnqGH+BuY/FdUeyEpq/DcJg+ystX6kaOkyRyFytQXVvOvA170bYm6MfpHsTS4ll
722z/IxHebeyfNVr4H5HxEjR7xUo+14kJ7/zoOWJzpTfac9EMWVUiUfchAIOpw8v
04xLj5IUxTScaTM7DnItp98HkYeFaqX3jB3W42jnrmuLYQFUUyI+qxC3VWJelKsO
r1rpAnLQLwuxd7TiFwoWYC1BU4f/ZKfjserVHjW7F5gdcmO7Vy1V3xcfzRj4flv4
cCR1wyqIwSwx0xyQRs9LPqJkWo+X07keTti+hBUr55aoo7aW9YdWFdbTlUSRSlQt
nYEDTtyoAM3nuta87r47KzZ2scCjRDBh9dX5mvWYr3ltfLUNVadJgDlNrjnVXCbX
oXJBRQcTIzUbtP+vAdbN6KqYpXJ1Ibuo3zpu0THmjeYUHIMTGqkJTnT1rlN6LUTn
LtbB8XKprd4jOu1uRxyyPdWu9W/goUS5oLVVroDe95fRQU0o2CWocFukn9Z0sfDG
pinV/Z4z1+4O1tShrfeJbscck66e84IjX/d+U07TRGL2i9aFsMqyFQQOGK6eEOQH
Q44b65PzEuJraBRgLfxUmRO2PQQBWVf+i/6pIobEytrLWWNnsUuHc9oCJFt0+bW+
d4KANhPZjqP1o6LF0WK9XEJr0ohsRwSGAVhq9JBf+sKVWXTPI0zNYu2vsZgXsTLR
Rb9PtSLuVnB1CrPLK9uNfOlnVLFVDmaWS01zoqciVpeIkmvrLepUyU5f7fKzsqW7
A+tC+fb2RqTM48UL+mxAVLdg3GzGHZe4Jcrp+jQ0znxjStQZiKdwVVk2agfd06HU
yf9ICMOSFMgHqjGNRVFHeXIXh3+km/SsBnLXK0IzW2rxmL3bgMyZIaWgWPmLIuZg
w30r6na8aNiHNE3K8hTN+IxMpNXtdLqDU63MB2N9auUJX8jWHkrVspU+b0+/bNrf
Dw80VWw2m1iBK2j6lUx86ao5BdjMP8ierGwlMQFP38DAVSeVJQX3ct4lkxw4Cbl1
Rb6Re6QEHqy3qB12Bnz+YBhQPLuixggvpoLSUNtuTYeTxKguaI5bvxlhHRAmqd4e
9SioR1eZvzxDHxrNLSUEh++11ddos1crWB69XBz2WiLTL73TFqQiHYcPQCQ3gtMz
PdQ0iqGO02Dx5XcpyFDO7exS1qylC0V86sTqT6kW8MSHZegaifobm0aENaqqeJ6g
3VGZ0veKHvaLGauaUqf7Spr6qdTc+j2N+LFks6WY5MFEce2LYUpHWz07byItXf1M
Y60iCkcDIjiECOP5jm25xKqpe3PEKXiBLeaRyPRRpFhByMhMDgGj/he03yebtx7W
OFleIck6vV16y3q1CoONVongqTcViJAysXqCLmLWB7JFo6TCP8cQszSQ39nuEnXo
aaM6GAxHTv938iQvINDjn9S9Km3GKziI2ZSivrOufz9lZtAd6wqKtcVGAOuTznZI
wmhJd+Pnrt7FDvmT3SLWk2yPOY0o/STgGKlYnen4xGbnaRiYqxxgD0Svbl3xL93O
LfXSOFHzX0H6Q36BWsRNrF1Jwif6JOrduPzGkB8CikmgbOCS0BdTb+3eMVHNHhjU
IKhYjheGCi7gXyWhKv/E703GBizQzFj5DHWoGqGhK+Z0ds/Fj8eIMJBKr4UWjW1q
772eeVulFyqXTBF+ZqP3PFktVHXpIL9aFOtXX2QhTYgDQzfB4kA4FoGKsTnXZ6Fh
JQpHzNNvyNJHDPaOg4CzXO5zsGWpKk1dzqZMcb/i49azV8QuXVIPRuUZwPVp07w7
Zw1Ty7vylHd8iD2z6/qrSVcV3zxQem7mvw7RQeA7/wN+Zltsb7o5/udbd4dxj+gL
zzUOaJl1aC/Xtancy4euo2KDNWWO5q6ml88R4ZxSTuMc5bwjcjD164OM4i+DqSqo
Avr9bYuGXto4NDaLwYxveoQUIGLroFKK2C4WkVvEy28JDdMgQnqbDRRDqvjcZ0AZ
ohTnCOFUFDNUO0zWuYRfnkAnn0W7/fhSh7S7yXp75kBkFP5CqDx84TrOv1eGSdBu
80O7KvEzkTM2bSiXMsi0dzk2aJNqiOTxutN9ypfniGsIiPv6QHgGZytW+Ynla40k
6U1P58dEKMP6Nl+jiuI0nKh760/s/EgHoNzPUCJEpnYGeZxqFDga+6eOE8HVdUxz
ZHbfinv6vTQ15cKTytO2x8D3CdUrHKkxAJVTKYNAxP4y60Do0A3I5jgDtuuABufC
FdO4ynMbEN2NaLDHT0oK9lGTBD3evM7TFQENx2W1g4JaqVuGHfvcF6ekmrymxuTg
UXekBIXkwLrodLzV10rJNx886vGwroYJiGV8/s01raAf97K+IPo9vTblOt6VBMmZ
DpOHfXLwXFnKDwi/anqYT6O6BWvtDkS07/2B+DCqnqJGXD0+k6TmfImXyzOIKzLU
br5eK0UQPnl8DI98ivgtNPaKAcgudX5bvmi/Qk2e6jpU1kuxe94wLUuI3Lz0GYG/
7Dres1BuCljzZtmGGWqG5Abwg74MSWlasx/VPLnfqKOq9SAdpRnF9qq4ZOui0H3u
m6OX7qh1UTWs6n+hquMHXX99h20pQeXrO1A8Jiz73mwL00S473HfoKQCwBBz3Nn7
5fV/fIRy/4jDXgQbSl84Cm2bY0CpNB698CLAzhwYdcmsbbXws+gzy7J+4xTO2NZt
gXnMb71A4LkWHX8OXL69N6AtC5nhTUNn6oUycSf997D2Ncj9iTZTUFxW2go/tZBc
gPt1atsXi9AgOcqIdDwIqS16eR8L/j/EMoo/u/6X6Pn56Am/fTPi6cTmmm30T9wy
uULDnJ5EhSF7Q4EMiQAjDnm3p3BQj8rG+9iXfkC8LUEtx98OZWLsjJgzM4S8y6gJ
rJgWBtVvQ+tbjud1t5bx+jKDYvTTlYwI8vlNCXf86472pGYRyEIXRo2JEa7sQ5oz
/ywtcwdXfr2QwDNRDIglq4s2Er06ghpnQVOds83e4110bpbL0Min/MhYu8NG77rq
xvgil0cImB/AgN5l3irAC/guPChaObDL/ENS/ptWwPRV+fWBdG7HheJzHAwancEV
2PvzvSGSH7+hmumLN63qKrTqUhRycb+h4TcTWHwj49RTdkPS0ckDby0kFJ2ydvRo
+/pOs4QNaTIEUiOg2nZBfZkgmr8kWnwlZEQISbUWP1MefpS6Ut6e5r430y7Chi5I
13QBon/Ok8jyx1V8pgI8HOe8ypd8Z56lPh6+Q48fYPVFM0gptadh0bsZznk1zmeU
audhPAhpTCpLlO4gNUcab+TNKI8LRtuPMt2C85FUb6fAVC7CEYETOZp8h4gUwsUU
fX440R6jeTHyOy+Ddbf0e53OcXr/Yly/LGP9BlbqrNkQt62KXwJY13+ds6xsmy4c
Zf6ZtHWTmX2r1oH6snEKeAUCI+6p/IyCZqplFkq23pEhn3Z+yQ9aCKXqFDmmX98l
psezDzSUR/kX0iXchdh2HFEkyWFNl0P4rckJChnkauYoO2BDNX4ox5vAvZkeu/tV
D+N+YvERJRr0+B1hZsJ+JiqnmuxN8yWPhVBCMNTQRrJbgKRsLM/DQBFYjk8myALr
V+fWSbJAco6jV1iFLeL7P4Vfs5+PKAjjyDDSbaoapLMlLGrd2JP7Iw48zESuspSw
hzbPN05cPzxldWZmN8ONYd6SR7Gz0/LSmCNzmtBt9TUb7HxbH77ye0mIzvCApi1p
NAcIr7iwgAwXVsgPJkyp7YALJ7I3JZtFABb8mpL3gn1+wY+Bpxxp8dM1q3gxRHRE
I1Owg8h+1J+DJY6dzawGgb0bME14pZfBcko01SxtCZUrOyJoYLalUsRWkZW3+82h
+7Vx1DqNG+PZ5GoXJUMwPMooXYZ0mzBrV1Kmyp+CU9wUYFpybaZBwWMgyfJ4pNgz
Yz9WBL6p7fJIa9SHHZufom7iFhshZb7JBbX8iMn/ZHwaxXfR0MCy/qVPWRLYIxa+
YsZ3AcLHZe+Uyb5SRfL77Inz+2xdA2t+bZ7JX2yVIJmdXEi60mv9TDj0hbgDlHKT
E6yiH1Zf9Ju3i+uy2dcz0aDqjh+odN9BqNWTXEuc0prAG3rnNYrhS5pB6pjpPX03
hZ+vn8SyW8hP0/kNL+ribGMA7KaDs2/VIXA3m3ExOUAkhYiu6PU4PWL3RW8jRoVb
Y/nJTJRdp9b5ng9Atn5YV8fJc+JP9gHEVzzLHKFkPJ0VfEucrmV1NPn/2sMdkrnS
HshXGbwfkL6RsQYSPlXAXiAotpg4QUcyyDTyTYVWMjgpO8IW9Hb4ayzfm0S+jw7z
SVe8bMWRVgTZpdWOzS/YjgEhRUXi1qkccVQbsEwgIFwcXQ8UIc5G3h6Fk4HhgSXk
Lx/qlrc225LM5Xj4uRxbRHZU4imM0cpxdc4ohjZePPN4VL3oyO2CxBfCykPKsYae
iaLPk1UZHcIZIU8H4/pbsSUHk1B75LJlkJzhRBHJr2mRaXSFTBdDrY5aTbQKxYs6
XtrEAAhZNvxCnBeqznL/2VeDFtU53+3j4wv9uJ0Fti0ngYRCLHu1/+ADQwyHyKYK
+IPBgK9zIDbEPiT2MVfpEOh9vQF1g03UTvQVirllwzzLc839m4tUOx8MCqlVnBZ0
rwrz3dmy3f44sR6/9fYqMTT73Xrk2Susi8i9hYL5szgTM4q7WSHuFYkL4wL8wUzp
8M0R7Tzk7BHZtocBtTAE2RbqBKhc+OzAihvMrE4p3ymNSGMi0zkV/7fP+Q1X7Y4h
5+WFlM3qzDFVAuXjgPM/kwNz6mFHFaP4S/zEpL8EdsyguGxBISp+m4DdkNaOFtW4
OJ8bn+BYfE3jok28w5i65n/PCComZBhWNk5CEkECB9pkJaBR4g01vm3D/fpn19TB
qEn9eryhhykqEyhIKBGhKo51xdtsQ8V+qVqRMNrAu29eys7ZWYzkbMPl4QfW4kCN
0wAExJHdWSOAOmFXErAJHGbA0r0KnstGQ4uBkQsG/ZJtxT1VCS/i1MuX/CKfBQ16
lobUs0TMNON4oHuyqOQGMYmVSDbGcjck3MRMcUMnAMfWxfVlfQpEYeC6gEOCdETJ
N2RNX5r6VXEr2FkT3DH2mJ/JaymmImSY9Pri8ZxgDehv71S3W6tcKE69lv1cQ93T
cDu+rxckbONe6kmIK1i226Xp07lmpAg9xqbkoLEkzJKyUTno9tquLPzztduHlF5n
Xf/gEDoh64hJB6Jf5uEk8mPy1MjeufQBejUi8OxvlR+CIUT6KxEg/xAeizHGsigo
VH3yU7g/OyBL9rgNEQsv/ihF83O+AVrqZZw+fKI9CMDY8uKNTyRJlxmJeZvGYRMC
FEDHSPH7ReiYG5aqBzZCS39oiFYKCD4y8tnCwF/4SFyyu8K/bHH86ZfYcu1i4kl1
HTow2lEpbVaQ5NtX/da3wLFkUjFwZBdymkv4Sz9vBo/GOe/jrT4GmS00PNvDN90T
avgB6bPurwEFeLtSHbryWDeKrdS7X3v31IncQJZaTIE1+BF6zhan0ZKT3MXGUAGK
YwBfAa2LFVFOJt5fMbcVkrztLiKRKURFW6cVLa0FeGKUYlgvPjNejj0QeJNlfUFG
7IdledPEYP+HCvq5i7AgUO7uwsZEylAH09FI7QtQiGTaNZD4tvoeNoODSdrg52Zj
uiipgH6UZ/C3dXLnoMnN1y1GnQ2LAhh2x1PS6ObHiKKDiuZDdiFSh9vnl3ZA3vmW
KootO7kNQxwJZUebLOV8nKJUgL/f6CF0bqwr87k8V3E=
--pragma protect end_data_block
--pragma protect digest_block
5DJ9d2ojCmateAWStXDJLc1Xg88=
--pragma protect end_digest_block
--pragma protect end_protected
