-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
a/OSvdh/pUtrnQGEpmwEiIiu09+Jn/JOlWvt2C/TtzXvMyCLITEK6QwhV890dmta
gtk8v0EuTeITY5clOLe/FGRES+J/3mXbyb9XA9v5RCZdbqh4Y4K1Zudzu7rB+Cbw
pp+6V4gzDLxE4nd+5lKc1grt3A4PA2QDzwIGVgQgxvs=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 42000)
`protect data_block
t87v4nOwrW5fPoNlZq3pDXj2ALHB1fVMBEUZX7llApOY7DmCAeBEztAjyvDjHbjc
xhhmJw21+uGkfEbfSIzLYfKHhz0lshtglKONHMcUsanMZdEDvva0hNf5j+1GshIQ
YfVavjgH0sj52fWAncjqpbVvoxvS1FEsf1gUAs0u7jklMh1a+R64OSw0+jkqhApG
IKOHm8oO+rZP2gXgDWYms1+RoICBHRT9+f8d36oWmG6T5Gj4ji9CXYSrR7oWH+g7
E+iWhicgiQ6JCCWFAlo3NGA9I9rbLUpeAzEVKbDu4hFc67WkJXC/Wic4fyhwvlm1
SK2VywxUJvpSrkxPmM3/xouzIaVKDLma3ySNjX2sXVOFd+iPO/cqDSZEHGuJTCVV
0cbv5U83SSYRqeWI4ZNqFkevuUCtNLH54RBOrp4Iq19ZK9ikYXdWo6OrMouSzMu2
gtcQ9bq6uAaICi0AnepOWUDvz2O6MgyGdMiCkSr+h+U2JxAnDCS9KvGtyerXtHYQ
YRlzhpVOHg7IlUi9qMfhh3fl/220ANmiSxn6yNC4CqWuYnKZGoBnl5ZTlUlBJ1lh
4XeKJ/REXy/PdoR3uz7SlcB+5Mw3q30I8Gj/qpEqwVVdZ26pioAoKAk2YNs6TWsX
HZbTvUp7Y4A3jakuQEMCn+MezDngWv01m4AphiQoiwAOUyONNlHXkMlF73mZry1+
y1NNmdidkWRcJvXW9GuamKbSZaHDJBqX2axgMpHNYw4KIYvuKsynuaqDoMT9rw9U
jq5nrjv/ts40PO5MNyjl7Py4YyNe27vRqK21h0y9XSL0nmvcMvGA/NDDe3J2pyWv
AtmBp4/2/FIg1Spv6VvrpDSToncWAkIcHn5L++yTLqRhtXITFW4e1jkrxspsevoq
aCa9cmqZi8PQFCw4qKVeA2b5Zqeqg+KGxHbYwhOrJypA5L/nqOgML5Ul2NkODhqz
7Io9E1TS1yqGOTizgc/iH4yaFDY5Py/ldflmQmSWJSvkUMO12JTmcq6EHo2mT8ig
RWm7tBmUaf1jMWoq2wkp53nhIiRUFxsuC8fsa44bvgCPVQNRbSRtaIt5xEjAdsOo
KRSJqJyWlcm86MbWuvI51kG+3G2PL2Up9jW51q4OU6XswF9ZpgZ7E1bsfasCtz3g
6PME7ohte6a1+A00SXC8u3A0oKQd/lNmnOdzdt4lV4ox6Il3JfU3NPOKqKMJ2qtT
xKs711zNqCafZqx6TyV50SRxP0xmzU0/m/eFFb8kC2F0oX7aWhJxeO2+A9N7LuKp
kHmVDWgzXRdz6X/+wyyQUtbpjS82IIx7HraiwTvZLzGul7qJx2OBTnn9rGQ+Yzha
ZVuxTcxRuDbJRISitLgtqopGJ7iy5WshnafjgyDbYBNWWbRAreCdkDMW7Ntr0dXD
KLtr0AsqgsnN4zbhI9BKpJIGiE6GpIZzb6L4u/LXtgUIW71ktWd8rqLu+qJBRRgA
bsls7jZn6uwDRIsPnfEYkzNz2X79I1W3T05iffwdgJO/wS81vTKe4gNZsSnrS12+
QLy2rZfCP3mAzmPB4jZHzY/8kq4fr8xuTWt00xI2AERIHTkfvNO3cMjEkuYygVYL
rv/uuBuqId3uzS/R9cwkz27HSoOIwLWZLZO9ir6a5tedQnbejD5kshbKmiLGLtd4
RUlrgyuMixVUhcigF1MlanQStKLVrdEijRaOZ+OKHJhHdaiM6zQKcI3IchNmNueo
cHoi/N5+AfLZrzbtQ6T6wdpoG5l810FG+/D49k/qYIooOOgHGCDu7EJcOEMdta3o
SG6oi8becvAdQWE8or01X2M6/4WeEY47V5qH//OR56T3yZTTNDKIVxa6hvqkLFAe
p0l3+YOJTs6kvMm42GUqktn6rwXHCaXEjqkVTbiAp3bAw0N0w1UrGB4B3Zn0jn3G
+qp0CKXMMCkAZBFGa+HXWDTdK28CW4+1z4fIurPaoZVoNOkOSPXrx6GSRnTch5M7
JFk3+1byWxPSZ/aEdB7C/toFK7d6EY3pqXxgsk2G7whvyFWKdB7jtBqix/jOtCLK
72IfMFX+aFHqBpbGfGLfqLtWG3DOPTSwTM5917BbvcvKM1/s9J34DOouFLvlzfyb
Dde5nV7+/Ol7JG9TCHenXAcbkfHllQhtzM0/f6O/uC/lr9GLIY1bLZzd6XaXwLn/
5FltngXQZwGTmo5bCmvb55Q6ed/fEXnchTUClSrWwi8OpKqon6kav4ES2ijXpu2n
MVnCKOLg8CAJaEWrENl8YOQxZA6Ac7IoOEbfpC3WA5FU3Xg46r/+3kkUx9E5H2gD
+pywaKi5i+x83QWvHBtZ3N9LSwo3KLsRZELeCRYHFVU+v7w1rM9pw9P9FDrXEq4P
TqGdTwZJDa8tTVDGrlJ8RAGgpeGXtP75CeH1NuF46smFjeGt8aUhtp0VLFX9o6Db
Cn11Tk3RiZKo1qXjdjTZlF2kradHGSgsv8XFY6irQVaDVy9LsiXk2Za3gPHB0itI
JJQBpWsXQw2C7tzQlKsTXNLbmk6pYYgqJs8hNbu9+AGsD8/Qa6ChOnJ6THwwmLUG
eEr//OthJDvYlw7tCRuzS4mJmrI1zJHwdwDvmfUfG6dpQWbuXfQ33B11En7guTuO
OQuGuJNVmiU3w06SinH/mkszYW9dTkmgrXiNIQJjdLk+3Mb+zEfDIGfIepHAyj+O
B/87dI6pjuHZymAGybt+CoEdkQaINsI46HnIC/Tdp3rg35WDnVR/qOedBKNQDIGX
rpuolFs9Q7s8PO3TgvHAcwgXQ5IP9fJkfpLYGQyA4MhM2HjmOP9deyE43buzq2r6
bdEZZxzCs31O9AIWMCG87NmH/6eEVtuvDpzcw4MRS/ARUGwGVtOU3VfCsTz6876Y
2W5w9uxojU7p1n8HuQR6WtwjeHk4J30t3rOzQc8tsXgoE0ULyB4EVYX3ikTKb+6T
cqnIHKA9FB+GJKFNPznKZR7gnXWazBaKKnRlgfhkUjgosBW1xyW9qL790S/j1Ij1
kQqSeugzh1a8vBX6+wF5OGDzb2gxM8BTu/2UHVEu50lzZZaSOoiG7USDol8BHwId
gG7cr9zML8fEJJUrQ+dvTDavPxkgU5rkhZpWcg0sw+ddHE1RuohZHahe3VUbjVi7
VbJBVcgLNaW+og+S6Y/27Dr6lOgN5+WNJviurG6nwY/h6suuBX7Fw6Jht78VptU0
Xi8ZhVQapsL9zE4Z1T6y7RnJm/7a5rvWTLDe8256tGMYiMgl1o+N6ZDgBvSjk99w
ssecD7K6di4JYtUHmztOq5EafMcEhO9EjVJB5Uxjn03l1MUM9053bGoVmanVxF+A
4rU+Mi8XzXbLmpholsk1ZyTYVwqI67Tud3HiDTynqlNqKgRnHeubtIxMUprqYZqL
kEJx2nEwikZQPIps5MIdcn3R8jgiIW1toVUO9kwqY9kjZOHYkGmtPE2/9vZxWBoE
kp/HlJwJgvESMdbp+jzr+MuoiW+k6uiiAzdjLJ0crED+YUqGSGyiip9WQ8xFIfmf
BojMFwfAh5zngLnqhG/IAK7ACIzqw4j5M4/t2MbwsMOo0c1ILRdpCdjaWG0Du+dj
elwBDs0cRvMheFq9rQT1Du5+Wv7ZMssHrZrSMUVRMs5joRhsiSMYfN57SliPCS0U
H/34jzF4pUBTMM5uCAn5WhHdwreEoiDLa8YGmnu8ci5m1G4i8ehPSA7BoJXYh075
vNy/YUlpTLglebW78rq6cpZ+xoJuzQDKH3hqgCZHclgyJAV7YGZJ+jIz8joy8RHX
eRqVLG09LtmSUO5MpOpOyekqdVUm69qqHIr0xXiyLNS6iBTZ4Y3W9IfuwAQMYFLn
pKK4ASleDOsXengY17050bHAksw0YxWbjS0Huu/OgJRg9ltfaz2yKJLfFtlsMCFN
PuLmZvvZn3KUUKdpnt/bu7hFUIi+YyEAArrn3W8R64+EWLNHqFgUpwuavnQQOOEG
fYdh0/tQIOrHgVQXKmPBOi+YATkNheKuHMZOc4tKFadvnP2aKWWkcm8EUcNXFcWb
54RwSW8Mu0g/+kPO6sjFejDeTWkSHbjf3PT3ySOFPJfyWRJWCF0MVPbtoQw+Tdw8
pgbJKdziOT6LRJiYVpXO15aif1azuIZD9aPy9+RFZxpBUgMw3J/17XnqVSU0Jzma
+6IVXfTe+BYbxfutSn2SJ33aa1rk5GEHYlvWRR415uFrCqhhHP5dodn5g0oKIRP2
jj2bSkBpILTp8mslTkXuvofIv/AGzSfcpPRT+Jf4ekhZbE4yiK4XQprjI+NYYhU4
q2arrQ9T3DfHdRJoIcZrKhSK5PRHNvpjvUKCSTjVdRjbL5Z7tPEoHgXueLwMCjkf
Uq3jkh3kHPm/Ao5nDc5G/MP7x5phWtgy4eodpE93NYrOAJAW2iH3fWSzaK1srAD/
DtsJBTkpE4Ga5ii5OBRJTweKhhmFVj0f9/5jYOZ2cNTxeQm2b6Nwyf+pnslqDV0k
fmazvbSxBdiUtv8u88yzpfXEPpc2TjTlMF6vp+Rs7edB5TKVkxLB+WwKNV+CDzSj
mSrQhyiRtlCf7nmph9dBNzzhMZE+xHZcd4VR02icY3BEvk2KgH4XqOtQykEWIHv2
URJTiP8S1n6HFkG6R4Ol19HqvOJ9+AgcN5Cm14vhxJnTG61wB3Kk5s3ybVwJeCie
l/7FTNIdN32gm3jYlzzWXofR+21JSJK1NdEyr2wjZtZiKVCYgQh1OstwEf+njU8o
hzdzXmmjseH9Irj3/tNiEoDyZFf1d95IPfpdO1hX5i9MkWk+Gke5/BOR1G+1VYiG
n5pfAfnzOmNXIgbgEYIJAyjteILB3Yk4s6onnNaiCwDg1HimippDz5gIJ3nBMRFT
VR6OKfJ6T+tB/2lZqYkzZtQ/C08h2NPgqEOWE7PRce4k7Cgw5DcLb/meBDnpHDL3
2kkYq1vGZS/a65CK76TQn9XxIv45G1ssY6WqZNbLokcih8fqMtJNZwMqICHX5eiF
9RBe/XAKXhhjpqXgzEAtoCrIfn52BmZU+V5SGM3kCy+RLGl9x6MngUN3GOzZ+ovp
WZ2iKaytn8diG3u7vZIJVDQEMaOdBUZN2W3i/0j5JycCilPdXmY0xqqRQy7SJVO2
TZD6yB9QpLp2ENZvYYBPJa5RstUTsnDWF/anmYPfb4pi+ojPt9BRD79Q0SoyGdee
VNnTjISUK0ZZ3z+9asE1ZK7h89gQeIO09g26m1WPcgenwxAYqboAU6o0dIVYUbcu
l88iZa3b7PL+0BJoUiBzTNPWUtGCI6MnqPBS37zv+3ECWatjZZDfIfJoABSs7xHD
peXemna1VxgIrnDlOMwS5HajrlNduedqo1SbPlQZXgh1HCrT7+E37oQl+vmv1Kos
8UXWmtXXWpFGet2SZakLHfJ84tCYTuNOJiJ5+LMeva872ZIhg8Vzrf/IJZbnSvkG
N5tBHPYeJTY/WP4UeVlQl0bxSXQUaj/mg0sVbTX5EsqCS6MEzp1VWNcdZDIs50hg
0iptYwcTPk3SQuY63kP0Q8JKs7KSqIiOB1M7ExHCGFDMXSjNHEaCc0CeFCovIdGF
pUyYMz6K92MnOfaFXoqGcFlitJz+nhcpINisR7lC2BLwvcisgui0Oz4iGzSCm4I0
Ug1UJ4yXVIZXcB9loZZy12ajoO8qFMYdYFHE7zNj3nLgc5Zy1ILa6Ga9ezi5Jk5A
ETfsq8QQ/5kVXv29AAt8menbWcpXomOm7Z9RkM+vffBH7SLsdp8sYYe/qfl49oth
BgzdtROC3IZ7Iq4CQTcFsQ+gHXLYcTqhuouOII6FiJCRB9gtYeyxKWuF1vKD8PgY
CfFBqOjUF0OIj5KJlQEf7mglvt/un8baZ4393kz+oFeuUnmUfcFzUgh0ccTn6B68
/igQOpEcp0Vv5Xr4sYYyYgv1xypgRJWVf/830tkk6Q8UMzYxIMsZDhO7jJgG9bn/
f2xWG2EvLLHRhr+cFZBrUjV6ifNtOE3erHVymUhMoqwlyGgy82HWWLJgD5Gorg2r
AH7VecAj3fmh+zuURYhlfoSeT/ca7IpclJ1tbNxTCofVelYms2Nh1ze2Wz0UrUeS
a9v2VVbNv+iUQTfUZrSR0oMHpM3palo1DoisQC/2B4TDv4YHh9zBdceMC/munKpS
M0p0hUtAmS9YzKRjiMSscTNj04ZYxyyTYHoeyi9CPXD1xuAQ10CU/92LGwEsdM43
VLgcO/T/dDNa94zg/VcovF8bJTnsukKB5xe2RFrMVVWr1lgeiijFbcDttOqG0qCr
lECVxM97UCeZYx8gih/jG+QGiXviD9kw4FyR+1fO/hLpAwx2ijEZYkDgxu/bTYNA
xbWSwfyLIJxy4Tk+p1K68dPkGyqLendhEYBP5m+XDw5aSopliIzy9oBlaa6RVIud
RWe61hbCIrQnBl1NQbGbeJo+Z688WEMkIUUxrIFG/GF7sn99VRl0F3akSnCY36Q6
KjGpnTamACjcgMfcFebX7ZZoRzf3SVCwygivaK4TC9wFiR3uV1jV9B+C2fQLKbx9
AC39P7m9Dt6M/+SXz+MrVvcy76eOUh7X3kmd71hv5KLrD9P6/trjbQmx56vst2Ih
zsF3DcMWvkdTwHDo4bPgSNM2RZ5bT6P9ftWkbaWi0s40wuxl5wftQxJf9u0h+xTw
/WcCd72STRFIKrkr2KTG6wI5byLRv5lX81h/DSUBuLwhfo+wqXcd9jI8ZFQvzCbD
YDJXYH91r3UvMuuTlK0SPMX0kfvXYs00ZwBnOuvVZUexPlEs6jIs+zBvuBPTvN8k
UCwBYQoFPQaEfBVmWN+SHgrXBSO0iLRkxFhEVeAoJc/a5D5yVJM4MbYpOaAFN9g1
WWsbRq/PnXhNaBqw6hFuplTPBeJXpIIsC7ZSJGKW12DHfm9lyffdzCUcfX+xWk9h
FLpgOMqfDvYrQuJqb1iuLxDqEwVCJxC7NcWR2aDA9IWk6ZjCb3EZNdyb3VSpQBLZ
lZgs9B4u2pBTrwBO1CeXOLA4JqLOzI4JwZXu2CH4eNFfs0cSvTf3n186C4ukqoyr
C2nYSoridlhsm4r3+YF0myQC6nQ08lG/BR2jGskM4Za/H2SJ/HxBv9dnPZFuD2nF
xMhZ6IPrQ1zzKay+JkVO9DP9Dc454OjOICXcWNVXfrKwWZYBHlNCYzVLycJPwZ4v
gJGua2n+R9wnylGPN2T+ccgah08HyEZhiXVQLRadjjyah4yjl6JnhZEJtLcMFUx/
TRlBTxmvUY8ASM7l7wZ/3EDEiFHgYoDtHwvt/elsjPZZilXHxDTuliFJ/OmNMR4g
oJt7cYtYJr5OD7eZYdvqpiqoib0FBZnZf3bRqOu+pG35jwoZdTrjRtTo00TKAmKi
LR0V4T4afdJFsCfI8iHDnvrb4f/exlTnN6COVR99jKX/YAWBPdMOfiiL/VMd+TJ+
sx6os3jBQhF1Mrstyj0yzyYjxpDedTFUz7yQNnN3pvoHSPvsTvAERU70FG+RuMR3
sRb5qaONiAT+U5V6otLQIgGDgu/hAbeup76OnYOY8HuDzNpOq6ealAyLDt+fPRfv
2x0C7JmFHn12rPWSVICdAyJFy/LeQVR+3jA0PYgHS+VgeYXCRTZm6/C6gvs1JFqD
0C/JC+9zluBs18WGNuNkb3lxpc1deYSSkLUAN5cBQUTmKfGy/T/hA7MfOgM4ZsvP
xDtt9L2o6nbk/vOBu+AidD0bFzmwgedSXuLJR8gZsfXropkqTbeUK2KdOIAgKaR7
M7ElGLENPIggn/l57TskwNM+Sbxlf4TZEIzivs1lyfKVoWYpaBIZA4mTw20QhbrM
mvx6/KI12ChIyDsPq2lET/h94XDDLNoxBkc8PBsJJhfCQHyz5V1Hga+FubD3aOQG
eSv06FyyrGo3MmBZYcDR8hldXKptEcaxYyJU0uy7uFHo+N29Ph87CE3uMaahHFfz
7QVilzR53EPZlyEBvrpJBskAZ+IzrbxBhbNNkM7sMYTmmVAjNh/Pg7dUCGrtt+i2
KK1QpOgMqXSJEi2HA2s+g+1WPC5havXsKrt2ZOeuVT/fkJDUr+aBQFkEadIsrpzz
8lU9hKKy291pX5a0o0g6OhQ2GpAbPMZPklfyqTSrKaGaLJf5P7a8VXQ5rSGWY32I
64v5WbER0P/veZHIq9hoPtLClZokQK0MbKy60q2rLQtTB86gnTqD1wm6zLjrlemr
oNjTU4pmUQ/8vOgzbWhYmpapXHCNiGZT/DNZu660W0/ISd3Q8q3O4isqsyyYVZ0t
whvvlfgq5XgwLKNjpyehqniwSmK+a/X57m5Zgm3uncwCEaHDE3lFxCGLr37b+HW3
2ZycRrKJ+lBJCJdc9DYNqarXeBvTlOsZJNRiIA5vN5UKw3n6ji7Irzdnt+gjj5zr
/1zjjdibr5gS1g3n+0RjCtqMOBWlnHB38JKjy0qfev9EsFFQJhCIHitVXJmhXFBC
QV8kzgNjC+oLv4vHyUS2A4OMr1+2Kf/0zhjOsoduhYNR+dmBwEkYTG9suh7e0TSF
h36qq9LCu41J52rpG5TLrTPwHoU+PSslrpAnD6lZ5yaiMN4cK3Pz/R0/SGfHtChi
Hmjlpdb9arHDuf+GBIVIyaLkFSzsxBoGKKtOjURgFTpWgfRM1NspSqPlOwlKG6IH
XhT/ULrh4v9FMXBPNMPBt8Qs156sl0KK258Q8qfJJdv9ZnsNKzx1JOj1tQGAwrIC
OD35tbMs5p2kkuAk6dvtFdRZ0OHgwj9o3ZDehhjFLL/jvSUJkFnlTxpqY3hbyaAX
IMQHLFTomoDcYHl+/wVmgSzW79OneQCkVp3bA81kkv9dgL0R4cs9nSmTOLuVM+/R
L+vWa9xnStz2fOdN3LYVv18Vzx7OKMjKEGTAUZSIkU05twbeIJQ6Ndu1EkqqR6Ot
LfN76+bTTACjxnGGlRpUI3So25t+yrSSUCLSp5w9uJyzntCIB5qw9kdcwIsbnOaG
uLmEdCieYXXqQRABAFDqhT08XDbQ1bJoruSpmV8+Y4xaKrXcaNRuChTAIKhGlg32
mwNMtmWNlKNYRvcT5ActMhFO/DnrlLmhprjVWleDRwC7+beR6WyRu8bgqqM9iloK
8Cffe5r422m+dx6fHq5bVbzLpptQnpCI2j1T75z7FOQwD7Rtz18MahQfeZoRZq96
QGteoXKSqYBBvqXKJ57c/2iiRXukbmZhAzOxGCyFG6Q/+cYXJNaO4atWe60zCKoQ
xVKZHffn7+0W02m3CNJf5FrvDWUQVQ+3pCQl2RRuUFR091eAuF1yKhQeBAs+Gvt2
LYuznRVhVEdgzR+08GOMC1KNRR86bDajbwTcpL6m7VJKLqjtCHVwhrxdCBghtmiL
uEPb6mq5QqxRS6JbsxYVRBnxeU7G2B4k8scKZocl21NAJ8Q22sCYbRUm92+tg7Px
W5wfBaRc8qRtPznGmVVAzvB7fhyKQXzXrZ7z0W7j9vAaUWup6Zxe1whJrEfIYsYu
/bjxto3Eiqv/2qnz7QCskSoDy2/VewUOplFo3oj5TWjokyREKREJYiQL2ax/jPbM
WeaGQvWyUKoGp1rW6GHqgQvBYPxWg/TuBfZWRG3//ebOnA8YxZKizXVQzmE0M12I
mdLffUXL/bWEpLR0iWganJcP/LTEAa1vSS9jJt38md1ZbxXh7tNWUb6Rlt7HGBc9
gqiSalh3ulFF2Asq/h+Y0ipzqq9gLLVFbdM3a0Uq3ZkxLcp2j5g6p2dubiOQd2su
m/Z2lNYLXCvsx1FXAOFEM3t2KYcnmUrCvCt2h+su4VXdZ9gcayFN5gWXClP6q2EE
lrb1KcafqZtjWIqBJJdNaNjBfTsA44g1BmtyJChtKEKXJ+hZ0v/lK5VyJZX3JVzu
A5wkTWoLOSPDFM0lwXUeIBbeLLG62sjcFb/7X4h63AtQH9ujIZAEg8f0WdLC9i6t
AEfRc7gOkfpyrP1oxTA5nZfOdBsNH8sRD4voh0QMpiD4fNtBXwjPv8wZ6RAltsOb
p+j8UFaLaImIvfmqwkWtyRL3S4l89Y/yN1GSaJ2KLqyJfRs0HzXMZR1RWcMWsbIc
TbByHqJFRyEULoxVDOrkJUZybhe5wqqS1WMaFX9a3tyD40V1TaUEzXTh4wZ7RHlO
/g5f5RRncYoPF4ouSy+0ML/mlmRZwXRexV7fYKRt2dC0QBEVGGDqFXmkYjNb8XlT
R6l1enesdo6Vps8EvFiaMrIL4v0VnaFv9QL+gODGrfll3VoUwDUWMUeurobAskai
a31ldQDpCds9VQjJBMMdwBhZNC1TsaOv01Pwjpcw7gPQAGEJmxa0+UGfN4oYlME/
UFo3Oi1oVskRcPdnfeJOw1VkXgxNtzbdBbxV+/0syfi8a49qQLKaAWVisjnWl4xE
iK4F8BS76fg58i5mVqJ/6gI5Blxu2FGLBTP3XcKtqtWUa7V5ciQrr9aJcZAaRt/9
p9SboI0rtth2lad2wRc5+Pm/uuSeZcUJBwMZaPewZqnIbyIygSc0q7V8+5EiW1ND
ttTjJPbdIzHSEACrf6hZE6ax7riqz4C0VWVM78erg/jG1h7Q3ZOp3MMnsyFeCgbY
fKvH6vaVeikNrWVNDJ/ngINw10ILwqto5pPSqTPbxUhP5u699FwMUK4FA1Ha/2n7
EkEqGSNcAz3A5nXnpyA4jk0sGE2HFMNHOKoEPKxFkVVhSS3cY0btDZa/MC4tsAvh
v5x9LRakmO4Epre9Urxbtkw+fHn/bPe3pxBCYg83q4wylgM67cqI5+5lEWre83qr
yWnIy+GzH5ieHseuM2oLKaAzz9o39CKhDaTr2XCFYKsTLo6WxJyqnEoFQyDg9ZjJ
oWb7WML6Ef41JRFhgYw6ITpvZjYmWV3HsRWjP78ewVcHpH9ltEeAm3nTmHPdOGY+
iNRSkg54bMDgswZEc5vFHtxH8UJUsj5jTsLxPpUGlxS2qXqwG2HDILBlFjiVp5Kt
Yhn3Cw4E3hFMZpiLLBsWVlhxCYHinR0oXcbTjMdM6HzGxk/PVY6ypt1bwZ7Jm/21
rjqGg0vv3nSKeQUSPwWhoZQ4syZTM4wM7pIf6HtPL2ObZamKVTakYPlYqp6rtTFF
SdpbVhrMCfZ4twEHuSLsV+tJ2q5HGwRJ4/4AElOqRcsS/rtl/O2gW4Ri+o8mxAAG
fi1ParhDoDR/DK+3EqBOkkMl63w0O8j3E5OsH6c+Kt6s985I08pKB913sAOdPo18
dCWIspelTTY285xw/vQhhtC4ySbVrhA6TiyLAhrn7DbBNcQ3ZRHcnRjqxaww4Hk5
7FxA9dVSRNZcz3TPlZwnW9g0hrQ97iCHDd0lkn279XeW1prhk4SKPy56vsASv6sY
OLTvpGGQ3nEXl76PRytwOT6BFxJXDu9j2QVWUOlWWJAIkwG63hG3XkFPUlpi3MWy
96gVifmnLVKNc19vj8MP8SimPfUyCclFhuEgnsfGQ59QoOpi+nVbJ6w1bT5r77Rs
jm4BbXARNYqK29AIJUVp9+p8n1I7e4+udfqZJ3ASdSP9DJXsG6fBSCJzEA9QpgiS
mbyvnQW/vqfwGbT3dq6f/EKSf/EAbdpmycX54VQpzp2KOgQU+dlEpsD36RyJcoXC
DuGesGl6K5ga6JkjcLZPyNIxjqb2wYQOoax9zpVZs/GmPUDOFEUrR3t4WySIEGu+
qz0daWV3iB/Ng3nvoMFShHrrlwjjxJsslCnWi5cZJEka14ITEu+xSW4xilx1J7Td
2tQ+tK0Hy7Chn4Gc+mdDxdw6lq4ERRxhJkkUafFVjZIG2OE9sGZb6KfdEdiP80ib
Hrx2/CI43pI11Ukb0bNSKbSGMpgIX98ttZcZTfefL/rF0gPs7BU90WcvFcdvhyev
7ynmOQ8WO/mxN06s/2qc8hIuiuBxfThU4nE2GlDu4KUBOPbQAR7+A+2Qorz1lc33
YmHWcej8vF6bW0cqVlbovKX8ETHeR48k2GEot/XsY2Gi4hmaxWpTQCKeukoyIvgB
3iysXpYCZrrnAcRp8W86W+DeQMp/UVCTD0KeedfLEFb6xL0d1kH4YRlv5QiQo0d+
wKH7CcZs/h43xBD87GMVzC175xddiuyJkICd4PQNFCwJ4DNFFN4QjlBM6pgfYH+V
YuyFJHXZk+YIPTs0LMXypWJ2EyQ/VhCo5QyozEzpm7o31pRY8AT7lZ08C0cnY/hM
HwbpnRnGwVzhTVye6ZJ9zr8tiAbGs/qJFVogfIh0+3SsQUev3MEEtRydCTiC6Bg5
50QeOEg0+SL36eN3+QzRgw0RuLXWn427pinQe5hCL26E2adl6zE2WpiDW6C/Uc4t
CuYhixfK8l5vn0s3vQfdUb5FnFjtpsi2wBUd4VNO4fuD43xePFs0cu2FEgqspNGV
NprPAXdPZkUZgf8w/goejOohWepjD0nYia0IlzYcAgtK05vhgif5n1zubJ2jLbql
QgeUUg71c4X+UII85XwJEJ75KN+SETz3NzxSIhx+tMXVIoysFCdCbYPCfLZr/mXp
m93C96PdDQjGvXbBKZ6keGP3IvpQpiVOnjm7nD36TkdeNcLHJQE96S7fHZRbMxpS
cBurxdfPf7YYHj886l21k/DVyMjYIrAgDu6BPXSh63m2hN3MqRGEQUpWwDbKjvFP
nDfRmBa0CbU4Er2yVOzGIdnYY37zsMAGs+9kNsZuI9axeiTptVEy5G77r0JxM3Nu
Oggmm6cI1U/NZk3WqDqKu5w+qN28bVobq8I3sMQlGdzV+kT5IfFGMGtDvX6VN/Xq
/Db4S9qXRWK/0SdAva105xFAwMENG9C8SMAB99Iu6tR9r6wm7kGXE/dGmgE0jmPt
CA5z7KSKgsZnLSzKXCtDEvkICDnS+pa+eo4pTtNwRnASemKaSK8cJn9LgsvOny8W
ECJ6KCXAzeJi/C8/UX/D+sVFII+yTJ3Q4BBw83EYDadcJ8aAMt55J28eQy/narVs
gNG6aei5FszK2t5kIwOLb2sVIDzfZq/xaTi4A/2S5+SHL0EIByNnh2JOqHtqKaZJ
nclbow0gAY865qbW0lxmxqbPMQ0Bu6snE35ezXCYgIMBh/aQG74i8lQHM3x51Duh
1sL35AI1jtTQWB4P1zFV1vpSiQRpSXedGHyGRdlE9w7ALp3yxAKCu5JthEgDNHim
57n1s7R2IJqqHeXpuBI10ClZz4fIaqjRx4kjK9VKtQ7kOGUdt1UCDsG/9tmhAs2+
4V6pkQffavs9A4xPId97NrsaD9KGhUVbGa1jvi+4hNx/WLYHshQH40UdsayanHEX
gcH9Ei6zRy2+/NmolB/04Ai9QGJr4fCftlLUkgl2hVGt43B4N1ihr0XBQrm5IqZl
fwEoMRsIknLGoJ80ZzU679oUEM5mv+NM3Krbrqt8hlvNmt40HIt27hduNf81Ry+m
poGFPcVCoa6NNdl9wyjlnunvCsMV6tJhuoVzO/HHKWBhL6Sq/LuM9anpfPWdUYGM
bXf/+eDqx1ss39WHgxk72MK0eB8swcdZ5LleZdWCAYPTU5GzJdhiwnVbnHdz0Qew
thKxSXK4p7CupOrJPCpcdzEnRivBt1F0wGIwt01sxOqbRGp+Hq4amVvPEZAkZJeg
MfFnVyhYyEYYWiBZ9Hblwzw7uzZz5mSU7jhVD2FT37ICEpcGfsjm0/dQOAz7yci2
3V7ye4E0/SaGdsbQgD00l6L7e8KdmojMLXIS5UJze2p5Ou0RZkAJ39/K6taFLahL
K2fO5dtQGimFk8QQQLF91IvPDOe4GOL/KTHFL+KrfLw0ztpG0rYjE2O9machE/fe
wJiSVGSNyk3PRzBOrWWSpD4D8U6zWMoktCUIWy1i6MNIEr2M34j8bMEOOPWYtria
htjGHk52dAcGCQkQKRKvKK8/aOJpLW/bgtz9aLNdgHiOnHNJyvaH+RH7GW7xEa1E
VpYW6VquZolJ4+MlsjzXUknilroCyAioxrds9pORNV7m0Y87gK6I8uYfhEgkZ+oy
6XBygpr2AkAQ2gm9xYrjMbQNW3uOJYlnj7uyGAiRrl3Ne/+9bVLRjhyNHVaHz2e9
NKy7i8mwDYmtaqYjkMeORSI3s1KzLCvjggifuh1EecwG0LtkMZsukuShLbQWssHR
r93Xwv+Mn416djcBxWHDdATFSm9j+F1EzLv9iR29uq7HAvBnYtw8Sc9R5XA0U7j+
oci4zexL9lk04wD5EiJK6+kHnbCVwWp8WfoMB/eDcdbid50MC8rOBOjk9HiBUmt2
XGIgtyciYwbsMDKllq3CEsMkaGMMheZeEbym01DfnBHaEuqu3XaPPx60/hyaFVaI
iPuwBidaqDboVnDqfPpmrQkCuA0O8S711Djop3exIcns1pzKhqyVL4FuNw3LtIsu
t5ts2WJf5RSxtoQ0/s7ekZjjHWqE34vuV0Z9zE0LOzWLPyK6ZMruDoiwzDluJuh3
k5xwm2A5+BrnhdWZBeemwWRYhFRcPqsfNakc0WfIrGZ2NK7s4aOcJeVbzBdzbjV6
x7Ff/b30jU57gkgRWPuGzeGoD+ZMwyywPTJJqCxUNE674mqbuK1+fJ3qF1tQNgif
oMKOvyIeYHWmdPnzFIj61ZApi0r2IDPmmwlrM+eeepL1D3nqcYsmau4Pw+T74hU4
0vA6IE70Nwzy2I4Lvr/1/xyYl3wTGUckyygPOKFjVONG75VbO8bJ9KFrPFg+8mmF
sKZz0LNiSIO6w6IsebpHHbfcmM4CADFOjVPoFhhnFwZNfrh8ft7ySmkxGt3vAC+i
ryM0UlxpvA+gtG2AVEvG2GxahzhXeG35VhcUHb+nY15UbGU+2EsyST3u5y0mlADS
v8cPq+Z/bUt0ruKrBVqXhHRt2dYjhHO+mS1JsfbKNjUnZYLK7bC8VoImVW6X+bhG
cA2w+GIjtwCOAKuyitQt78uyD3SpUc6c0uqdJVhKdoIwOo9Mp98sof+0HxGMEOux
Rnvydp5aXtdIDs/btZ1KT4mBSFhR8c8a80syfXLxrjhfce/8b7w4HtHFe4rfu5C+
p8xAt0JhwoNY/m0RDcNLdAMmDrZy/taKkmW20NAhUQja5H15YPoxV1noye6RnfW8
cqP3ihPGd9aZHCxZ9g+tgv3UbrASciDisym6EvjqCidj+A2ixPa6usnvmwLC5uBi
5SqScB32edevSKsYfWqbzqqInUAbrD+JsDXRooN/A5iS0V6z1T3JPW3FJ7MZoTs8
FhLEKM1LRtfTknDUiA7Tqs+1vtcPjhJW5/teDTLQNeQzwK1cbec0ZmbQu4pZbeck
hUoWELQuRFu50Pw4FYeAVLLO9+2rR/ckozYPTzIX6PXxu0rx2JfFz4d3XmzLkQ/F
ycOZYLnzaCczsbI0+VEBiQDoKzW/uXynG+i4ECZ+Q6LEYdgagQSCZ5w7ecxw7h0V
X+ddXfuzy9W3TnXHl+vCvgDoLwvZn4JSrZLcRIO/7Wlz82nIMQtOsFjlJOvj0CLp
Ct3J+uOdsH1IN1Sn1lK4DZ3Y7agC6u8uqrPWGbh0bsWcq0l+jYCpw7fgHQcOwWHk
6ekExwTKcvjuFIFfBsAodt2QiqXZMZ7pLib/rMzR32CoYaLqW60Ug+unqLzdgn/P
4NKfPFVg0c5qOdWbdaX9QQUq749tcNGXqtAsAr3P/tWdHXWou4u0Ejh19L9P5YSx
mlLCXANhuleG9w0vRGQ5GWtdsop4GEjwu6QzUoUsG3M+FMX6yCPiApo9PwJmkLzd
JlA853sf3/k0XgGswz++2jyGf+/81+Uj9kiT00fg4c+IFClDWaf/6ei5ch/eE8rA
aEZ+kJwV9MrH+j0K0oYsrGDZebwLZ2x8LnbNHoytxUpw4qMNh+pnqRGYwJLH1e6A
veejrWVsYQkkVIYwrtgvpuwSnEBgZLLEEX9THfMPlOXyjznCrYW+lNUlojVuxvXo
uhPKRopKxWgp8zad3R2/Lf4d9FAsskPsK06bFMrOt9/vo/FyyxHG/EeRnNeDiJyJ
vrme4dM5VGyt+EfPFIVeIwj62D9YkmXOr/xn4DCYGHnFjLj8a3uhCga6Se1tMOZU
hqgIqAlTzsAvddRIFptsqelItnKIId4osTNDiuAPycGY1uTYKui25f3Z8TPFugbG
zYnY151ZzzWXMabqHuy7okQgUKnqZRwQued44LFohJwfwUHO7Wumc8w3K8ESG7aP
UoMjKEiYiIy6eIj1q8cAgr9tZ3XkQUWQbAST+r7AmJLai6v+cO8Y7V0goLTIxnZf
V79u82ipA/NgAfCsvNBN+Dk7BSr/AifC1NrI2fbQEbJ1JUhAoNQC9eM+NiT7CPJv
oGBOgTpw+OziwTYvMoexP9n/CBmkAEwWuUakxdyjHh2vZdRbzOmrsOPlLsy2Arry
F5D4oPT9JcpG6SOFFafIrn0bkDu3/cjMC6KnAdlDaguVSo5gUwaEYl/91SfEU4Ch
bVR2XVQKzwCeENrNeoN/M23MiNoo9FWWPN0s+XBBpV+Yvw+tl7sf58dFuYZ2AxgS
AYmezu+TlegYmlTY2natqZssTevsmQf2dod3nZOgBa+be2nxYw+Zh/mWMTbKWSAo
U0THELA+4PJpeViKRVfTn+8G0KabNpshztjXKn7CxyiofZ+nSyQGm8D39quFmh+0
uAPgNah8zu/wnepe9j73UrH1FQBdhGJhEjqhZYwZsIUytfllHy8Be/iVCCSQgAUy
ZCyE3OiL1wVRjHZYkATmLqDjcELQsT4SRLfsS7BNbX9PJh25jr0BZ2mHVngEqjnz
cz6WQnzVjQGT1H2x85UdalfGoszPt9tu2KfUU0n2dMyXLESS7c1MtoC8Mym+oUYj
8S2veIi8Rpp2MnuRZceUpRJ137N/XzhBo/Se4wU9n0gFS52SKTqFHIjvK46OnJ2O
WdQKv7QSd/6C3DXXJreLO4y6lhAUSruVNL3DwQ/2Bj7ZBqHFYFWqVLLJmZ8b2GHd
H0ICuOa+mug8m9Yp5qMT1DB7S7xWw1cpIeG2xC0DBBVHl3eymu0aUx2vXBwr02zx
vhuVURG4Fjyrxbx8GvXsohgCrxKG2ck/6AzDsTefozHBitbH72ZClE34X28fYU2y
yumOtNsko1MKGjCn/NuJksDUoLvHly6p4AMk9aOGPtnUXFew8ZTxHzLwIzLOLmgO
pwnQO6BRPaBID4Dlyi1/dl9DaTyj9sAW2QPAFT+UZVpwkwe5qpE6uy/mjiJpFcAo
h0Ze0igrlbCT3CloCGPEg1fYj1LNmTWejn7V5lBF9cvf8C+IlAzHWZPeXHh3pgSh
B835FMNcl7aSbapXPVlMYEDwkhNAs55dHKnv+8Ujen8DxjfvUZJX6dc61LOeBUI3
PjwjqqiZ49ikcBEcUHCMdJZI6bz9wYv70lgT2NRPp/VSOYsAFcglMpKA/5qBCqsN
iLdb0YdiatjD252AspcmInAmaUJS+pAZ2mELh70AvMR183BjvvLjgURGelBDfdiE
GWMaHUy44+joBAMENj10uQMvkab7xytGRGWep7rkysLrj4i2XkVXbPBLY9/bcJVh
Bw6jNBCpa7V642H6KDg8UfI4sTWO3RwbNSTGDl8U573Nen9puvuB0okxqj9252Ye
haTycK7B3MgjIkM39OMNyWLYwiZNgA1Ni8vbiY7YPCQyYI7i2VSe+zTSWaHjp3Q8
LwZEgPTWuduFnvZdsHMXza59u71vpXPN1V6yUKzCNPO8N6tAasNrpNw05Mh8zmhc
v/sD1KA5CmaszQ2WsppEtA2I8uMhw3SRkWgazhJFfwHm99xahefEjCjv59vuZqcF
QNMqboqp5uMbpk37rUeOzKNyK6XdFlBVuhDPVf3lnhFZNtMcnzwenWL+S1tthDKL
gXvVNu0egoERCoJay4JtNqIgW0YTqnzuDjnrDs5HQ0aAtyn9Zafnkn0Vb7pEfOzt
mY70Th18BBq9C3FT4MGBdSs63lhPC8VyJ+jAztjtKMlc13uuRjGD00qkp49Dd0eN
8VXuWtBRGmKsDRF1pxfDU598kkIWbDAQSjz0dJXg6qLjidglCICZegPtgf3AdaDO
vey5E8u/Jwex2cECf5CN9/7EMKrYusuF7ou2mMt6fcakDJVmt+IP8qcKnxdm4sIQ
jzBHiLBgjzFNe22arjpxqj9J7dp7VHMJupivb48IppbUyVQO9iaNC9Ph/Udv6HTa
GuXpnORWi+7urOwNnCGzeFDZM40fI5VouH1pSkZ5YSSoou3oZJRy1nPpNTrUfR+z
4rtjp6Cb/H65gbD6ezFsLI5BvsGftEu4ZaEKjx0qBKZ/NVdDQVduFCqk5OKWOvmZ
m43yJpGSLhRS/QeV/yhkOQShpDsyjEJPjzELkFzaHAQrTJD/zr+i/y5ZzuWs2tdN
RNbfOY6skediQhlns2Qy2EFY6+o47Y7gHysZ2F0FPvex1ytTatHxoqXErx+zI/4L
AJSf1Fi2BA8zvNR6OotM7WegHsqb9moLv5omIjf9Itzj6PNPTYFoxedRk5I97O6s
+x3tsZdcUJ92vlP0jd3EUfnPv9ov0K4wFj2shZZpaP91g6qHFWNJGbeE8aIyRijG
W/SwoSGwygk0VDxuwjBMaCpzznCoU4PRS27QrF3eFDX7F6fH9x9F0nLL0k7RGF8b
HW3nZ4NwuhfBWbN38sYRIPBgeM2++z2jWhfy+jzxB9Wf3TJg76LSgVe+ewRxPfzu
pY/3frjrhyCwoZgyqX229osqlX8ifIXkiRddYQTXh3p3DI+bPhf12+/Hcu7LvTOn
TNUFmc0HY+Esk0NzVfteNaNewo8nHKuVcy69dOf/yZ8yQOSZryUs2vjmUruFngMB
AsnTGx3pVPzh9b5N5kKCMejy/qanfw5O/MzqCWuAWoEEueECy7bAEo3lIwn73BQs
BA9mJKQPjvV9tzZSuLn/gRo6y8k/POX10x+jWSY7akBqx3ykRQe0AQ8YMFFmcqgC
E+RNKPMJbiMyUHLlEZ9PBwxh63/XlgD8wcCudtS74tZ7/lyJ8c/OgdTtkbUXIUKn
yLHV3+Nu6JQRcShAWRoH2bSxFIUSjhtUU37DZaFrQDYtQ+nSKfrIlZBmt1pboF/Y
Cn5GDtoPm/y8GXPpqcINFB07IBknazfhPCshZ15C52nOR+eMW95va1gRiOJ0kM0E
OQXJcnJ8iVcjLen1TtdRqpXgiEjbpCERhWY+n5rhwmoo+1DRR8gc+Deb+SneI/NZ
K9/Hxj4YZXy9eB5CvFjgt2P+8J/fEmbVidCR5X827CPdB2aVRju7/GZoQTlXfI9I
Gk4BqRsXORldmPvdS1af2pcDkurX4mM1mSqDJQyzMS2NPSRQt9IvjTX8A2GyDSIv
kxGfioujHHB0hHe2duy36K5zJUbtlF5NaBl5JZuTqM5cKajKHGiRFpUx1IgUrj4+
IvZHSCe1c31kzCl2WvcHzQlz1k6dfx/mjTjsnTnbbzasYI43S1nsKr9Z8kOh7G9L
/D9EYlLkCh8BUfSuz0SH0p3GVPOH+xnTHCc2Cmv4GvxrYPUhly7zjHHqC8ntp1aj
62mBQj5f+/XpXOqy2leVzuwQR3UYONIi5cPrSf7d+SEH29zQrYr3E7rD5qca289u
7DBPeZ7fBOuUSGNrgYGWLSBCEqrrS+ZJW4xXhTAFvGW8E4h3cpEGoL8CVo6LrkTq
jvsmgzEzagLA8jC1rvycjcQP58Tt7jkn8zTi7jBU11oXSBN5908kMxyPTWQn5DDr
5BX02F4hxhINzP4pV2SzsWKn3ITr7FMSK9D/i8LYGdFeYu029TJ2wiF4mH5rUFzt
UAXeRZ5Ldjv37gQuJ64H+edwZvHfTP3AoYasmBFiU5KvNKcsuCT4xqDLIvfxIIpy
moLJEC+1Zd8LoWGbtG2lCm6b8UXt3OBVNPmUVxeDQxoLvL9E1LpYnlrhkqLPksPV
vZxTwx6JNEqcRWR42F4sy2FX29xI1h8SDeV/hXmR1o6N9dG0xPwXzBo9awLbS+NV
MxpIVtuOM+WETZ1dpAW0RkDdqxnPbdwornLxHn8Isoc+bzbLTIYk8YUPLGY/lljz
y/uSoJ6sMjjiP5bcS+otZsLhoEHq5FXILcYtXeGC4m7LxD2fXvuc71AMIpHQUKAP
ZJQVkY0pRxK0Ldn2/l1p5gu82xdZmbhY+cq/mB2dg359yYo3Ja0mU0VlpfIf/EHL
TvolB7Nd17v9rp06sWC4+ExWvsm505oLFjI1CQEItlNMkEionFgntd6BIDzo0HZ+
YIgd+dMO+lvgrDoeMbu0RHAmq2tgVWhSaUBG63MIhDNk4++CF5YDgL3W1hZEzJw+
D3Nq/Uf+5zdgyxEVj3JrOleQiSx+za3yFmB9Air5g4oqE6Bj35GTq72wL1EbLGMt
p5F3pdSMRvtv56ssjwn1u7tFbRiQ7vzDZjo1tpr556Hn+AnDeLS1M1NtFi6bQPCk
7ClqDllCDlsOh4zoFplF6fwo4XPcmY0v1qaoLj7KaLFnLXOR+rkj+LwiYSA1Ydnz
pE+YZb4msxTujzG8fnS+cB/YjFEfViurNjCprOPcWxp2yoGyFQ3KxAxEMa5WmUV4
UOYT7M5nTGsox0DUJiwyosI0119ap0jcNnCuvjL89v4UQ6QTrxQIRYhW5GdZdiy2
R4JRHnozoLq8ywHQau4AkV0vJ6QtW/XmdIEvHdJtRKIXJQw2crlcCeKudWV4Bkjt
F+nTE4JPSmstEhrdDV4Ptl9O368VApE+v2wWIv5t0eVV04u/mdC4VBZ9rrw2lza8
qi48uxMTuXw1EWovsj6dBmN61k2hH2eXWm+06EgsICOmHwvkhmMJwN2i4/lGiVlL
ZNEyG/RJCj8PUbRJvcRdOcC8J25Qdms54za1zUl48Thn1mVEkVOslesT3pY8Lu+4
mo1B87/HKg4Stxr035eu6BjYVh1kWk1CxGjhqkantUJpEbNrH/NzK8WudNudtIen
cG5u0os2oArqwtKBLlowFnLRjzuHQjbQC5VNBZBW5VlZvDvQrlxarAzSHaYP9gr+
8CgFrhul1AMa5lyFPxAB/XNo7EqCVe2QUv7jGHh4V9DJ6crgdkOyUjPuXhB6QdSM
0hDXeYJQdGH4bwEh9UlRgvxaQa+qckVou0oivvzg8BmKpKN4jcv89M7hE1CGzkum
vicl3Iju1HyyiRKULbifI10XVWDh5Ydr8I1ougp5jkawavaeUqxW5q81dPG0wBgE
WGTPyIX82M5dUGDeRBNBesfZLOoGODSrlYi+spuxLnCEBniDnBPIiYGvaPsB12z/
IE6Pl6yKU4Jr6hnktGFSkIoA3W7UmXs8TAqKj8Cj0gDTZEoyn/KZvETe2xllC6JF
QF6EIEUPFNtzc3YmM7DQbCZi3rdcHS8yhmRYR+LPZG+SQTKk0ykyc2yMYCZ0Fj0j
kgihpX8Rtrq+Co29Z8KsxeqcwfnK2tKdSn8ubpXvHRKHUGsXqBl4GsRwyfjSMIfi
Cnc36QKmjvB7UiBjTK6Rc232xRQ4xmgekFC20fA2kguguqzLCX0cdHt2ZIHQ+WmP
pWI5KF4ZxP3rCi50rzAnbqOOVJ9s+wt6d9LW8YCGa7ydjR7bnt4CDN8e5f2HTObJ
eY5H3BM2m8AjTyGjA6iFCgyWBnbfdXHDS41dIaEdU2hnCkafQstWN5lya+tE6WZt
8rXxLEQ2oxmHu59/M2mDZjYemqluQDyyoIVq6ovdrg8dDyk1qVSEpNv9pXEXVJ7q
Mll54iILoNp44s+1tjEF2EgzTrFD7wIl4YYvvd6tIE9l2lMUaLKypd8cqdQ4XM+j
YK9nU1gsJyThpO0kIgg1jfJvwmobGd3VJiAQsVF65cNajyvjUoaALfe5rJoRbePu
fihzgTG+YUbW97jdJJrgg5ZmfBdcPX5A1+v+UdrGs7Slsc3ddB/g25upfzAjaMvB
qS6GFadouJ6AvzWmwpabKOIxvaomJUU7XZtKr2zmJ8MNQj2Ff3u+fhKCFX9ikstr
Q1xbk3FSak56ILl/jE7i8epSGFdNPkqU5fC5RaBi5gTE22rpG19NXz1w7NkG8YEz
5VrxPDL9bxUyxIhwl5iW8r2GZC+MQH1YdAcHPP/LRIUyZy825NhyjouRVMCEmOJ2
Artv34JsKZ7CWm4h0Aux9jJIxiJcQljHWqEhmrJsPNMJJVOIeLVfoXjdQR35uHMI
01Ozm1LJ2dYclioprwUEypMg90R9Q2OiMfVqOUvGi490kZL0x8UCr/z6GveRvuOj
rs40SWUbD6kW9jhbV9rwXSiaNZ8tkzZEAFgTqtjsF/JXeTcb9eTzl9DXUjsFJQ/7
9HrhX7BGeQj2Fpk5pgpDol3fbmWopzKf79EVR4+TwnAroy/wjTMDgqgqB57bQeEY
Hjo97BQaifabgBvikD3DtrkNBX6oE2UQQRi9Ax8kEFETgPIxSGMKHWHtwfjE7orU
4v3+wjVqiQwWzKIWh1iK6xp+Q/pVi+DymVZXMYC2lOn/0xWpqTcX/OjLM8mKYYXD
lsTMrlprmh3mPJGjdeBOXy0bYhTRCFot5W7vkWORrvQu590nXCiP6i/A0qK7OUDn
fDTb8Qp3Op57IdGEFhBmjq2FfdRY+X+QirXgoDGrFtq5sFRpRcGVnCISKZofz5XC
tAcSLkSwaHPNwiM+L1d6KWzCq/zIZdSFR9EzCVQjjNVrFS87Hp+U+GoO56QOOD9C
/xy+W4E1fbonGR/BRWbMjuZd9zDp9L7rppwu5OnXQWqpWmrPvpZQBOL2YJ02H/jH
OWl+KNA+3jMtkZevHLCxpeN+llDaWcXYSC9w+kwCsf8A+B7WjmD8QZVQfLjgP+9+
9blMOlOleEVQ4PZbLTJalV7t2yRqtNsZrnBHoSiYizNya1gSZU0M9+svAR88pLM1
vBeeb4dskTR6JdZgKNmrcFIC5mLmS6FlIr+NFzQFz4aUaorSq3yAU8a94TTG1VX7
oiGqpe/3FOVOg7mroz+LkBg3IUC2fPT9PRU/kYWS4KHUo9KdA84qnKU/U4DaUZ1i
CK+APXIhV1DI1zZXSyI4pvAcr5fO3vmpd0IJ8dV2U3LSYnwmqke2f2dAft4fqAgQ
wg8v6eAtUX2Ij0HfEAP6C0KPVFNjOSJi7Wqx5+guE6DebgX8ftjhccjYPUbycjxL
3VDDX1Psu7wF8tBCRAI8l+sj1RaLFGYls66n27cq28Fk64IELrsHDZOxxiH9NKWV
KHZaWZNeoNOyi4xbTFmhu1tpDdUBmaErMku2EEsdi6GKtAhJK+sKlYzAVHv2teKs
i0tfxMcOyuXEWQHB8TyZ7sauAHd1JoWVgm/2QK4o1ih/wWB/iHONVda+ZrZM7Z5c
A5ClgTxVqnn4qsYu52P31SGjOqw9RGAcIXZfIhB7PRPgf9DgIxtOBSge+BTI2Mah
4jXh0rNsIPmil3IzwsbHxYPjrQf+LcJjzJpTMEbzpNKhTPRCtda4QecWZXhEc/W7
+KjPubJYMpBInyIoWCfnaizp8gnFxdl7Q+a33ZtJJpnEZK4Yy0AHG6IC/IvvvGpY
yCUgTsalFgL76pv3NM+RQPrL13LtruAZtOwUP+Qlomne72GxX9uSjDCw78kpVdSD
HT5ep1Bn+RrTFsiKKmvtV2Q8/Yj9UYar6JKpn9eaFoMsMq0VcmzYrxusgBLrP20f
cbjvwdc8YVCplRA9lnpO4bHCiDKHuSh/L3U4iURcB1NLj+M3R+1vq9vP8P1h13da
oswXHzZXDKwAA5tZOpPBoRyB4v7s/A4xZeET0W3tzOBARiQ8eFPyQT5LxlsTkVKR
fBZ+mlrzkRoplY2D7mIiMIvfLZGnSYRPVfIAF03O+YVeIVJBKecUJAempw2seQtU
a3kwKSHZczAavA/FPCpgDLDZSdyTKN+GXlbxbhOB0TS9sNmISsfOfHys2DYgWoHe
wx7HzYRddLfBrrlbngadeuG0dNPhduxQwaWuFvHubDNy/iuqVK/lrWQKiOWaPyDF
s4d6clo0B4y9Oh3Pf9vl3XyyQiR9tiCTXk/gdTa3NkQ5bAk+XRVo9++hGef0uflc
k7n5G40nKWZoVf1CTxJNRGEHHPpiziRexggkQF8uPPz0IAi6lQBRvluMJ3O1ZIYd
1sBM6nqlTM6yN65FvDqKPZp1w9QfVzBudY3HBsVthUSk9bQzpIZtGjdlSfJ7JiWp
ig+n2+XGqjjmSQA8AWLBrFCYhJhXAjrXPLICaQFIAkFO81NhPJ9m/8tQ4Py8nwMf
qj1tq1+SIWS06UJttHF63dfhK+ZIloJhOs597aNYfTRi5rTYw0IOZZtQuhx1tQl0
TvJ9VFY0wJdjA9UgrS3vabAPTdH+MLMaITWSYZ692DPazZPa7B1m9HgVcIbQF5hd
nLGoi3MPZqtqTpdQZ0xhacBSb81cI4/dGERoO6pJGEk6v+Wcb8FpRJKtaNX6vTRy
wh2fol9QML4U/0zukXnBDcOarvF5/zYHLfhN7jDVZbgPivPg0Fu8xiffn/v9jgyl
soDcHn4DWjJbriclUQ9a+SQsFlchtQRtWVcep8wTEIBhs22bIjsU0hxWGAPmBWy+
ubO8QOiLncdOEcrYuY+ej0Wg0ShNCZy51GNcNxcRezHBzuTuNw7iV6BpMA92SRQI
3Oz0nPf7hMrf5HDqBoa+ANxa3d1aHtsgUUc4sWQdYzUzXJ6RgcGlXClPFRabohFp
nqZppX+LIgEmiIPKK7P9sXbX1gUubQnf8iQ/KAiH1Uyx69lPGHYm2O/mGboQQI71
wy96NZ2LNzWCmET4HUgX63HRqlwmHEBjfu54Nmv7i8tzowyEPl+lDup55ByXgLcR
NawZJhlpanuOCMR1E5MxzfPDDcfH3VQjjm4xCD9+YuPmPitUX4FGLYwFfRdPP5wE
aiD9GYRhoLn56RcH6FHPvopbjVeGbwl5wR9NFLCliR5TGpEBvUtGN5XG6BKEof15
Bw5U4jd4OU7qeInMa+7gP6EcOrsf6Ne+qm6xos0zHnIAxQmnZABZGhqgeKkLGvWU
hkuUV0szFkRcvBfKwbjVVVnXK8HzPPuPyXTV7IC/vrOVuOr+y7Y7NfV2NayGpPve
qqS+gejUItwEydzdsxCL4HStC4DqcdE1AgIWm14DITrnvKUWRYE4e29o6t5acPdn
z/5hRpXG+qW/F2mGjFv9//hql9UMuYW2/II/u1bR1UUL7YUpChPy+PsvLIN90Rc+
REmNouUZfY90eLz3bLVDfyUuF5burobqd82BKlebpG32Vaky37JAcXdFrCpZ6zfU
HwmuB2WfcyYAbXFLORrtyPMLSHsbqR+iu4xrDspeqpIj+EuDeKD5kJ69cVWdr//8
Lq+7mG5xn8PzdUI2vTpPZGsGYLFGtt+CcZOWm+6uygAartKMIMM3OsON8ySRtKUH
5R6MLA4LsVs/rGlE6GjuiFdlF9VWvI5XseEmw8pNIERSv48uFUPsrBZrBc5eHNfz
hXKCTxqc0pUznJ0+UfGgHNO+cH9LoZ4Lzb7t/tiRsIA/Ylsy7uMOCK0wb9AMKnpu
Arn5wyF/+1sD2L7naVqc9EeVO9sDZSSlsEUNlBXoAUaQkrQiGb2szHOXBbqITXSB
WEZ84mB7y5cZ6qf8U7x8cB33lr58R0+sWVNjPYd/WfVdK8GuFIImASC+avp86AMK
XLlJOL7rvHOZidT8g1BeGkm95lJ9NSJkG49wjbu6d3jLDw8SG8aoOQyynUQycUL2
JnW6MvF5LcW6zFaAiu5kBqRFuI1rPxzrja/1VVHgr+iab7s14LDnCalRQsR8Q+Ot
0j8hpoyPXWMa7KHZaqKMcyHmKNiWGmVRMSNT2ZkqkwFbLohz820BXhPj+yxpPFPE
gfJRsoluUj/mKzmQAK6QbdL0Pma6+TyR8l7LKguUvs2sH0EBkj/IG1Bse06qIFW6
J7wrQkii5/UK2GI/qfABZZY9wWcXg3LEWUSPAOyXUN3O5yIQbBtcwuB601CLlVb9
ZReaEJF7B2HGEubdM6wF3OxhYFiFDNolPIUcCfUbGBKoJFkpbrcQHihsJg/RKCwX
y+jLGTbmeP6dCuQxJSV/JzlrhNlVf2lZjnBTkosHuw1OtJE2EVCsd26N6Hixe76h
RDdAAkZbzjh8LOhiHhmAMtdx1qRQe9tOoNOHV0DJ2LMt8kXdPChNOu1mi6MMWbNf
fHgrNCms6SNC51V8GHgEDFxA9wUVAuh9BpLP//TaOg9t3rRH1bBNWy2X/Ra+Iok/
/IDwHjySQR09OgIbkRxvhEvN6pSBb0ydiYgBy62iSuDGFJFT09Ha3NGX8ZhwWyzO
mipSiDET4k51j8Fp1d3EiQW9B35k6oMcT+UQ5FroCwgWnzSvE6cyNVmIT4R+Ce+r
9QZZabzxMLwqXPkunD7b+5bsYMt/ZggO1pK/0QlSMsVCGTcF9GzeeLm2UDgAcfI+
eGr2YLjH2kHeW3PcouilKgcdeKjM2mz1ai8byxMEPfnWw+D3SaGE9U7tkUqqinwC
cracLHNW1Na7Sb+I67+3ew9D+FsdFNO5zRC+DBr82oqX49LdEuQpp/oilhnJP38H
PJUkdgbb8yKBnfKu+7YdwAcFblmqwDNJKB08/Jh5TTS4+bUTH6pMu8ECJhrTfev2
Zx4y8s7WfU7jKYiQ5ZEljFz82VbI46G/MXP/fqRZUIo3p/IwyTSq5jl2vDe0QQix
B9yKUXOF8TSwevE7FI5QmP35gG8J6pcU5z3fKqaCfx3TDlUTvZl34UmtM81RTK9m
ZN8+Yj4pqJJ1sVb1ZyTDtySqTUBobravAl3hNXWR/C2wcz8WgDHocFqaafNH4GOV
2/1L5MwG5DsOQtFhxjVyXvs+jVM5LLA2O+fDxqTnjeYTOn7TxXiZBkdqMww0esC+
YxPGoS/bkSr1GLirF0Y3HAaQGDdui4aypUs+N/ASIwh7lkix6xKxQDF0aXCtODIc
yiVbQmHPjYni0iXBbvlZSVkZMcUdewe1BWaFL+3XQZPbW0ZbCRGEG5yZoK3zUedQ
7gqPqFvrb4AsVVzuot4FcCIHxIVM0QIIB6gdharfzJ3NIPMe6v2TUyN6hXzUej8v
hzKPsWqyPOeQpGnBDZpUCDzRTvT2XQVxGhNqs4eBQY0t+FI3fzB8n2LR+ik76uxO
EybSC3fY0imWiP4dgsTq3LaNKq4dyFkdTW1FnXs1i1ItGfjJxL49HAYFDDfVOepi
j+cpJHkcPFihxmf+k/XTZTK7lh5wRqrec8ldQ0wPDxtiiqYgY/ETXIBxpYYvoLnB
IjavdizWiVS7aFMtadm49cJnOHnQYbFDQvs2FbOplJV64kRMsY/wpbOjzXZq69aD
9ppbAUWTMovHNvmlENToywSTkpK+RtTCFBCTXmVlIo0aA25xtoOLePIpAxZhODCR
I6+iXfkCVuK/ftDHI/W1CwtyE2+b4XdAFG6oqmE7mbNbUYjP4pVPkWWnOUOlmwx+
i2BgOvXk3swekWqdLmg8p7+T8FKC+mbEpJp0BRvSbE6VaVWZESZjDFQvN8az7GDx
Ttqu5Lrn9j/H0H3IRL1a1YAeevQ1Ql1tY9qLIgmr5BAvx+epRuXOAzRAm5LuBqDG
sqj5Y3VrOkWEKDh7VhulgWecSW28+WuGCkTJYrLt1qhuRbMmimYMNCj287ORgOCB
kTKMIYLlQOSpCNMB4JrpgcXwwBXriGtt51kqzQ0OTsNWFs7T/3OD5H0Ul5rekR14
SsadM+MeAZN0jnSUZ3ztf/huPt1RZJlvZYaqD3Euza98BEBC5Ies78DKapsgj4Yd
4gYhN7hZpZ9HDipHa+XwmcxViCjuaycQ57592Ro8tMiuGmBBhfudZMoA5rCmk5NO
ZJAPrBY1X8M49BcBuw70hhJSRMBNHeKMVApmk6MtBYfgvX0KzRvTLySZz5xRFgs/
IwpBRXdod+PP00RzrBIQHq2qNxIPlrFOLScjhaFGNY7WrBP3Sm8zLA5jrMALmtN+
EvF/M3PYsEFTa81RG3ozd0WnS1zdkmjEbTY/W5wZmEuMS5uxHrh2peEKctzGSaJo
UooWdNp0+JVARdW9wLotpZ4o95NKFu5OIEJlxUfwhjIARNGgRLSTF9JT8VkJ9T5g
1VaHJN0em2vlVc9BO/baUN1esp4+k+pe4s1Sz4mNqhQ1ttchn3opc50/a7eGKUy9
NTZ/uEJhr2rP5Az0HaqcReJFOzwdQ2kpQGWsnJv47mvJCoN5Fk4/WBuyZKvYlmFy
exPYDnEMY8svT13AvioCuO9JZmW+Io0eQq9YFcuZ/NTVh1pj2ODI38SbcjBCoz93
Sjn7Tc7GsoezeRTyDhaEX1QAbPnbdb5X7Pbjn5FX6iZpn6mYIUSJzlnv0ndjVUDM
Qov7cCpO20uQLOjScVbFv0f/4fBo5HTXh/A3uD9NZywdPOvsxNrlufaKWL3TSxoV
Jm62hklfxFB+NR0pBWfexSXTmHfZaBa9UII8f0rBOJNCLfa1cWfC53AiNKg3Mkzi
J/jkVmESv2OUujxP4JFu/HUyDVVYxRbaEUuCB7WL5Gf+Dm3zeEtrIrQJQ5/Q37H7
P9sLrZTmrawcOU0l4UA61YU5ITa3yRYCBiE3yaxWnybzuw+Upi1G+oBuVJblPJdZ
wc59XzcGR5GEmEEMWllFcGKTYyfWpbeFUzuFlDH4iqqaK4XdgRnyI6gDEQMbJey2
IfxvOe6uF6Vjs7OUDxmJJ4beyJDIi0B+M8ZZaj1IB6WgLBIAc6cxtBcLN91XByZY
f16PTDar86+t0ALy/4rx1g+FGqW8q+Z0VuJiZXRP3X3E29b6ANeFG0YW4KZ7ZeIy
1/is2MjupwoTwp0q/uw3z7EXrOUhc3RoBNtU1HjY3xAyvz3xIMhdKL/YTgjEXsRG
7CX5VSaQI/TNowDzNd/kMgL1RrQ2HzFgHT/xmhlc5t24G2h7BIuc3DMuuTpDll5Z
FiZbaq7NY8hvIGbShVm6Df5ClAtgi0QewCOeCeBVXiZ1dseQ9INKgZkpSGSUz0OE
5c0YZo53KTxr1Qws2VB9oODKMibLAcoe+okjsi7KWFYJTR60OUkwJFuo/HIcpI68
HyBVZM4FR6sJG2A00w0U6s5eFf/Av/Fw1IO7xYsynDIfXHQ9/0Le6Ggu+Jq10Ajs
KvLa2IqX33gJRwUlL9yEi3j5NQgeSoc9oysNnaViD4S8tgLXe7WWMZJSUcLXWSuX
Xq+a8YMabK06B1xrf8np/PFME8kQjI5vtbqBx0C5c3dV8/MCSU+am0LEp+brZr83
kgp5ITV7jecnirQ2icXuMH3ok+a3QWP/x4ER/ZA/xxh70WIBAINgS1tsn8YFXLS3
KqH4pjQVRDwfdgMyRCrJYicnCqSPBP9ViEGDeDzqFZNMx4T13fgJUAK8YQ+Y4zGR
skRBVzgkNDeA7lNapeH5ajFRwSsCREewAaHosj635fFLnunDJlcVe28zVVJ4dPWg
seKxqKub9s24F/9wS9oPEY4wGysOAPyprYfWF/Lm45D2lh1z2yk1m2qPITQxHAcL
1YLpkuP0qc7z/WJFFQvC5+RwMpH4rkih1g+2UK4MZ+o07ayLJ5nPbFizXJbomnRK
wvZHoO/13WmwT5r2HAwp46vpp0Q+i0fQOdzD9jUGCzOipa8zddby2vwEx9B+mClC
TI5a39HUTIKnYDo/g9Km6JaxWfC57YbPAqZu7169k/CfurC5T/FqhF4eZbP8W0sK
6QcbVPOZVzJCRYpQuFkM1VzSc5hAYkgJ0fk5pS3pIWyKQsUHKv3O/q63NBcUCxRg
zhJ/I/CR1XTbqRw93Z++5Qt9T1GOn5vAoBiorlwXpixwdOkZT3z/W+sKqoz7c0Ty
3Q8B+L636MyK/ITLOzbCadHXmu+70o6MIqwwEYJTsANj3S3h1PDlUtQWPTFhmGQn
p0quU5vD3wbAJtoh8gEVqKHHQOolnTM93n2s0veYBlQ8bQM3h0EsDxjnYhuEZSZp
STLkTP7SWl9ZmCASYXH7+rzaPfgcjkGqMgtQH8R0d5rqLN3hLVP9FayUx7rEgJA6
GU5ybkWX0Iq7V2ydpymI4/Iq0uwmV9vl7t7T0XGGT/hyNsNZskR+V6qo2agFuA9+
4RzDVRIEWI5jomj/BvBgEbvqwdKqQt7OrZMAtifryslz4onMqBKR2oklKGLCJd/O
oMRM/VP1FWryej/H8bMVOfdJogyHqOZfAP+jIW5b5akFaT9FfE2PswiXc5O6mUCJ
qnrUv/HYzy0wghHsd25nVRvsl6VyftCN9NlXPG4a7B1kan1Zx7idHPRrMyt4T4us
KHtIozBn0xXjNtZfGROoszQ7LIIC/Y++Isl+9bstWrQe38sh1mWkC6OBnVZbCFd0
FHKv8Ez+i1qMynHuSgX7xuTSeWau6r4NYBn/s64OZ9Y72coLv6InSPaPnK/JuQmD
HwJN608OvGPxXvopdvln0conokAiEVMOdt/4HwKxvjDkFJ0WA3YktiPE1WQdeKLk
H2T8gmJUFj3fPaFtLaafRIIv46vfNkeMw/sZp/HayUEbjAYFWYjfLkeXRebNnjCO
/jaoi/EglMTX7A1WapS351YnHs+fcdXG2ZxatGIUmvufeSHT0ZFj+g4mNQig+5ke
Go5ldG5yON8/07EeYMbhlvdeu42S0aojSC0FAmM2MKeNIdS1Hdv13PoqWXpHk8Ad
AbNf6i3/gaYst9RK4qEh+6llRUs81qAQPseeyLEDib/5tTm+jz/F52tCoPj8T0D7
jDKk5KML+ILwyLj50P+a7kB+YiMwPaFycYSxubFMEfcuL0nTv34BNcy1+WNOI+cD
2HlW4pePkuTS0f48QG7ZxWmSLRJ0bhgl2m2KDEr8PDNOkrIJ+DUFQXduNJB9W4XF
ZsYtHDOql8HFBeuprxbwr5YNB4UhIz0sByzIGWtUGGV8QG75pKhJce3SoyDrpN5c
zxRrcaoCNAgKZIXdfz7xEnbCi3d5hUduBn4cDdCorrNhxH+GDPV9sfnUPBx/7dZc
MgbYW24d+xlf0u/KNRo5zizFqDXxptw/koOuKbnHxJLjt9pza3NUXMW/dY8OHVVb
A9G7hbGIt9GPHzzllOlIh5GpF4KvG5foqollTrxE2/MtxlE6NLHNwfTGIj+CC+HF
VB5e/s/FvAQJ5+jxr3RwQfRbqTNQRYQQS8YHz4v65w/vCiPOhGlPzLMOBl16Hxvz
hQducAHwY9o+M/k/JkAPGOYxeuugpAy4ixSDkRoq4xs3Fc/XRSmOHQR54ofsw6Rp
sUMHKZ091OxTwUbNYZ1m7ZtiHEibB3H7OJyyQf1WwKH/dscOwWHVHoHcnf/FiIiL
cAW3MHY3QdkvJdO2I6XfsEpKgL2VaTUa4Uk0/bwTOsb2RANxafyU5/Y6CiibLkNw
IAZIxcwEcgQPTqx7Ok5qJc6v5BT61d/+nUuQAB38fhldg25X6oOujqsa/CctST6h
IW2IoxUuXqjZBaMjb2pGIUamfpc5EmuWzayWuGKj8ZuT0GwHBcRhWD5NO0cXs1bm
oYZb9ZSyGtdImL6n3wwEeTySt61dvivb/1cUTPBb5IPu73iMCDifjPu1tnN3ppa8
2ntxVjcHGGQMsdGzkbfqqjCDFXC+PZwXJ8OW8HZl2ih+aHjP48DLpXUiRLABkoIs
GiYHLyFSbq1WvidIC1D0JoThc5IqdE1Q/86Capw3lMTSweGSL3q9ZazIixLSIOHN
L1sP+LnoKogdix+cFmXysJX4vyh0GdbI2gwjmQZdRYmR70gi+U8hGzXY725ZdbV+
OFPtzTtUD7yUOr+wagTwWr+4uIwOZBY46JvHWlIWzoEI6fidrwFpiQ/reGj2INXA
9bkaNHzEA+rfYKnU9Uq3o7OV9lRTvs0VKbQdqUETHcO84SgpBE2bjpaxc3oCrQ2L
6GHmFDvuWIHKVOr0gYd7nGdMMWf0uoT8rVLvuEHxYGHkCuJ3L0V7A9DsQBoqDL4e
KDHgmMQGx5W3LJh8V/WtCuCqzf5V067NAQmQZCCCq7UzlqRKm4RLouFzPpO7FfWD
G4/Z4nCL7l2568bmv2zBVjsERWBM4/2BCRxNFL3a6yhGkLIDpBJb2vfaNjD8GaaD
Q0hv/6edPFsWrtOLehocH57eae6wdp5Qay/ousbdeI9JG/iSBHh24UBf9TpvMjqm
GndScmiJ+X7nWWgGU7iZhQhqXmKHH8VJ8Q48ZUjxGreQv44sPDrfqMLRruRLlQE8
zcgjvGB8PGf5dJ4Q72vwSVxBAM9Bypc2XyAhwG331UC6RVAFmL5w9pfIAM/DrYjQ
qbJ/1M428RvzkDEzD01z33qIma6FDHHdOC1JFPuOSt7pk+A4qM3hDUBKtwBz6day
9RNrn97zFm0T4RQfqH03V4fJXcFUCdlaQd8mAFR8EX5vJ+pZm2Be7aw1QPywolYf
OJwtBFhRbINIBdLKC+fhVza7uf5XqlGAve+xWG87YXFbaDg3MmwIiMMncxyPvkVT
aCVSWVHUB6M49rc6UdtIC18g0XwkN9CK7rx5Ue3JJwBpSRQfWqCwsJFATys8SW/j
ngBo80bPUoY4lVoW4W5M53yDaTRd6G3dgYBtVrbcJLi4sdLd2RWV5xrUx5GgAfR7
PR9ywiVBtE1kaylPKV9K9SlPHH/jHNG2i3Zl9b3Tvir1WC0Jq8a2P5/jzW73CUd9
sbsq8cwSKLtIR1DEDvCNaelMH/CPtUpzhyDZLnlBsX+a3ewf7ILbrxdrzjgEda4e
DAnTqbhJvT4Pu0YSbCyDxKSQHBhJrBbYUG+t8e2T+1UVLHgyLUHVdRg4clGK00gL
ria+Ut9ITcc3UeE6VGv9VqwVbF3tSftuLSG5rZMuP3rAB0zwF+H1lVpIHVdqPy6f
CeoVGTXnK0od7BIedgUHlbTtNGYCK/QTiDDMOy8r1PqSSwuS1KTXMVsC0f4zN+5S
0WzAN+12/3Q6OyGAboUG9MRe+/d+Q2YEpXD0MD5OkJKENgl07pR0hV66PkNm8w9O
psJgwnzh7LYRG6XrmAqUkL9LMscQrZ+WtGPkD+/Ru+ZhwOOsMzWclBFRxO1oEu76
jwrXOATC2bvynAUeOxqNWasZq8HT4YQKNWSgIEU7/XnlB93ygcZsxwNHMsBgYelg
0XU67+rMUF1Yg/XYU/6rV8JOemNniQsKAkyCYdS1BbTALZcCvicThh5eSpq1+06e
AqskSKFq748pFV8hFCh2yGWAulFfj/TOKar1aX9H1KvXQiVdQgbjIGX9vs/eaT9I
E2Y7Bl+/Qm86EgnxfyonwWTpXy8NWe5iIMriEuJpEYhYs06XoOjFThDK/Msf3cl3
H+9oxx2bSBWVg87DjBMvFETw7LXOQV9kQCKkzCDdr5borR9kgui2FCcQO4k0oW/y
pGHAxtt3OUFMPY7xRicPYMnD6a4owiqBA1FZULVkS+BZwzDWqscUl71W6bItRuZT
20zYHI7oKjmN23F/+5uwwRLJkzTuViN63cAbx/3Yk5AYFWXNzhTARTpSfrEsMnHu
Kg4ID41TAmMpBATTSDA9ev1JCXKz0rT0bxYc4Y2+Wj7sN2Tab0hZMyCEy4ExWmb9
0iXuJZ7r43Rd+D6BywDhgQmo4TETxP/zCCOz70IPndmiNYvEvmWGtkenU6VmDG7G
278LFKMZKw8tbYPanUuBesSiFSdheYGRdOoksgrJ8GpgUBu8xsxgS7JdqSBPs9Gt
sxjMPa5kdEKAOVacczha/zvHPt+Nif9Yib01N3G45qm+/RoMXZ4S23XDAUYRc9jK
/BwypjnddeqoAVcAXwPqdMf6aUx0tSodMf8mECGxzwHrO7BPqti6kK6RyROTPkq+
nMA0Y6/juMhsaq6NIkkeaA57eCBdnSB+FIBIJ8f9NsdPL7uM7iwKN2bnGnA80iFG
FbCa+AjKz/LV+wpCE8wizGCUaJz5mptzAKouC3EZ308/2oJ51CoX9IjrpW+kXcBp
xwY4TbykAXymixbi98mwTF4ZgXOmK7E6whwRvoDHhV6J+8unc/bjqCNVk8c8A+hf
FzPNo7k9+Xw49lpoYBfpdJTUDqw0s0WmFHxn+TMxGVsP8uAWlPUgwgiu5g73jIdG
3LTvRxbr2VEDEfreMwCrJ2bte0nv7spKELuHwxX3E84bpn7N29PmgLn0Qdva/RuG
EWN+NH6hbW07CsRMPkTSEqTbjPfX8w2c2pAqcRmPqeycyvDB9VJPTvHKsIgrqwzk
ADASsriCwrxCa320wlbCJ21ySG76Da46+3/2eD4u+HtOHZFLRCp9ths+Mtrtszsu
iBtbOQouisEpNresvXq3pnMNCNfnJlv2q3r5U6ANsleH1I0QY1J1ssp+jomZA6Oy
FSskBbft0gLI4bDGpVxbhQS+5Zo7GAV2nyu2CoZTYIf+GFgwHZK0KaMmVUs8NIO3
Nvyj1F12Az3t4CZ05sofw7INJejeiXcIX5CcfOuJEV1Iktl28fqWa+T0j4UKe30l
hOzMz7Fpzr1OCBew3AVD4Vn1AB30dndCx8jChff78IrC6dFgn5+SS2qtknAP21my
BkLH1Da+rjqxLkMuR5ObZHkOllXxNAoOVIxRRgX3dXkROVCUOc95EW7EaeC9zvxX
2OJbFEr6rRbpTQoOy9FzYPjY/dBGFibJpkZINzHeUacuTQNYDQoIl2MfC+RyOcFw
v14FZ8GeTdauoA0pA6VO20iWTxyFG8/jCvqm+y/MSaKfuDLWLrtafHAsJ+sUF6R4
T2RjUOdturaMJRD231fgG1mTMpp9OyYXaH435km4aHKynN+6voiKbBtdWfTjS732
os4qlFJBgIAJzbgxxnEZTO7xJOciifne4MDqeyriQGzhdXW+UuUJ4vJhhNq4WPt8
EnNq9CXvNNAUX7kclZDjy8B7F9Ljh5M4ptUkyHzPbRPeSkmeTFu7jwE9qaGimWgw
49CiipeYyoWCZocy7o2NELGm+JO9/NlO/lmnd5u305fdywIRj1AzIzc12ylOIwVb
LbNlQvbVKi867MFS3NUjdehGObdlHzo8yt+KDOCxWF7m1baEWCOOtiCRMiAwPaYD
Hj9GIprIli2kkv6oX6MvtYYLoX1dXuji2gdT402wWEV0XAtM1WmNdLnn3KDdHlkm
oJP1ksggSpzOMsZSK03NkhUavoVMyf7uLuVfY9YVu30781W0Y417aQM0TAERt2WM
153KFMHyaj4jgwzo6TOmwcpgN2MPu9frm/mliOat0JxM1GZVj1enZjCz2gBC5pTi
Sux0o71QPjFkasBHjKLanE3RhY87u1aX4x3gOGygAWjKOVIQ2Oq4otYsh5LSe+dI
RnKxbrG1nL5SaqSiPXjUzGwAz79Ptr1LzlyIrQWwSmUDZJRMP8hMrTO9Z3d84y5k
VT5r/GgGlPDhZP4SV7PGR1FuYiuR3F1GRVQje8p2KKKk6RzG/3JTvSYGfq+IaozG
Bsg6Ntn3WAhkHF5bkP08ER375BhTRW4ZqY7RonH5ZKUn49mUG/lnDPzIKVGUo/rB
rd+wQpkmlzGEDgUKg8kitObWRj4ar0a/h7uk1D3Ke9oKhGsGebx16Zke8xzjNT4Q
Rd1tgLjcheKjRJ8acxog3RoR28PnqeRHwtjHJcnLLT5SQaTk8BC7yyVMYfJalAV1
g398YyndauXRhrG/s3jdvGgPnrvGtkJ5XqJHuk1ew/FKOF1rksZoYHQfbRuj1p+Z
5XzdT2namiQibGdsCGCTRE8TaraX4Ew4aHHPjtTKmf+b01jnHXBEaSLDneq4+biD
GxkCNS41cV6C2uOyzXt8EZYw7U+n50nW6oS30AemYS/soUWNbwJmMIt0zLGIsDEW
4OGu/z5ANC2B5/zOTDPmlUyDUnr24148Ht/5d0528xb/pUMlBv1EeMeSwjZlPlTg
I8Sbv0Zd/IemXPIeck/YCrPI63LHfxVkqAKsayUodUUz+8KXnosFx9gB4kDWt8g+
cTTX3K/TGQBuC//gMHfc37j1VniAxNQ4Aunj/WDu492JSPrt2SljpnHYscY1cwlQ
MZ9V57J4d/SdgVXSrKONqrevC1zhqpkKr4X6CKgY9dGbRJoyaAP4FnLG0/A7Rhp3
VhYFDKH6prVmaTuabyU6vG2Xi+D3whpZrsr/cVAXBFwJVuwmZ2eMUChlbgYsgJC+
cWi6MpeFNtewIyw3mhBka+nnR8V1SGPK9tpMQTrb79XLBUOGLabc88Y0Nenbfs5T
Voa7jqYhHIV8yrKyflIWjro8x5bfDTSVjXqHwqTE+4CffNZAaWJ9p5jbnu8l6yVF
C2Dlnbd30MNeiGLp6fypkohh/I/2ByCW2LtumiwIG20r44TSlgTIQB1D2elvjZ+5
0ec8NawYj/Cp7QvJLUQpL1lk00Zu8Tk/vh0/i+jLRAZdNu0kQvvEWWMYhDS+bgiC
SXtB4WVb/OWwDy0KP1AjAGdhUCZgrA9B6+1Cbog4qVo2P8H7UJ1PfjqQX0JBBVK/
HAoiiOd+GMd2usSNgIqAQTuJHaiaU/HvGOXBpDyjrIx1yF6/VAb84SYaJPJtsAqz
Z0rIha62MSFrgdb+UkUhbLl8MDDXv9Euy2pD1lKjFT4OL3W4uz5QjbWjgsku2V/X
QrTsliGdhC9cFTPEDkjqV9n/C1+92XRJ0QvwY+yMdpd7mgmefGOLA0muh+iGOAJi
1R3sGKRmHz+k3Jfxn872P6Vy2FU8PRRMBIKqbjz1y/ELC8mWygNuns8JF9ZqMvM2
yE65H0t4yFisAkLy1NwTbPwa9h4/IVZ78ZwM/04HQXO0n0G2pVnplN1+m47roxKm
HqwWPUuZmzamjTldFDscP2l/0TDFo4gtVJ+Z+vE/uyEGNK2neCO9vcbOSmayoNyr
3/NRtc9aFV6chkx4hP8prspblG1XZNOoLWFZlB9WqPn2fy9Pr/Gq4EHj8Kf5TU+X
0By3dO2FCDEFkOjo/rN6RB1v6crgjFjjzZ1VNSKxLxonFPn3zHKiXEqzhjAxMtx+
2cQPCTBKQ2ozL3AQHZFnEVNokQPE0optZXHQcD1PnvHRu3d5W/1+0E3BaR33J1Zr
Y1k/iwStvAqGsl6s4D1+qpfVCkq546+Ct4tRzaKrPIwyQAB5CNbBDKuJOlYkPb1R
T4dkbPvGpUA2QlUcSXi/OShxkAQEby2phoffBZPRpsgqN83pE+SWv+QqFfsK8WE9
/DlK3Q1vaXhHjMQCArd3CAebBvOCEnXDhVqSN9Q1+WFDJad5T/bvmQ+hIlkjqsua
XBXFOR7IbOWPynbbTh9Yv5LcjIllebjEVc327mJoEVwY4gsxH1I3D190TvLo5O3z
iPEQnglRi59ROxTHJwMLewSKqchGT9AEiYJZPlbO9tr43YazXt9GdC9P4YpmcFH9
EaW+YerEWPuhCqgsuB9o100jEKKclxUgwGv6JPaK/7QhpSoQ/5FWne8Z4IlXVDVY
TdRSpVQcfIwE3n9k7t3unS+usAXsKDw3ocbQDpTvjv6is/fgAv6+9yXSV+HodaJN
IXItuV+K2lkNwcMYkL4Fcj2PULnnAbg9hH6LnVwYDMu6Z3povy9m6l34kElsDgwX
5W4C+pMYc5NwUCuCF4nHgRyViqhcuujpQIlC84jdqOA1Fe9gIIQTIc1y54Etkyj1
a/0Oq3zBgm8KNFHDxv7Y9nV5VRD4vfHh6sc8yHRiIys2njNnaqi8RHl7FQC57e2h
U16JkHX8WvYGB1M6EqjbzBXANfmytnAa3iNqdTZIEJP+SFmFKY5SypD8Hy33Kf3N
7pmMs2Xj3w33rad9WJAUwL2+XkPZylNJFV5rC7sLzrb0QdvVHCZJeePSiDTm2BR9
fvNBMPGEleLOIl66niUp+DSNhz5MdHNVK5YLzzwzGJrw1SQlVK3lBRx77HvxRqc4
Cus6NwI15irRlP8WKyaDSuGpn7ZvFQbUiQ72Mg9w78vvv6F45F/vz5EXOQeDTxoj
4bFtNCAg5qLlk5CXD6ehwkZwo18IUABQLniOenPS1K7p+nlfBjfL1DeDbAfc38ZV
NxV3mcA0U4HPaM6WE2bRKQBsYeoW5JO7t0KE7SkRIAlZ6vsK8Qy35j2rhNeGGngf
VY1unLkSGiSM+Ksu0oKz6hg7F5NYH4M3NSZl20jbOUvx2VKNiEY8wvijSVUb15Ob
Sugw+oxCAcFT+LPbr6EuJFRMwuJQQGTCBwoQYdRFseI4arNVDcE2C+h2htcBb+js
WlRxQnx2nbKaf/EMoud+v+F7iTRp7lYZBmlRD8osuAB1JP/y629mNLsAvtVoyM/W
XrUHy3brts1HbIXjkJWdgNZYFVtz5lirPdD+qCxo4Ll/F3XuYcCnQQWcWryO5ReC
TJpNJNFukVEGKdaCpIL/weoCCK/JO/chsYczkqlMtiERUlMoW/h9TmuV2X8LkBCn
140lrDKNK5/u/jXgq0kwuk+dUvpE6D3gsNYbum3qwJnqr+MeKCnnOZNs0ghYgou2
lze2znZ7Gv6PBGco6Fn8b4E1o186evtkdxAo+PBSgjWZzTnKUyClHolE73NUrM5N
W5UY3C9oex2UcaMQ8iDjtkkjHeFbhwTwvcz0CbvLWMlmIzvRMaucuaws7oPX5hqo
mwiI5BTvWEHigcpjyGFbL4qTmJxegxIdPj84DAer4ucQNjRnOjtzULYLhiq/j9KU
Q2ST70ZQEdmW52i458ceI35jqo43hJGXWd+WoVovh6ReeFAMPTlixcy1ylry+Lhg
iYLQ2LdZkaLoBXKqaXV3UFGIiforfn+TzlDuyYxkt9w/yOC34B9v1DNA6O+b7Ko9
pDJGtx1GgNu307ZAWkV7iaCqaaU4HUEpgEViP3U48n2C8Pl7uKodQPSpMQrXun8V
ieUEF1GvOP/R/+2wtHPFKJAmxjdTOWJmqbujC/okoxnx73X522c8a/1ffGFcvRGm
kHIpYz5i+R5EOU4QQKG8reS+RQhNtjXBnOqbZhAW3BMxsMDIQXvFhUslIEik4PoG
orpp7JWRKfEkVgYtg9my8Zj2rMEdiXOEJfbBmoz3JjKLCU3dv5jseHhd2r66jPQ9
lT8TMbs4qog5VQjGap98Ml9WfjpmT3P3ImGVr6G0M+rU34IVyhFSlMavhTW5EjGv
XG88jkPP1QIPcToDZMd59E7GehvJlIe2DnQKjk1/d1ROOvppSVYk/+dVDHnN18x+
UTnrEBpY6JNAsX7hGzeOX8z30LJH8LxzyZh7H56CR3aQA6n6A+uwZ6owjv92VGVn
5h7itTC777oM9sXZbb7unMbjuxxFDZ4Dasai247hWGAPZZcNP0Ye2gH0+NaKPs9r
VBhH7moQ/K7azSXRe5AXFx9/nafi5NrDVhERCnX623LrFdbsvZyQBw8+fYS6+ytu
Y4Q8sJBsXjWyxyV0FazbV7hyP/rJPCUItz/plUqqgryfghRr+7D4qkYMm4g3ygEb
nzXx/RloiiWoUJaZRIcUNAAszmzeabF++vB7jG/b87FWBgtwdXC6r9fNJea5BrEj
OnudnYvvunkr/YIhqMFYz7s2ildsjlzxnYL2fh8kW/l+E5+5i61M/kKqwBBCMvgY
zY1BmxX64E4hXjimlZ/g7RwbpKTvfQnQPl5I0T0eWU5rzLkG5jcvxzYkhkVB6GMa
xGyIB7A0z9jUbmJyNDAwWm0akBhavDFJ+yAnyhiQ+kzdHRHbm7GGg2auqCLijjyl
s+1TSG7RnwekaDBRMJofHwujGoGeVMr3nIQy5vdlzB2bNgW8p5o53FCa7XPATLwd
XN4ezK8o4o2yLBcgLnZ9kwYoJ0OPpCnrTOOQ7Tf6mm/ePFrd2cm6jOWrIyhbX+at
MiR112CbJzIM9yfHPJwExNjv7+RqvLOqVYaG3ywBUDmEpON3BhVVv/k+1RfbnhkA
3gpCRsiXg4YdUDM8sgyDVYCtG6arOfuq5rETJAqx1O+1UvMAtRGR/ibDCKzYOsvq
r8Pk/rNAWxq7NMBY3b0Xzm2uKYE9DO62rxEHOOGKcF/pJN9JmwR/lTNKux6nAE6m
a4/FadGstDeOfmg1mywu/By+J2hQ3YtxzlVoWH+q6GM6JIVzYMl7Z6xE7K7IPqND
EKweb4bRMtspLzck2xjb70c35xDToRlR5/tV4bmWLfnWbDakLyebK0LNw1IJ3nKp
j9R6fwEsU2sUxZUaPcPMkoX4sUEYZHEIqKbiSwPrRMzjRcsgLUFhpdChT6ZEUxSK
tIsYLBurGyNf+jQtGZ9oRSjl6fiGhDktdxzXh8ZLIw7brJ2qDus75qhWGDhK+u1h
LiRfgSxzi0MTpFLI8mpvD5Vb7xgQcnLX0WL7/9jQhOFH486+EJJK0/v2y96sXmxC
u34CF65cW4jE49iWGgCtWd2cy6ZhtrXo7/coBFC/BA6DPgSQ/9TRf4QAP0PoNGbR
0j5iNlszVE9kjTYNpiGO42m5CUnD541oCqD34LflyV0oanIy4Q5357NKkUByYEYk
E6YiZuGeTiAy5FPBgZ8hKqveIn5v9OPizWoSZ1Sv6K6bzJvedtqVmgHBBi0ajSKD
Qg3wsWmT01vU2p+u/VJ+8q/0XyM/n0sIqvlIyyi22p8pdxPWeNxlGW6/DPjzh6Hu
kz4VKqmKJlkohfR5ETEoviYmjNg2ct5q9DGgpHz36AyOG/oHRIPhXrYppIlhWQS2
RgdVCTtmVqvNbJcV6zO6G8/NBWe2ozIPRJkKulqo9PhOtsRJW6tkgGZB091dtVzc
gcwlwzosozNKTalcePFQiJBE7cwpBAd3KzrMdsoLSufM01zfrAKrRCCeh3+Ob3CP
++sxhDC4L/+3XqEaz8vrnJyRRK3Y9siy4xs6YXhkwgVFE9IuIwMA3vJJ/UqczwG/
gDAAvHxUqnqD4+zhByKrEND7pNBdYHBEq9ghEGINHglkn/4u2bUGPaVh4uM9BhAm
97NhqZ854WA+hBS08KczQ1IR/agmKeDXYdFMb5H1oSnDn4OEJhO00XZSnnZyCV83
XCNrH6j8OqYbMuXtU4fdNhzejHH1aF8S7ofeUMbc0spzOZjFJuIAZ36uOrgN7CLc
WdbM9y8Wp4hzTqeyU8ByWQ5ta63HGP6dJBBAD61ieIzFAUS/YGV5pCs/COiX9Wsn
769mljQFvS32PuWw/LZPCEOFY0hQRKly9hxLQ5/9Y4MOesXLIJjAZnuaM9kNBR+1
UIEvJoEM2PJkCLvKPpF2a5QKtfChoMnbA/EhOSBLwSegtRR0gU0CP+5GGLRs5hMG
fMef5mS8QIGKxzaYjo3pXxm5GOFLArPznKdkqslLiruEAnHgy0wv/0arD/ufKJZE
eJMXhwjqS3v4oxjW3iH7jBnpjZp9tFWMga4yoaMZfBzlZmMit0kV4gquKBys+bqW
NMjFiYvu+RRS4iwaWJkx5soZKf0TfHK4WhKZTyf6w2uc0u9qut6827XN/QEqtZml
/F4n0P84nvTVajDy4iRj298hso1QQBqTzSb4r5ITIi6o97VVG0dndHt+UvNkaSVU
+QiRHmEOwdqp5cck7zNVFVlYs6AHSJLcoLQadz+6U1vGi5XW/s/X5TEYxFv1xWcj
AyPfA2Eop5MiP/uLWF8bP9gGJ4FhK4LKPLPB5emYdGfqfnFUewLZYKUb9Ze/Cgg0
NX2oErrkr+jfKaT+jTwosGM2hZs+WMB0DHSFPMx7g/rdhY+t5BrKsFEVSAc4fFiJ
qorHuPVhJiauTwk/SR98Oxh/ooghuhiy/T7vSnAosRXQrefwiQCw56Q8zbW125Nx
8UlaLf/L/TWFn/jqG+3stl+a5D2/6ooV25chGUJjVnY/BR9Z9T8nqG4PChGK+Zh1
2tD0o8mXQi4PfggghZzjAUFjCj/WVCzsCREXOGMBXwmUyz9tFQVywQ2J4OGEBknh
PmBbb9qz87t52OMtzq8qsGTc9OHSIqK0GkM1KBBuq7OBH988rE/l7TFEmY8UZ/Wq
lsMBQL3LWQUSzuXhYEoyrXEoVIl2GImrM1Rx1M8+/2Z4aF9+AZZEQOHSP/3PdJ2o
l2mcmGdi3A7XpW/a3aLas+ytQrALup2f4JhsGgXMQaibFJ025ZSeh6NB6JTOan7P
kHe5JmXxyqyoWRrwvfcNImPrsSLBkcMw2qKVHYUYEO+4dBjlGF6dbpTlZub+8MoY
wBaAt+clVd9KkEb9kKGpY5xXOZaHYfkqYtrhtWequM54HEBEgQQZVh2kbm0TgJyd
e2XM9W1v8YmIMG92PQchHvmW6jJNWQcLaZy6HgaX5zDFnjWW0Iteahtc6t2P/E8g
aUY8zZqzoHmurwiLr9K3949r0vhp7NmLGg5BWRZi29Sr1u5r5nj3mZL99D0ppt1+
NWoQ2Ok7RtMggjbzUp6wtJSGZvj4Y13q4SjiurxQ9o9bb0PSupqEoCj+eDw/w8Om
R2Pz3pTwHO/n45ExIiHC7yCCaUQpOzfuehX1Ya2Swdn16KYGeIlEfYNhJwQXwjBu
kZZxZKeeRtr2WLy+rNqHjofflNRYwfLM41Khf8nEDZ164CI+NF5/ou3xHPafgl/9
TkDp2DSrsEwpP2k7DI2FEdpOzOeMeLTrklzE68BKPyZCwfL5D0Z+0FT5pKLglgD5
R/YS1RYc4BVEHkjoRM+HtBr6QKTsIW511l+xqsf6Y4Yl68QzHf/ZZzBB2Ek+o75k
dOZqogP1ximJkOHcwy69M0WO9FjYdy/5L8/7t6T5xRKsUvJA5PfbbwwqkyKmCsGw
ljit1sUGzuuxKP7Xb1fdutdbZvAndlf4T6HlYGvYK3dM5Q9fBRbHuIhLKLvIgOsU
350WdqH9eqKukdoXmgqshVrJGkbwCwp6fy0SaA+0PtBE/iEyMhNRZxqq1YuCw+9Y
j6FZSvzwTuo6ppuWsq+gkRYHYL9Vg6RajDZ1rl+cY9eV6fUhgIQCI+C5zNlTp/Xc
uzQuoZjQmI93PLii1siV8OiiSPdfrHWpQ4u7IG6DuKs3LDACIDx4dJ6UIpBp+o2n
ENkYZtryddrdj3fZA7kywltQPE0zOQKDiWop4MUKrwCLihuuSKg9x0wJz+8frRi3
Do5q57YzMYTNKX4jxdH9rOjPTbrcWoPOKPRXWm2W78uD8yBTFrfiLVVenvU0dkMb
TJ4A/UaNSFV+zhz5tNiu/OcIRB/5BlQ6KbNbsdIRvbOTndthxR28BORE1nmhPIAg
uuKa9HLNyYdkWtsW1THalLQDoIUehPCXdpBH0JPdMRx6apVZUg0Uz81wS+DHe4qQ
n75qcmjuNourDODL5S/rDD8Iak72xXvAZ9ItBMV/7msMiMF8tQIRMNJYTRKAyLX8
LzE5G5GqjPuaijjVBbdb7ZpHlQSVuXjr2k6CbXLfT3avNbuI6/BJSdeK16vcmZvc
5J5wSDaEr+91xupz87e3hZNGbSBd0O0h+dQYkN9ZxfiwWi476SeS+0HikqoqIk5a
rIbxykRAxr8XfGef+AfT2qHSzwLfzcu2fnJdnw65yqeeAeP4J4llmE6iLkK+Koth
2LMq0i3S/JUTSvNpyMkXpAXSPP3s4blL9StwskVUr5NO+DrkOk+FEmo/1tLUKPus
Ia4a4SYFYLUUrE8sLWWMMB3RSWkb9B+UGRvq9J/FGkNLFHso5s0TVv49AJiLWH95
yTomvxYzewxRIytVws7SG6Dj1U1FZ9Y4yF8Juhj4oVz06/Zy1t+vlOpVA+fsqZJC
xTCgKtM+bLysAXVxLsTJ6JiYKlZDxKiRtv9g2kkwdJkSFvfbNpxeu9MmFu4WCXGq
Md4Gmcjx5j+c/pIN21kQ3oc9+5SP7myujCwrNJZxTqD9W4iBiHbiDLRm9nHg1AcD
fRT4NqsoMAG3z3ewMy5DYk9rB7PhqAtqe/kW0PI2BSFGaBbnvcUA1HXwQspu4xii
COv5qP2OoBJPSnZpIFVgwhVJ9Ig4bE4WpmaQZ0Mjqe/734Fxga4QlF8uXGJWKUEf
4SUd6U+6x0ZN65V7yyYOijTmvSTRGSJqats1fGg5aL5r7ZNMUjofYbcNOD/FJadu
I0bTCuZ8ukUmQJfDRzsWbRjo3STysktAUMfL87oBjArZskmTFIOhRDEkOsWAwqr0
4LzVCEvX7ZxhtV57ja+6CMTT7ivghwHkmkfHg4rkEIkGs62x30p9tcLyswfgcSxO
XS0Cmm73gb+OpdJlQJUkP1chis54UtZhBK1FdOO9sDtk569Hytdy43dFnerlfMsK
SAkkXyn+hr01TuBM5aOB/tNt/peRFy2wcFvgJYWniye4k/5XGChprHgFfXy7mRvw
VHRWp2XHyPMoW7CB29pUT3vWVx1HKlG1LVPeFRl0cIEi4koz7CCbBvxI2ef16/jb
gH/UKa2vV+G/P/6QmNiogRAZoT7WAfQ0T03i31g3vcWHci1Gae7yLXaGZIUnBV3E
TkMr041GI87jZP+T7ayTjNncwqsaV8gidEqEDCOn4ywO9dJRMcpmeqtPpYLtbHIU
Iw4KVC2Zp4bLwm0fPXMTal7Oo6V2wXR2lO8+V+repg0LStWdY/xcZrdQNiM6OxHV
496PBVfwMXbkpkJK46BB1s8t86hCCdCEEp+obJYaJxwLUzHiSxFzNPOhfqCNXws6
GL92dJ2dk2wcZabGC2xKD4gPSqRz1MfTZ7k9KbQ6qDBYs5uLzgJxA2d6N5eHImSq
c6BLZtizd/9VmBUJ8gC5+j9y23UYuEDCCkOGftZF1sJ8QtrqWGoa6/kMcqa5DorX
9m5bYHlmdg4/q8CFxZPv2WWzA/ZF2ypVOX2cEiuV6prWPfHO9gxCWxGDETpnc8No
2djNLHs7WE9zH1VSdEo8mNsYV9SRM1NBakMkVYdiyznfCZsSOC0Ohr2X9YIIcaIS
7YLgw2v7Hq/YS7EGCsDuFwAjlDxRx7tnqsk8MvI3LgJPxkCpREFo+B/FCso7WS/N
nfZjzyCW6iE4Gd/KuYuURKyIgKAnZPxuh5Q8cnCu6s7JBqDYN9iWtC2EYiNB287q
iAFbUo79i6IwL0OnyXs7OBlD4ClUYAq3xMypbIT1lDsFVLWKwBAKK36ol4xOd5y/
oGvB8mnPPa+OGdX6NBEpbG7X5AmOGypzQBhK+F31fRK03hueCPMRBIcNUG3AIfFQ
+kacbBFJEE6yeOUAnaEiSrgcHBINgfNQ71cEiNwKP5SfxG4uZernZCW3PmL/Igxg
QkbfmWTZG5NJDzm35aZWmyqeOUk2JuCbgfSzdydGxsWB9ypg8JTmeOZecwYX4FJR
6pbTTgBJ8/xPI8fV6u+pGFLusLrZxyzWo1cb1wl3fuIjbVQn6Zq/oOFU0gHkYIRc
91Lhe2Se39sf285zScNeC6EbTa8IaECg/eEUD3ABogOkg9rzWpXAqfcQy/eGWCDf
xjYTd00HSsZ+qFEMJpIw9cOlx6zo8cxD+bYDTN9dSKjDgcg5Z1A1bCPTCXhLecG5
yb8HEwbesLVj1mIWYpUBjZkGk6gvWIcjf11kZYPcf3soaI7NvKLo1KFidToK925A
XLWYaWeThbEKQY2AIxHToVHGlJD4sPv0TF+zfxJjOVOARRQJ9zf/esgC4+TCqxOQ
+6vnXHYOHYe6JT8kLfp4XxkNJu3Lzv/YBaw26eYFgmHCjUGUhKIL7lFr0VhYWxM4
rXAfd3UDh88ufZHa51A9S4UtQnlfY++x0WhfLs27kK3MewKLBBiZZLzNBSExMkiD
Rh8lnMRkGR1B4CBV+kFKaAq1fMSd+rlT0oeBcJaX3oRKJa1raryAmPg0FY6sbwaJ
hateQ35yMw5a/wOGJNQyh25UChkjrODbMnYe0oYQkFecVdRg/5lR3dTPmlDE9yRU
HOfjtuet3GsEWPtwzt2Y/MSpexwa+GecpPV9N3hz+YuOCVVRDBUEIflLZmjsY/FL
uq4KKj5bvxQPe0FC6VhdeftoDf5Fc8AhueuS00XM6WYgkvPxiB43pc9kCLu4dW8K
p5TrayfPSxbMNCtoK8lQvKsRT+FQmMLBI3tRLVOhSiOMGUdsrRoafZVYkifx5xRv
o0d8mpUrtFQbNYxcmHuJF69oqUecSyltbyphFHZm/zNLPk+S+daY9OCrAWVRRaLi
RYcFw9BAwPfASbx/3RLUTYMfCyVvc8bDrvPMedSLSl0CGjF1VZC06AsUXCcP4ibZ
0xV3pwRDIcwZgS/vUp8cussSaMu5fVvNMm4AvwKzEhd2sxXTCmAyUR7y7c8XCPUB
bpulI0X8+uW8Isel61wekcdterfJbyNE9AMfVnwxzn4Dy2enIMr+9sOx85aPoe/Z
ZV1QFgNHgxdeGH3HwyIpL6osDodCYXEhu7JoIpzvwURWregBo1AnD0ehtRWvMw5X
Bh2ZDLvZ/LttkOKx4hwNizeW5d3dRqLE648XwV35HNVL0mA2maazCa+9BMdnAKSW
nqAFRHB7rXLtLyQuXgff+oUobth5i1mXZzAEnDxkeCHW8r6eqEkhZdHIbvvahE1U
Cjf1sMyFhl3ZzyYUsSEoNG34aIoiWX4pPUWTYtzWYoKE53fJ2DCBlLn+8IkQOsCd
MZUtXd8Z8VqN8VCESyORUxGRA+bJ7P19SFyzlj1JwxxWi9Owuoh+bKTSO7LeEmcS
/njL7ORTVHDH1kAONvhQnIsNu+HZ4kejVWx9qglgQe5JrgwjQa8qlpUgw4ZKna6u
HKYl0k6l6YrM/ZvGAeEE357BKWVgzFxYC9gRe9kC4rUM0rs6Z+oizszLHzkGrE7T
uRno9jd3pD5K0nYdBCV61uQBoPMrlaaGTS+Fsw/QEdolARgMDODIwPgs5aDjq7us
zT8V664J3JWc6CIJu1IhUQ0SyhZHt7334EjSVSkSU+cf0gsH9NITw01eShXavb/T
oEYkYLeKXHmlcUdWMt0PNh4BeSIvDEz4BNnnmKabtUL5ASwoxGK4+Lpw3TstodmX
viyGPpqTB9iX7DSLgfHqCXqdXk5j/2e2F/ggnPRvbqiQxEIKCpS2WwrQC2y5k4Lp
WAzB23SybF6kK/Thno8IpVI3CqeIXd0X+dQgtIO3Aup+QFtlUWqlbHLcFkmLxy4p
LRVHJU6KQwTgG/1AM73lerHCzJo5/9xHOJow8vsRgMNMdIupV2d+w11MPdHOJ7wa
DJ7vnW0HlqPqgxZfqRYtL4WCNHLCny094eITEdb0JkEYUBZrTZfQQmurOf40Dwpu
vBA5+IrgxYMYFrbCBauQyBQewqFbY6n2zjxOijqzdnH9whTiLINHe5xQ23WiJHx1
a/Nmx22L52SGppvL4GetqZ5LohIXCeoAV9VE4M4OHuFvK8FvItl6G9unHXWWNx3c
P0bjYj+IRKUTzgE33YhbwlX9F4ZDXTHjHoCrk4s33g30Slto2tE7RPoee7w3H7Mj
hswKnMLsRdTnkkua/GWsLupDNvi/oynR/+MNWNa4BbKKesarVKYKvMHJAGBCTFE8
ABcirJ+Zq2Ap3EDoWQLgG2WQdvtB2+awMtAjjYRC2WVEr60U/1RpnKbF2TmaV+CM
5AhC/NxuVsXTxZDPta2LF2zzXW/d26Ts/sNCXyHf2r/8+UBrZA9Vp3ewguimg5ik
W/GmjH79PsAEjkNce/MjF2ThYwMAPCHzBZpV6Lvt7eXN2G5DSGdAbn8IpNoIKC+Q
zrWpBB9FvTJi4nFPunMd7faJMQOGCBEIRegFLqcMWxCuH2PBViwm16TwVvhv5/TV
0bn8wKZ+wSNw8OTx8vg+xRhbt/eiiz6gqtLPSgKlMSN2RDHzpjPszXg2pHbBugXA
n/BzuUokn/JOWyfLRjyG1ZPIETzfzl+0H15AELIKVnOuCG+r+Oe+KNkk0PUoec7R
pGaUB033njh3afy2qNBWcy+pc3iZ9dm5Uz+xWakfaxqUqVqzN70anVzFCrxORyO3
ZS1GAm1diJd0ftSoXCFLthwQm02DQZaVFOGCSoq2LPO2DXVEbktEqroYwgHeCnhN
G1q7UbY0SDCv3dYvtsSEw6go71FzRLDT+tF8JDNmyYqIaAgk85jSFpRqPtbyC+NA
T6dcHtx1zJpBahJ2kx00yYlsOq3nxBbv3A1hqkrn0dGH9Tw6fSD0fYowoziq0DpJ
GohJS0nzAZpCqCy6T9iqpTUeYUg8TLdrXBHrwdFiH18WVSx5EF5vSlrmhl8ch4h+
q82Fj8/pvryWKOEdmRzp1Y9eQZLmjn55wvOQX9k5O+yxM9v/ZpWVOmlfeV8tHY5H
KcUzm/itBQeg18srthBwlkiqc7FYbRdMPjfo8iwBHkiC7y61YfvgqkSFYwPF9Gh3
Eh9/1Kr09V1G20LnrkSUYYrh1a7/oWxsriGSYqdy2jXoajpocPm3r3WCl/cb+B7N
Tuw2nIxFCk8SV8y/GPUm/Nh36hRPZra9vjnlAtbZo6fd9wGIt6vQGxFSYGAbVGBD
djmpTIiT4wI1nhn7R7fJ22TH3eJqdG+oA1lOVM4lV86MpuQzrJEEkJdw8qlXKK2f
wh5NUztRYc0nV4TW37UmYginqJl4sq5WV02hYxusCiiFflFpJ8au/d32yaJd/ylO
o9hw6Jpruw95rPA9Mz2oVjW7yLABWfANvfCk1L1MOZ/zzYTwCYzxnwjXaRPq2SLs
dpfepckdix2NLzuLXrMcRmd5fLpVEZulh9sSSP6cCTJ3IiyETlm67Zd/DY20ZDVa
ckzpEdlJ5muqDq1us+qj4b0H7Q+F0t5qGPRMSm6MVA5T7TAtOw/V4I91asF38bfF
K6rwEK800/T1OgDYc7X0YIIIRwWzzF9v5Z0LFRZ5L58hf1h91EOaXvRy6xRRyNJW
wpoE7R9ThoFXYnwWaw7n85VzgYIj0BJuga/DtK4O4VPIgoHDtADqi6HoXp7m1R6l
03QYXVfh33y6ZQ8BPKqRg2/r1Amfkz2j6TAjUoT1wnAPZVyQ3BLqeQIlsz1jkw30
IfaWWArv9MwTkmSU9vLmVI3+EoAbooUhXJdWoDRqjE7ajkhjmbFCG+H5eqArcQef
kXpXSTXL0mGr3CBaPQXxBw3xk1iO2jUFBhINGqlbU3kmio4DB2mf7A6/Z4OlEOwR
rbpB8xEodH1dteBvoZMKsQ1MAIXEvEA6XFkd9NsJpmH5YPUm1FQvaU3dV1zNCw2t
58jJeSMPIq7L9GtIANxJeEpuqhJzco9fZFKlQYwRxQHimDuRDoYRQJ6xyxQGer73
KJ/rFrk6fZ1V7cbufjjccu+6YjJMcWSevNFbFrI4UiD41I8Zq1javzejAQluB9GF
1jKKuLjMmizDNvuHIv3aGedvvDCwzaAntCUpnOw1dAbCMgGUaYsFGJ5Mom/2/xTJ
AUDkLr3ObGmK6oNpjMBs4VjsSERda+8PUEj073WbldikSQpqrjaBqIpj3UPzeK6I
rKnaacZXZ590x62+WEPwldXM+wBGMnnz3C3VLkEXhwMmaHFjoxLC7KoqKE85+0fJ
pJCE6Codfzodm57NddPxpHd6gASAm1wA+Mp2eJG+MHeCOGLt4m7M4d/zvMDTeI0G
3z1hOmJ2Pd/MYUcp9rlU4tLaIQfncluPXPgY3mUVf5gMNczmWRlzNxiXJJnpVgK1
aLmCqVpw4bELd0RAxi2hYh2t3elMKwnS5ird5xIKXMq/GmY7v/2JFPE+PEWkiTd3
VQdUleXo2a8oNml2DZEXnWDHwboBxnlsPasEwuaU4DsRlD2h8vY2Jh1+G+zr84xE
bhP0i6tzdRa5/T/WrOD7l45RzHj99VTe9XKISnnJ0DJcDTXoJSSMHXMQgpvv5XX2
lLq3n9gIS3L6/oFJ5wRFkRRPbtlmA4nST2f0oIJSTLUAv6x/lkKfUFs/BjtCQcbW
SHQBlBs+TMlLD/ZOeXeI1mZQtZK3kf4IZITEo3Anbd+8i/ZrTrY5TqHHgs9sYGRd
Kuhgs86X18pH41ln3D2jIKXV8dysTEuHy2zi4yxCRL2A8wOMVVQi3lQlvNjSHUJq
AtuwoTT/9hT7eax7uKuhlT/ZhVPR25s9xQBh/KNC7Y+ZkdjXp64BKuMRYmDlshC7
g308YJGaOIebufT/nO15yO8wzC8XtxqT+ocbiKQkZhLrDSoZdF7Hj49vve4JO5Ch
RX9ZSTEI+p8f88RFg1b2AVBvqlJKz/iNJdFCkRzF0SG+DPXsfqdTpD6E1dGFXHnt
NEpa+KzLFJEDQF/VPRIL+rA0NMdMIltu1Hgj6xiAF5gYBA+ZAeF8maBGtDYl7PjR
fLDzjLVOSfSQqA9hEqoHpk17ejKmKrn13FP/P3ySJCEUnsssZT5Z6d1QTgHS6waA
gFHD8oRwl6VM5PaFtAo+Ab4EgXXWhl3o1+aVxGkDEc2p1FWCVyME2rUO0nmHGaRA
S+5grF3E3wEvKByrjfOuzaHnbbNvWUgg4y4fWqPdziPSTKNK131I0oEPhddAyUoT
q6zr1f6EFj79wZSOYyznThnMM4o/a1RcSNCaXAscCpXC/GpmvrQadiXkVzTdyvji
CahgCX57JzSIzVth2gNLI8ujnyhxVi6N8saUSo6OBmFTp4WlE0LyQ2sZCIdbU5+a
g6He6JG+9wXnH1/qrjSf6qITD8hTFbtW4B3yw6bBiaCWfuhP9Knivnm0FJxTtor0
iGN7bYlmhPVbjdnXhmP9wBmsjLB+f/wIn8UyTGqOioiFWSBjv4c717ZLG7oSUr+S
fyMwksn8/dQ8u9YLk2M1PCphZHK+imoty3SfPZScZtzOQsbqyzmj3vIB67zWjDdL
mj8kHs2q8C3fBOvUV2Y09XbSOGi3Q/BxX4XZRIv/omqmzERYsKq/UWp/x1JedAVE
c0bkF+Or66n4WvVZ7bnZvo1gMlSEp8vStYyoHaXqYfKSeGcquTxy+Rj4hrbhMyE/
+uKaYa7Emy+yNPR5fd88yi0r8yEW9DdQUOy5VJT+FqZCvqpemyqozAa0iYDJgEQs
4XfrgqjPr7pUiUwDOQMowsYF3kU/IM5yX0yb5695mpE2F7tkgbfRaEf5AR7meJBZ
eCsfYOoD5Q7gc5E/lPLbG9iVcTLU30pHOZX0aHcVY4AtY98dwh+5E8ugEVgfSAzC
iAfi4afRvxqW10BvZBSfvdazI1XRJjjLpASpGyaNYdY2PYBYxTWMR6D3T1RtAtij
VxQaYTQ2O+tA60X2K8XmdudhryBvDSKRhGSgqvrs68LA8SmubVjqpVTYH0GBdi1i
OlMGZkThzu7CA8HkCGYmBnQxPu9H5NN2mhQ/HdOHsPVZ6AXY1Sr1OWEi4JpaaXWW
m2PtQMcJGVux6zFT8nK/XLY+MQyRUM7BX57ep4nTv0buSSI2nhkKdZIFx9PjIcvh
MP9W+U/BNxv3wlgPQ+Whz4obRXATmMY51qy5bUMEfV/YlY6J7orcx5m2EotsDai0
xV6LQBMzyZd8q/SwHpU51UHg8JDXaUcToM+s8AYv8Rye+g5tinGajbFUogIePnoG
8kmpdyXvyYAJgD0eAor8qo4yOabEU6Uuuj/ytgnZclN+ujn3aOFwcYV6lCzhLSkU
HZCNk0VX2vDyuw862L6XlxA6TsUot9XrQBAvQFhE+hRncDjT6Byq6tr8ronkueHu
zxxf1mjr6LC/8hAY3HtggwsfuoDWY8LFA25vOcbIM26ajR+yL0FZ6dJP+kLUoxxX
z7zWKzIjJhG7tDNHQph8KE5hJ8h/XB+tkuo6b2C3LTw/f2/isCzYL/OtTPR68BEM
u0R+Wg5Idzn0tkYLvNY/5cAPhO0dAyTdLsbgHImsde0KlM6VMvX6aVMhFjLxHBSk
HW6sA6Y/+oTmrl5eAjNo2cwj60kENpuetBijUygPWSDKXyMJ50LO0wINQIBagJ9G
yHXtrYbtWkpsBfewHMmVtvCK0FDSNRfw/5TEqbiTu2JzwvEb6GYzG7qSzpeecyxM
EqIt0UafYNwrMVJLQzpNqNkllCnDwDePpFUCc1eq84JNA/cpgr/1FjFBKIAatlbs
jHzeEAmEph+sGv+syAoj6u2skhDwPQWC8/jB0wl2iXO6YODsEETJCHxDuZYLswS+
+syRwL+qC8EcGG5DbvPGBPbrbxYoVBg+18FzrdpH84HDYtt6BHvuwcyK1PBvgeUD
1XemBngZtaVTPXKRJmylpyIz02S9rFNUTxFUbprVE6tW9bY0PkVKYpo9t7QxxM04
IIrxtcgh8XK4XRSWW34YJJ2VgRGY2PjK1aVGFTWOBrZafeZ/l/tUygEH6FHzRVdO
SnNkqT02Ktw3MjyzxxlaP3IkVDIuY9CjxKUiJKgn1H9PUDfbnMPJhmjp6xQqjl9F
5pvhPtMfPZmL548hOzSwofABfCCRU8nhD4d9lXk+diI382gIqagAv6YY9GMTRxDQ
calhcnzrU85t+FEJzo6VTgmcjPnis+9zZROq30JJLjgsPIxB3OWNJDM7gbKE7Y0d
68XglZ/waG4Vk/VyfZ5766Jl8JHNZP6ZC7zEe4nVg4Tmemlr8Lks5nLKzqkQp5TU
KkyIvXO2RD+ORRbSmfOE7xyscN/0DJlrvpUGmhov3duX0zfZCZ9RIYTCbqY03i1U
7hF1IWif95w0BWDWkEhxKCN4r8bP3DUHQ2gbBRkmYp6/B8ACu/VpL2HcmANhf/Sd
WfBuUX3StmrhH51QFMfWQYlIgHSMyG8FhhEOjStxkrfiVwxcsBn1ceuREhgg9jbT
2mDip0606x+5WjFCRKENm2ydoaEpFIacQuXn9tu/f1v022PzhTNS9IdQevoNhMkp
tGK7ut2CEi+EWjI/zQ5rTWBuK2sX+A089ZRYa4LnBqj/sq7ti7P+S9jXVXFXnyYd
ivmRSMx3x3iHVVX9HuUe6ynSVSVAUBeWDqgMJFYeJ+bB1ycK3Sdvqhc5CA0WefSJ
imsUlt2eHSy7E5mgdYiwiltSb+8fd6kXA6kMCRNWon6NJeBuPpryFg8shWOmGwGE
lq3xoVSsChuUPFj9UcrvzVo3XYZYb1DHqBhofv79pTf/DjAD2zNYdlDbiWOyF7IG
59QyVamrM48pVCnLtjGVX3Ubr3y0fKYldSQPv9iK/5fxGwksFSaHiws8Wcfa6RtH
sdafSTZKUe1zhu0HydTm8ATqLiOeA9tkwSBI+OEgMpAMAq9rhak3JVcpWuc6YvYD
X0aKjpAHbN7kSLCicy7v5aKHMcg2m97PxVzvj1oj4UDUYJQzE2ejPOOF1QZqsWXk
xAG9OUyqP37jGPH0sZ9PGPWqDzDd1WuuvgIpQgrr8iRMMr8C3dlWkGBFRzOGTXrr
SIqkATEIM6Yb+26FaFyQuu3qbxxg3uqFvNnPu75SWFrENKZ9uXFCj86tFvYqtuqk
JEZP+CHwMKWOhJBiiDhAT8Xtk6fxLb3kvA9S3xC9FjzEOym5QENq9+0bCZ60TbvO
bGwSRPjl53Voo7fvQAzvQvovoR7FJGn6Q7qsq5VogQIRusFPVymfV2Lh37YHe621
5tKOTkF0qCujYAN0MdhqfhesSVnCFH7CnK1zhj+FzSb3APCTaHE/hVquLbn+7H8J
p82lv2Y7gYZqEeP4vdliZDTODDhNUZz13/Kky1sPEqNeF7o81SBryyFdsY5SKCuJ
hrMU6ESPuiP4qp37U8oz8wO17iR2ghq463r29FRuDVE64SyIXSm0JmEW3dux44Mi
wLPyL7hrS0+NUtK5C4QMEVK133t3DmQaCYYR+yz6r3tNmQ9WIrbZk1XyPFSo+EPm
EQjYhLnhTCLZBxQ3e987JbpFoISW3XCjnNEATlPB0ghxOvlH29FYbp2+Ecq7A142
ywfmzLHeQ5vqWKf0TFUHHFoEg3Q3uaVVCSTwEDE9o+RDaNIbGnYb68g3F/1DL5eY
I9oop7qedjZTZbTjwrNx1rVQBbuoGKab5gfSckdcneEeUXmHMMF1cxFUyYsPiDX/
YySdUKz1beOXR31SHT5q9CZz8UGj26bWKx2e/4f9W7w0Tk7Ey5G/2PIb+f6jaiSo
ZIhvazQo4uJBefKcWLPmC2UpT2QLKpZF1/pGPFTd0//bpQl2dPIWQxec8qdz0WOi
nzGR7mdCaGchppmdhqpQGJqSrgt9h2zdD+AzVDMkAc8TMybANy62lhQF6/0yARL5
HgktiKZVio3qfheXKQ+GjP2qyE/6W6WDnApo+r6TfGvvmYX6s4jsg8rglxuNJudc
BA6UBJ/xoQwWZaJ0p7qf7iLpwv/s6dEXpOSR9J8vJ8h1Isic2bTwnZN4MkWsWfrq
l/AR12KIo0oYb4nAJMK+wyDGiLHlu1iQYteo3Dn2IcT+tznna2+afZz4qq9YLEB+
dtQgFLtmr4COq2EWhuVSmSRVD9HpU2yek+PELLAknaDckHWdJAsvg8XgsWwUVNzt
F+YRF70JC7PGPtsvpfTQCz4LwjWLX2o9qo/kI3iff1Y9cCPy8c0tsAjeX/E+p6h2
TRY4VbbPnCMN0oH8bAHQot7DEJ1rwf2tGbtwCwisubKojiXfEpy6SqgCDNx+zlhR
hlFo0VpQ1LT5ELfHEfGdAnAtFuB7mdphrEDlsN+P+XFzGjvU9BzSA+feBGEUKg4d
6JrCESHdQVs4oi3Jxw+scMZ2v5fa+8uzRgbzMUWEOYOifnfhY4weyl2jDH1XURIA
As0lpNfjIGQyx4bnF0JewBqlyUAlgYjy3J1YNG0PBtpesxlhE4PCp74zlUJmi5jx
Pp4tboj2Sqrum3iJ2Bshgkc7FgTsIXk7eUwQUftrQb+WWKSRJrn/81rZ407Ffz1V
ol6H8HXom6Wvx0vD6L/9SDrJbRK2e1Luua1gSgRxHJ67rtShK/oOxcv9z14Dx2mA
v1mvhUQR4nvnC7qQL+9QfTRiIUohZmaHQQyzyqEiFNqxx3nWLH9UW6yQfdxDle9x
Hgb1YItv35Qo8uduoVfXnaRomwQPXb7F1eeY4uYBe00fJeDsYhlhVAMUND+hQEhd
T7SG0iCdekGQfgJJLukB/MbdB5hUnrMOi/4IY2zOQTqydZB575rNtNoc9vEJ3+32
c4A623j5z5fZjlZ8VRwqGrG8Jv68K0a7jrcXFMurxdL3kWEekmguzJIILw5tvenU
L1hl59NbJQcdmTP+VsZKVSz5QTysLpAmCj2Fl/Yf2MdO+5xjRGUWFLIfefqmFDXp
IuqOp5Jj7R1wZvI4gSr8AbVeakdpzbl8VvzYsVU60XvoksPv+9hQ1PU95UMC1jBo
sgCoQLG/NsLpKbwlE/1n3sRXn5Jw8Jf9lWPae9JI7+61zfSKUY6RjzkfgDrKzh7e
28DFhxSnsDQfSi5+5Kcsx9EWTIq/lDVOEaqlNHPPXJ9w+HBvatBgl0J+Egp8U4c8
v1JfQP/su29WTA3TlFY57T45/N+9/VXU0Qvy/fRg/1TC9IrRaKlGsHAAMqrctp+O
RRe0oZIs/0ujA34Te/eRRNlYY/YFdmDaeYIRPfVWX4Kikvav/0DE5Dfb5/g7jzA2
uyej8llJMrdJrfnSfsMi6JDaIGGOnl2df0FiDZicoWFkNbx1JwVO09cQ62mR9yOf
JHBKXmD76GvbL1aTWvXbEqelRItD4l5Aok6aorgGOq2kmQrLmQmaBpgPbtfdF7UZ
7WkieR3riAqLlErUqTN0WpuDxAbUfuuhzt+AyKhJgMw/2UqPwK9hOgDoxP2VrEPF
3yDwswfBcaroPja+qxyNlX1sLUJnNrmlHTq5BejEtHoJOhnyWn0L4+lxfVWimKDA
2ObeC+VCX6r1tAfUhmLEj07s7VIAu5jIa+euN3tDvvr+kaoOJ64IzCJoPoF0s0bG
CXoBlo6RzedPwcvGDIXCfOHCElZf6rn2TDdUkVC4RwtCDL7wA7rhcwdlCxrNulv/
Tikl2ZjAeHmEUjKEbL4xqO8on4y2qXud5uCsDj6p7btJhwRDf7OpQzE0eQdx3mCc
kmQtdszC1PsD9YY5cNFcCExuLuYUcCbTwT32Vq4H2pBBPupG3iV+5unKuUhizOOG
B76+n+o7dXs8JFsD5znoeE026o0DU+lbH6843fJ/Ipq897fh3UraliCKrE7pzjzF
Ulr9ofiMmSXCt4/Pmpk0TuVZ1dpWCVmzBzR6OB2Smrgg8LsOxvZz+9kchr1Wgapj
UGRE1yrpjTChck8V+j+vrD/4dgMkoX588/NcS2soavP0TEXWi8+98hhHW55Qdgsn
dQZv0E96v59DosGcNc8Sh18tGpdgyZ29II+fX+1ZHngk9rBU+1H8SMlmt2dk4FLm
X+NbhV8J15Ww2xPEygKSKj5858D3+kZqQznCF21Uihs/6OcYr2FMKaI+3F+c2c1W
xa/qd9nGbnaerNRU/Nv1JZ6eTyp8G6j9AVLFFStiGj+Q5fdTBwNghQvmO0qQQEKi
`protect end_protected
