-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
WY/Jv66A9IG8s74nW9fBdIF7TjmOcYWLVrvF7iPwkP0yZvXO0cevV7FY47tQNycAmEU2H2t1YpKK
t9Ymm8cRsk4fLBwb6NSPjQt/YV+z7el2rmV2mID+INPMvtZzNo5D7F0U1c5FuMMwtJ89t/r0CJKG
YUA9nlJk5+K4EvSaB5eniBh/QCRkwlXEtKV/PX8/jB0b8Fq18j6uutC7vr6lkbU83L6Jq8tMfcYF
8O3CisCfrx3ZvMW/jM8VGTgfYo0exmMDNeEagvmyq/k0x4cMgBLYf36wTyuN5FFXiGu1sxx1loJH
J1BWbIdyzWtWLuYj39IboZGcoEtT2ZvpsitTrA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24944)
`protect data_block
cQbnYyo6bw+uSJX7Tn7kxlboQDjhsjZtpFyZsTsjmg3pJITZy7sajB6wFL9VC/n+ly0DFTZOhSRm
LvBI4gWNnbOUnhql0rJEYl6F861Okw4aq3eBYrgmP+FLwOJOQb5njFMHdnz2HajB8mWY77oH7WC8
J/ZaPq7GSEEeY0VZc+TazzoKEoDJb2OuK55JLqES2eMJFflSw2JJ5mQwkMFCvk9suwbbxDAG9XMf
9+9Wxl8LBEPwJH2VZTbUh8LSKwuEcdMYQCS0xjEsj0vrXaHYDy9GnAaU25f5C6PeG6vYxqXfca0S
bklOe6h49X2xdc+5bP97+IKU/U0nGSnG4ZQdB+imNUewaLAIiBQcRnDgvMRoY/ZNodznO0hEEANu
oYZ2cF6vkU4jv7EA+1QShE3gDUaE3/WUjIU67SFMzJIh0oOD+Vf5+WiC8w4xmYXH4R6FVeabglDF
sJeJQYz5JtAmQMJt9VqmBC61SNnw7N4W0Sow2JBxL0vRcRuSjGZa4QSBqwZNNfCPSHXNeZzvVAEz
yeWd+KAHHXM+VpPDvr6Pm6XuVpqrQqfik9te+vROzBvZW1z0pTi+Rqeu/dya6Ug7rWccHbGsEuwV
pRlYH1piS/dHpR7p0yaOFyhalYAOC76jWVVIzFtmOptQsxmNe0ywhn2bH6Xm3eWHeEtNd2RmAM7B
CFqi6kM9pygUVQ3a5UljH5aPlV8+hgkNQqN49kF8RhNhv1VdY0AsAI8wY3f158QuX6jkqp21SOay
q3JYYlJ4iHolyJmohSDlg+bRZcE0cCOcVWjSbs7s8LO7Xhz6zpfzss0jkQ4OjuG53O90FYXoQabj
3E2Tff1JvA8zPcT/JveF6XNHUj/IhVkkl6N/7ZeZJtmlJtfQEx8phLscNRBQOisDmKxm5ft8SxCR
KkmO0fecvqq7brZbIi8+nsR50euF91LBcgMbV5oi1K0dQzKZ2o+NGeINmW0WgxMwH7dBhSwPPz0p
eG3gLDtSH8g59O+JjFmSvEkHVmIkjDAhZc242tCl0VrDGtfwMPHiox8zStPyb43bxvnuBKH0pf8X
cx+GAfwdo+dLkjISS2JXR53mhfynXHm2LI/lCYRttSHTbADh9iozNodr3jHHU7zvts9oKaChy83U
S0zxEprPtveZA5Oe7PgIlmlqmvjUkrDVpSwRqrF6GvK7OgHjng1/BD/HFGdd7a2pnfrq7FWk/ysC
uRWK14S2CHjBG64rTZhIRYCIwMh0qZDTQZxHKd6fTc6R3GsWoQOkjTXLzDwEF9THCRuXxlaK2zQZ
THeBpMC5GOQgQFMbPBnqU+zdeX9dk0rDF+DmmH+s9QAVuD04aEtpEh1OK6GvvfBfHN6fmvUKvEIV
aA7Af9w+9oAwai7+8ovTFLrNhIUosuu6OpIkGnbmsKscFcz2GcC6e2bniwt+6hG6UkuogAw9Dbm0
VcR+VMpA+7IFtYUaNKBfbnl91MxUqEXPuA4VdWwdzTULfyREjMeYrDM498ft/92pNYbt6FkiMsbr
I01gBejEUdUJgX2w7RWqdfX3EM0JrBxdMIzAtVsLMBb7T6l78qxCk1/h5K/ZxRtV5FBDX/i6WD15
qhkUawR2J8FH219q4gU+fv5V4hdCoJT0KjBB16KThfj71hnNdkA0uNK1d48WVPinfSVEQdYzGYQp
ZYYqR+ESX8FSjjvpCTENHhSHSrwLc4dw3HiNkdGnXemISGKj/j3xsYNq5wBbJnw91RMgHqgzR1U5
k0UVC/c53KYBbM1VUKeIc8WlHF+w1KjZHtUSw0sYfbChL0B1lGKi6A2gkOY7syYBdK57+KbGdGE7
fPutCuUoBN6kzCJY3hnBMXA0mLjyDltbyUs+JpgNoFpQKcBy7Cd0eSFH7qKiF6OK9lpe7DG6qUcG
COU95SNCPQAOrPnsSqGVEAEG21WMx22GG//SB1syig950s5EoS5SMYjUqFBxUikxZrXQL+tFzRhn
DAxtxgQAn7POsXXpprQjelHkUxxE4Y7jnak2RyYoJoAqPjVg7nYwRDVZ+1UgFIgWCe+4wKmiafUe
PtKN6aZ+npqNzweeD4Onx2CSUaEDq8ar7gY+x/1aFKA8E73YWpAj+k3Go+6YZTl08MbMckXO1HlU
Gs9IBSUjJ5ek34Qhc5DXkW15J6YwtAO6ICbBxvBiEDMOYXL3XqWvHB/NAlhYddqeRL3VUgioCdhs
3Rmt1drMXSeD/DWpND0rUS4dsXzaoWVrSXmivFqm84CS/8TZrcBq3Mib4x3B0dx8jMEAfCViD7DJ
QQF083bHfO2tJQurOloCDtHEZL0WxwGqxf8vc3sy6ALmMxvluJzUbQcl8txV+xzROWnVKfgBIAEC
WEip5PleIa3RWPvRIFHqMVzR8H7zM87J/OopqEyd73PJJ0fHLFHDeV5XJ5qR0nhpvSA4QSoRsDOU
LhQAnSV7GONNU5kXoAFK+6QjcgfVYUckYmSE/9suLegFzOKvHhII0JWq5NilZb+4vYHRlNWPDHNy
UoNbt4aoBz3/ENjZmTpLwO7yTFxg+yEMvy/d6aUSMNPiCDDt7iFaUmQst0ukJyl72+437Ssm6tgr
v7PnBIQMMuArpKUR7lc2Aw4gjwY0ZmH3ELQj1Wqu/0Oa+jtaTIh7E6DgCaUJgzO9/YFoay/88fwN
ReEBCWBv+HNtdG6BVXz/juTzJlMsJM1w14i5dI3aOl+zEhyzmHPy9UelCu4xRaMJZkG9Bd3BSXBd
ZYpM89wdJVCTr6GH2IN/C0mE5UI6tPlELeEfVjrLJixYIwvAjw33FzKJrxnLW11FdZgCogTpkTsv
GuNItzwJQENCEMMDAJkah/h+ubw6tnFfaZHsB/qCCsvuGxdCo8+LRUlY/D59pmqDgMIcdqxpPxon
ouZ99NBU0WwWpZS28ApWKEu6Tem+FFyBmt03VETB0OF3dAtGTJiyIeXHcUrWamRNrd17dog5+5sL
0+LXo7KTATWt802BkFHNNBsc+NgiwNhulo2ezTsnTRex3BW2C6DKGoHWbQ+fd6/G8KA/h+KZi4d4
jSCnf5HuqUHr+a/Z/0+MUkab9I3f8PlmshWEnH5r8n7if4m1APHMcenwkn59ZxHjaP8amnszmTDA
Jb94M2WnUStwMxXP45s9OwWLI0iDg1AM/MtfChm3XMDg7PW9F8fCU8BEbr/8+RJSVygrvfH+mrsy
P9dMe4YJ5EMSBT0sZK2FOCa7atUgVWeqORop7Fictyh/w7QYvS9EfgzU3EHEqxVjF5dik+yTOwJJ
E6UUEXykSvR+wztxyPu1HaG225fLnqr5QkNfpNSPrMGevVZKL2OR2AKfRsJzDxAwpVbjoyarYvU7
pPef0w4Gg389UKXJEI60aEmh1hsZBBEUcqjksCcMG5cqqrpBEThpm4Q+q9OGD5VMhPJOOL/y0J7w
guCyzrHYVTxxR9YMBx/KP68Zr96Qw7vWF3jIY2aFxsUooBUMzmQjyFnwojC+aVnD154QhFZLij3N
532FnQ++nNm+8HHoWvSP0iIdE5tGDM8XvHG1akAgpO2rNcs6AtoegZc2TjLDbP4q3mw/fQ+xYngx
BekjjNjND7v7i+O17WhUbptTpL5bIBHTcZOiJK32woBWl9wBo5SP/+z1cTXiE42vrQ3En+amD5dm
EUZMl4a/LITX9iI3DLYaG4vE54rXqqUuETAG0qh1xO/HY13Mgs3KsnES8GhtR5Qqxpk8RfljMpy2
BltgA2BUYV9c1X/SrUd3Q3Iu8gG7r3ZFbU663mLwFUJ5MBQpr1zOoxe5+i/KrrHa0WHufesTKPss
FvFNtY66grSb8TBDUezYD3tUV8jurpx1+aR+mHpnJZALe8PkNW+I+Wlj1ZpGbF0WMCDdH/l0uIqE
GaTZyGjPhm7YOrznPkQeVTk2ILOqwXhRZbabOY3V0UB1A/omUQSpHjS1oW7Ls5hcPQXLWd/SSErI
OEDJiuHOYpMqkLdTzE+t1vMH8efnSCp2/bRLy/MJ1opW5kRVRXcPQIg52Qd9L7TeKVVt8ympqHTz
ajo2xQjApi5xU+9xVimDe7x8onIgI0aj48CB7SfB9W59dW0Ei7XV7TY2gCm65YZez1ZTSXstdsOe
ZZq2eHXZHwLtk0igDkOBe1uVAFQyXGtSmxd3/Ip9xaTt6AqS4cVTnLdzZhZ54A8+CwrxtAyO+aCI
CaKJXhg8qKo9zp48TirXENHv/BiC5Rby1Pb6RnWbTmC2E2n1pXlYLgHXneg/y3MKAA+NH1GiS9/l
ofHsU70nNyNmhre7U0XHTePUlW61Tq0f+xskHhwit1POSzRMOVACb5PS2wRYedGkQWZrBIv4BY3M
8eCoonCxAdsRpx8+raITzJS7AIqlul5ZSybDidyQiGxRFRMprMjzZ6tFmYl2M4Wnl8DMQCOlW0Di
AiP6XRtAV9NfcRA0lC2bxhphlt2sKddFSSbWmtmDwor0se9g3AW8Z4HPJ6rXxpj14k77Kfwx6451
mFrKUJS3LvPsS7TNHdkLnHOZf1GtTNVbC5+fO6SWckfiMbIaIhUEqDxotxCvddPLmsLQ/7ufDVBW
RgVZMrtXNVM7w76K0vI0jyqnrJXPdnV0mQpnv6Hl5PpJFdgZv3wPJnVowbgx2NibA3lGM+e+klzC
JDTC+de+LN+zs0OnyVEkCoBpBavuwUEfGzJhO9gDDLJukElBni8+4OPh6utoqAlpvBIHWbF8WILm
4f5pxli54+HpgtpU083ppuZa5yuCbHxMoxROtgYjuJfm3qJhk1H4rF3zJWB+4aD8XY55XHtqoOQJ
WwREaPJns8OAEMg8OY4wxcwNTlDtFfG9eg7I0DalJ/HlkADSShDTJNtCNm+5RbZO3lHFoOk7vsCf
wm4D6OSyeHXy2oRT60sCz43Yt/NB/AqK6C76+ZT9Ha/c7FuRJ4uPzTbA3cRvNhuGEDLneMc6C1Cb
U7kBxZELG4aedjbZPv3nyaUeQWEdPiDJ4ArTx3h9K0grlzBlzElyS5xDVzc8qAmzaOnS5VzmnUcE
l5BhhRWx+Bi0zGG77HZgYEIg9ADnQUe8+F7ppkD3W/mOKnZtiGCvYpERISNFtJmEhxvbSi8n3P5p
nWMcMeriphvuCDBf4u4QULOhqUk4JC7/EUwCTvhT4XULK0cvx/1164FOZwyvEBr2SXWobT+RG0/j
ZKA9U3kp5bzJ5aDFXqNZKCSoNTwjLcVukYXm/O51Fc/op8JDnyB2Bmu8AVvood1wPVrE8HdLIPS/
ZkvEg5bE/X1gXhu6iQoISK1cmOAf09p0Lu5OOyml9335PRJZHYi2JXmYK13LNsOzcZjYco7ffYLl
887GMLvEDLa1vRKdGO2NVjDoFWQd+qazpRVG6EnuqbzcpbL0x4AFqxAGF3uFyFy00r6AGo4K1MZa
K57WmBhEfq1IoyXNAue+e28g4KUhqL3yJXimmfx8yXFtJvjBmFTzuj3z99RGi0ritS/a4P8Mj8vn
RHyRAeMNoPMhEdIstifn3aoBPamGkwc/4Og7X5qIkPkVadiJWg3gxonkw3+/ha0icYILOCXW9e30
f+eIlC4EIUPbe9VdpWQfwyNmx+q3aJOJf4m5J3Aky+fP9FHAEkdxkoCc0UkpBE9Yp0Z7jlNy12bE
LhCfeBQQs0GY2PTh9gSy9ANWKkCkXaeivwwfopNQdPTHgk70b4euotlDUr3mMTfA04RzBTu1B9jT
GbSh16ISmyc/2UFtUpxCraBsvyJB4nBJTwrNCRczWS56Hj5/MjB8s/z1M7yjUoZEelDjg6Yj1dPi
SRgbR5OjpWwOe6xhXklAn30oHEZdhp7Rk0LdUfr58hFSfZdYj5Qu3HZF8xWh4pJLJqA6x1YRGVn1
/YXAtqCZHmT/njibHO/ABLyP+yTF5OMu7Y33NxzddMHHLokl8gYVkQu1DQAKMsWQEpniMEFfsoRh
Cxv7dh2iAwfn9GzLMpP0d/fDYtUXP0YR2WJMbYtAVK+yDJWUpp0/d1sK6WblD3zSXPNQRSr8pnPU
ZsVp1SCBLm3zyT1d27460WJtYghh/wscB1OUfO4osNDEvGJolDk8FSmfz+pydtDqixpZrtoqkpRQ
Holu2YV+WAaPQmC6f4u1RJCTluWtaE+tbR2l5VQL0v/GaRX6POumvGdgrKcc+McKsRP9JVzfh/JF
JHbLr6NrZ1CwOjmxWjBw38mzo16WBpQZmCfZFE2JVXbHKTDW8sFDWXkpx7qjJcGGNRvDb7BxrUWY
vx8FJOuEijPheOGmABw6K6jRohiD0AG2amokstm7LOe+uwYsx89dCAj/aeDm2om/6mDewVbNbdTu
DlgyLLVq9kEeO9uBz0zlaaCMHLB0ef68BzECwUO8zE+WnsSX7LrYv1BjQOmahGf3qfAQFTW8iA1o
C1QiCYmdC7ifJUee7ZpsBt5By4OS/7LG3tDH0iuGyrzvIReKgQCuIj4U5VP9zW8ZyH3FibhrxT8F
sR3bnd7JhBgVgHkoTqCTDs9RBS41/PY5fnUCvN4qLj79oILQCCnw62HVXcw+gbEzsuZ7Bf2x79BG
0BU1LmQdA42c/pfreQUkPEYLiBZHzpDmlbjP20zjnywraUJYcSvG8LyXas0W//clzeDV1+x2m26Z
bZfAHpGZOliQPRL1mJH5kMg3qBndLJPaT5WCeHV/75Z4wh6jUKynuGihVrBb8eMO3bBD2w0Co1tg
KA09yAMkU01tpBlSsAo0JsIsavcC+/c37cQ/8h5l6lNpgQyzXbmTmobisLnL3PbTn7BHWsrDXajL
ND9LgYGU2s3HOYfmCOMHf0Yc5PJ2gprGS9NN+Ar2ooSMsGoD2hKkIa222AyK/erSCSZHcw3WUJoo
OOEVKelXRoppKIy+BqsXo3kCSEDJqFaohUAftAMggzjwkKFZGwjb2PrtsAywKPmom7MSnVxATu6Q
UCgiaEDCUBxhncsdgj7p9aGmFGm1aTvzoy99e+NFuTZfxhR+Uf3ZOvX2NQzGJ1ajM/wx53EU5B9H
j29Tw31z0htVtuuC77mhWtTFw9ZQTnNecxQ4ztldoD9clbN91wQbWdRKy1qzTjTQka0LMjfTHOvC
POLfzkNGCudYjTzJ39wVEW31OiP4aNJyGMjuYd3Ql9f/EQOVN5M7Qxk9Ufl6S8WSFHRDVjMRHPGH
IsKr73J7+QNZ3gzG9G5MLHJPyPyFxg7vQeMYNNApuH0/GPEZpiT9PMwAZr+2CuSGUV88++iQbyzi
/vVcGK7GhhFJvPvU/0W6kb8WFkFPTIrmmhmJwBU/DsYbjX/sztvXk0nDsz60Xq/8/d3T9EIUb0Pa
zVU+55QqJbMK1U96curX3iWjkUGEW3lZm6pRTh0Ql/1wdFRGexysoJpugYz/Qg4ULTBS8z2X2kDo
KoUMZUYuhv0HM1JcQPJypIlK8p/NKwQJZXLOTE9lADBTkAM7g345KDvyD83Ox7b/R5WxB2juyPop
f+g6WFVGqPcUpO86EWNroY2icLqASEM5Tw34NXFYJh6P7WBKJpsXz8uLlbABHna3ltc5tA0NOxV/
bRbZ6VlfyW4c8d5huFOvU9PVe0xjwimIz3O+J47oF3WQqXsi9UU+MSkCFVGN9aQmEyhYb2xyuUqt
y798xixPRuab0hUwJK0IvnZyw+uePxs7iT3DmhJlIy/m8pCA40Po7MY64GF6iis+Gn90f9D5DmrL
Q8/ongj+50Bk5+x83eNB6bi4Qq5lv2EYnkMtibDl/n0FdHHp0TuUhmnhnyfFalvfisT0AmD1u635
2TyBMsmGV0eskqnb4FFIvD2/AOA56/JMfPSvGltFgg0CaV8LATOQbiwQDlrcC9WooK18z5NbVgII
RYvwyfdMVWzBw/KiI+quSA2npP7/n5ADDK8wJUk+q1u61vbPS1VkUNL5P/jvUIasGx5xh/1htsyS
L5pcTE/dmu7hUQjrSs2+ebEwq/yOgDYP27SbK1xUSDUxqo1hTvCE9HzAxdje8eiCqCsb9tI3kZJd
4EnFIhRfFY/JsEVkzmmpJs7aWyJnwGo/aZuAX7uDNVjzT36GxuXxQZPEV3psmu8zuGABfFrDxL02
z4Oj9wMr0q0cxZfuRRt/UD3nSWPjtf7ofUoRJsWL7kl+gj2CHEjJrzV+7AjK7Yv8Q5Kxtw7c07hu
LXj6QdDuzmrZ485X+zdK0Z3bvwMylSy4FjUW698Ak2K5AHDV7AyoEoaaA4Bosqqj+tM12dMMM9DX
1NfEXGQHdfSZ+6wVlYk7vwsDPP2v44gYXU7NlVu9V+az9fXZYJZpeCKrIUzmbbO0W7HfrPOIGh2u
cSBFH/lEL3lgRp+sqejxMYsAAjhDTY7ob2L6aKLkT1TRSut8b+TLx3wpo96ekNIrcBFoMBfi8Lib
ahSa+yv4awg5d5rTmmn8bHjwacAjn5vMzHTfchgNKyYYtbMNv5xRwAoHe/lVR1PGicXVKYfr3auM
b+7mMQezsePSLmZlJO6ik82RFzhh5uD+lwBWubPzfyvaqFL/r5mldVGno6uvgTv9I4oB8XVToR1k
7qVYxDgZLOQFJ4msLe39IyopqaFmOx++zUn0T8+UYqiuFZ+4dJAaGGG0WgNIgVF5kueWhbBDa+jg
prOQPvZTJosDRdUbpX9M7JxcSD7oETPnoDucNMm04UuscqN1IQONF8xyMZndLfGWQyzQIqW71ZX1
8jUpTqL2REzkPm3HDmj7GhefwuGqFMJXJrpVyiZ4eDgvjdnifqP69bWwjEHAEc1AZGAKEb66774L
QKzpllNuF/OqMeI9XRg6L88kQQsVw9gVhd+eQHM+2VEOppHjcFBbbnXhi6omNr+cBNhJLkKt4BcY
P/tn1sS/2dKofwGZxwWD1v5JhPfVK/7sV+JNclsNKr9RowXZwpfv0F6VV6cALzrr56l46KiE+26c
HoLZ6KfVkV6tx3IR5iGpqUi7laahst6G55zs2ToEQiMjnHNC5JG1TiR2eRuHB/22sVW0HPs2oPh9
qc8vZMOZQWI7uwIJLXtEOLAfbUO6QPqsFhmJBNNCaJXsi2LluuCUXWrdFGe+Nhto5mnmxNZfSdEn
Tx05GxlZ+7Le3keP5pP+4hyLPXhHoUzuBwDZYhX3lBxVLuD0ojykgv8hilDZKl/Q9zqGf7DognXH
fKYTcFqlG4Akt8YlPiolEKefWN3MoTyGsGbwaGL/7OGi/M0OeUI/6C80bEorb5tUN4y4xDIvHde7
PC8McknGN/D9qR8FXlIemjpbW82lj7r0QgEWZbEeK/JgtD+MWLAKPDlRGVcKV8ttvUt+ZCIHlWzB
Swx83pD/0ghXeC5vVA6A7DPabzYzwLb1YTTvJVdme17IzTm8xAqRkckswEMKTTtneH7Y6UOBM6sM
3RSJdSlAdqJ8PO73pqbk4L82fD8UtKb5wYzUxIS8oFn63lAOp5Uc646DOuP7CjRZkIhrjeLQPFwO
f/z7yMEtaud5U7bqtnEz3iaolXvlZcFbSyAnv1seo3u47FY78zeWmPrcQFUY+R2LGOvwiN7fpcwT
olJeaatbr0IIT51d+3YPqtzEu8AbJYlPHv3da/o+06tq4Z+TD1i58Aj6LJnV7wY3SxQdHC1/VWYh
KEyUrcJHeBwh0xSpxBwwkjO8JvTyWoqaT0bjLlaMJ3DbO5PI/zmtNVVjvH8BSkM6ExnxuMAGs1m3
hEicYk26vxVkHavYZD/+ID4dwVeVHZmnVrDejRW4ny/K3jSl2dDj9xFC1vyw5PMdlzdZYFM96hQw
M96FaNkV7Ys7WORKp0idhkEVyaizfhK5Ptp67HyuLTRnudUB5Gvu7bcwPOYiP0wkzn9rvPO9CDA8
H6fzVTGWF21OTeOTD3A9CmSrH83Ll8yaiUifhdtNJ2IUZKr3h8VICddmm9znkDzWrj1MxIA+jy/Q
Sgsr7pgQ8RkPZGMWO82ALR0EC4PztDf1fnvQ/HrW2T8MEV719TAG1kpon3ep7fVCfaM/a+wwgqTr
80G9+ufCXsuL9yWdpG9/5zE+PCubN7bh1VvWqHCUswZtcVrwS+ArBNvwaoIY+ybIhm6NOwby6fBn
SvkIGYdQ4eYf6buLZ76UZm2eZo1otbIWaeFHqbBMH2o3PSOXd+ee9tnd+rk17+RI+EzQAPO+Aka+
UIqk2Q5TckB0TzdIOR88pMS5SK6nvQsUZ22Y2QSihllEwKCb9YsTsnp7XvsNC7gc9sdOJstgQBNH
msAib7fXDQZlNRzFCOV8XJ7VWY9hIsPbmVBgeqHbmua2lC2ksep0fvbGp6UfJJcHFFMPUE4dZVo/
5EK1a8B8MZtOf8cLFgOIjR13dhVGoZBvnkRWQuXmrCRnjeFgj9vKLZMxnwvBCPcipsaPnDG3ZIda
9k1Pgpw956Szjke4tpckkH9KU3kRHLUT0Dc0pNeUoP5hGXJQI1y4DfyHtmz0N/Y0inf2Nol835cV
K9Fq3x5EO0OADexCrLalxtWzZ7wvKti2bCXQ14QeFfb0YCsN6tdGETp8cFv8qAbisYwTRKnVqclc
44Om9Q6sg5Nq/nciQBZkLP6Gif6aKQ+sqcp4Qmsb+3ob3LKEqTdhAaZJ8qJlxtA6gXeZy6LGTNJJ
jBALEOuEi9S+Jf14FTuRkxgdhM6tqn7qDh8FWFjlcATQrBscabCG6C4KRzl8dKy7trdyFlXJi1Y7
rxYOMrjANXj8L9oM77CSIlpmyky3jZGP/acSgFyVUbJXDCQJ4rol3OozF5fvO1x1pV9eOavj0+Da
4vx0ebvIi0P+PcggWbOnS7pfXJbCrSrxf3iXKhNEXUAUWz+QDZta1KZL+VMpdUJvSUYsPOxywBMu
sGxdC1cx7B+0ZoMbKQSrVna9fQFfvcVISWo2GNTgbwrsnV0ICvwEuI6kDVTwMzKeDHIPhQfZafW/
rIh+qzfwv8TdDZLH7hiz/vzHXIu/7k71bL4LEh6NJy2Yv1Br/IoDvy1xeh/IGKAB2YaZ1vVNHnpd
TJ8zb9ZY7FDO6gRJCVTGzEhLOj6bRm8uoeaSfZYOE2A1bBCFm0juX3UqJ3IcIew6PQf2f89K6QIF
G40hjq26fKbKAtHqwlXfzRNui9i1K/thD0tg2kLXGLz/ScEEOWmmbDIQ9pViYrW5y32cF4dIFeBQ
SphTF9LXMxCTUaK3Lup7AlPSHqc4pMum3L6Hw0Dhd8uAA+RFBAyXzSSfKeRiYFD9RZWEo5koI1U+
QSIPiD4QNFyVBoGe9nOnv2zfkwDXHFCMoklSqQqYqb3hH8QtQYJJ1edCRgXod3aDn88DCnLe2sYj
9+fTUfGCLZJ5DyPw1wL/xvl9M5vEmlIBQEBJS0JUZv123WXYbWKmDakDLyb2Q4E491q7L2Zlyl6g
qDXO9sppwmGmXi6KxlSdofDc4wnwnezWXnNGOtC6BJnghDw1k8FfVBXxqNGMIlXyrN7J5akuToL2
ZbPEeLw1m4tnY0k5x+ZT5s7SNRziaiS0J3GT4MsmWxq37w7JtrlSMuok0BLQsrinVIxDJjkObp18
Pf/Zb9HvXO8AV27SLlzt7NTTwX71eKhVi9NhgbOry01ozdIzYm1uIvoSxi1qNemU+uItxRPuu5yD
ur2ZcE1RfKMCzdemCLwrVJiF/Ta0fCcSCUjpsnXOqNCpJZk7l+dVzz6fErQNroqjFyPEBt3x4rok
QOAtcdvwWLkttgFS+rbGO56o2H2Br0AuziSUHW4iEpId/lsgicjhdMpDow/89NIsLzv7le5jYkvY
+2R0gKkuF1yNhbtg3/xmP7BAbuJnL0w1C7L5d48vSigYMxZZgOAT2GgD7Vu/wOqM4ue0mfKu9IWU
/7/aN8Dao3tG68p1YftkF5hJihtX/vP6x8uMEhGLFOGmn5LDOHpYR8vBW7blP8SBG2fwEHGp6p++
CMC/g2G3/NsJKgh8owfDk1rcezuYWAlq/J+clzAg4FRezBUk1nQljipr+KO2cDCM8dGzyx1VFRRw
NiZLmiOfxBzMg35sVWu90jC6C051oLQhpRfmHDKRJoSlpwm+gHCjiLxQMnSsr+ovDiTGyKo+5vz5
8HdYmdJQXQPOjhJYlemcCyyOjc8jDsbyFlw4VGTXnoO19vdsuoWavX3HO83oTigh7SmHM9Ini+RB
YJyL04fn/GL6JPMAE732QIfm8BxXDQbxyA5cGMNbrEGabtkkSwWRs+nN+vGvw9K4tUwYdzILgVlF
NDRb8zFiuhWewiZAwdy984BYRxYQlAaixL8cM54bCWiQCPrKQ/Yb2UFurevyQ+Xh+YSEq5GfgQ/S
zFArXXR33xCyOnTrDzHg5uZ5FZfosOBvkJryAy3W/cH0qYqWfGDnCwO6BkkbY2pCs+aNvNatJLXZ
lvPISiqd2fMtdoJbq8qy1EuPGc+bEAc/hGpkFjgpzmYEp0NAukZxUTWqzs5n3GBp2cZJ3mjzHu0H
bXiTsclrTHYPLPKK/9TO/dKLPYA1npxE1DVAtc2opLMuXBYBzam9ogMkrXg2grLMNYdpxK2sP8nD
moRjIb8+XW0UkP1CH6TxcnYU9fmK1IfbZwdERV9I5J+8yYefAjihXhV5X1p6/8KOoI3FKhrVnIo5
FcH3u8oVwNqIN7hkNzMf3j/Pkq98mecwaUfuee9Fs6b6KQYfGRnEUcFBkjQKCI+bilVGRmlUDSyx
5y6dnKNVu/EE16TaSRVOE1AL5YYsLHjMnLjzrfbrYio1mTutrWrXwuh+A6ovpMITIAXS7hGPA+ju
J75sZMbjBmF4gr4oiaB1o0Dn3/C1AyhR+PegIuQUTxRoJbfotn/nEnzK+sNQ3U58ttNS4hRUZjlu
lbmF9GV0763LGJl29FQVM0Bgvd+zJCZtisEdGLHRCWmCrXADTELtF4crQOuwK2eBEzMRvFPRV+9j
RvC/5hpJSrnEEDlR3trLQrvpA0L6t6WNiohduAKSSaxFt85YoFjFL0ktSYT2J/eGFE4E4shB+9wY
pJSUVYsGv33HHrqv2F2p2c2n7Yyrn0nXcfnGbS7gqoYWwl+NHcilNU9fV5KSCHgNXhJp9fw1zH8c
abYR667nEzo6dICV5tEF9ey/CNDjWh8MzPdD4h2hq2izbHPUa/XpEK2fWG9SBYkfvgau40jzsbBF
iiSzep+sYKZLTA/VroG6SQBc8dFHmLnejc+5VS3npI7u9uOxCtuHU257+3orLFi5CjrCzJIc7YTc
IdcitzCspGZrHCY+xCLsmB3EPLYgQLh3/CFWgXf3iAvFOqczl45meGkwrCkSk5BxDrQiDifl3hbD
ucNq5W615qdDu87aXnKA9yDWUE5hqX9pkpxtI5pDMJI8+QYjvcV5B5fiYw6bE55DTuC2fEoqOLmv
uwMigst3Byqgfd3IU5Z/rDoGtieQFb926nW0jbmg0K4R6CnSU5lcgcz8urMLuGjwlL8PgAkZynYv
uHZ87fMB71oEjG9MyKJHXvuqKsO5YGkzmzHRbI+cGKZfJhi0Dqpror1LDDjYRr2ElbDgPL0Q4VQ/
zl5C9+YfFerD+ZoVyrzLhCWSMuvUzud3d9mkb7txI85KXDWY1lSwCc9xJoDiJQeiNJxcUTEE7Nse
+TRGEMFW8utzqE17/Bf4RWr9WZMzVs1G6WU7eQPVvIQt85hOm2Zf28R4lbSyKx7o3QxveCIH3vsJ
rbUewHYF5Bgyd9bhLEja4VN5rr2rnvVSUZa2SznWtpvcp+AF2OyANF9vFaPHK03gsfEmafZOp4zS
yc5J/vaAwoMnUBvOYtrpK0sSzzR1QIEAK1jfh2gwtAfW+xThLCbKCVej74fUNorlKEuFtnPdz9xT
ZwcRU9EhHW1mOe2KBGxwrT5DwYfL8CADzYeYrFCPgOynzz/tiDb8/X+vbRSd4Msz7bco4JPFAxPy
jzU4DZgFj3ywnNJ0VA+O+f9P840QW0i9h7v1E9Mnv8fBxC+Bun/QNREzxRPXNz3cgM8+pX8Y/Ktb
uqwFh+gebEyjZi+Jm2V2X2ESUQ506z0PS25RuvOTJRAdScnJNMri4x5/kJQzxInreepfo6TXqAGz
rJNqVm67wKT44ZD2VwKK80ABXjaREPs21TQuZ49/69ioJZpOO7HFwXMo4VgsLXt3nVCoWnsCvV50
isJCFtcnaLR6Lb+qkkPj/X7gQ4oLyNuoIJTxhq/cQad2OHOjRX2UhdRslFNS4XMscOga/YSdK0ym
LWZ9Q5IohG2QaTHT6eYqMvPY5zPzHVQAlIQPql5c8xa2StuLH67RZKX0FCKkgqQclixYtaDYGmOi
lz8NRj2b9zSztf1SD6oNlOMNrWjPs5XnWGeaUF+7fjs465OFy1nqqPAs5uUEVeq2rDm81Czz9vVj
lsyH0FYZCmRHBWH+cPV8WjAx2Rm1zUeN2peky+awSivi6I8JbPglrLsao+NaFeep39mDngVq84Kk
0WrRpyxt46T+0ig/szi838mYoMPMHDOiW9XuUdz1IFnPU2u8E2mM8uLqVM3UNTogC/quRCVTxUpK
XxhqgaQJ1OXhC3U/Vz8v68ZqxVt1kjZT2y9VmKS+8H5EvwNrIBk3wZhTfcqHfGmNfITi14m75EZw
a8ESc8LXGxMqTCBz85ivC3LS0XD2kouAPHfsRbPqsKAEAhYCk1C4f38gE85J7cNIt02o78e9Dt54
rNgUW7rWWc16fpLcrj4Noncp+MV801CPgjC71pafomo4smrySzgs53cfcFb4HzviSmwKNLRayLrd
wklLj5MGxXeP2sNr7T1S5YKNoL4QB51exL/GDNr2U2GplHcz3udwiX+OS9WJkRxdOsxfBaNKkW1i
8MQUywJyAOiCEofamChGTXApHFuE5NYNFum5jVL6p4pHXkbtCGA3z1X7gd0X27QQWsPawE95dPoU
yee9hVbHBeAiUUzfieLKi788rWyZuYC8Kg9qjz1Ij8DHVvfb7M3X6MSXQsGPV1287WK+ViCYN/jy
YCtrE37kFJeEkS5MwKOUqRm/MqhqfjeHN8rZrD1Tp4j1xqSQXFpOsIUkCJJjTnlgB5WW+nq+ibRq
xNcex8WUCCKhfYAVhWL9rwWMGbVkF6dVhWJ0sxlQGv6vl52f9sl23nOcW3znZvS+CZUehs+2wBlK
OWxu6uIDmzv25GBbthj3x2BJjbHdJjbUmRB4hqZZ6zcVIc+qxzj2uivQFytU161A+pCu9CIsrqso
BkIagoioiy72/XFPylKhcFm4O/T38ZZmtPFfFQQ4qlKEZo4XGRpMiKm8XUVoOFpsVsAe4/tgaQ1j
oPTBon2SAx4CwrNH75Hc7+EpeKrWtniocvqdaGL2yMk1HV1JSiVr+/inPRLdNUTOuJHasx7DNb80
SV+l9m+4BhsTdBHKY7fzlSWsS68qmjVIyv7Jy+09JXOOVdPjJA4nu7KznPllqkZLskl9AyPc5TVb
bzFw0D2DHBvPcGY1PozAij7siuL+SIISosBf9fBFVfzxw52+BFb8FG/ITGP97APoEFNJb1oS1jw2
lUxLo52dsCTevP0NIglagRvbianjSG3wUDrQT0bgxSiH3zfePGKS6knAu8qH8dxuT8MQca34IRSR
l8Gp91MIh0A4d+RU6GiZCa6KhKxZmnwE3vwQgooDFsH/fzVXv1rsmpzV5fkW5etoSw5Y8M/oEuB1
0pEa1k31D+VunR3SO/vakLLezdEwBAlN4e3PSplOFWiNysIcbdB6RSB73Qfh1oUFxe8eHHMCTIqe
3fFdiSc6WkoPyxJ0l1VNn193EgBMSCE/GhYIAXUMMPYA77XZySV8hWpZnfIogVnO4VRJQOdJw2Zy
LUsp8Y3nzJ58lsYFHP8QGnD2+1JI7509ob6mShDQiUxAkJeEldbNNq9PC30KRjfa54i1bn858Gqf
vx/gAbifLLa/51WWH9J0TYh/IIumBGalXqJI2pI+sXFgq8IlYg5qqbMA93pcdA1+iVmzkrLMFPza
Fbp/zn7hUQ+t5qoRlWQF/2di3D1rlKgzZn2MnQUUH7ZKL30YtH083fglztULmZKOhAO0kFCeW/mK
7c8KPw3kwPSWaAH0vETA8M8Q1vjI+YHG2caz0IG3uBB3GGm8jX7wJda/VOjn2klbQi4dVmWwiGYt
bJnkLCNPJtGRNwzGODrYCyhEzMSk/EFP3yovl9ife3lo5NkK46YfTjlspJAECgGzHBdP3tY+hD0V
zMs4uK/NK04IuO+Uoei7U41dgMtKEpydEbYJ5RKT57Px70Rj4cKXdo4qeJsR89DLmvi7EMHO0TeH
OEyYwKrQkTMWSQpqzQhOJ89R6I+JE+B2vy1SeCq2OXqY0Nf/uznkPgGrBNdd82s8GUnRgkGLav7w
ZF8kz7u+lg759OrpptHMfRO3kA/BnsMXw0JayFJX7Y4yAB/41Ctoc67/hc19okWXujhzqBaulE2P
kMRKSl0HJA88HjIpfKtSOaFVhRnB43RluJawlK+ewfk2k5ajqv2C4uCewEktD5DWTks7zYJIAeNw
B1h3l2b4LFVvOnzCJjzFXQX9IaV5mzKAGjsNhDhXoUGZLGIN4wbi92gRI3OwHigIrlhN4TfSClHp
7+mQvcJkIQcA7kMF6ZjSHpVamfFX3RWr8nKBDTRgzMSgFcamMMD4GyV9+b5jnQpvoz2FxqAXNtrB
GlkVSTPAEle17S6ITcfJQhd5j/q9D6AWZzpizaImcsALtpFRNbWO1imT4BYVAjnhJFixJbCV2T9+
gbnbGMWB9F4WeH/T8LkpRESzhtGuCfANEvmuJYSUtXPjtwI+D4S3ezo8zAJ56hQtI8qVKJMDRE2e
uSZemvxs+xAhLZVV2LcxFCjApcFI2guOIh2LuokJDe8hbrLpQ63BJIiV6Kn7OIelW2IIcFpLLjND
op4kGEKVuytwdP5XkUTbKx/Sns6xBuVrykvXqNje7kOeIWEwJN1m3qAf+s7NvqOdRJkMJlStFIdr
GYhh9ivOUtiOWFR/3adeqdZE841Ig+1KEpgkj3GW1idr+vlSfqKiwlV/wuZB81oJtJ+FZu5UPzvf
+lHMYMAfwIEk9UsgbJcsRtQahczynuit46s1tT47SVz2KAsQ5pXZuIZ15e4uekGyH6wTBq7hYHr+
vO30jba6hkyxHAdr90cBn5Za3hy6G7chRJovFkuhxrZRlkiAWs0KzWkKuyLBEKod0A9MCcr/hFFc
2webOxmlK0buLUY/zxiuTqgs+QHCq4inr1EuEPCxBN4WW0tS6XwLEFSqq3OUQUcBusxkRSOw5nJW
BOcRVa+Y7dfO7oPZuLuX31lXM1CmOYAFVCxogH8ZgTczXCkc8lzsgyL6p5uru4rV9qBEQKKWB7fL
PAsiEAfmGYhJC6QCgWl7oL6m8GxIkLGCgNOGGEpu7Cv85gVa7fj+miQaFp2jXD3FyQc3wayKrK+G
7aNXAACgB1BZIMKeYDl1ZNF0IICodmPiEuYqC+KRKwXfAJkOGO+fA1j07Lqkegy2aykJORUtOMKi
tZKYxOlqwICi7WI0M79SeDeJ/WfNsNN4dO+sgLbbws3NK6WjpuEDKrYVW7viWz+QerCxGVS+TtGC
XfnZrKMYdfTBx4fTU2IJmJ4jEmoQfEjToQU9LA5QWJL//Sio3wJPm8OI9IuaJ2G2mHtjWYOnjCcf
UWk9r9OUc2zDs/zMgcYmjJ4fbdBhA7vqMv2anzl1nmMYjrlTYLlsrcl1GEb0TQc19UwaFGyRgIUT
MxGcdD/iMosY+VBwYAicHb5kZQW5i+evvcZFWjRxx4Tdg+94w2sCh1oIYLIuMMrEabcEUvBF7HJs
Mg6SMeh22bfjz85OBzLxKGSYc9F2nlLmuGhMGnsiMyqq0AAFO3K+cgHgXX3ke7eMJ9cQ+AieR9iL
t/RID04mtVX25yv8Tz2BKsU1cGUQofdZHTm0c6ZwZkWa+k1zJePs7U50QqP5RKMJvgDFCJZGT3aU
x2SzvU2Lpu6O+SUWKekMKOKgNitHraH2rxIp56eYqIjhoZz1oefE9g4to/iUTeq1iMhIBGx1Pipo
W+tgWt9JcVQd9i4Kcpr1SftyjJwyKL5+xuzOj9712fz/L4SwgHsQ6xWDSL6rteRnBANufmqpvB5o
Pc7sSSg9VuK/8h+deAhd+U6CyeqBD8idho3MeW9PJ/1n6I/weCbABvCA0rTpN+083ZAogE2hZl3p
8xgJ4z8bdqKSGe6J+J65fyCpN82FOD3e94LlBB89MZcHweF8ezrBhWu4qaivakIeHWL1aFSAmCBC
XGSW8Rw++QPNePfCdexSjdoPTvPLgOptsRJVKYrtQQetEYjymNhP1rjL75VUR1u1IjUSo0ZEOTiP
7d+DXkPG9mMTOivj78M5CdNuwLkQc81BgG7H3829uV625SrtlgibbDwEzeW0z+/GEc4S90Fk0u1s
YMgvSosI50KpzcxBafDkpDKGjSdi/31Rb4sO0+2Al3kUZcL/Fcc8/xrZRwlzQAFJge7D1FL2Knzg
FyJPCIVjOPdliBuinUSq7k97DNAkL07NQ/P8K7XVMVF8PR3bdHP0WvcfHcgrMEB/pyL6iGTjykzP
cmvAXZwSSSAK8A79laHAyHmsqvuZgev9y88hJiylo6x7vpuDr6oA8J5rXcNuRGKJfZBR2Fu+i+1w
GVzhJx2UaMjbGsTAz3EtnLRJNqQTzqs/ZU6Bw5zjZDFnd6MJ1r4HnHbPGgseOOEfr3Pc1+d8DRkd
dPvjh8vCnXzIJ7wRuEMosjmjI+1SSmuOTfTp/SBByzx8M6/JPERX7rSL9XIyuJdzdp/pNq7QlswA
2FO7gOWHQRtyGJe48FkybcE4U3MI0oUv4NMr5gV4TFuA/B2i+VRIuMGu3JawbqeuZ4WG3ihr7Dn3
Uc3i4c8C6v2dyQ7pCZ/JqkqemWxEBN3D1+fT9WW+weSJlpMmgvByb/5x/ji1Q5m6hh2q1B3NMnMB
a4k0OtidLP0nbLzRetBSmdWaQpq3zrfd7W2NP83ivRM+ORUhkBUTag2/yNwVuCzYlAoHLHYS43cs
4RPhNZM2eQkSpumlilf44lB9ID4jepGxdov2CDF2xFtY5X3DOSrKFLldT4bp8OKt/Zh3pc/h/Gwu
/poyiqZLt7+CCOpnizfYM/NULP1mRYe+5nhGj6cj2vBgJvoUSEU/Mk82Uh2PofqXUiRCGWs6SGi1
BlGtZUdurmeYvFGgovJlz3Ll/j75Y1LvkGSuyVAvDLI+iHng2aDQ+YJ1kY5waY+VHMIn2ny5+PoP
tQdmLRhidV7Jk6KoQj/SsryKFAlKyGoCF14gsfIQ7pbw3A6ool9RO4mt3A9dE6F2qS4cr8YX4W5b
X1uYVFEw8RBlWrwzANeN3PeYwq/XhClYvKwdjETiheq3SxdzBmXTCCZoRO8nZlktmEjmoU0PGjRV
TJPy/Dp9KsB+61FTBf7b8bY7DBcjI8FPUkjiqV93v0oljdHpu8obnUOPT7nKVhVoshVSFj5i19HB
32KUY2CdK7Smox4eNZF6BYxcqo34aOrKoTKwwCanG2zjGGS2jD2tDDpycXscaDKnnNW7zDvyLyHK
C66Te4RUW9IPjq5pv8DVq4qCwZUte6CHat1N8pSFDKluowhd7A/W17/KXW43zgu7V0xXw5c8xNUb
f1h6euQGwrBXsaqT56Q3BjYyZo49v7m3KLYTVwO1ZuqGf6R/d98xvroJ67T/+UWAY6h/uxokgMrY
RDm9lSjJrDh+ktraPeDNEeNMY7Z8qDMajgJvAxceNfqER/H0I/CQTJ7WaPCRsJEHGn8q1Pegnlv0
ebocabOVdrr9mqNzOqs94hAG5Xr/vqUCeFZyiCEwaGlogKvN5Ubbugv60KsxEPg+IaEQWFwgRrPl
/dzy+HLOUysM0nRGG+sqjvlp8VoI+Cyleh4ekggyWOP71B8SUdUVam4hNByw+avvcjgAgnjFwugv
cFblFVahM4fWMFRQ8Gf3tkdePgON3WJF1KesPJ9dLOrMtv1GM7jNtUrzMxD8L+3ZZX4JqaqZAhr7
Q7SjO4aEIrmi3ODO2DgT1i/3jN1sIl+17F4MMPjgCjFy0UC6gTL56VEnVhW/iDK3L8ZI+ow27Wai
exNtT19T6N7lTcEArH4JoyFu2e8BjZrcoMI5VsuIvO089U1nDJovAB6RwU7yw1/hWJzO/uLFbR0M
t6Rvgjzor03iT23ihZ0O8Det8Ph4GRKk7HYMKf5TSuhw7YL5kZf4xHDpy6e6U+cy2vJrKfOSxxgR
tXjF86mntz+2DGnZJpDKoo9xGP+CwY25N2f7KUyOgRQUjD2HqNVNqEFCwm8BQoXPAHlsurSxFBHn
eAUpoIOjnTo6bLRuA6zav7Z+mjkCQi8GzaP/WC0n4TB6jSRBETQP3gi5FVxL3xTR1RJKsjqzVs82
UskaoPI04cV+P/Tjl1eXxjhIyQvkhgf+55P2Z+nvlvdFGXsIpKR6oh804I1upCdVfB6T1etVdfgm
qIWVHiURQCywllM0dQOTnwzkYlp6hvOC37A8liS1QbiOnXv1c5tDLhRCjBX87ANy+fKF4F94P16w
nmNjRcbYg/d+b8E8kz730HNHG6plNNyR2Lr6hSMezdxKbhdUe2IeEh0VlQz0KVI8eMpFzyLS9G8O
AXSVGW5iG4Dt6hZzKacDiG7ItPfBBELActg5ugc8oBx6fjxa7dQSujeyd1EwAvx+yILExavaRLuC
QhJJ2j2SLcfxNbvwgdhPeIbAnD6LqDToMNaqOLRegYrNyWKeuv/M90IcDZK6/pgVIM5AKuu7lJiQ
FK1NbQXTpOxKJCJ/LvaOFPfCLsPuzDH7liwwt3I3THgxEoeREVv+aS2ET77RkTKSqLgCky05lYeA
IsN7L2njfM9Es86qLAo2TI0/ahv+iAYRiEDA/NvyswRqwO7fAmB0hshTacKualf/mT2VkIV8xhkn
47HQ0qzJOL3tR0G+sBiWh6CJstVUgYSgN++707csCCYxoS4BWieL8bzI4wd7KB48OaBmMFn+W37M
6Y7ARDTwj7FGus9b+r0zbz+jzjjQL1Gcu5itXe9T/xjbKM/o9LTy64ZFEslVPkSCSo5tsqKOFAGA
AE+0JPSv57Wq7pgCQeuPBnjlW6Y7aaJKUaNL33+hKoEs+MOLcG4JXXeV06yjyWeBA9h28I9okj9o
9Yt6tS9Dhq6NzwPtwBLzWQ1ybAhBM39zva7n2/K3PJvuIz+ZU7m7AL+dy7dG860GfHa1d8JFei2A
uAyLypS553cY2Fbp3fxwwGQM34Ivue5fOHOQkSfSOfw+QYYzudNkH+6wtJmuuFPGLvBwxsF6jdbo
D05S7CHOqAQmg8/ewdfFIVTgHmA9fcZEAZubpj2SI58T8g9BQbDDYywzm0+0l6l8KRgz3/B9JIZp
ktf/jxLny0FqF0a7xvwb94eDJe7Pf8jxyubvjxNeOjwee+pW2rbdk3y0UYLdZqqCOInVJpia+bCq
4ZVrUW6DCSYg8WO3WYMEfXAaUiqciuMd1Dp788bOzWiqcFX/Y/DJIVG46MoJvkeeUYmc+rUu4jSN
90SIfj8NOhHILIg16WN5VYb7f74YLvQ4ywea253dHa4CXqZ8M30KUvoIoV+xYKwpoXJdy2d6AvdT
d9RjyN5PD5Z0BHASeSQTFGpt5z0V2bjkeFQrQHLuH2DGHmdmUAD6EiFxXDeGliLNmt7y3RUwHWec
MR+q3K91CDi64wI26aVYeUxSqpWKWsuIYCfYN6VgAXFm6PU/yuS8gpDXpcKHaSmVEnrp5EBr+HQ4
HEOmexX620QGn/gdrYP79ZJzfmvmPxsownx0mgKPDonziRftaaH6LD9CzyK1Kyt7S5OhXjW6wrt7
XxOXXvuLkc5k4XF7HiaD2xj+6aASO4FMsaoiOaaEwXWJp4Z9M5VX/BlyHOIoBqu9tGDDTjH/XDhE
fjIL3SzZKp7YFURRNofY01QuPcntX6kwsOUeNpbCzrK9oZYjNFyCPoEMz/t2nksVQ701JCCFAN1T
XKIrmawna9XH5mC2beMBJc8K6HbAF1S/HTqIeHWLmXmr9O6hVAw0JBYiyEk5il69HaS66AjpAu+M
BV8Z5ylvAjtCZSvHBV+rTMWAG//l0YTXRE0D5cgTmm8rKuQp4zKBbiD+VL+DKi1d8XtrpvmeoBoA
3VX8TukZwUmpr/zvQ1oehaESDQF+GJetjIVai0KPoHFfBSFqUKiegEWeLQ6To/bIRmTYbDYd30EJ
X1lQI1XHgH5YwCfJzr4GzXX+YxIqk6GJWhvhaGsEZ2CWYO08A+HtCTpFlVjqYzyDyVCi1c4GyKTc
Aw7+SFXd9BbuJgKTeEuz1LWXAeOlrCsH9GNDafVsUuWmG6A0VukHcvelbwH3gsT8VMRLcg51E08b
qbIbZaasIMIHPmTtv8P7mGaAE9VRa5uJG2bZH6jSNzzqum6EZS65WjpMZ9sRxR8jTRWM27Luctxk
69KhaWG5mBH3NrdjsqYd+58lj69W1EFyX4qlGxDRttBQt5hojiCPbpsgsRpCWTPTSN9ditOgM1dm
2bxABgfdbDk6aDizcVZw05sdzprWDwL379zVM3cijS20sKlMQlJPTsbZu7qcy3mcT1dxQx2YtpQB
dcTkL6yGVNOpUuw3YovJWixz7bwzCLFO8BAsbgBnDWwXHXStsjulaOGk2DenShHlPed8NIRvIBGF
M3P8HSiFSwHJPZyifU5KLz/2O5vhPDxdoDEjAyKGj0aW+RNE+z4HJUBinY4/gZj1x0zT/+/j7TuU
ADd92pklCU8GyZBUkIPb3olg5kjGEQtSZa71A/D/RCSVvbM17j5uQ9LAsu7ZGKgIogZaN6dW5OaC
GfVeiiJ9uFP7TDRrQzn3Bod/Aml6UAar66tgOajVx8/sLyDa3VbB0TKLNo1PsCvkmRYXC5r7O+Qa
gBSIecjn4kHE0pXIsoNA6LEVXUGISw3M9qqrmHVxgPJylt5hVE1Ptj2owl1/JU4nX9SX5FVlCsdt
0Wi6ms46DesxnK9k4ZadsMPG16AGQZUMRXpyWZ+vYPhMBkhDN5ZcOg0AJWoZXdzXFWvHo4R/v/Eg
NuyDSDYt3ypKgFYUW/u+bl0++ga1jw/UJnbyCmh2rFHP/XJ0J+1bUFPPLAD2QJLdCIZ/1ZHh/GSQ
XhTKOsMHAcJpp1UTQlc1lOcm0dLf619/a6zI0PifVO6lWD2pqT0w+JyvyyHrDJGuThbM7JfG3TyN
gK/+Uk7nAjrEDkJT+KruX6qxS0IUBh9XWeak54wJBjuV8U6qxY5QK+vd1J0Wt4e1gYrQFeuqWdvu
psxTXtlBuTcGkimyqsUInad8H8Vkfy+XAko/Qcdi1yusUgg6HnBBtmYZ8mlYPVEuHjRVRB/r/KAh
EHqVl0UWwwDhksdRR7IuXMcWcdTs0UnF1SCcYZ24ItvaeWOQa0mJSBxrtvhopQoK023U3jq3BzYs
yhvIjiS6NDR8C6mNacZw9WGKJybEzUzcNhVbia4VUtC81ieaz/x6npxgXvaz6Xm9OX3s49ix03Eu
c29dr00ayaWCInvcA9bkTmyehdpBHbqQdKCbZoevJGFBIwT9yn0b6zNN/it/a7Uwl2Ntv73anWgl
WIBBIRtdzsFLI3CmghiwKpcWfSfxNMM2C74XkEaG/qPLRL2DCyAswt8fnVM3pWMYh42UayWifKEo
0pz4/EMhnldIyh8a6rF7qwLd+PE7NW9ES10rwYUnzjrgK08uZawNRfyY9P/tDfeS7wgb1Z5Ctp2U
qfiKm30MjygDhlw1CNh6+XhEfTamu+xP6VkgAqNhmPDVwPrWtLf1rMjnt89M86okNSOhA8qkcafg
4yZfqP0u775dKO4mqj/+qvVWJz5+m2LbIoDqZW7yr4zWxzGHMxDlSLIBCUyrvQCVZoXfzhwFQgjs
sOdF9zFOlIukhImE8cZ3yAe2GVBZ93Yyi0unjH8KTI+1eOWz/xZf/vLl/So/1gTLUxQhhiyD2UxX
7TcKdteAba3HXgRMg4GcezJZQwe1DpL+2i7IUec2xPJGa+5Jf+SmHPV/mC9ormscgX6C5rIkAnlM
eewbsWn/kjbRu6G93HjF3FI4tlPLhXo/ZgS98oxVq+tyX47dPrH0Fid77Ps7js7rEqQRzaK5VQvt
MeFLLKlyjeuIi5OVMp//BnHcAx1yGSEjwLiXbKSXyw8duvX3EgbQek1vbv+0sgkLNp/gBH1UlcEb
3dDMvWF7KY0NvR9EjP546yfQQ9bOL9B4POVqyvbLeBMK8iW0wK89c8Qg4ybK8sOLGisi/F/lzoDR
CEqGdM8XymVvyYQ/F5GQ0OmKPcHoCC6wgYEH04ZzovtGnKN1eUDaAT9u6NWuKTkHBe4vIWshUjSO
8OWVMGvNa1ud6UyzmC4NgZp1qYsJlVUP+C1/ssOkwN4hRfSXlPeBaJE0Iz1ZNKRbWygeZjqs9ZSV
GW3jLQP7ofOwjsJztyhDFj1DYfxJPvDJ5oaQlbzUCqbHnk/OLd88r914TPYRyXoRhUaJiuN97Inm
rf2QVKpa+ZfhpeJd+h6/4YXIFVtOc1bLJB2wpa/HojEw1zASjgopcEuSFsDuHw2HVWFXN7JBMlTm
FmA0qBy5rnfjTsU35TbHv6fcqsSnWWP1NbUzm5KlhQ0fkC/YS6WmAZjwQuBrsYIkixk56SIYDJPk
JpnDmME9KcDPXsO/9YDLFm+jeMkrciXBkFCUQORT1CtffM1738vtbqQOw+R7k7gP7M4h7x3EmBSC
hcfXe4wn6fPij6vu9ieU5Ua70+RTHyP1xq/egzpc1CLCGPYU7GkEi7XTjkTD3BoA9sdRbT6PR96G
OSDpFUW2bcc2MqwShGb97leciCTqnWRExTTHxVzYznvh4N41CEZLHiUTmDc7Bhxn2t2ltbOoW23X
L/fz9o7/HwPRDr96Omzkxm+RTeks/Mcdd5BCxagBhLaOEqasBAoIOCp9WI7o8hvrJ5W92dmO46JM
hjTnCO9B1i65txaO/Da9ZSZWfDOA7dlusP5RY2YCQfgrUd2RbjJorbtcpy4RaOiGhSeq85ItoDPh
yl6NW4gwqbOhfTeRznuME32p5VNd56iBgwKrwoLc+Lh8Y2PO6bA5M3Pd8Nq6A9+noKXTYw0o7Acu
KlPhfFfE6yCAXrIgxxb2/ztMWru1B+LI1EKfNLKt6AUPeWNN0fIiOaxmIhno0gl6wzqxh5x0ZC8I
DrpKmFVRermBkn1QQ0BjR75PtPeS3wNo9qnWZtO8kmbIPu/ys44mZ5QKnRt3VJl0XY+YnV3YGNSj
XkES8sVDt/9shuVRGeM+/b64w1WhTfHx94e1spfZFYJPJ+oX1cKbzuVruf5z1DvOl5VGQUNfTngA
44+SwWuYBOV3O99jMWwzre4QjJhtMZWZsE9waRKxj2h5e4pMsPDZtJKkTSz1cou9zFUF4xuCIYkY
yzon/D6Vai/gnyUBHM3o1e/lC3b49bjICtFHIFW/DcT02tlF12gjNigR43R6rfY+dLdAZygZJANF
sXF61B2ZlQoEjJPTPlu5oRWctp0Te2C6bWSgBKn2EKgi707iy6PYMzxsXMdckWd4V3+BJCgVNNmC
A/v2D5zUn4PfE4OgyB/ywd8MKbl6hZLnZRhZKyHpuOgTpbsvWJ3PstXosnKl5ivjw4spwjPqQMCb
BY5jCYguZ+r71PlY5X67YGj8ZaFTFf6ARSmrZTufTrooqT4a3CeoHcwrW/ymSz8nuKqXUeKUM1br
LI2wE7VFzgzwKJNM86NGeAB3FWk3jM7dvy+6tXRg9saCUQEYfC/jxQSSYjzGkpKqk7xshEhTch+r
zQCD5ecLZsYJ9fDPuLVn9LlQ2Hp9q6x7A1w5vgeNYVHnU8UjRqvc1FZ1QUOSWwGNuGEH8xUwzcpJ
JVc/TKFWlLzeMhAIzzyuNQNzad+wK4cWSyySIfN4dtxTBw6gKXVZ8ECFJuVcyZk+yKjivyN8AbBj
Z7GRG+mj1RtR/rib4dMxl0nObZmfzHqiU5iF9XJjJLVs9Ay8s0WpOm726MJhYaDyWEPTecgPDqoV
YEd+wDPR2xfBKR+ZQp7dnlthACjjZQhfK8/Abl3Si5DkUDRfMuPEYfgqdhJ3MMj9hQb3cdhYQisY
yJ9sHNAfXP4g0emh6MnQGDmfiojxf/o/DoPl6eEmGKeom6wuM4Xm5LhrlMbnnSdYHkLhWyesCN+A
Xv7rfPs3zFJyfyoz/EqNaZNmSCJMY02eRkIeGWwXFrL0POn+QRHB1gsdYl70quoJdOLu+jpvfuzs
A/s5jvvEDV4IvZp0Q6PKAdIw6olY6+ZteeSB+7cSozhGPGOe7YGFlVELSc00mTUHhhN3xqKn41km
lAKXi9UVnbCmaJcpLGdeQ0Cz8EKX+X+/Kr0E+ySjGt9xXxmdz0ibEy7YXT6U/7jJ19wjQwHlutW7
6L5J0Ad8LkIosI1ccAOd690Jn+/YnuejTzWsbUvbPRm/TiQA+o6tJJP3cg2xc167bH3vP+0FTHsu
KRcw7owkhk+xOLwjY1qyG1nhUlXqq3WGPbQ6uxqcau5xaJoVaL43GTRy2xFvwP1Bm8NDP9QDZnA6
qfP9k4I7cvOTwXv2LmGoihSDsv1zToox5ziLgg3v7AX61O2vtorBnU1GIZqNMBWe3z2eOdRa5bzF
BDeIEwf+2yb8jacHe9rvb174wUE9Gno3YMbCAqNQoBrJw5oA8gcFgiAUKUIyeR/ZBy0N9shR9zt7
AjqwtNDgAsGd9OxZf9PNse9jQgrufTcSwNeK5ZqxZfNcEDai5/rxyx5tLkENPsYBkxuzeQv9srG+
aTl1YeD/IyXCGMB1FQUZlNWM9I7ZdyPhkUaTNhpmpk4NwX27hk1Hvono3hKfoZk1qOTfWsz0wEuf
ZsI6sHh5YKgQXuV+5T5mix0EJFe0BDdq1tyRzISnvemRZr5VWe+q/ceK96UHeOtFtt0d2JKonbdB
KdqIqI4CQc1Uvna1iQvR3ZtmtkjX8T1dskONEEb03apXba4JKg+GwHq7fpVGI8VJg5y2RJCjZPTY
qZGiQCG5b8kRedgsqS2q3UQFj+KlqvtXuPy7ou+QQkzLX0qpFtD3/t7qDFm/ITUqWNHCXWxfY0w4
DJbAo7lsQSlEZaiTwnDmAU9+oCVM0mAxQO7gdNBXDMWiGLJCrC6Ih07xyqvYeLjSROSHLYHo/qxI
BiFtJuE+5uxUqAPy+9KIlgqADXnt0PspEYnCcFzLJIfrveYZPlB9iLrEOtajqTc1NPEvPfBz3v7l
2b0F4pfnXc6wjjeUojpwLFc9E6wjISAdZ/mbDnmkuXbTOnk+unzhLGdk5zaysohLe7l/wyJPkAAN
9AzESORaCFHiIrv2j3nRXDkmnlWqxJnIS+4B8P9/KdKMha+1Exuq/IZxgBB+ZFK2Cw8zsSsyTgUU
MYf4VvHzfJFMUJiFC/E0tlCSI2AWiG0Ticp211zn/5VnoVVVLJhhYivhM0dmgWDw3h11PZ6BiYH0
iM12qlDp67yOO2XaGASpnO5w9OUnDKNZdxjSs1NBJNnEVSmStE04rIj7+fw6haP/F49todLDoz1p
RUu3A1pKFuD+mVAvtkyxv4B4oL3nzaHK8f8KK6162glDxqetEgYTkXYQgxQmu+a/uf3Y8iqgqrOr
rXBynpfxuPCPW0yt3i6zFXIwYHSqacXTFKCLEvJP1p3I+f5UXEmvaoUxHxZ7i9z/qUPAPajdnc7H
v2Qs48VmHwHJw9BHouh7HvCn/bIIGgsRls53ivqDsPCwOfPWxYRNEWdkTRsWEzGTJeCg8RutNUkw
07xLFChj7yzrETsDX+85q0jdSI8AK/Gek+FSmc8tu9XA9krXo+sgqdoWcgGefLhd6//OF7i1cN7b
Srem+Xx/rnPLA+vKqOW4SJYZEqcEJonj3W4amAxtRYd/4oADHr7ekw0YoYtKVdT2VuDgwsHP3zrT
YLNGdwaaSCSUp0eenJVd5MzQq9499pxUrwi8vJSR4fAuz00NSMXIQBfsEpNctNRObtXlktPVWka0
zhmuNivUDwQVAqnHaIw6Hgpe404draEoN43Z4ak9dRkqdGAtuTjoXMLyZKxEGq7DKZRotMB0JNnm
7ak6NUpwLGLC3w/QOOVQE4AzUzJ/+ouZK7LySSU+J0yLwb2fW341T/QCz0gad4F28CPhpHQH/Jy+
U3roM7idSOEjWjL4m+2wMXZs+nFlFhVkN1L/U3dko6uXPIHBbEGzaKHzpRCAtqF3cV1igftlnqb8
RxDrpCGFlKYAqw7qIiSbnKnaa2DaIBxfuEChqJ3MZO+nk5HegeNGsATXqdA6/Xq18qYhnHURwBpf
Q+wHGlJL2G1NOw1Tsbga2MeBUqRAxSYSLvz7QmP9ssCfCLUbiurBW5pTcdr26vUFFZkBjdhsOusi
GIAynyWbgKaokinyf8vSRNM9Uj5W1xWjWxzdIwHJZZsXKu0sW9MMQ1g2Wg3BZmoGrSoXQ+cBytfd
uuKRFxEyXHxWV1gxHwbHWPXX+0RLMV9BLk/jDmij97qbW1aLR0rES77KzisgQ3Cc/Fpl34aTlx+r
8+eQo5uuOBBvuzi0AgFYFh8V3J3iEbCdozxfmnEimSKb2/AsVnS/tb5KkaJ6m5sCsvj6oaqTMpl6
1qN9GeRvbyZT78GIDhfM1+PJ03Fd7incfj8gv1pKzH5AhZZozhs3sK635Dvhtc65knfq7yOsTk3p
AjhVENyZITKgxi61/MJY7FUA3xZalmENTd7nPJVBSEliKjdqe0ane9NevhKAflq9atOkynUbOGA/
6mngXXJuDab39drc5N0VP651ERdMOuNEpa7bM42eeBeIWeA6M4hWZeuN5ACrBn/rB05yEHvOgqho
jAhF/80VN7K4rVjInpEYHixtOAFz2Zc0P0YJJRC9VNCCkqhVMg/m0k+pzDL45Igpv94j7xxfdySp
K/TO4Hv9XbRrogq75awoo7sr3TbgrrkT5bqZxmvNiNlP572vdgsXpVKg0K++JkSw6JWVGx5AlJJb
IdeBYX90v+ZYNxR1NkYunAxgDN+SWcgNtdbczaRmFKBgT/mI9yBKDexD+SAAhhVyPvcPZhFg5Ttv
NHbPPSdjoL241JTZf/6TXzjTZpddgqQ6lOEi/h/vb3STqmgXxGoB59DeM2rbJByw+OI8CDRzqAQ4
XEsjkI21YrSD1/ZuzoxZ/+l66ixgWMTZDSt+HfJnG+EW41C52xLaJlImrZw9WuBQaiN0tys9oGbu
/qS22m42hp3BPZfZ/etfUTMMXsjxe9CmCCtQGpOd/3704bkPr2TbagqGLBzB/56hZ4ePQIqZBGU4
nN84WR5oQAG+6DlunlkfC+sytDePevvj7aUNZtvGq7VdhIVrrGiAzgs9Jy7R9yVZL/48NGzMFrUt
0vxfm4JaEC4x2FZ5dmnNolLYbGIzrY5dV+tplRCro1YTBhHB1MQbdmJ6rLczefK9LOec3WwkCmA+
T+1DqS2ISPSXvrrvHS7ArnVyKeGMIxRshsleivE3SJb7zl6tHyTe2pMUBHPEP3yAqXW4iWGtxmci
8O/EqUPGNfOC6lN5E0EtTLz9l6GUxG9E1tmKVzOLovEuAbi1zw2ewfrHPxaZY7ROdNZQpEZt7Ztz
CiTjCsCcyTBm0RB34hSxrH4edL2MxegV4XqYAm/0POUrQJJIKWgOfI+wMqS3mZ/DD/EhRRs9eTZ5
/p2e3fMaJ8vH1/pN/1wkvnj9ZXzs0a10hI8/hkXZemUH1SrcbfyfJHMnJSVcvATZpjitM2KRubgU
x6dYssACnlEBcBhQGhusOqjYbwWj93LVb2OCfv+NHWf5ak07Nx/aS0/qG896v+gGes4FfOQa/2pl
n7jJYSQpGCWZJLy4CgMWpb8/0Ldwnv7XsI8dpeAkOMOCkHAuIEuBmwOGqXenZRlOyFxVL43rf2O9
nvWHCjWQAoLSBm/G+TIRT069rTs/Nkk63XbW0Z7OYXw1OI/2emtqOtNMKXmcc8RCxV6LMsbxpID3
bztrUpWhWP4cHiK4CfTGcYTzAFrUIzWGQRDRkoDpAysMjPjTYPZxRtWSRlLKrHIezvvKDJ2TwBcS
4ZL4Dl+SqN+9D6GpzN6+yxVnQOs03l4+LKdI1G1AJ8NCrotVRClHIpni9HbXmLvSIroQy90y4U7Q
GL9tNxAGHKJiId5Geo/zC4gjFq7KVTsuuzApu4v7Uadcd+SrOO9RmBle70nLxPYVjttO+TFcMiWU
GFM8MXyt5OiotIIWxKR8z2owamjKTbnqlD2uIfahzfa9cmlXgjIeHOvai7YYMlk93zi0MQV481xJ
I0wCZz/hSlc2Q0G+J8k65sfcHtX2iw7REZ3GTIkhU2szNVeRXPzzxrXbMf9xNj3gLwVfzH2C3tv5
+tfAAmAP0/lbAvMetHSHvnpxKiHJxheuPoXjJDTxVjWOro2F2eY8f+bGZicppFnQUPDM8/qZ4gx3
zaDwxWNLOFCquBUZxzA7beUAksmvcrnfDYqXw2Tpcn8SVNyKHa/ctJsvS90M4lUNFPJfyLNcThNm
W7R4KC4lpB9yfvwBt4cBo5vOYVVYkJo5n6N9+eo4FgqtLN3rI+95Ic++YAYf6tqphNwq7Z5X1bnV
KndLZEnOPevkb9TMnOE89TASuaeCDfqGuOLS1OxrieTanhftvGG77kdnnrqOrrHmyA9EUQYAVz6P
bT8kCHhhV9/PvozKVgPjqsUBzfwJAvyjQyqhG6kQiXxEltx2/ZBMwsa9LeKx8IsPinFU9/oPCap5
PZneXnd5HUAfHmt4YxB0fnltqWrTzevmY87uW9bdJQc/6H7Zo4vsDJvVTUZCf7RxA02rs5EsvJiQ
cdUQ/yyTdCsPaGtheoMxMbSCAgAoCLq1rUj8s6hiGFv2iNJMqAE5oiKeB1wn46aqonERwrYIJZdv
QolB2KxDXYt5+WLdY4UDFcLFCvpYg+/KYocrhyysMkKk7Ne5kfunubheya2ZCiA7HAMhh1iGiAd3
nQQnise7zCn4vPuambWJy6uZbQxz1KH/xHRB9TEs8WGiwZn21L+iRbGzd2Z7E/HPM4Z3jjhXgDp3
KRMpwfKyMMed8SBhaQvRF7Ydh83NGFG9Nvf3c9Pm02ede24jcrkKpklBDgSRf3JQqFGVxRQBpA4w
yqiJZHMcxBeo95nBta/P05R5qip3vQKe+mTVGSUyqKGJU7n8f7c2cj9ruCXc6WS9/UeYBGxzp8lg
jy+HJ5uCCB9iaTDhYhoKKcCOHoINhfcWbNJFC7xsDrjtvUtHqEkwtcq2dlIXGYwPU/ch0s20fDQd
o6ynjZCTkCcP0zMImGomFIBN235MqA0cutGww7GPumHdoyzVuYpXeXqjYvECvsXqq6j+BIBLzRD9
GCNgNQQ+XyhbKLzODhog3tjqSoFMMbN/BMQj/0HPFYIIu1D8ShtLk82kVGnMHV6blnpwi6RKzZ4H
QbbdKNtj52pFmbuq21zAieOlKjlT4LC1TeW1v80V4YrRoRRMoEdp0gTlYQbHjhbp46bThsEjIc3H
mGBOw3szDVHiIVLWeWk5xBBWXktJ591GQMUULdvWARMvx0uy7TGoJeuu5Kcspr94iM6bATK3YEvs
JJ7rZbT27PSmHwC7aI1ugb7QLFt25XjsKvq5obHoRjxtfJPdHbjXwZoj9q+pTzxX8r2AMpDCXgAP
q4vjIQf0OduVqCqfBb3gU8xuOTOEAj1gkLSU8uzrRnGrwTcw/jiRfSajcOnFNe6nczPPxTUBz7er
7R7qEXiEHRu7CT4EgqhL7aEWAq1rA3DRKOIRQo7LAqZ4H6f4/LLyutUNxN1ndzwHISnj7KzLff+f
Fi0HOCle7yW+fXFbY7kyrvnmLQPVH3eSLqxxwJTHkEgDXiDl7wqwi4QcnWzos79SfblOi6T5lbfK
NM4WPD4Ckc6+q2ii+HIXqa88tj6T9d2JeVTkuq9BuRCz5CB0Z1FYnW0asQlnL3AdgutkPEAiHEkp
CRw02vsmYgfVqI6MCtDLHUDwh4dXdJoaBsOhM/Num5pX1+8+pdtJcuTGbZoBvuRbf+QpkcJTreCM
P9pm2xlQjiPQqDdHxd+I69olWf4Ncta7t6IsJGmKwE/ne/IW3K26h5bP+3ciMgbFdF1KpCJqhfsC
UdRvGvaKqw55+E+5Or2/7Y6jVhFlRSTlIdk4rshGgkl/lNZEhn+Tv3F5/ViBiAjORjlSs37Xj0Tm
85lBIZvqjJq2WHTWkMd9UpUMSOpoaun/mOVkvm3B0rgBBMSGzhZwMDCdtQKX7wFrTet8xCEOe61r
RuQ8sMwcZXv2nLO3PFKE38gSwIyrBSENCTMZE/Lc1Fe2kK4z7gEGBAD4TsLt9LtwhgcA/7VL/iWo
ZY2EED8LaFLoMW0sVoiq/pHywGbdt05ER+pB93yAuRbEIbdoaFoyT2BqP1TD/qt1LWwCheWZmNjQ
az8kasf4ShAkd9gvk2BqxCtVD/fE/Tdp9ICFpXL3GtzphF1gxuDmhZhuE0ZGLsgXijMwHM25Yarz
b0LxOi3AuEJWhYA95kD3KuPfwvHjYCLgBPt9Mfo6A4grl0E0onHFLeyImE0m75m0VgQUArX5jYbD
gYDB9kxQaD6/U+eFdjRvuaMVoJMo7EuNC34VqOiXJQP+aXJmMk7B7Gqp7cMDn+sGTjrWIiacN5vC
V0459IHE/uWgjmKfZ18fWyB2JmoTX02Nd7v6Wlb/ErhiznRxaCTW+ruqtuznnG482OoRkFZo69oq
x8xnEdPosoTwmlKJ5/TuCEd1SJZX/C5yxCpVVPNRpBGh2yEzxO6fyA6KqgvF7dUMyYp6UeZIrhjc
SXyeqxs5xDkiVQKR8W5vb8h9nWSSCpXroj1Z/6Z9kqVC41Zhs3vq50yymuA7Po4YA2ew/1f7RliS
jsPC8Mfa+lucShookxJMlqhgnik+kc6B3yo+ATDRXBIE0Vfq0l20a6bmIWccYoiRm3dUpGDGhQyr
F8m57MYStjrTIwaSu8XusDXs52kOM6bYpnaRVLPca6cmpBJ/U4IxqIlzZr1H8O0kkPr76TVgZVCQ
Y5JkDE5q7P7/UyxXAN3+/y8cuW2fKMKW7hoJLwlmauZ/n3+8/35Y5IzAh9Z8vxP/1BG0myUh/rhC
3u4evLQge3OW9xGelxYmUACgfg6afTuYyyyAbFhDDGbEAsndFUIzS6Z67DRoISeg3k8gSdi6nAhx
A3AaUSBKriUyxIyQYNM7gTqtiIBIFqGvVnuH/NEoOhVbjnKTWYJ2gCOyFGiybjgVwOff3tnuFAkt
ccjku2S8hy+jgfwqk0lXecaQUNAIbU6CpNxTrLBPGoonChazCk6VgHttlGGNwukOcmkBWZuVo1QX
loV3gttrnbLNT8V76Dkzen/pH5CCcfGvNqpBE4vocFqcuL4=
`protect end_protected
