-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
0UK0lPwNYix3Iu2Xovg30yMiDmWUhJoFLgtTVAZXw/nQycLeQ1fmlqMVfZqliQfF
7jupSRFx9ybFIiIE21bqU2DxHdvSkzJ3p/Sck5F2/5SQEGDk2OwJd3St3Et3c6z1
oWO8oLFrHYv2713yy7q3arFYvEkeldAxBrCY0wWasaY=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13248)
`protect data_block
YJ9/QNWVOvOYSROGp3CbIHPq5xSvGLUaT21CiFTZGB63CYC8sltJ0DX7ydGYG36R
yzI43K6+t3D2d0vRbw1oEcPWDEVuCt5wzca/d+FrKUdOzIDhmqdHdJ1GSuxB4pIy
fOY+ZdxccftziNc1rawqrheNBZLvpJbPBm14paYellfccIbHuVYfDfPTA2Bh0Mt9
hm24m8idoVXjb42FOrdC7tZyf+trcmT/3Mxax38Zu8sEwy9p0eY/PcQ4Mt8X7yDW
YJTHhEl1GpvXRwDSWEB4oRng8FqvGvC8L/MzcozCPnX4CQoPFNlCEmORufpnM8qi
RcXzY7nclUhLdTdnTczZrmjb7w2rqqhjW3vlzVo+0H5MXvlKBQsEBlJhsKe0fMZA
/8aiiAfQf2eAxtCJHCdgLlbUzjiibDjWfv9ellb9b1Ea2vc+9+e7V8neS7QSmSSm
rhEAd5c2QDhNtR6GbuRAWvArOma81dBmUgEpFwDwuzBkdexGCWR4IAd/m1Jx4yfb
lyYqLL5vwf5RdXOdq+bL2Q0xpNiO0Sdt9y9ktSHkSlc8W65wA9W1zz7dtPBCneCY
TbtstE/tRwaGWmnAEf/6YyLpsTeUKYPMG2Rg3EluyWh3rEtGPrtUrl00czyZhJsa
dDaCb1oKDt8CmzD1qbw8LTxsc2GsRme9JAQ6fUb2QtnJUcVd1zIKpTaxyk4EBXIC
6wzXFFTz0EnR5mcuZgjcNI/yHJH8sohGYtJlUj896YyJG9zPUidvoKjPSEw+tqsC
5xy9q09YUxoVcvmfEsTEzPJrhN8Dwc6nFRVjanJp2Q2ZXZMA2VtK5D8tl/WvSg5o
+C5zXAjovVorU2GaeaG9w5a6HLUQbHzhLoHkoB3f5v4kFQRdzLvIIIA2y1BVE5Yd
IeFIht8M74dto7kHuylmjUxsCtAwUkg2fpqK4qi9wmilVEvjEqpGSyTU3tAeC8BD
4mHqn/doCzFKKTsn3lzgCuyZyE66kFfTT1xr8iGyWh2z9kUgm9ETEXZzkwjP+sBl
+4fDYU3zpd2joMNlwql8eot8yBHVXcrEzmiTSjrFPHdmK35pT8y+SAfEe9UKv7gS
S7b3+gsoMWhEPKiB0+WP3NqmqZzwz1AW6cliBpqmUPlQ7D5M5OIKSvIe/Xpl6Iwi
Mpksexi1kH+5Lg9/SC1yWKII/QrUt4wCHDUKZrPhxT7EFoQ3xas90yuLWS3YVlJT
JW7Qu7hzOboqskjWXFFVa+JrVq8rkh1scSVCjbm70IZYQoBpfPZ+VNrQbgQNBogA
n3Ja/aljS9oyUZEuP1SwbEFaMHZb3ZSN+aqmAH0vWfy9Y+w6X842keEuKPsRrEKt
WBCryZWp+8T2r462E/xzAzpMnvGbfI9n8pNkxa2TYRYqUbQwxa25BhXDIFFscawA
vwL4i70+FgTLiV7v5n2FvfEw3arvqkLtsHtvC8hN3PTTuYrdigZG3iwuDjCu3+BZ
Db/ERzf81j4ZjDVBqFuiXKNAN5IvvXlJOQgQIiguOPZsvMBhUQlNqJvWludWTUfU
vuvndNZ097Xm51Tp7UYSIIALFq/Sq5GWfCas5CortmRCPpcd3F5rx38gMAqPBGRs
kUGzsjx42I7G5CKhJCoQZF9IN0RUj7Iq/k9Nk3vpfaOtkKsnjH96tNWJ8PSgP16K
qOHO3rarzHmjbUkuc9aS5gdpeNOTT0UqSw1YA2fVaEO2HOLMiCCmu6od0KKw+ZlR
1vVo9G4QnczuoF1yD+q9oJIrqR3aWG2DbAU0MLVglYwH27HwT2JG44sa476cqtmy
KZwcG4BTbxaJkDGbYwWwQF0fAnPmUBX2kn77xYCAuBwYnEpyAzpAsiAr64cRSIhg
AAh+vAtXXcei96CyDnmpOIhwrfsZQ7M80Ef/HK8wyWGevKVp5ZusA0W+NS2eMR6F
T8C9+mYygy83gHdaPM0g4+VFBZW7Ss8xrAN8NtAyg6gtoped0QbcyrCX4YgT02Gj
LVDl07deTxhiaYjRzmwmxN69tlGics8udvdIVyiM62804oT4N3tjNq3hoVufyLsg
FsLZ5pdTh3WGWE9Iwz/B8fQHT1DacDDXSrJFM3K0gZB+OAIvo4VoREQtR/iy9TmD
s38hfYHRHx0K2WwCUha9zaLY0ZliAjue0J9ZzothemFg115wfMZscsxUzlytAqWZ
GZtTDRVFhEsIXK/EeuqpbiONBBduwm43cOiLjZzN+01iKFNbShyJUEL/cOmu6fQx
Pjz/p6pcpvhTW36hHs+0Nw+l1BIQCIDQ6G3F7hGTAFX+kEg/i0B2/owCn5Mpq81h
pZtDsvob1KAung2CRKMljAWwLv0RD1vmPa3gUE1UsWcukmJ70plLI2h/Nq6KseO7
7ff5cAzISkPOu9kDZSk7VSnlA65BzU7qWNODTVqW8849dfppZCWpBZWSMixg7eXx
9DbNAHrRsc74mA2/JjYHcAwE14JgQ2XRdQT+6yAbgJaSVyYPhBWnjHMFkSb+sXAC
wBXKSBssGVjN0qSNIpj2183mWvV4DkBddT1DSLHFOLoViSuCDkxspiflnb82ptR6
KcTKOdiPEifJzM6qTOV6cQGgS1xNoJaidibEXjb0zT+Nxi9j+HSIdlugqqhNpcHG
GI3jR9Gf+/s+fIDc5x8pCdaF50VKFhrOP74vI0vVLvl7jo2jIxWhMynQWO2G2dlT
8Fs0OhD+nIdK1Ky3g8R2/ks+ZjWkM4Keq6/n+mGKsEZsSD8kS/ZVXTyXGIsqq9k+
idN8ZpoRqZMs07Zi1VpOTvy6oTnidJPO3v6w2WT7bU3GTQSPFfdGKqKAAEiVoW0q
lk26u5/pz4hhOOiOH+S+rOayRNc5XikKTYYfi8FjfS2DSNHabEIgZos9ZhloETvW
keB6PHkZTkwpNqQ5qfZe0fIFmgWXzggWCXxz2aNMPhCw+dQ7DGRSwSc8iVIxjlKP
D8i4dtCm+dNigp0hkhgUmoXvmf+cNyxIvrWwd7QrKXJZng5Pg9s6xjNygQ8TunYT
5kZ1k9RtpuNhN9Ccye9ZhkCwqmWPnswcL3z+7kqHyJxXaERAW6jyfW5rwQVytf6y
LVclsLKiKwlPFz+NLSvE2zsbSJfSZ3aRf6vXD2ipobrOb0VYP8wEZDW4bk71wHHN
gEt7La6ChJL7mIFWvxRAVvE2ydZ5FkeGRoVDPXjgnrb6kBdqspvOqTICbyyI2tUz
HSqAkPF+WgTSh6lX5BqcrlzBZERvjJ33yQ4PeBrBAWhv6cPfDyFRa0avX9p3ojJt
Fc/7R+cFum6wbKs89C9+FScqNOeUqVBECVnVIAEWSH7rekhA55ezyYRi4xTlGyaT
wsUqOr4eWhFwO6TGl3BojuA4xbOrdGZNJReUXW8Hazh1zPBz1RajDKYHEJ/2OlT3
bXMwfdt2yn4c29wSN43Ddx/ZSoeeLAhC8eNnRcwPnZ3Bf0QJ7GITyOJfDcmBOy3q
at9CPGWjDQmcej+ncgaY75btARPo2xJhfWQXBqZJ8AXyIfK8Ip4G7KfOd83QyjPP
WQbmPelnKLqxuSAEHFWmt3woKmmjFOV+60+8HUJk2xXsQUX74oCEA7iKWuhbFF7c
tWIVgzZvNLWuYBo7Ve0Nl22JmUhtoSZMV+2Agdem90kOE+MR/xl4NA5OVE/0Nqxf
VsaLy4f4+goMwq/WvkEi7QqlOc4A8I8s4034rpI98YvJlPS9ZnPJ4iA1u+oZSXkL
v17pxch2LVAWEPeWSsByRJLL4uAy+VGv8BBQto1ARTuCQyqGIsdO/YDDv5n5XkjP
hBwvhJQuE2GP2jQI9AUSo9UCTu5Vbz1CXNfCoNhYBcXCjujJPDGbpmJz/e5FxS6z
higXBpP3TRmihZr8sM1ljiMKAuxxEx+DIJ1bvxJN5M40zWllBB1Dhjg5P2GKBb3Z
72G3dgLBU/7OyZVUL0zW1RL1NkKh6yojNdqDRJ3Az+Fr65/T5+aQfVVob9Stmx58
Gh5ctSqT0qtI9CxQs4vhep/48KYBqU57P7SGdbaJMXZPAUCt4sISnxw7f1hMkDmf
4wyAUFS8CYFXM4Dve4oUukK0zBPMQtfp4cz7nRGDbFOaF8XBnkPIPpb/HBgZyJPj
PVqmR/jZcFdmIn7Ao6eijtNDs6YzzPJBt7q4US0IMogaNgEHJaRztRweOWTPYXTm
L7k3Ohdz8K9qJbG4/VQRH3EC0lOI8LqfSruRJcltvA5lHea5HfAtNBNqAAgDWIDd
syMmvcH74JDD0BqhfuQ1kn5bTrTUL09I6iygijiDgvmMlMkhNeCHMx8OF+NEoU8O
VsW5lnVBWqUQFicW84gow0y7OfzbXYeFntz8wYhY9qF+4PiZ9cZoUT6g9N4fj6iq
YXUPXO2puDUeKU0DzNOd6Na8ZV5YXuWiDoUk7DCWJSu5dfWA3/015zdEZ4qPBzQM
wgxGBrYS52zVUTZAYKPGAbqHYDlRy0E1oT0tpufGZ9y6VBwrqLJt2ODzcJdZNNra
sq88H9EF2jLe0vG4iub6AbfhR0VDOHg6IbMjXXe8wEKx4TNVhqHfVgkm8FLaDivS
p/FZPnYV2B6zQuMKVEbYVzUXBhjG/AfpDI4N+waXXOYcjvtNdh5os3OFLxOuD0J6
qR2QHo2Ayo7rTTa3nIXyoCRwiXJonZBwBFV353TW0B+VAC0bXdgsFTZki5PQcYzK
6cISU0PuaHTZfLOyrFpS0MViLbNRtIlSD73l7/VFG881dgo6mkVeoW6Xsv6XYJJp
7DqOwTobYCuPcfVeCTtl1O9Z4tfceUZt1hsZSg9+XzPbIL6aCWleHoFH1Eo4jln3
VhnjJhBZXZxKf1nQO/+LQG5ka4fl7RRf1BisU9kcytcS0wO+VmM8fOYQuH2KJOpK
EryFPvAjyYUbzBCiW+NpkIP+iNHEQ2WVbyEhF/PNVxClFgHgFVtmbXVjctDm3mhX
XvvtdMObASKWXO3aIaYK0XsWcV/HuYUGQIxqoBMazkL+miLg/uDGTL4gH/3tCH9Z
QBqrYcx68xI9DhVR/J8ennlsHYbJby7HgCl1HxS2oZO9QcSKvkQmrTUdad4nTMMS
Qkpz7Db8BKnapun6ltsg2TU1AGQc4YeicJqnYZNQZkvdQjrfazjsF4klLAOxYODQ
7yizFXtSISoEEoRlC85K/KKFYHcGzv3qVuuW7RWxRDj7H9lkQzcU8b10CNVOpLbp
zqGXro7Fn+Zk/9hVZx4tCDTvYsXGdAv1t5CyHaMY18fSPLQ5Ihbry0oRmNs2yoy8
CwpLD7KnBLCZQWlvlhF5vDpW1WK2qALr3/6Y8KlcZfrPy3MrGyQb5YDz213IlXAr
hmMZX7szdXM1Jw/So/IVZeBW4uSLK9gWcLL7gvuudlHeKrqAYXEuOJNCl/Gs12ki
S8NFzzYahyW+ONieCiBcIsS3NWiHGN7u2VzBFNnKedJsk2fFWRzDTgu2Opl0e1iS
xPp2DY+uxDHKwNS+aOtwjEfSFgl0LJ67fynLOSPGitwfVER/PA/dbI31jwLnQjyD
+SNr0wkWXoZtbj3reWBrDaR4kovA9KQaXy69rSYZksXQkzCCqy9LCS0Cog+7UqyR
SrUiC0x+yClfvciLToDeEu8rodpj5bip7f0ep7wV/vE98VUfiO7kQwK5yh9qsVdk
bmPuOpgKwlB+w4+4tXcPDZmRyjv3V1A0ZYUsJOdXr5/Ch8PkpijKVmiy+IEqUx83
gDVw4JfUp3iQ6Krx5yxxse7FWHi0mRN2qd1u1HpGzZhRHE0tlZYZNr2y4lqhYlMO
et6isqxUWZgAANtmewd4sO+5zBNWipE7pwYOgX4IByOMFAyjwY9hXQFeLOehkgwT
WZSvKNLEJ00NII4jxbBSwIFKmJj4sKOMONakhWu+e3sdCGYD9Zgy0aW+gnwra8OQ
jqRdi/vUzA7j8rHqhTGAW1TImIrKROKNj4RQOOsdL/k4MwbSXupo7OvqfAPXRbNN
+cO9n4FtGv3RHZR3y4EXBTAFTwHHTTxejCv52xT1UAh+WWmaK0YoUZ5eQOap7ulu
b0UwnFdrjSjD5OKSUBK0Xk5fml8D2FJUXE1gPmMo8Ydj8U89oIvc7B9tGh3aBKTV
KIutT+RKWa78BBhmpa3embAWXd3Nu2735FyZjm3BCRJmoLBuzoc4V9jsAu1TjH8m
OTDXGn50SdN4uxsCeBcCM7ulOmeo3McyzrRkBhvGBybFEiAOnl+gpj98HtVrPLtI
kGJ+/oTauoLgAYT6B9SOOYHkKekvtYrdo/sFefLnlGFD6EpVh8AHmyFMJgea0ZOY
ulaSWj2/dssacnJn+eivb8LwhM/PbWCmXRdCGsyPWZXDZrbGrNSGeBWCV4tQKC/u
PJ2rGPSDtM210nnYiJWJV/pJN6+ykQp+GM3fWTKXOY91unQ9DyoA8xk2dPX1VS6S
DAvjsM2B0/z1krpsQzoojP9zZ1DIWFhPUoW1GQCxUW9Iw7TNfnCI4lfEhHp9Ufed
rY3Va4JSMoyokcmIcT5UGGDPQqxuYS57YuAWgfRoSIaO7dP7fsFDkpggzk+tDsY2
zBiRpBjdF3Z/byVp+PtVb493Y7uw0PhnERFL6lE9qLUESGeShFT0lEneuPo+PM3r
m3/fPJhabX/hDkliVXeIw2F24UPerffcZG4uWAihMLDAt+fk9J4HkTUJrGdCnfRA
5pny+wpl7KG7ui7Z/vIRU+X+UezU8XnD7+mPyymD0dHVGygbKkqkl1u1Lel++5qS
/wCb+INWM6uiQhGJRA87zVkvBKaaz8XqO8vlr2kRfhI42USJYCIr15I1uaMBOQ8w
LGbkqyzGN+Ft2O7IEh5J2llmv2rDCB4ttGKBMXp6Pc4c5UAWqyWu86sPpPdVCvFB
G+13+tortwa+NOiWCOqZj0xsn2/mhQDw74qJgtA7CLxXs7zzpF1VMS0FehrmPHjF
r+ncUp6CpywNvyvXnWPqE0yrCzmKotTWhGFrOLvnGb/AN3ZAEY4ocuSeWxi+GhuM
2xikOzrdarpJSIExqn1xeZD6p7OiclG1aH8DrjsCSG58EPAxYBCofe48tUpqlIb3
ndoqwcMOr7v1im2936bI9IKFiFp1ImpuJSgeS3hAIQ1+bk0PPleT/lnOqTOvLPoK
/xTq7dqAatVjoKs8z+CJJbrLASSe7tc+F4DvlDYXmiQblf/mUenDrHv4awwcxmGu
iaSP97O9wrh+p2nQnWDhuVqUk9HEY/EPpzNYdyKqE/CpN729MO0vS+r8PHQ0IoXm
YxDrdNLt3/72z+eHRX+rbNMatqH1GOHEGHZ4dA0HDkA5Ukgs6ddeqcc9AAeevGGp
OAOhKSGcrHZAP2ShdgBvan4HgpRFUEZzurMDUrjKVxB13YtKdb58hl9fYh6v6RoW
lG6Je2A84RCJc8dgWRHUYhRBeWQinNbz/aDSo0JfJLzE5rOh/hNgUIyNahbSyZ2h
aJYaZtLQfpbgFTQFYRf3Pe+Jp28YXqRgBpblR7o0Gv6kqM4m0Z3DmQAAZjLGGram
TMiB3iTop3u3S0ejZqRcGW3haP6t5jcx9xR8Q9woEIzeIn/YXvoKQbRuOm05k0H5
2XKSiuPQLwOhzCI85afzbZrEu70RuAMnP/RORvj7b3oWPaw0OuAMMnDKC/3UZlCC
wc2gv2fhYcr4LqM5eImRGkumXV8V0d3hQcxKUO0xQt08n9IEdkPCXcbiM1U+rnHO
sg0Sn3UW7pIX2Gub7/FePcpKFIuwPBvqo+LHhLrD+vlL8h/PHxp0Qp6O8qkPlNF1
Ja/jDghNHsPMTserUoR/9k4WdupgSGDSoWQt79tXni0IlPowJQCgl89aqMZymcBB
sFDvgLuH6uFZrP3eg9bluGlJFA97OMFqtNO3KBNCUW7C7jMSxu3SmqWZ6OyMC1ph
Hruj7Cir/+X7VjJmlp9Gh3UmeyK36rP4HlQ1CzYnRU7/b9qhHzy9WES0ksOLs1I+
9ewOA8Kc4qa4BSF/gGlWknuLW1gheZCzYy6LlPKU9w3E8oJhjzoCTUcXjKmc7shF
DKLvnMdv5y3H6X/ox9T392yFUhqKPkYEPoXQEEWN1FUrid7xpDOq3PI3ejhiXAZh
BvUqav8r7zXQ+ICNqLRAMMnoz5eZuCqVUKpsEZbEtvPuj7HRZpqw9oYvj0LEjIsm
rU0cvdlNYhoEyhkCixZPWR4Kq6Dl5CxjuWJ43l6k1pnxGYODs3kdyD1F+NsCrSfS
KbotyZSJrxPFYc8Tsl6QPDLIfp4EudZ25YjB1QMsQAPZ2m8owzSfV4rgM/XLNJfP
+tI6ZstLKT5E/dYoQbqhYtsaHycJLKQRj3Lm6QDQSflXESD9IjHjGrGjGyEo6g0Q
/D5tZpQ6Gxh8FGzS1FcMTpCP5E373k1UXrOEAN5gYXV0eduYlYr872X1Jq/2bIFc
+U9D9cl9azx2wz/XLQ4OcSK845QAQp9lLeZtspMga6w2sZ/XNn4bgWAH4PQudc5J
S1lHEl3MmuGFBKkYFjfbJhoschzQ09qI/Te/rwPVVnGOn3qBNa4OWntXhlspvgAd
9yAP3X2XTVVcAdRCVSclIXmBBfXbCtO5LCk2yN7PlAavOOV8V3ZBBtLTn9ls+MOk
koOp90Ud2Nib7u8z993k+wn0d5dVCmEe9cmbcEq3AW12xI/JQqbo0iv9Z3iE97fe
Hgp2L3zsamSxNtnRs9kKcgbaoIdBTdi7f4m/GmxySk2xP4SSKnfJNUK2S2S4f7tm
sTK+ynJVu95MjzZ0KwjWvKglwTjwOmTG9fZArAI1p33VfDHQpOXRd1Pkc23tTO/l
PwNKX1qK4ds3bRiou5ULO11Z/HEKLCeQIbHbpmbP2e/TLJaV5/oTIfvoCBcIrukM
3Um4jc/fGzIDnPUdG5Hx+wxZy4XpJeRb9R1/PwNBIZ+Yl8Ru7OvXpn+QH6N5KaYT
2evWk616Uw6vh5x5XesJU+OfDpsCQQNOZoXu3FetbG8GTs1LAodAc2bcirPX8tzk
kMd2/4rbkJ1739MP/NjYCu0sYvxJ38+zjZtZzLqoHfG0/ZtfugxFhzoLQeOAyivE
zPCh6pgo8yl7ujF4qpGl/Kw4nXVyxIl+9JQiXmsh5uOG8PYMH3BCrkfPcum3FN9y
EO+9ZLepBKFxjTiplPRhmlg8eFQqYcIE4npHkonJHJE2VCVfYuVW8uaEnVW1RXCE
ZHxs5kH78tBv3UZDtP9+BpsCH2RxS508vEH04ipKNl4yv5If7xiDns3pyZnA7ta+
oxEwIbQ+EwESwc7QCKm60F8QJW4PfFjLqu6e6ZDOpJWUT2JBBVeB2G9ddyFv4068
UNi+UPVRIt9rpkBvfdFg/LxE5rFPAlqFM2uWmMto5PNoZ5/X3RAHt0wVS+DfCx51
Cl22AqrsTNjbVI1exm/Zx7pHUBw4yNJaBOBZPE1OA28EVi66w9cik2Q0y/NhcJkP
WyMG+9eoIYqE0Lf1FfWBCAo2xAcVLMwSL4vgTdoU5md6pTX6a3q9RiKogp4SQu3C
0Pkr+KaenmoRfNoyIuwXeZg5yTXPa9wxuhuNmzTRqujPt/4TwNGNG/2UJyxeWAuK
mldnwcXAGqBRJnWd/zfNvF1ZzwkIiDo7IbHcR/1jduIqYxJ3cpiIG8lmcBWx6dvY
3s8m7TMAGlXPtrjcLcdjOmwhVl0UyNBHcuZYSR8xe7QF8wnVOjalp5dwuKPoVuBo
u00ys7n+c9jM3ewPBwMOpwWDCwh0+qX/tA/ewcB4fd3gZwG7ELpybul5cf/GgPgA
+fhdnpHtJ/oKWUcdwTfttyTPzmiLE8k9ooIA+wTFyeAycUB8w+yiSoM1EwWMlIEW
TsCzzqVqNflURJA/EUgdioESCvzoX4g4kI7hiOimPq5dp6ASVzxUWo/5sYc1KXZv
vn39ll7Nwa+EawMncUmPcVK6miL2FWOHyYwaL6SdJMq4ViLX6zY5hyfsEfX5i4QC
rMiz7bYM67CoSah+lKFr5YI07bIpteRoEzTzyJFJPN/7rQf8bwkSWV+HYznXFwXo
U2bEuqe7vV3W/sShIU7ENroa7CY8hLCuGRY84tS8eKqpCs52Mlm3GNPP1KvOiv8Y
S2foE0lr5sBCO1vTzrlZ9IfJH/yn9xUR+gwdI79aBOAOt0MFbw+XnpA/qCvPM3jR
HgPF6RLd7oqW+J8GP6+E/G9YdspStJt6cBt4ixsRP8gcjKvo46PevQEk9pzR3XCK
l/b0ba2Wpg4Smh2j5Fc1hwNXY8h949MLgdf26QX1MNisS0/nWeCZyLsY9oM8jaWg
Tq/UFb5nMhnQH6rrehLgS2L4bdayLqcZ0xaPuARkrMKyxXZt8NInq86o2cuZjnEM
lUbg/BvonGa6ZfYfVV3eIpYKSk1jn2CeKMH4HEkqo76JkHx8mrTplrbWgjjGs0fV
P/usl8gy5rszN+CwPAVTtNGa4kMR6s1Q9k5K3gZqBkmAuBzApfZ4QYbObsZNCB/Q
ffWgT1tJQ39oyEoswiCkCF7O0TGpyDkh1xz5AZBZOqzUy5mnDhNEUcdeOAGpV2zc
ABSz4BCA/QeEdtRCS5IFDZIWnXZhjnrxJ1vYd3uGyNWBC6H7Pa2mpfCMQ9HCF+4y
yPkTmK2k6CpeXnT4+xxW02PZLP5arGpsDRt0t0RILVli9cjxoLWXtZDM00RSfEbg
yfAOAM0qpOHjSOdMNxKJ7BMJFD7imZl7jeusC89RuGPy8benkTTr1N2lhgVOiSzJ
/pM/MYaIcfPIiea6qffkM1Mf27QUDd9hSw76E+PDIYUit3WqTl1OyhUnvUdNCOMc
NXtjhnytqFgovBJLRCCOJlLr3p/MTFcWX9g1th5Cm1lZ5IMxCmLns0SLbpi0OKQy
Ls/mwV1ACwjLQrg078WV/+dfzJjDYyp76WU/MZQEYfeQ9e3LnA387yI4bD1AcnQ9
k9LqYEwqWR5GugXuxK/MPQh4sFQNKmFyfj+t1zo3HgTSqARbs+ES37rTptndegI2
xvv3fIXNWi/NxId3T9NhGKlyIGk6OMPwKxwuQigQ1rJKoNMom/5/V57Wx7wWMW/H
fHhbroxUkFA7kJsPFFpAhOowTw8iGSeEQ0PAapNjMAkUTuWIyTcfAtdtIn2keSf7
wl69ZOfqCwOQ2eyH2/IExKb0qQlO7YAm/DuKKJ4yxp+GSRgEMm6nELV8cjwv3Rsy
A+Wh9ImFXkXDLVcn1bhExDcckTP3KIPdGnwniYRjx7H/9PTcqLW3gpcvLm3yrtLF
ZkkBOAfemyAWgDSZwW95x+SUiIivaNU94AVKTMmJk0SwAw71AR5SWQ4A1fMstZ7o
9lt1dWKzj0pipi30maqcEOlQA8pNYCnblMDoVziZh/pQeUJJYoIrXMMrJKYSNKK+
mWYNzigfVNHyQbhcY3g286cdqf7jKzPFU/xmLdcL/bsISzHpKqDS7cUnDJjt2p4/
sRC/xMZMo3HlYX1oyNziHVN0C/nzxb+ODJ4XL2g3zMryRYUdbZDaw7Wsq9x6IkxU
V5oevt2/pGO5Joq+uFq+nAtK9HMgMh/lTK4A/OtvDDUDF1ldCB4oiL1PO9DjWXv0
ARJcHiJ5nObr5a/LofKGVthWmyWxFAY8DiRmcAs4Yk6mNDiSa48T2mTLhMQ7K8MZ
cJt0WzYnFOSlrqw6HY4zQTCPkdkzua8m4F5Oc7iexm1XJmkPkQT52zSlJEDozhB2
WCeKAQcxNyP6X+ufHfniWmJyltTbLZ1y1fGmqNyp9qNx1N9B14goGGdO9lF7xTST
amEkbo3ED9cJrk3V9iesoC0SFG1BTNxHlE98rLwyQOZVl11ve6ox6l5HRGXR9/Tg
Enn35K2wDaRvHLb8Hgx6ywusek9HpwJMttGFN2xYtgqpMvrE5DO2hjq31ZvMx6O4
gWMUO//DZCABJFKS9HgQshyQQ/bUTXc+hXF3p6V81Vv490HSC3cMWgd8J3uKBIqJ
+4WbCAtQIkENqBmtU+cT15tGKwdtct/88taQ+1G6kWQ//Mwjeamg5g8r3ZcEGq6T
EcL3mutTz9pAXfmj8pA1irXaPreYyqtuKbtepuKDBLRVMM/1ZjjJX502DRR6zngk
JdquaqPjtEMz+uLRqrRiiXt8LExNYuGRIAa/kC3n6djUMO7JqLQtclbXnNKOTQA/
A+Ua2d3jCthewduHTyM9MAH6e/7rKaAodNBW2OT+3ArU7W6FL9efdDLfG0fuGux2
EX4PyC9is/XDGrJXgQojfPJrGBgZ+hAH7zQ2LhT1wGEzHmtX2SlJbUp550UTScjK
mbwrGx+1f5+Tw/xLZ4WV9E1NZsOBIzH80IAK4/kmDLpG5L+HuH5KfNXanh8KkERp
V7obj4LixolCOEROl9g/+Lx1Y8p4ZR7ZKnp3yGwznzBN5l2Xxq2NYTm5odIoLGvW
n8LC2uGqTvEIL9r+SRLOCt4SFBdqxefATkvJJLBCFuq1Xxt01n106ihpkBmOyTiP
Wke2pYlWRW+DisUqqucFQ0N3lgeDhoRDMnaMVI17tzzlL7+6K4QbFPZoom0vht+k
mDunF19d8IceRdIzNW1AKRaADdHxL+HGPzMdOf3b4XAQogz0O7o2Ysj8ioN7yoEx
YY766WRyYkn7KwG7cbZtwFFHmaed3VrLJ27BqLUL+HYxEhwR+exBkTxZ08JIHY5c
pjeIftsa4kwlTghiyQ7Hy5In/ng4wRuDftu7i41AZZFffDQJK8rcP4KuIX3/v/X/
I6KanOP8wDVSVAK6O7dr4yEXWFud8blUTzIhT3RMi2oqKC0R/0Q8+A+xdIgiQne1
giGxlMCEMcpY6cI1onSEsm4iifMy07N/4xRGVqcEjnkQ6fHTRrDDCO6bzF4pc96I
Mie+c3dYhpa5K2uPFv9zat04xsGgGxQDQ/TXg1DHvj2tnPiN7YH3oGx/CrJP3rt7
6YVuwK7w9B3f2LGf3YnAdxrcOBxjDcwDbtL4tM8qt1ShzxismG4+QC2yEfinBKIA
qg+FgngXlLLIPqx9I7lLxv+cfRLT+pBALG2kfAP5C82oMPCT4cfRlSAr8pNHTFmr
hKHvWn2uSN/tR6CH5D0O6oeSXO5b36Qe7FWYKodUY2uKXdgCMIJE8YgohAMWob89
b270FzZNnCnZkz3sB75NEGHmCr/NZTc7o3csFd9ksogMuKTKN9B7VwOz7BNwIpD6
dFR12Tovy3j5rT4JtvwOChMkB6DO7qlaSM+NU3nyLKuGVgXmJS1uIJRMFc8hB8YR
D7akqSHNr4rS6NOI9FOSW1dkkKOQOeHVaDGd6RPZA+h0lb8k7DG9/lukEF07LKsa
k1mmX2uhFSXDwvx0OY+1m4UfTQFX1JhwHSo39DYEdJz9V7putbq61bn0Rc4EmdMi
EjWqkvrdIJsYb2mw8gmImHQxpQxNx3KExM6QrdTvFJv3UbnidxYYcI4N0nI0VkNk
GIJ8eBtp7KC9wtkp3tTWXwLjO+0ue98bVZ67+/TR8yoq8zXlLEsPlRJf2ugEnld6
ZH2HGaORq2qUNxQFxBbnjlAKQEoSMywDtrYxJxMWTZtzfM5oT20VNYyDdOIXq4kc
JnRpX7Bq1xBS8juyk5bFWobvEHZbSsxRufc9FlMgvrUnv1Wpn0cQsufPkz2EHPcA
XGhzJSEnPkF1LCEQLpRPF+vLORUq35vFMG/Gujcd5BVWa8/ZaJtStWp17rTMEw7u
uxH8c+rfV+f+8/TG+AncAN6/TxlG+WkStsR3CH+j6mgQtoFxcoh8maI/0/x31qY4
E8cO2QbMjR6DO3BQi7iJsf2IExcODouhChWnEl/QOWxGDQGCnE1xP/CSsb/9nU9J
AhK675FYhBrDB9ezihBangx2xpTBM0Y7DZgZjPjX0LLQ3EDJOyTUui4kPFlxKeiU
y2/8Lk9E0wnMw2d1Bd+Ii/6A32siP09855nBzb8WF2RIN6o8Vz/C2308OZNj79wt
G+l1B2+L8dHUGbsySHsNypHMg76VJjD4OErT4gxTBKVRaZ4Z/3jdR52BdbNm39wD
7/fHjJeASA0zWCw0HMrbmZpbuUE1xTfPeulBP6/4RDfqyWqTF9cFxE/gKhcNCks8
tK4SzcgWe5d2y6iSoR7v/qsalC2ITF+cfxkc1q2XS/Gc1n9aduyerKzQDRYXuTCH
8/TWHuRYzHEUdM4rRMj2DFT6qZrf2hZmgvsH6jG1H8liL3I4y9Lx99h5eB2iS/K1
6vZobKsm+YCEhAfv4UGFr7PFleT+g1bCdjY0DMyQwWRgDIQpQ/ojJPMybIyxPGm9
dYdOhIU2PU0x9KE2Q0xi9f9iSZdgPamGTo8ZBRSSJfuj+yCsjzCe2b5z0N2DYq6U
N0Vc5YI2SLRGii72ZOFJcLgChPOeM1XZ5WbRusIzT2baxxiVu1THsT2+Wi9PZ/z/
DgryxSb52fmCIvBATUceIfLBGVL+vAyjLR71TzRE+6xbZbF2kT+NAAFW1SXJH8HG
P6ZOPGjyyn+x3swBrcVpcrzVXEwikcgQGWlelIbp5Tqby5va0i3GARQyadWJ0QzK
xTiKrZDBD8BNlvHzbu5ICbjVp19zfTlzxzeKRN+1VHZQ3o3kc+LMYCpYY+mHhrGS
25f1AdB3CeHYE3WLLso5QbNLG+YdRlXLYodBl7VAHN0uj7XdfDMkkFSNlUwuMVwV
/YecbcdwVT9I+PHCg+NnCL2DwL1XRENc+FBvH796CfZg3FJghL1hVlfWGXMYgSbg
RUzXJgFPryygH/ftOFa8gec+tmpr/wHHno67nLVvL2HNpy7/KX0+GCEvV8fVVurm
/zQ2kfwaWvpWH/q/pOW/WkbfwBFZ9bddra815THVuRlfFASLvGeqwhK9WYQFvGwY
Kiidy15DkdBFuh3ku7ZsoXa4rVvRrAWSnrlMb40w+7bDFxKerXXTVx+t8BQr55uM
dap/AVSYfugMyOhfjZGGC4CJTGOKNt20+7hstFDeSUD044ov/tCjJXUKY3zEzeu1
gkW0ictt+uyToLqN/CCdotOojFqr+ffPPIVQC5JIDqh868HqIz8MEvrvonybybhN
azAbjBNISezwcVWwNFI4x+gsuOK92jBIL5YAG737UTPv0RzAHME10Mnfj92UQVua
Xsr5cylNdnedUOprdYoq+NzKoXulHWIQbAcMEqGdWr0mEzg4TC9jvi0jc4PZYZzT
C+Op4KMczb9x5ssx1QYSrHjUvfIhyKkJTHZPAT5zURAk6cj1MlNjTHAZ7tbFr7Ha
oSMt3gJp/Qz2vyS5g058IogEVKwiKsijSdM8UpuwD21yspS9vvxt2B2vQB3IXdB5
zrz556gAZWTBgzXqi7bfcRuhtF60Hx6M5rRODcYeER5oEsaQz3IJ/sLcGrZU4WWV
R8Y3o1mPP8rJLpBj6f0CE5Hc+AD4X78ZTu0spOEAQQhT/3Bkypz2aC77qO8U9AWB
0LtADH8zYiEGvZCic1uHri850vqZvOJueuKb5n9rP2voUeAdqlPqBaeFPBC4CBBk
VGszju97xrV9rtuky4c1VPKnlbS5KSnmuyigionDIh82yAF49/N63mWzokYvCHCz
xEMv/ZoQY30abZTmzqDFcLK0zAAvYgZ9UMaz6hDkOosnkd3x9Q0hGXctLTvYoYFn
Z3zmYxmZyhpz8iU9LbHBN2u9iNKve28+WhVWNUSWifefRNJTUifGQ/fzjgtrGZsR
/d6VZu9wxODZWUPawMza9Sm8W13haOc9vceQWnQ1alrCsXU3uz+S4DRcYpoAUrAC
31KlzNDjbAfKeyZamfPROptF4npZxT/M+vL6nUO6xey9uNcv+SRXS1mP3/juVsdY
5RAajEGLCyBkz8UnptN3zAOR+Fd8lE11TpL2q1XjNwfJwkE1wtaT5fJ+q6oH97fc
cTu0nY02CAm/ph9oOoRmYMfP51mq3EueSuI+AJFrsZz80zkfzfy5Esu5qE345ThS
pld+1weG9xU/QVq7w3k3w/fycJg9CR7mqYw1kP+OvJHx5L33OkuTctvxx9oNdKOo
pfEZXgM7U6nTCgZKjlxIWP4eHNWF7PIjFblcdjG90jUwlz0tXiCKOy3yzon1TNBQ
toxxR9sCjefqyXAqxmleyvedgGDssAV1wFQmZW9e4tVap/FX/I7pbgoXR8WDvemH
H8zNACjLuzr6dI8v8gvphBreiln694xZfKw1QaVwoanFVxaSLvASdDq3+lGpu6KW
bU7lX3xlhayOd5XC55b1i/juQEXLtwZssVxsXceTuH9gamUUAfcQ+hXfxLLvPsLc
ICxNJwgiVZHVfkshFCLuWx65KTn+YSNngKM2X84Xgl6jwHBk/87kEb5iSBAiNktP
ldmbnVOs9Zqgc75yuxQpYy7Ye2LiDFUTQ7gJRj7uLwo+MxfRbBoe3oFEaPdfkT60
DXPh8G5dStybKS0KqkqFgZ3NkbKvmXvEl5civ1GA0N5mX2dKDJbUAj08O16onQcC
ZkN9wSOVrwRAkB9/gSdLRKnXj77u0aUtG2Y0WxyiWk/d8KtB39ttoPE8qaslB2uD
v3Wco1nYFVQbJa6RzCoWz5+kdsFBd5lUjE3XQoCQu2Oo5q8ICqkCwVEWuLSDLsYi
mIlbEif1qBT3p8a0QogG2/lIc2O8pEvbKJ3k49BXQ6BGbPzlJFvNMsBzUDSFiKw2
4HLaXvYGFlY3fLYXwUN+6FuyTNqO3XsweWwuJ6ownFRwLzPYdABsVr0RZ0/5qXGa
wXzm1RU2H14lwPE4uwkng+6NH277UqsEYZND9RJ/yZzxeWBKQGA59qHRcHxKr9Ya
IgpFWYYSNXpuKIkS7L7LzTQVpNRnUmjjw2ln59z9twP3xDPMS9LhvL+uOK99yHWb
AbONO720rISE3zowJ1zICvvAkSVvvSTQ6B/EArKtZB11AeYV1dFcQ/baKU5lREWM
ZnTHs8qK1cPK+lEpN9s0HyW4CzaHWWkL670FsrglpYRoqTMYApCpTAFYesDSV84g
FBRRB7QbTFFlijXyM3U/egQ+y32hjLdhSB0TofcdFNP1GkOWSmGVvIWy5V1ssD0q
ZW85ZHooPMip9qxeeInKG7bAqvM8ZjPKzg1m+dkBhlozGPOuVAxaVk//UZGWY4sL
nJbgTGOdnH5eXSbYA0RoJNNTYfwAngYnVHpYWv3m1Rm6mocjanvomCkFhHu95TJI
HU5IZ5bkZxeTVeR7ce+3DgkdK2cRwuCR4wny/KS7wXw02FhzCZf3yMcngB7DUMi6
5Xlo1BGQFM3gymROr5URl4cRAmq60TPQNfRl5lNZun8iLoohcqUi4ehR9VhlRWX7
UsWqfz/l3CwXQXMZgXU0XC208SrGsGAeZvJ4FqrxoaIP9t0RyJnxIc2ZvjLrT0ep
XLqTbHIeVz15xtBxQorNiNyJaaoyemys9hpmO9KS7TDknw7xf5Q/wTA9j/eOrpeJ
NKH4Nn9gi2u5nuT/9pORZmqZ3ZREQsB6iXZfpAFXGyisB0mVvUiGRekFvCYwtYHI
gqhd8UqCOoPNFNaKOB6q6n1sYo7zXWVFJKZMU7hvNEilLlwJPQaZtnOHoloX1NCK
Gcd64xaldJrsZERP1oCF41AFUNGQrFH/U6dJn23QEpN6J6BdLRkMiA1SQvEWnqVD
B92nhuEJsipwSaFVFf8X6iejX/bSYjDckUJX0pTLhSR3xLIb+F+JvDQuh5AYvAHp
4vkvrnkcAoQXHXoEI4+T9iR+3L5zu6UJe4ilTnszDJ5QF+sNDP1hkiH5zZp558vS
`protect end_protected
