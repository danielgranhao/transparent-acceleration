-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
xsB7DcLX8LlcCGj/bodM4FqPssH31L7C8UmDU2ZmFnGa9EJhE9JP79siG3oSi0lz
7Tj7zP95N7GEaqWNLxuM8T7rEI+DZoinw2OyQ6zZRKLonOOlqrTBGMAfH7Lo0i7e
6G/Sj7UhJVQlNWDdGypEOoZnF18eoDWUpU8nHJCX7Ls=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 49792)
`protect data_block
Yt76/WVXGnkX392Z7CKHyCnQcBxL1hKvKMszjXO3ZnEH8cTat7mVFz7FzsAFDqg6
eQorSTt09iky3QULV6UnQZc5T/QsdgtKdywAsc4KRxs5bLzQXBv1PlWESK6jm71A
To5M7jT+m+LsqWltKSWIUuMt/+2g4zZ3PMHJMiH8lW7FiNfVBihjfsd1Jj0i+Hkn
cIJwx3UIoS2q8wX7GMPf17l2o9xi2ckOxEn+r2sFEUoOuxJoWsPZ0qdL11Jk6MLc
90HSEZnQTfRsAgzY7VLbzWF7bwER4k7L1yLLsZah/9TfGgfwLCI1OG00M2CIrRsC
WZelpHVq6XMg7z0i/6hwihPOPMIt1e5cxxGhfoBiKvM4paVPJtgLltGbhUfxZapr
9SIP6WcBnXPkHtJnZwgaGaKkQex76E73Iw62JzZkCryxBKGF0wa03p5iHdeRfupF
kRmIz7yhu9eTtijfK+Q2ej6RHOPxpC+c+QqZ53fOnHHdYFDwOVjUzYkFDpVBCHSf
c0hCg1dmPd2tHmR4GKH8tbJQTIMXBBogWVOKFu2leobVxKjxIgRx1sEkyqfA73+s
Y1YrG1erriMzCpMDVQkqf/dPr/Y1rWni7APK9P4GaY3ub+z+LW9z75iZaB7ga1Ns
IEKpveQlY4I0ozgJwaSLRz1eYLhgh8vDdVQzVwbOumAiwNhOQM0B8cDwTMiESSoL
pbDvVoB0BbWPzM/EhYDBngzwn/6Jp2BojSARu2tuM8Gri5C2VQc+NDzzd7AwSZvp
yQpqVwgrsGFCB2uLOl7kbzMbNF8KpxbHCiV9nNYdxtXlSG7TTsFejuxTI7ExPTev
phZq4ywT/QB1Vu0NBynJVqnID0CCa+AVOFTfDOEe7FGy9/r8mpVevlSpqseT45bM
n1LrTQdvkIidFunN9yh+2C3FyQfAc6luvtain+EyCwURUxBiKO3MFS3ZNXPQ4o6a
rEg5XzNjhZ8eZ3cZibRKMP49slTY28CqHxgujB3MfcGO5sOsdzDiFIS3bW1YQbfU
I+CHl90gXMIV3lSkvO5MnyqaSR74BjEWkYX7FS4Z+B8qcccJQmEBoJP9sI7qOVIG
1XGF3suTbPUSP4QstOEsPbmLDXTAbIWFjELt6yB6KFJy3pSSWj2bkf5gwJ44a5HF
/hyJaaSx/OwJ0CCBfPyhSmXP/vhonVO8400I8Gc7QnYJjVHDrLY72lKnCEd4mDzm
VpOfKO6k9X9r5LWeEYjzWF3B8/eAARydzalYNdMUyon47YNfN2hh6UqedLl8qCNa
GinhsfZZ9d//r6DKt8ogfzhL/DUKhazdRDn9kZfN7+qBfUxPQpS0X97G64x0EL4h
/Pfv+or7zw1rA0zFE50tn1gNx8NvxzQcIaSIB84Gp4dkeKzW0QFlTg8LhWMWSNE2
4dKIBzZphtyBtZhy+52zKkiZJoBddpa7SH53+yZHfH6IQ5rblldvHSOsCnGbeyOx
Qwwd0CO3tocxMXu0oATEfBBZJY5PjqH+VCy19kT6hmXD91VLTN0QLw/TVj4aPyBs
Dkw62/mvuAN8S2QOeU4tKc32xktw0hTHdrz474X6njaKYmQSbY2ko5ulDTzuq+YZ
Kp+IA42cr87BGIRJeVXw68ycv3EsA2nCGy762UFh4p0TNSnrO8y3Y9uNNeJ2ibge
qdzlGDN8ypEAHAX79NIcs5NZvGXsg0Cm9Bj5KH32rG+qUOGzE394HEyGP2NS6aVL
Dml78brDyYNfYCL4/DPsUmkgK0I4VS0pRAaKXXrt+7UUo/VSieiX7KN/ARi58js9
KOCq613YAeAoO8pWhyELHhkYol5EDgUmfSFXeydLiE+eP5+Hpw2MNSk3VZisPwYQ
GH+be94UaQzcY/fSeO1dHX1tktgZh6o2PWL2CD9JdCPxdS1s0Rw2xHi7fpzJ0+TI
TxpUKklmyvD2pmXdBe0GLe1xb+3wOgxnpBvxveFBhCHr2ePw0LSWDp6un5oK/qXe
ZvN14xoBjtd1odHsoI/f2wHba/21XBMPj8CQPRO1VTc8yhVUE156zCP4BmYSWHC0
A4wGJ2Uzx787H6J3rcP51Bz1v542pI+oEutWrStP+iCRapNYGJ2Zn6TLqwdEdk+4
V+yl3TQs0Ia8ijJMAup2WNFWy+alEecSI78hPYSjGzP09iX+e+0Y7Bedx5CYw8SX
Yo98l+bx4mtz7iN9xrl+qghTC2Hl+X//u19J6ra2weR3I6JyXvojeqGyxLdRLums
4xa+Q9FCovzIyW6HNbG48ag/GsQFZZAdXNlN1A7omO/59l2/+1AV9tkH7tiz54E4
WukG/eswLJf/l6bBv4FtwvaZD3MjUqVbfioFGPSy2zP6PBDBA8TorXnDwTyoodNM
gUKiMxd/EY4Eh2n8Y15IckJxEjaUM0HBtemUW4yYmaNX1RKWA72MYV/e+MMkQ2WT
JjdvxZC9K1yOH/fGbJilWZcETfTZb3qD2rejNWu+zu9fuGW+W4CbO3OJe7vOFkxo
7DpftDKFzUqVym207RrdI6MWyhW7oGaZFJly+msh55biXisVFdTsIfMob+0oS9Ts
Qo+cY6zGvtX242TG+eE+h7ynmwrVPXTArO6xcfNGnKaUA1NGqhrsr27Bm31+Kiit
NifMT7+DwFI+NcJzeb3s9B23JQxJJG9nKQDHthXPtjs8Dy2LSTgVJ/eP/7uxq1oX
HYwlZL5/isJxVUkRykzLvNWNFSmcaEpcbUlfTPAq39+wzOTgWHYgzwhOt+QVFPu1
m6AvhMzPpZwH+DubrSuLBqE92grfZxCquMo3m2OGO5V77cZICRh4+75PPK+0dZbb
trV1o/rbygMfchu3Qh2h+ELbs/+N47NaGFR65yYvE00+zHVhN5PlF/mui4LLio+V
Ms/wRE7aCSTR/jaGTvrAaKHlnxlkqOqbj/qJGHPNcL8v3EFxhvBECLhdcwsXGofD
FO80o3sptQ5GHBS7OlyCQfUCycyGMDpdPHEyBALIAncP/Gw5I5MKjOu0YBWb5uhd
vdL41X21H5wMfudblbl31ZK66qF7b9oVciHeJ0MpMoL2gU5O26RGYWKqIwCPzWib
0gUckCQq9Ony4N4/oIn4EH1z21ZOy7QyaStPDM5LgMXnpbg8F404CeTl6UNIX25Y
cWCacBjxXBsBDiUHN4fowNWh3+pIC3HVP23232tLdArHpJMhRqhVta+OVkfiNOr4
55Fi22ayYYos18vY13K6hE0z/AgsBQuA3CyU4Cu3snNqlREvF8TbCAbMuti0f6Sa
qOrE5aLiQeTBQrwk4YKG6/cmmSDpM70Zds1TlZ55uSMdNxVjIGybV6LGNCrIkRMf
FikfTzNem0Y8je8ROSvYSMsJPPKEjq9SiSGhPa5qcMIeJCqExmzQQiOy94+EBKMr
eZtk7Xb5FsiZq+PoryNAJ4b6AUDwKFC5nXm9scnK6oh50UBj+9AFKekj3l3l5mWx
DCXLH8fAANAM8kRKtrsvBAElU13QHm6sCg3ev6l4t2dZceK3tU3nXXChRhGe+wvx
k1eYEXJgPSr5nrXg66T4hZ/NegyWeyvCfxDY5QWqos72bWWPwzI4eKMxDLh6+R9X
skrUW0uXikOc+qHWfQcgg5jr46rGCHfVFxdsjO9roVIYernUn2Hft9/gEU512LpQ
NBH8eHLVURv/7RAv2Di/takUnKTypYfAd66gzliXT+NekhH++cjWn9CwRSCKAFKK
5lLs5szZvLTm3Dp2769LSkswBLp8PFpCRBzBPmkZeQhhcGt9/EfkfvXcHYxRcFyn
XDeKUfU93xIiRPSlCGUErYPLBxR0JLegCEbn7uDVab8AkImgCQbN+IlcoaP71q0d
4mSomc13XaiMf/5n6ipgtZ+3CbZO/2LVHf1Wzbk1sqnVJ40gNxR8mC2KyzGOsl7j
gPG67nGcBQKucDc3HyJhgj0V5qenN3WkR35Woyl3KIu9xmmO8cD7MaNzSzJTPzPq
gFvStXi/ajmPgtOoMBooQZZ/tCMTdNQeEjzEckr8aacOpOduJZLX/DaiJV0mzgre
diYvDgE3eJfQo4v7PLhkpwIt3X1RNQhsm5KB1VD0UWMmIx/aFZhZGngoXgwaQIsn
WAMkd42EwD1IzSD3afWJkpstwy/iY8ftdwMhU0XvBIlCZecarLbJg5bUXAz8Vc3q
SI1KxCvAfL8LHkjh2XfYgD6s1Eyvk6TyaEIuFi8ju6Upd1yF8yA1zNLXk7hRJ4w2
CuQFZskz7FlwIrJZ9tz7xvEdQWxmQJT1oVDU5Cyo+q3LG/ltqnTdaWVMsrpoMDnt
7i1bC+fqGv7N8HYJAdCzmcUDT6QcybDjY55XtL/IQli7I6Zz4jhvxkFJ6REO7fRB
MkY6bPfSoFBfcM1QdCf7wCFLXbzVmvkshGlapCc4Vha+/KJniwwId0AtKYn6AyZZ
bBPp6wfZppNVjoNm73P/RzlsXA2XWN+mWj9TBIokR4P6YUcp4G7JFjYJsCr+vy4g
YVKS+ba8cAbmq5P2Vl+PzH3BV7QXPfUKWSWQG47Fet64mnNpJCbG92ZfRp7rm9z9
agSAwmz7JqFOa0OgUVwJvbk3s+v7Ow/KRizrXQiDhJ2glYubF9OhSELU7mXfVm7d
1wlYCPRwDeRRvZIbAkRhnpoyC6oU7oP70Pwvjto9mjgemJvDI6iG6CnSvfkTSies
TQ+gOwMdguIqmdqIVgZDhh9yST6StKftfyVo16/xmPvr8ifJmPMS4olKy3uJHvU0
ygz3QTiWHTasp7PT71yA74H4vhpIULsGEEef0hMcE7ZDBGk9KXhamEfB1ZkmS/95
p/EF0EOk6s61prWIGysq3Mw6PLFt3vSt0IMeEFzy8gE+bleVfgjvTSOsPSSiy602
tJA3SMYcdLWp9/ZT8GzDEaGpLpBHBSv1CHNAy7JIrkWK5/6YPYaBd2auCawCtnF9
3HSI/03VrLXloVhWB2mF+D49lc33uMCtH8x0GImj+3VJ8+b98YU4F1zzx9sNnc04
39ovhmycIe9ZqvdW2AFIMgAGY06taLPSz+VR1qLx/SVp9odDv+F6WSjlivEE9wWK
tQ0NhZ5ZJF5oL7tv5c8LY1xnsUwNOufKlfcxAfWLL6dJxyqZTu98I0cGhaNmuojK
tH8GxdBBV5nOcC+e+XPofZ+1D0jLP/e3QTetzox4OcD4Qpm/cp+f5I3/UX5FVgmn
HWy7iMBHUefdzAZo/xtpZjS/f72DtQasOYa1q9Nb/t/Z/Q/o0VN2FBf6XGUyehs2
FcDH/sNOA3l4DX0TtA1yMyQBe+P4IbaQOs0KbILw+tjPyLKz9Vhqw5VSd/zTB5ef
NWJo8cXMpe4Cre7474xazpXTl6cCbIokjtaBUxZ7pB5GUlP0YcDNrR369xg3DQMW
h88CFs3RJD00UZJSVZpnJVrg5BekVXVAGrtnTp1SoaCI4oIZGJcvEGsbP2ZeWEMm
HEPXCLYeg+gE9U5sJnkc5iJywUFQQgq7f+KvTRIfTpXYNsIQjCdYppj6tdloQBw4
tc9/Edx1ec9jmjbtkcJsk6ubPx+V4Y2NMLjfO+CCgPVPFORdadYQbYTFDXfS3lzS
EctkgShDmsZZujpwJ92Szq6vbFt3tU3UuFii+1ZiCS4pS5uYvBTn0/0K9P2wc9m0
Zq9jQT5wqJUHaft+qsJFFxZNkhyuTIrtwDkMzO6w1KwcwlDqx9bYOT8H6JaBh3G2
OXrD0tcCTYfErp1ipWQ/8bIVCRmfHftfRysvVhfUUQv3+43eDv+Acuec9Iz40Sfs
IxWMO5Ziae/ZUAOGfbPujL2qPDeQtLevKDF3KFR4g01e68ZW89j6MN3lKAJR/JaZ
n6Um/fJ4ZTcLIEDidH0YZUlA3QhH5bcdvvSo3rLCM0Fx8q10Lr0TsOTWeyR+BDvZ
KtwshFa+HTTqGm1A4rQ7TYmXJ+9K+F0Dxz60opWpkSZ1q7/w7DbDvw5bg/PnpdRg
1flPaygOB3N9YwsDGxeHEoTr1Qlzc50L5pkoZyHguOJxS9uatNP92yZdgAlBm85n
9Q6Howfw+LhJG2tv9Rf4hD3zcpp52nvf3dUy9Du2X7Z31mXBpoDezIuBWxdManFa
MMoWiTyvQH8zRHqxgTjtzFHgcZR/eYXEOhsWIWBJ8hv5xnBm8W5F4z2AjzR6AIMI
lPrAKWVhCxW4VneRHgBOsLn/x4I8HK8AEvIJHf+zQthDO03h01Z21PJRvkwca5Pt
bumHe93YZ0CTtW2xqTA0a9xcBMpqngVymqxE0WStvfjCwqjpIXZBwsRx5cvA4FCp
rnD14rWqbdsiwlD4KwhGpJAgzXGNjuBMen6ArEQWfRdma9XieyxN9AdEQv37q2du
lNS+YQCCgbdaMPLB+pO6JUZkRIwUKon33TJ7BBYWWeB7RHJ0YXN8RzV0APxWEe/e
F2VonxfAaGsG7fdAsSQ0eWWlIJGYFWfNQZvfMWTIz/faeUgT+VueA+cq1PrJzRLJ
FUpMNDb6w4Qm0tlAif44tFb+HGi9TE/YSMPLboKE5+HQpwmIfYBxwXgEanrgLG0E
7Cp66FuwxWTl4YE6AAHBd6Ysi64AVhuEuhDHe+05tOePWD3sjQt13xOBO3qAmWPd
tRiWggUFXy646YCYdrvrDcykdPRwq3jOmG2o6VRl4LBXrMMMz16z3UOoV/UQiQzu
r5SszsjEdzsolgaDwyF3wE4Cd6FXEJ3ea8jatEMhwyLW6i6QRPM7lRWhwIYkK4Rv
AYA+Gy9l+MxHrcsB9UaLsJRomEkP/+rN+cuBeTX+AxrKTnHBd3238TjZW6834tgZ
wU0MYRciP/jML2bIn7O0NuAOuneqpFMvP1UE/bkXxMkHcqRerfSy6CsALjNhe9Z2
wRumt0Rsu93leENbHJ3ppdllPEV33UxD9ATjfaSIIsCf4Cquf/Hl08nN3Qi898ox
Xr3aFcwReYxDQpHf/c7NZu1d4AQiajqqzRtlXQqUDgiW7bCRyxb72nKSUktsznoh
XLObl1qc946qP63xYp418uUQOVuRGp03sxbw/4xRp5Z1miK/Y3T5Af/53NGUpYjp
nlNbrfoUCI10G3SLFjgQGZqXQNQFGHMyjYibQWFXXcMgoSu4B8vvSJ6BWUImlL2Z
+KsgzXJNZuTam1L7J4feyMAL9qnKvqNQlcOz8/GSA4Vrcc5YPl8yj6UsjjSHpi58
d/+/EnxMotPQCAjP2EEpedBI83VGX15j7ApYDD6wMhtAjWcCBKAsvjCi/u/8TRvs
jrBlQoKKnV0vFVdKveHFAgcfnmXYfLzdYf/ya43qxMrpN8/gCh26MKEYIQ4puehR
PN5V9R2/jql05DQd329IsY/HxXuAUdjqNZJ5e/+mt/p5BQZqeBLV7R2dXcGNVyUF
9AxJBpQW6nn1vL0cEHOMwV/gHzzqfqTuAiGqaDizGobkeyEOahGNX07AjLb/j21y
GDGSUeKJhZoNFWt4X/bdPlAi9xdpRp5k8tddZ5kunIoUAb1QBs6ed539PvmDuR/E
2tT8I54ki8l/sHFnnbmZ+z9jIOgq6F70mGAo183lSyZu5Pw9GPreEJYjZIGMGSrQ
ewJ4btKdWfV3f7rMHlTwfJm4dy2AhgcMNmQfa5nxpeGG+Xohjl6/ExsV976wX9zI
uxphE5kjPFEuKzOiJGHw6vPN3AevtqhwJn2JOZb9BsMScVpO+8aRwHXNIuSNYyRy
8D1mRyesWcol682Ff5/Sw4vIqyvplboAJbPcBd++4XjtIgeJfq3ydevm/2YhAZDx
db5kMyNVWUjI7yoBVbp2BRvbP6DNt+kJF5i6bhi3m5F4iSG4Has5VO+2KhI0vT79
ke/z854qq7kLTVvdsTiE7eJTeDh5+aPgZPEM3F7X/mWMH8U5okDn34cLXSUQmob1
NSWj6bkbc1HtuC5COze/DHfQ+1hJ4qhI7B1Wzv/0n+xAXXBtH/cNG2lZMaB8c6kn
7LQVOr1l4yupm4rFGyUvTsEw5RAQ/CUdDkWoI5YJbXEN7TfywXnpH4AkMJhxfp7u
NQPYty8+5zvrtKB6wvxNXv18Ykre1zdmrHpTIIzfXjs9udc6IclIM1rWVuGwzTuE
lUegOFDiOsyq9LXFbmXWR5CFTXexEJh2I9/XyKsJy8pZUz26xQ6/S18mFjRESXoT
IZI60R6J2IJjXvrMNNQ2NFeEJyxFw97/0A2N31lin/y0kqjjb18wn9Qb24P+8fFp
qfCjp0B1jlrGo0YmwoZka61O62VbqoxKsDoPweSI3GgK5Nqnra1xlUlCSEdTQlC8
RzlMYwwo3WooIQeXpLJj79MMdgKDYLkR5kGHtjDX129Zq98X/zZB9aEilVOV4ahx
vDY2yPujIlwA4Iv+Xa0wwYubroxBpQp0gl8skWF8mf4tMOmEt4eljD3SALdhODti
dqxUM6kDoaojcnQ7OU89IbCAdKDqi9tIqKrcJCj9GrZixlV9g65OMFqxRouoEKAd
rvrGmajy1KMAKTT9i8dUj9iU5h+7ZSgfEHV5nwnIAIQKZlPLu22ppEoLxYvP+/cz
tLMzTcZdyqm8NBXmd54XSi3v8iLGjgx0NvgCeM27BrgJ5/QUABFhqFi2WLty1R9J
D6py4fi4SQ4ylECoez4QHH+5rvoD8Mg4WL5aagrkZKqXg3UErR5M5IJ6OQlQqcj4
UnVXrpJBRAa33fpgCxjwozkUbJK/v9XUyiOx+/YBYwPd89kTSm34cX+7blGAwQNb
HwQNpGqIbuIe6n1EnUOeKWVYiyZXP2DAxsBSej0Fcq7F30Z+UbI490ES7tILt5Sx
EU/xAf6DaEPMD6dLsxn7JzjibW1e6T+bRifPTGHwdi7IsxqOs4KeZvtX5jENcZ0T
EhYgtb1qUBkbjZc6afKFDlPfMDiQWjZS9pyWVQawtLmUbtI6VaakasFsVzzs5Rnf
98OKzIX7OazjmR774Q/kh2t3LvgY9aGoMAFiWyCPBhsekab53I/7iuWfdf/g3C9E
3aZaee0GF5wqxWX68MLbx0UbOguaEEOnVbJ0/pTL9+N03JNZeM4pHnW/mllac2Bt
o0ne1J6T0tpIgNZ3SS8M0NV7MC9gsdE8ZfqZI6KByA1lYeKnb0bb2UVC414Jib0j
Bz+6SHB+9dZhxXUc3hPWtstP7WoOskUBJxES8Dwl52n+qJl7hUEnDW98uTg9ZXDi
sVPd6I1vl/XRKgC4iTrNHU6gVqZ/lstRF74i+ulumgbCUqXDQo8YAXJ5jSns9d63
FwKnLJlZnu0MxCY3Orgxm7X6OjZ5CawjvFU8ix/Y4DY8BIh4dlPbjPjfPNnYwC18
NAgWzS07P5U+PctfTTUSyNoMskHX3NlmF58TOMr6/LvSvDQgk9rnLCEJA33lNU86
JLb/gzwFzYFcf46Gj9DPvns0wDr1Uo5qbT2Q8al17BzPdP//WOcLUvsY7aaiPtJh
6HTb29T9GFoYT0tA3W1T5KTIzDMK9kuvK0Qmd4wWmLqTTSf0pitIAU55k7Z0tsPa
RSaE+03TmAKsldIEvZPUoVr/6eczJHbX45+Z/5hsDGJSwGLlvmEUureKaTRx4J9n
hHcNphKGOF/L8xobOxQl8/5ChsQd+HkxJIn8v7MW8hlWussoTx9x4fS9UbVy7OnG
PLAvFzBdP5e9ie3MidNuPQ5ASdaTq1SoDtJK2+xgRslN1+ayhcfbqedh5O1GfSaS
ovjmoISZ/5svhrZXG7P44N8FcES35YI6tdMvdUw0dk9yY6ssnkJaWKhf+te9FBfE
WiN34UcB+JiJtN7YNHg+QpfR+/HgfLlLtgDp4l9ELri4RXR7iYaRIqA25PFbjyJc
dXlU5ntZ72880Zt3YeQgaFajQ12ZsUyfzbDmdc42iN6COfXR6Fph3hQKn5Hh6rYz
60E0bpFKVOWK9NtCS6ESfVZRDFu2sKMN6/AmrqO7tg52pLYiKQKXlJzG7N3RjnJo
/67itTdZEFfUrzs3HjsDaNTn0FS+8KsoE+bjB71bGWv/M/V94xqvyNaoeo96xo/z
+QxHhgFdPR3eyCmoltgPpzHdHUgNLA0rMtZDJBfuGOKbJ23f6Y8+J48cpSMIuOea
NfsXyIoQ+C4BT0Og0B6mfvnRpukQBDpplhZCIUNIZDd4SKYEnrNHnjp8RMI6qvbp
WDbEreJgxn0n7lHd6DF6A5DJBAUX9kgilIqbiqgAPJIKCSuah0y5PFuSJXhQuXNj
2m7WUdhpN/ibUaQxLa4UgUeOvIEdxqZaWu6oanzVjqWOUTDsrswe+bq+CsgMhlQ/
bVBJRPpB2bCT32gkMMJuF9qVW6Q7QEaGz4qnL4eJBOOD93hzaPjMDwtHasMg6C0B
Qw20G4QHDHwwLSgaIIEbHxFsCZixt1CFdpLEZH9K6HGMFw2VzRzdkcRR+CmCSlHe
HBEP1kxjxXaOW/Hy7oiDuhlHtcQg0LIeVTxikWIz+XDAs7NX3Bh6zj4g1IjJQuZA
+YIfVSxPQo6QDiTgOtDfCEJpDQIdQsmJSadNxLNqSwVPVJJMLJoBBbHaQGgGwwiz
bBMNwgH37Uw08mW701sobgd6BHFzT98wxwB3ktMQrrLbkwzcfrm3OiInR/Sv5GsJ
aFqY8MrIl2ge0eyYu8Am6jY9+h0yvbVLTCjgjmpAnBBjOFj+D3UdknE64g3rQL7X
h3wwnUinc9mOtyfJWS6j7Wp8+8nem6i25RpRD6QjMtdEd0tYmRYSoKLgznh0/keV
msXjbJOByo6yXU4SvX8m1tLBkuZvQpZ95bCDQa4XxZlu3faZs3ZKbch4FjWLfDr2
XzQ2I6ab72WTZwjZG0gEIlztmP8xA8z5pINqPHeAoTINnjExc52tKbLmUqWEanVm
CnxP4aZGR31A8/TzhG0o7LHaLJDgh9ro08fU3JZghlAovG0g8nwlm+99yc6yhk1U
aehONP1v8Lk6me08NsDebj7Id8A5dzfXh527MOCRIUmY+tJ5hZ7eMfcdF7Yg8jWk
/UdpdRrW0JGrzQN7BQMMC/ggn+ozjqQlgg9MGylOXlInWI9AX2TGaleuaj+5Yqou
HyZ9SfWtnLEZahC0/k89SkcEJJ5a4np/yvdk/bljFuRSpchgmHQmmLb2YASoELcx
rsw0vJBm3j2N0RA/iFqszQx4jNrg/CmTegaaKQRvV2aY2GzWRtllUVa7JEjjAZxz
zrBTDe3LBnFwTKvIJ2BM/Exs9OOtmkH/HiPbxQIralzbtyajERpsqAoTXh7ANDYb
BR3cD8IVJvsnOqiZVCI8OdNwQGmfFXOA2mK6KypLUVov+8UPxVyX+wYojnz5DAfJ
qBsD7wrhg3iRjttzPXIdVMSWVEWsAzi1Pdmk/GrV/39Suc+VHpIxDm7diGZy763A
CfFgiH+ZI961xT7ksdsxzG5mNsZwhOZ0LWZ+CoNtFEYTjOrMUvylCAIehdmqxXZo
IYvNLFkl3oQkhshKNqOhdq/P/ZE8KWg/UjmNsXzB0f5NhSu2h/sDZSzjPXgyCu63
OfUQQptikcoJQKk91vPU8BotPWYLP2QRBDpAU4IfFIyxXcCWt8kZiDDwGgt5+adL
dnoGNXA+iWvvcT/MWz/K4CT8++Kd81MNwvz2yCpLdS1aIFNR9yaKRRbapq4FkRcL
YTxq2xUt6pFGsILhpyw9r21kzTs6etCtlZR/DsFi3NjK7Qv/nMeL/hd0mgn5uUk3
nLNMLb1eCtLa7pl9pdIOdkS+3Xg89IHk/RCXjAL6npsV9+Vq+9G/CQNNYEetK8iN
6/ftrsQcicToYFqy+bt9ccHOTFrST27CeB6Gleo5AJMmmpOW30+EWiXNc1JCofC7
YhyiMGxW17LviPA54KBm0QuBeqzNMj6zlWVCC2+AjJnQOWN03291UlAwPf5CTAZR
XRfqy6rYaAklH8TOGUlFAj1BrDpnDnbVvACqrurFn2YnlsW3YfcmZkfiKVgXxOe8
EHXQsel3ui2ujbkeCp8b8gKhURChqXKomHC5dEU6kwzfxMpnSVsjm3wsXRledXzW
BwNpAJxtrFTvIYkPABze+Ayc8BuzCyUSiKhZwxvXe6Jo/4oCnjkdH51Bh01CcMU+
7YFwSLnB/xwIHT0HsX1sJw8oMS7ywsSV5obNRMnfhkGDqxBZXDBfBGeiQunG7TB0
eo88RKqlhQTfI7EHmo+TNH9QUF3uus/MOpxFswY2SAIi8oqtBlCTLYNzqUePZjjt
hQXmogwf2r5RgtFgHbtp6uKuujgAHDD+vX8sWTkOTsmStKzNGdJex5JAKmCUy1HM
Mq9x57F5aQFYaaKfNxD2a35FYxbn7MxSEnsAhP46XyDxmeHU60bkjw7zepQWpKBA
5vLh1p8G1JNTi0oR58MRivUuDcGPsUkmC8xS4kxctWcyvjZwZzcO3ufcHNaZTayJ
Io8uXbMsMBtU6ryYzTy/p+yGFexP929SBRqHzXUDZdBYZHdiMWT6AMEhHf+sMGsB
9d8jfq10wehITa1IavdnPloslV9D2EpeUl0aaetuTHr5GGOSNWFHDsgeJTAJlAHq
CqGcIAwXERvqymRP3m36vCCeEmhrr9Yc15/yjI1/+PDMyFB/V3bpK6reYNfMIVZD
pcrTazR8R/ICa0zpUSHzWCZKHjP+r5gyyBtYSO9amBb5Po4a7In0Ebt5AwI6apJE
g2nKlY4m3BGQlkb72JvRj2Gus9U7QOjjIozhgA5bTAYqW+SN2GGU+VR4SjgbMCKC
HIkFePDayPTQyYpcNpFGMWiwevXuymRnRpOAqD4iwxQiRk8voG6MY526npeqUi08
hYi4rffz7tlMJnl/EK1GniQbXHw8l8HrFKmR4/FbxmTT9FNGVbce9cMtGvQpilPx
Zg4xmGMmXFmaJ+931mT7SSu667qY7LPNUWZ1qbOfXBNYygiLJ/aREbEdpZPAngKC
FXAfxir50/54ImbIaf8q/hUu5M2Q31H7Ft84pdG69CfoY7rEcpk/0PkKpgr4ISR6
7I9VreSJ+GguPLb2SDaTwE4tVgOvR/BqKBX9TtEOSE1xuxwX49pPEhh+y32y/pCU
wl38hhRT6w3YoODM3sZ4PfxbiraQWoPef6m+Fr6t//d9fxrsLaJ8EJ88Q74E6/eu
Xq4CoRucMOPzEtTbe3m0RWdWUQ9Is6r5DgAEgyGoIUmv7APpWtjz0NhuW/cEFpKl
XIWBMx7GNXmxlEfgmCaFdYsZyfn4uIhENpUad1gr685551kCIXcXNQyhG9OLOjKL
kwtUJ2mOOcAW3QbWalWRj9UdbIIt2jSqa0GOMOZxHfG4s/iF4yOwzeHKJo54fpQb
JYp06t4lH8Rn1qf63kHspn2nG2vKXMFrbPI1lfC5DOQeM6vlqRa61SgbSquM/zOi
ti7M5MEE5fwLgllV+zK/heDqqwkHKffbjWuysZakFBEQYw+SGihRS/qXTONeIzZo
IP2qD0v3piIpVPO5zrD2boOClKFo6VGLG3kzXTTtRckaT9HCZJJreHUdHnxhqmAc
11qEr1FPjSEHCU7/axxHILLSucHwFVPRa3PMSUzplOLEs2+9TOg2dB/m0rgTwWAi
tbnfoTxTtPJNNmk5x+Evk74PKFh7sR0rluvGHI/v0TLuewqrneHDC6sdM6ExfiEY
9dPZ+axLm6GEXTH+kvZ+cYiTAMPb0MT/Qg2sRTFRJF4PoAdKvpaCUto4jnB5jIvD
t67LUQ4W4zNGBjkGjJBWSmJ9auKKTrvO3MNHhPfBGp6tV9cXGoqaQZ3E07Z5XpSU
vbe0xNRw/IWXeoUZAgvfJppYQQZuTZ/mU8VqJWdmQsuPT4AcW6lJRCYN8s6yULf5
R7Z6EdtuYRgWT5jpF5rY48YCiMSZLflbjSEMAbOHvcW2NG/Sblq4CW9FjXHyP/r6
YQnFhyqmGe5ntRp4p9YmAEOmWzfKXjhmx/GzgAZLo0DeN+T95C+/0j738UmMt52n
swPhdJigRbuHkt2Lp35fZLgrPW2RdvP/sbWhORTZ3R6pAFOMC1GycOGGwoP//vzk
oe39wlPJjUXuup2bdrBkV8W1/ripVACcUPnI0Yk0VfUVW2W22cGKcXjbSKekorH3
+9zvR3Bp1WIj0GgMGIetNceE7qje8YaypY+YsTNrRRmVURIkqzWiC99DSdVhBRSA
HlPamuSzrMbMaEgbe/wMbWljIhfkDtsouy28jbuzHA5OCY9zyrw6PS6Ebh31DCfy
GpMPwDg4nprFcBJRlqEczOE1pRqw2J5YHWX7rN0w4D5Zo8T2cnQkP40ydQ5xjbc2
hcQFzI8CProZDJ06omwKWcJ93JrC6f59DPv6jtMuekjOOIKhhQJjOjPM1KbqngSH
8H4ZuaBjydwRcGxWO/lcMF1dQTRLl/3qC3iH3LRWhzWIfkioBtdUEtsbwjFTVAQS
HklpoVegpZGdTFxtP+eZaLv3RuOdvq5Ubu2/0PawAEZhobER+19WI0z+PzFqoO1E
yW1o5vO73JmR3DUBUecNSzeB7Va547kE4iVIasbWle3Dci6u1Z8IC8Jhvzk3ko71
AiYBoW43OxJXJEcvhh1h4gdRBTDJ0khKqV+3hLZRnTI2uFhIl+yurh3p/ilQepmC
4i3Widxg9USmWyQx+F808Z+VW2JAhBELJmqtq7Qg7xQY2OUcntuJYT8X68LsWyDA
dUWyi336jbu6JlvH1ggOZbG0KR7oGQ5rWQMQEgkuxhWAcZWR5rdAD8DfgtMz/ZIu
cNF0tiuKI9Awg+MhkTpdVJBmZP3P61/duRP/FojhGQbmpLEkeDRFfgWltoe5F7Ub
6LUlCH9mhx+l3gXzI4u+LZRValn1UTR0LKYXCEW/gX81W/G5D/N9sPFsJf8Wz3T1
vHq27tjfLsmsoF1TYrAo1UJjGZHMwVxCte5Q3phOPALvvqSEzFqWF5HmE7Hs7pCl
NB4ABQbbiWYHRKiba3YgKlSq5uJRC6WDoc4i/TzMRCmvS91BJzJxcfnUUgv/BQbQ
qj79MqzQARYMqNnNX4AR9bVN/YzEQdXamBgRECc6iXswZk5iTmkxjydm8EIDHd3S
kG3nftwxMMx9mayNNMkA0UPA0bQqCho3CarEhe0H1O+OogolXAJ44TDXIKcJEm/e
rtwqAgpRkwAv6ReKvNRwmaYamfcTjo0tjLdS5259cH5wBDon9QqFhRh1XnjTlw9o
nrqgxmicJQNSeoIeccoYRCYQ/pgvnkthmAWI0W573fRjpnZwtHuJOVzl+uGcy+gn
t0RDPZsLKzSRmn78QszuABm+Y9rbB+qhsr2rYW8b/4tFsQgM4cs11wwro31ceX4o
aNM46W6t30pDF+vTNWWbJdgCjG/T/P+xR+8Xo9uR12Q+hseBt4cyBKfc05NOLzPR
wcKQJElKrEwbO7+e/+fTxoZKJ/e4s39iCgIvDlOrCbDdWrXy9O2P3INuoQpxOezD
FTL3pDDwC36oyU47ErmS1Wpm9zk1cn+SGKaYDGRLOH13GFsBPMCf8MuQ93/4MiMF
lC/juyOwoWM3BgJgK2aVzeII7Z1xxqCYgbFR/UAousHPAbWV9v2qSONlmht93z3O
/2Mpl9KBNBimMoi3f7dXMvvkDqPKztZa6sIkpAiSBBWqCjXsu9pSOpaIbiNaj1Pk
rsTF/N697v9tYbdj+anWZ6OYuytIvjuqLemGlOE8/SYVVyk1YuHEL9H1XkUN+l8Z
DguTxKgvecq6lCYbeOkCtXhBxgbxP88NSNktPBfL/EMo503lBdbXt7vxiWdS3W01
aJpuDrLE4wcLa0ERp2ZhADxHdL9XbaOpAIN/t9wkIB1s9fuLFYkeKEMIaZqMBHQl
2mU2s+AvCnuiJurwNlE21hCNju79OKrDswgeW4hOXZajRDWFG4TmnfW7xtP/aKls
yedg06YhfcLhimfGlFrJH9lk80Am5YiHXsoFh+dZeWXH1kpBnE0kiRB+aOnxlPM0
klKoBJLSjl4TIEypWeIqrhyfDFqT52deNriUq3WyASpfComSTt3/QNTYqD27V9eL
yGpmiCd1+EfRA3LXxKL4AZOM8zBJa7bOkd+/atkuoECILMMOeMXnNB2EYGEp8wEG
7mQOe3pezMwSHGrGKz+JYwiSmZQk1bLLtIiO29wrpCqpN3JV5fIujWPF5ormq2I3
x1CS/BYGObjt1CQUpWkaExdrn6UNf4jD+gC7eii0KlhUgvaxHrirRU8/8dc1i8Ph
jEc7c26wItAK5zYnGk7S91d1Kkmtw7/FllnS2rPCNP/DdVuD9iag3dmgP/72Dx/+
/vBT9gFg+mT+hd2pe3EOoVBO6yICTSBvccjyMbw6cejR2f/zjDgch+hgO7/ONhNl
K6nAjM78YxCgwyoSPJ+kYlwAYFcPJmdOIv7cYfJ5pv9pBX/bB40o2vLoPhZlE8Ne
c/8MWXAdykQi3uDxOV/lBRvmR05isny2XmrMznSTiOh1tMb8e8AnjQWDbwPVDd1o
fV3BXIo3o1tbNlbLGenLAIqMU5d8rMHMYDoh3y/1XPP2p+Ua5w5BecMNogshibGV
2UPZrbSJuVdKaLagCV1uDBEXSL2KZvXTUNFabYidSt6u4M6fn9cOf5/2jCzvZg2s
d69vA83GJ7pIHQFi3kYMt3ZVXxDZGu3zbu5mQKDz/a07OLLi9Mi3f8Oo/EM8mmVI
NCKh+w5Y2n5LGZT3Kad2dn6388aidGcxrasEo9a2kTYI3UulfYKAMV9OJYs3cRxe
u5suYIqxUvoDY66XaoUUWg8IaWh3cAwgqrYdXEB7GM+Hn01SmjuTiX9u0GCbfMGf
bpeXjyu0Gm1JVEEykaG/rCIUsyHIdyXRaOldCtVAOC0I/Ktl/hpHYWpFD+R+PmJt
ZpFUUJiC6dKhQ/vorCMk+gbCteB6uMSQ27KQB61/IgGuDMjxt9LvTDJs348+GUmT
gK8RHSTi4kHj6xjsh7kjEglgfu3FIu8W/VqzgU2uTnTdxWSlJiYAYUsBmd2WBpVp
Vm0Ulfn3tEOleu1f8vY4Oie6px9qOAEVyxyDbSauJdgGIaAAWNPOTIjjIDSunzCf
fgrOruEpCrstinVeZDyxOwuu0zjoNtjv4cYz2wg6e8P58HR2KqJe5LNyRDxc1DdG
fm49aOpt8pTJXXKA0x9SGsQfSaYHpuCUpR6WwtXv0DKNj38hAB5fXh2eiizTn1A9
6qCEod7juAJOpr9S74fiaWeoqstEnwXCNrfGxyfbokwKkPk4+WEbr8fu9oaBFwiL
CnVV5Ej3WCIwwiOP7npo3aH+GvF5deLGhRLyOiAdFePMvxGf1WWYvSReIP1ly9Xq
IJNK5q0GZurRzHorSqIuJm1nIlMzbQchcD33tagJsSs6JzU8Y81KBLvjvGAEz/WI
xnvFXThcqcdvcjkGRfgnvcIfSjkBLJaIae40V+t3zCotamayJ7q6JCXSdjGUMb6P
niaNS+makHx6QYZ4SxEJmWLgGs9r0k0SBPuJgxUQX6yLU3lw6CaHNp36lFyDebSb
ccd83MkkxdJkNz+crEiepYCtOPE2JopB185J+l3m1aJ2GEp9lG8eb4pLAW2Yfi/r
lMJIUMDP7wXYUBFQkg0uz9y2tG43xjDi4LX9TVDojr0CPgryWsawCvLI9no5Ge8F
mALWibbo49//o75UtGL2V9XmWw+aVyUdGDXBDoHJWtybBmzf9D0ehkB4hUfpQhmH
ZZluLWvtPu+0j/z8LX1zDWYnbeMyraP/Tpmt47MLLypGRJS2yphvSdIezLg4Wx7j
9fejSfzDXblZovDQltyrRV1SjC+XxgS2CDsvUlrk7lnXy3x5DrU1+lnR0Jx575XW
g1pjSO6ubYbYpN7ylqCmgPOtunk5SfnJPdLCxvHC/R4r+wtUSUGSpmKY9iIEG32c
3dYI2iseXBDVB6dg5XncMhkdwkhpM9O+tuCCckF4wxmC7k5XtqDLQIB2xq1h1+Fv
rKpUo0Le64nNCgdPemdH2UxYXJ+J+QZCQCFZ2CAuCqJH54SMrf6A+9b5AhhCxd26
mfZNx2LpQtX9tCCaRuGN3X1Rsi+3qoV4K26CA47rWfbq6xtg5jnJf3O+3loLqVwc
/QpvlClabhMXQE3skHAv5/Rw1js9xIbA5wYWq12Jov2uD/TpYl5eFbqA93I9anv1
iHrAVlY49Bt7Lyh0/8KRbqendx3lhDfmjXPEqEdMAOXReKqk5XUAHJNqconbGG7t
F2C0pH9uBq1EDoKKWHRaysnpX7PU+R1kzfx91/AUE2fd0bmlOuG7udDnvP3lFM9R
QTmW/9q3WMChW9zFdtqXzVDZJTzpTgcPenJEXtHcEb/yQX2kWRHziJ5HjHYBV+qp
ghkKTJ4Hq0zX6O/mCFu4viQYAYKtolgn9K28xx0B5XLV1tWJXD6utSLJen1aK23N
FjO6zCidQKQcO8Y1jV/dSj3PJuUHdVES4ivXSrCeY+t6Eg8WOXzcsJq8PyXJznqJ
UY3Nv0frXrR3v2POd+99lIT8SPq/4V0yf3AsMm0ZtVZV23nz4nksMWOeI42qaIFt
EE3kbq97fzG524QZCk2GvjvaXIFndypnoieFzORRvT15UQaX4Bh23/NmDN7nnrHI
NNo2dpk3kzglYtVYMjGcmpVsx0eMYjPJu2A368op9NTwDOPbt6g4JRcM3PHfH6PU
IQLhOwsYfzQQ0rzTb5shLNaWLjDhmAli4cYYn4OyDZH1qdutZveFp0qGYElRoeAW
5pQC4n+7lCZlf6uqO6slntPtArJW6BifefpmyLZGpvCUOj/ZeaNlenv0CmATfrEW
0oGGG4fyJlF54Mlsu+PwQUyXfCzE/urCI6mo/u2eOz5oREBFAPSHed+XWazmfNL9
jRWA/bP85Nyb54o9I1Ljm4J/xK0fEhBIA+Om9f8P+2ceoZ0oezTadoGdS0lckV9t
qUThryoHoUWDlLGyB6YkQN6R2SzcsP85sMhMksuYjMXJqhKUv4t0T8hWLSmwscub
TJq8ImsMJi20Yw1Skj3BjHWuPRYTZvWdScRornAdRsFbLatcOKngqsTgZm6V91gH
Pj/IEPHiXVIA4c8Y09XfULseY4MnUBxJH+9XKLVyuUhqbHR0/sdPm3ijICxKGcBk
f6g5WDZK/JiubRlKANXleaVrzgSRWP7lxZR3CQD1BeP0flvKsGgPHTRabSX1kn0J
uiYQAAssfFEGgzwpoVqu9cIYuEcIHcYk8w27d0L6+9nHt9mREplDu4uzoRax2+1T
V7mULBhTRNCgISLFhasbnP3GcjG5dfbJmAll8+T9VFSkTyKe5RpPh2Ys3H4DJFCa
mKgyH+fALjk2/Qe/a2N/BWXs1Mf+gsBe4RpDsf8/rvmq8XYZLwL/jfzxHodxVerb
Am0ZpVLTpSIzGhO4AWQqGk5lIhx5+aBr/KIIpN5kxARTq4kykoOw6UAFauaAoSQO
rhLxMgKFjoVFh3a9282BDI5p26H1QcO8NqV0eJL2BzwELc6n2Y6vQeM5DH8nOd1v
frHuaZJ/J2HmNCJvk+zioYLMR3c5XdQR8x0lXHA5OqK86x4/9G4yT3leNUveMUup
BvGKsSEYbvBF6JpGFbX6UUouvseqCJxIKBWHiBVKA4YvoN3umMmX31Fdq9mZqOYh
x/n1fJwFrcrcKoWwFEQanTL5n1hKl6R+6NOSBdZNdCeP0bQNzezr2gOmBGtlNKpJ
18jY5OTjejiun7ydEuXfdczWd6OXulJ4xC9ca6XowIb9/lHBGeXObtEoQW1Hoip1
Wy68/R+CELo8pkrAhX/iQ+BCTCKoixleqe520HFxwPaBE9Ox+NvYEusORwqa5k1y
12ryiP4TIJCJ2WayJnnOC/aSz7IvTL8mD++CMnSdvytLxrV+M0OgxyiGMmrDnVIq
IhsV6jgfGuU+XB3B7LifrWR1X6KlTFwY1sUqFSjSjZoTPqHyMCDTPCRYmyZwrG87
QJ0iBiHKsT7NR/ELorzQIwKCQ4+zD7yvecP/V7B28pOEInfJvUO+uAAnF31WiVgb
R7wETFkSapMG5vlC2xrZkzudcsNEAD7iS7mAC1rFr7jHn0imLsgxNIoAR3CV0QSd
E+FTYr7aQkkCTIfBBL14Dy/eJ5JEj2gvHFwS8OAUm0r9Uh6DwOopPEtB2mcjASG7
jSyE/uLKa7I2WRFo3Kg3D9C6IFSIxKsblqr7D8GOeOc4R4wuij72hkGfGnSBHrhy
OdYrd5kJ+HWDT4/78JgvaOp2LK7wfq+8or1snLdyKyF7fQVRzxkUOpvjE/LEJ/AZ
E/zPmXdDXQgf2kgLmSEKDvQfcgBuPMd1szRG4fwnap7p2n++Pz0tp92dVjgeT6xW
8q7ylbSmk+3x2VbwXH2NPLu2rt8FyDqrqVWsgYkTn/dEKUXF15ioCKRtFKykVPI7
aN2AhLyAUHApelwlMPjq1FuYuQjgPYj+GR8aEbTOAciHLNBOqTTL6IGY0LCnBC32
GaaA9f9XSk68zz56wOkjF5KZ+mYc99e7IvJ6xH5Qua3SFN4aqJ7LCxiVV2RCjCN7
WWTa1b8QwwvZg2Jg6HNnhYehllt/Q89urDITW7q7BM7hs0GrR5WtsOiU/raZuBE3
/2g9QvtCo2+HLiDM0LGJR77Ux9hY0CGhISnZKoc5Fsh0/94gcf+tG1TH3V/XMDN2
m6yYbwTE7+psVUxaNfVKFU8QOhPRNO0kospqnBTuxzHc7W3D+GTt3zUwzw3mfKjG
yr5nvr03W5rbcdO6ZIJ1FOvcxvQUxA3KK4hv8r8VBx4Pp9e5/GmxY2Nn11Jy7++J
c50x4KC5q2ugue47S376cF0yZjlZpLRZNCSGWgm+1wx+X7ZnqUfbpwvgDKT9w1hi
3RjJ1ImDQb0UkQlKdRJN5FDtxyANEwQaYCz0P1iB0m2+8sD7XmhrVv16EeVC+vTD
nw/h/VRGDYuAwM6bb1r/zek4f803zt4QuSd63ohAVpTpIt1C4XM1gtwaUcjNUNPM
UrPhL1jqmYtrNhGgVlzykxlyIyz8BvKKP8ottLPsjvq8zbKn8BABSI5GH82XqpyF
O6CoCug8I5tSph/3hhiCbIP+1iifviptTiSkfD59eIX1NuMdUQoFdM19JXwf9N0J
J2f4aki3CMlRnUz0SL3U2tZ1zEWSjJlCKYDOXT7ulTVbApCLUVb8a/jwqL28nD0Q
dbJbvoNY3hulDCzq+tt8cJ9m/aMKuvnOmdRDk4RfWtq5OonydAvLBtbfiNgH9vKb
1cqDcCqt3XvIrdwatIgvqV1t35//H4dKqRgH2Fb9FIVC9CrsiYJtFXvsmJTJ1STk
aF3LBUvXf+D3OOwhLvXWb65PFcoTmaGczECGeY1e1Dmo1ztOZ0OADzg5/SA3Sas1
SNhuN7f/NjvAgudvGCGlNnMMKrK8dnKFBliWCsSK3rlXWTmZTF9GVPWwm/y0uCSl
iQCI9uOpe77jjTqb9vuOl+T8kc5JTttl8DSFsaKzB+fh6P7QkxJBhiUDLerhCntV
hYDYsX2gla8j4A/6gOewDhdwtyn6ucbn5cteFY2QJSnUFHdoYhBtNBu6HCVr6gv/
fk1b5famVFsE1kMAjhLebJeS0sYr98kIpZ0e2eDQlz/yBbKaiEzYqf6dkVlUhL3E
v8qopg5ieRUmfW0EWievzXddO7EfipPDVP4GsjRvd3LGgTSp5Y1MnuqyB/rxju5u
k+7FEve/hPWGX11Be2We8FD3UXV+saaPR3Oo22zrTTrscsANnPveZ+TdUAFpaiT5
AxtEkf5UG324Hnt4sFAMX3aRW3sLU51dcs5jrGVE/QjB6lsUZECJ+D6LSLVuGHk/
LqtXvZFtaqqZKUH1HY216eKYrKh8btPay5tWduLMCshl7LRKAoxywTg/9n+/RLpG
NnzOJF31pQQ/pG1A674wLh0427bHnESbaHESv2JHpcbZEAx61UkoNlbugWk9PXld
jcHNAh6XvfmIfND6PpAFHiXFJg5Ve4FuCueRlje5ppc9BTdPHq/5nmANCC2TZn+c
mhQlKmr/Kwfm4ATqwPR7Vu9qmAYYswlsWi9tXpnhoKwrH8/8g4djFpYu4eBQYaaT
brNxJU7evUg9gCQnzJanoOcvXr8KcREqALtTnH8RRHfPJp4uDnuDrbye55Ry+w7/
91nUkGnW7Bxfpc93LnYgkshUHs29g3wp0WVkU5pYFeFCwfzkMd/uEbKkWpyH8tsv
D4gPqfVxNZ23DSa+qHPJUXTZITERpyr6qE+PPbTWciDI0mPLKvu0t7Zk+08Lozhn
0pGNKDg0ePsMYc5R2ica+DVMOuRrpTzImu3NF8aKFpvKQQb+RMTuCujK5yPRzj8u
ZegzloMl0p1v44nHZnsnjaEdxND6CqmqH4ukEEopaN3/8a8Qf5bC+MS6rn+u/9qf
RRu8q7oZ4nE2+sKOt4i/Ow1e1d6SDOXzWtPRQo9mIRXoHHV8wKM4ylJJ9zy5J3ts
O8BYz34+txfnSVAOjKvMlzQCyhfaPNwehIpznHFknbfnCQBjLEF1JD1lW86cZ/dk
CMzVmSO475v/6XbIjf5wUb5xomLZ4qrguDDoFyfHxd88gPdrufhLggofSE2MJX9+
GkUOykycTVG3qgApc1xvh06t6pPdRChR/G9kKviIDrtLiw7rimQB9SS9n/2dnkcJ
CbLt2ixsjqfKiErTVu0qdtcQVZ315oDU9tryVaf0j1vZVxUfUDCUTGRshFf/x7ct
MhGxv7Q3fhnesCMu+VzOqIn7BWvlO3rG/Ml9pCsZhqTa/3teGIcv4QQI3BeMOiDQ
/E/ZQWh2DRZBE7vRcCc3naaGsp8IRNoEwp//ODolOO/OPv5CKck5qqDx3jCuZeTM
eZsaPwHMeHCaWw09oHlgJ6N+yfu9aEk/Bo8AHIAHmyYTxhg95fNxzv3XFOXD8p01
VOaNDBb5wcY7USXJOE3otP49CBld98yUfAZWJ2wPETrD9shDPetqE1BJfEK90I85
EQ6qAHiMNc7j5BSNDAaIM96vTrPMx+9MBrHCj/OOc+Bwt7kqSS0Oc4TC2FotbYGp
P0NxP91PAkln7v9oNcBOPu3IpU/mDjAEpXzxuGNbfIx9h+EnevHNsgDiStE13DyU
lTwmIwrRLNYOjHwpQiQlgn++WAW6yIFHeQqTQxw2PJInRNOyY6kEXhbO5V1YOFut
MvyO8YFDdWutmAbmsYLWSLZ5cyODMdADd5jbu7UOlEu21JUWG6ucCncrnQT1QZUe
3B3HWSTWQ6UfKvohUQMVAFXgwhIFcxIIAk+xlWaCTjuGTUZ0bB2ZwJL5Bc+Dhth2
L0JyN9aGdihfSdyGsgFuYZYelfXbUZmsTkgacJrg17ij+aIUwWFRBDMPpj9L6lOh
oK8xWZRqSU75/tX02DcmZzDVdUEOCWmR0uKfwZ0xKYdcfsHnnN2pqpvS/ExbTGNE
XIo7D8DQVJ34BLEORe+TraDt6Y/D6TtX835Qn5Ta5QzTqenkSBQ0i6lxUIOZ1Vic
ca2TXjfAIOwGVDUtXTfvZ7vpY4P1tmU3l6TL56yrVlR6T83XpJBpJjr5GczTwdOT
aUhHTAzajis/GE88SIb2hNnHWPTBBaW4vpoA/RJzQ0owiRr7WJ2vfngxi6y5QpHG
S+NnlzVj5ZzfhB0ggeF3mDMUm992C6quq0NatP7OKprBZDpBTI9xLrL2Ae+IJiez
86qtmr7EAEgW8RIG8jf1TbEvf99BuAsCcWfUAN4br+8x2eWiv38JCN7DhRrh6ARV
GLM7rAKjj2i4eWBXDQxafkISE+gWfhSpptrHar7sVaFaZZhTLjaA4xhgXwSLCXHv
y5Nh/ol6PzEKen5Dd8jCDAargfotYQksQxeYUwaUoK26ysavhTsHQ/SJOloVbHhU
xECOX8z/CS3T0ndZxn1urJCHCJ72+XgRB4u8E9kFsHEEp0j+3YcmAP0BUS6PaXuM
PLqeDcV+u0wVth0zMWqwz2wHvFYDvPdntkPMYdZD04VzIdxAcxuwI3bii5rIG1Ys
59FFa8zwS0c2Z6OU5BYTkq9pIGDmPjEjmATRtPBhX6/4CKMujPLB3ZxSFyvFeA8g
70Sub7G7VaJey23+P37x8U7iJ5B59fSUraBzcbyAYJfE49Ia1Uedh8s6kU1RsPNr
dK7JATcO0ucGepMTTBC39y+iAikSVonT5zEhxctFzCVqNQeyWIb+11tw3y2XMm2W
p+WRG5Ql8yIbJhLTnnEq6D3rZm3oNKH/vFklc3D5CgdZJJhHhxkJnwfXNJitVbfN
TeLRn/DHJStAV6QOz6g23MwBkrmFE84CXICKGrD2IfhIxGnhcX8kwJbePfgw3EQd
MJyZfx6frOkx/u/vlohIRk8dEgDZB5YydDc49vgjuw80K4DTj9JOHq+Lwxr6grR6
v4mm0MbAc6cO0ewxFjfvAtUljsy8LgXkiGpSlLZCpuDk+C51soM1FXxdn5oDYgPi
JifggwKjEEI9Myz86Z773RX7QADZrDNfBWPaLqv+ilFQWGrveY+H7232eF4oOf7d
YUGShjO1YeoMGxOv28cYj92+v5/TfRFex32/TuHP/lXzkXInp1pWNv+FGtgO4SRG
Z/f5qTyR2tK+ynQqDS/lhGorWqHmtyp/T/i7jSKhHY5hfFDO4gpiMjn0GBeaasa1
NQLbWkyhmrk/7sjXImXVHyPwSkK5BcoDpx2YeDQ/WU43fJ2GBibfPIUX79rT9qRI
CYGm+N6sR+3NRrQPtnenrV0TQ/53ulrURiaY7+9xmbimw8yeOriZma+MaPl6k+Z0
JaPklXqgmVVxoP9PUNzJCpDC6Xm/SysRuuFkRYgLyjYFIMZLVj3SDJwWTwuoysBH
Z4z7GTwNipJZqwmhvDZa7pZ+hs/rKKNerEJanWWmKDtMdKbG4DW9dzQKOr7sf+IL
pDPfYeHFJeT9xyc/LxlTxsJ2+FF4jYb4TgKkQCgTMO68/g9Ze4VvyI9TsOhBJ0OV
nDzLA2VG3QxDOKC5Ga3qhHetEJX2enO1uQ5OG7aDzseqy6u17aOYbnLCJ0THyiqO
DP8hkBdOzWHO9DrdFPdfMiuwIEVgOmEv7gtKJ5Oo/kSbObI97KqIP8CkNuCTtfp8
IiPG0sDyVH52IuAfbFmup/fBDjCvByZczBH1+OoRjoTprpWXrqYZ9/VgFn+OCzuS
cjhnNHvmlEQvx9X2su+w0q/zknANKgUMtSyWJiMAF0TKTjs0OprzPteGTh4SVavZ
ZjhBbWcRtd+32hJ0cafeJhYOBjmHiVrmppTIoCKOwfvM8FJgukot6U5fqogp+fs/
F1e+cNYapIykHZ0jfwl1FnKKIGA5DsoxM/KM2apY4MAFJLz7r15/qpnPNT/35hHS
/WqPgkgrW4mZ13dr5aZcZBuPhHPogEST2rFGkACTD21Qn/mEZx9gDK6EQTEXPmHv
CWEvevSZhHka68sCMP5Dto58Lrc5P0wKo5hKFeC8j3pBgjWxC/GxVXXUbExA4uzm
MvCtNXtK0K55kI4hTUTbx+5ZbvcM22GzcGvUSlxNvKwY32fZqX5wbe8Nq1wVO2x2
HYjtXryq8TGnIuQci1x2fS9ymLfgGmbbGoVCa+aeb0nBL107yPoV+DTEob+rV+5a
8CZs1r9kOYv/B27k1pr7b0Zt2lV3PkfpimSvTuwoVKn1jAGn8LSICCCaB3x91WbZ
dl63A2Xv9gf+xgeMXIz1rtnntsygsChJRtoO2wDktWwrmKUBu1UrpVCQT2ZXF917
matLhXO0ZlD0brtE5uVfTod2K3bc5N9BW8uQAd7iuRWWNJzcqFGBCXUCWX+IAtRv
aX2sTbNi6rmETs3xOtiv4tGnVUQnu+p2vWJlauQIBV7XbQVU2uax71+R+EW3JabI
Ht/ktuQY5ZDfWVNXCtaDxoaTNE3G+Kg3Kpn/AKv6z1oLj4u0TZhtFJZX0Jo7wakh
4TXONTNPQFtCj+suWhCzZu8TKXach+XESuBSrZGqbcOD5z235MKs/EO/ujDyXGYj
XiHdcyq65Yo+b2quW0DA2Ey4kInyF5fZOlwaRiM5jlKmvaxKsgAHLPiqf2/3wUOu
8kRM2q9ifjO4VbsfNO5zG/Tucz5uarzt15vCcWNdlEOiX4A9B9JZwWcDoU0w/vVG
RaJx8GzkDfWMAboO4511mbYXi/eRwEmZM3p9ns+OxJv2VPuRn5w96aNLz99ND1lz
7X/BPazlXfVYt6h9G8HjDrTNSPqSlO7tAz8SJFdSRJ+jZDD/eWv+uPid3B4d36Qz
qD5zF5bA2Jv4RdT13cfUNvN15Q4ALqlOrEU0FX666fGYYvO4bpsSfNhWTX9pUn+j
fL2t3RmcUxWLCADzXO9vs0dQW6/SV6I2RxuliO0FJLThoU2iUKyhDKPIBBKdz6rz
ge+tpaPRPwkNzJlVMo9wEd13loNK0X3//FWGocpkciTpYQCBUzJQmA+lKWLiJchz
YMMHoDERoXFhh1dX4uqhW7faEOsNdhO3ch1hsocNgkkbxG9nLriq59xSA3Kl3VwY
hU4t97GnwXCnb1PQBlK0g1DTBFPmE65hItKvxjT1rbHc56EUqyX+t0eAcVRXaqnk
tWUmt+dTVYAUR4vB7AR3vycqrpNbVV3YiX/QTOGhv/ND14+27xSwt+gFt+vhFZbP
3c8L3cUSXWhTGlslXrLket/VdKT+zUIEAjrAWttyxqNic1nSxrgiRkV2BayNWyQr
mTpCgXG+/CiMOWoTSenid03VyDBadSzHTs8nRxsaE2VRyY/qTIzkKsZOdzQbAIAu
3a35coHto3UDSVIWILn3HFemWWEmU9apbOayZDq/1Y26Z5paaALp+RNE9MgOl8b+
qE4ccYvuGla2XBRDCesI+buqC9J26wJEqBk05W6LsftTGvtSSwGTB95a9npJ57sy
YdtyKbfY8TriOINbPPjArfdMbq5iazmVDPJFbuyDIUcn6/KyRngE9d+kmJs7xdpM
WtSBerUOO/VaT/UDayJPcuausOFYYziYOrnfGEy4UOkJKlyUlTFuYKAi1AEsEBz4
kCZ32MIMJJmXu4rRAa2GD7dJnfD1QjCEFBv0QdJN32c6jJ+MelSt6W8urw/u1tgT
Gx13ExNsEbpsTOzv6i4AGWWkD/qHV4lWGr1uzewbpn8NNl5jaPIFkot+qgkjRVjy
8X2SnWe90UAczB9ZzJyp2tCJ+A8UsKTYLsmMFifkJJdTTLoYhGSrb+HkH/ba5nLg
wo98lOtME6u/mBOvuCNLQiRqk9gm71hsgyRAjdytXGFmBwAWsdN5bgLUyJU8amRi
LAx9JJxYK5ySttZgvJd+eaFym9cnR1rAnx8i2Tka8/Jczvj3k33OxTz2Qm701z7P
GFY6X+PE2XSD4Qvprax1KQG1kxbn0wW2FkfpOMV82bqRCEUCK+LFyxpEtNwo/bjr
W5RHvg0MVl2AxNTpq6nIrFKafmgi0k6QajFH7aWvU1PMrx9BKeH9hakIPK2Nf+9M
qgeuC3LAdTYHcxg3kq5a1rUTCbXa0cRkbOkDU9ASCMaOY1lO1z79RJT4DD2wBHpy
N39n1J5xeepSlzYwb/DxU0H5XSoPwufjuDKzlUO4YTvkY2s4UF8C3I062aYCsmzR
WtNCZbOFf4v5UXMnW2XRvjqz2Diz2nXcDEF8aGpfHmKZ4EwuXiXpdzEb/NbsmYrU
53s9hkOyqd5CWlE//lYjzwN9HcsUw01nat+CcbnY3AVG4Xo8Nc7W73kDOeXIDLl0
1OjkxuDRTROT26QRajdcP+TNtR+Uby9dzOZxOuC93IqRP0DLlHVchsXNwe4YZxZ2
YDOvk/H8Kw3DoTNd5sBYOl7AmAOgIE6OPmRpojcr/0zRO01srFD7u6zIybWBcNGp
UVM7h07HOU8b9oj0J798QsVJJ42/hFXgOaIu8Q1iqyQYLrIcEy8CNJhIEfMMoX3Q
8Pv1f/pfIQDjTQbeTv2l4UuPfs/IL5qJpzameVe8me3P4u8rKpreNjhktNZy5VdI
AFni6zMTVY3kpbr3/Jchuq6Ha22N5XSX922lE1LyKBq7n95eM8VKzFPFA7CRyEki
C6WAddMZ3n3EYMMXwGnCim/6DHqNfL5lZirjQov7JHA12MuhaXKfW6v4BaWGjsZR
EwQAf6u7cpROlMxtuoTuXsStMLsN3pTU+gWQFs/hloSSK2A1FPfw/1e7n5NeMV51
ykdy1HbSCeRAlqvXJJnyK15aNJ8kmsi0l6Nv8/ojNsdrQ4lV/qUVxRwmjFrw+KIe
RqC1NaeE5H2riSC4O42QUQE220lnkILtlZKrqzZDIlGsyPGlMfDhyj60NVAFGlXG
zQpg75ZANtmI2J/UKpjd9f5PUETr6DFwwSsU52GWuRir7OCy86rK9TmXrmzdrJRC
ZHQfrpIz11hawlCmRmrntndhAvWDQndn1E3zdVJEeq+SpZh4znj5JwzhXblEGk6u
dN+98TsbW5AUWuE8ZNykZORJDc6vP44V/4vOyPvAgBol9PsLazZ0RqdMJTVbRXGq
ww0Ze0HII7vJo6AxGbxLUgkVHYxN771JYfO6WquGdRzYa0HvI2BGbyCM7Z8lxlI+
4tFUqQwlpChcc8VnGDwWsPoN4gKEa95BbqF/Jd17havqLTeezA0A5etDE9f/+zbK
2J7SX/pgpVyPZlKL6GF1NoGI2uWxXQkbithQn0WfFxqWZQK6vfE93h1125OTU+f4
KrjXeicDTGdHOykT5aOgCsyMgRm51H1GQalBNP2lJWyRajritLIlLxvSEpkN+ZOa
Jp7PPA4o66+ji+jefhuD2Dp9sXWX61B2o9etcuMlvhfQw3d9fTf6R1UphB+TQjl7
AO9hVFE3QG+kr9z76puWEcDL0farLSD45cFEWt6pnUCogSq+Kpa7KtJrT5tH2u98
JAdTRiQbrEROXl5ym3eIhm2vU9LCLNGRkUkCJ9zL3EGT27IqJ8Y3D5/qXBiHZW2s
tT19FLezDJqJpYnaBJU8sfqADe1sp+BZsP8gV+xxUyXKa2Gcm36TrTM47Fo5q2rm
7MInHI1/OEg9KSEsQKCRTDD8FLwciNu7yzDsFP1olz22bvdGZizxck1cfQZP5nyi
PLLMs2VdXKuD52RUvBGzoBab8uSnr7tdKVsZzKcdX6aDu6RSq038w599TOufwU5C
EQWYVqtx0E0tWJVZRiYMUpLlY5eOFfg+VoYFtmVBjAPIxk0SqzVEql/UiuH5gMBi
9dyDiZuAp9R41NG417TRcL6qBHbx9CbVCkkzNrFoBpCQCDhwYaCsD30vYlCv8NW+
yVL7vQcrtmWm+eLmNVHgERbxH0481C4+kBxUOkcd/1kPP3avLJ6rxc0cZD3UBFsp
F9HEbCFyF/BsEQSowApI5WPSm63YcQbvcUHXgb+r05D9mmDz70rmZyi0dhOV+FjQ
FZQdZyJbPowla/9dgJee930JruBd9oliGUiJEwLysYgk6ECWFKoDDD2LubVCtuLv
fvDLTf2r1I0V4pT07tw+nQSEN5+7z9WourqPjbE5N16y5HIQ6P9JWiXadfZ0K5Jd
X/C+keLc3OFtSTViVJrpGk/2iz3ZYT2jeLK7V4GoL7mgIa1lHw+UQRJvH4Yz04/b
x686aQggzPA2OrymtU1TYKFHhfcycyOCiZdSxy5+Q4y98Ud5aN66KAfR13zP7sGU
1pniSvNet0ZLz9vNWQnXpgXau3jIf8bVR7dQJjIk602iLwiLhM/za3e/x2ybBtf0
DeRODAauzm2+v1cIacOhkGfO1asryctxnC7KC5YyRh7tZ6DHWH2zKtQg1Up1zyuZ
qWJ5pr3Hr3YgrYqOpM9k9+U/+Cpf6rnKIukyrs3VjLiip6SuvJDd0y/9atCwRR4Y
J+pHmMFDWVBnBkXLtzrjo1IdBhVe34f5PNkmBPlP8bqRFmCgLuK+m/8XSivYDFKy
b1f1ybB+3vLzbGLZEtc69emSivYVfFxcjLLFoYDapCcv3iazb/7bU9Z2Nh8lYDoF
+Lik0nSesI3tXe13n8U/QEZEOMZ0FdPjzRkDW2SFjxtN3IABe6Vw/K3WI3s8oBfQ
r1aEWb6/DW4cBm9vH752gFknaOLyAyZ4w1FFc7xZG/T3rfYKEqF/mh1BN3BSFc3F
w7wijJb2GKPlXdmtBPvidwyZEnI6vES7W+vebRwHLN5uXRqFVV9M54zGrWSYtqOQ
uBT5Fw2+e/eSUXmwhkdOVqIh5rZvS88NR+/XfMm9waZzSctCP0riicxKIzvlvbgS
f4yjP/GskzJybmKAsXqy/kdoo9lIMKDnzFkMIZeUU4RBz5sW4K7y6yILD2h1zjOS
daUeQMrOd71yQPOMvMjye62zp5NO8yTOHJ2Ly6GFmOubqmJQKxiyoqMcU9DNbKS1
+a5hOB1NY09m9Ozm41yj9rw8PTw11BoGGVI3XgtipJF0KY6zRQdvMWy3bPr7fEwO
8XCsDZ0VhgjX/M9sd+iu2dWHUBCxc9hS28JCSSH/VqFS0IHhPhE1Qu4D59PUCvjV
bNj9YIiGs8yfpFZ63xqcM/07huYeO68hr0J1J7bNe+7BEUZjETK72o7c57hq/lJn
u/0a9qcBUjQtHf++vpSqetkrbGP7CCdcc+3wmYielzK16QKv6h16j2/UqSYaTX5W
viW0ErxujgIWoHjV6OXQnpTaQU2ve7jALvLid7t/LdISaeMykI73HjJwgauxitX4
j4qaDPmuxRyQztSN5GiBhEAAcrpkHfH+PUMzP4DhGQEw+rhWJtsQCN1o05/h3ALa
xWM7wA3vIjHsEhsuDcj+Rw67WeinZ8EEhXGueV5q04Y6AbyJwHTCWqCcwo96Imh+
DrNeHwydETVabhNpoLRSfTtDRPYDyvhb8kquV3/3M/dr1F58SCq1W/7CbG/Cv32N
DGJ764T1pDCXvTVdvBnE+9ET5Ce8hqeK84ioG6teZa8ZvIKYS3U8bQIQDGJfryBY
WLOfiC0DcMnZIaBoAjTQfhqsklaSqEG3GQY1zLFmhUaKLCwV5MXcYan21D9K9fDS
3LboxhFWA6nnPnIrKks9bwV3YoIHgNjUgBoLDtat+xuR/ZxiyyEYHhLmnpnQs90A
GrzpmT5L0oh4V8vsZ7lHY7Y4Cs4zSK37vapie37BY9R1d+W9deKlmlw9kyp3pr2s
GpjAkQ8PjUvANfaQClJ8PP4DQgJPCBD/rVUAdqYZKR97DDY6QkT2xgAxVBujGeQg
ztFSO1s6FoNJDK22ccvVk33lQTXv1anQujO758asZG4JqinBJbLwHhNo8rkRo2nr
LsqAmTK57bJHvk6rB74Vx+vIhBBOe7i7Ppqmq8ZiLYXeWh/fR6UpYzwy/5irht/s
fu14KOzE7/KNVxgTcONj0cJX8wTtf6p3QxV1Q3P4BjSQjr6ah7TBkJmptT5Pn19s
7rdNoi/Va2h1pHcm2GVSW+FaxAM6Gw9WqrJPsG6zFO0i1Ll1SgLnh/ic/P671AAw
iIYJYmfcmx8ocj7pNAQBSrTS4P4n2K1YGUjjxhLS2JQ+NTdE4OyNMBW/IsEFpUtA
x/sihT0+IsZlEP/yEhEbI75p0cZqs9AxXg8oEj/m6/cyVocM5xlY3DxCKtbe/RsM
9ajET8iFkEXkfSw4PdvdWDTl64D09+KoqpPSHiXACQjj+ESaEk1A5ORYlGAx4kta
sAD1N3zpBRuy3Ae6B+IvHmUKuLgcHPG2mTQTPC99RiWQcd+lCSsvmcCpwEOC2nwk
+OEAYgJD0SSrBRI1sBBF8BEfNLv7bZ2KkJAbPCAbld7/wmR9h63hAO7P+l7S/5JH
mMMi3F+HYolPbwoqhLaCiBsOMGE5pS1r36UVnAY2yZX222DNAIbbXjC61HF2Aji2
AhCgNChV+ahFr1QXvzjQuIo0s22Gft2A1W9l6HGIL1h5tyGzpWWW37dFV9Z9Sm2j
FlsUqHV178VVtn2F6cOWZ4JjbLyJLdXR/FtKGW3ymPLNLdp/W6dRolWRPzPGx66Q
lWw5XXLrCf2g/j7q57nQ1xnThVduxKx+dxgwnDfWFWo0wdd1oqt1iaq5Z5Q7z79z
YOzjNyLO2Lqz66kDM4o1FYWgKQ9IDyGzkkbh5l5glzvWlCGkq/PjhuRXk5/X4n82
jTb1RXcSJVIkhu6MyFryszgxAO1/tkagUV5joIalpFVcUZ5BMKrrDRb9psl2LGA0
wl0cKJ0Y/4BCp5OT5skZtazrDaccfp5pA1IS7YIiJxJcJEAC5KLUD4m03c8w3ZnZ
Te4RS+VUVPcV+iOdrXFQeRV5QO0nSJl22g8DBBwckWKYStJFrbG0E69qe06zp8K4
6PRZbJe9XSfC3A2kgeUg5I00XfM5/vEmI0D89wLEnNSTnFc3wdDWR55JeJOLQ3Y9
ffYpSFMPtpPq/G/X/Y+Llt3Z/AzzwyXLkZvFZoUHwepl05/H0jKCWJLNjql/RSlG
MfzgHVE35DUH6g8Lh/EJogIvs+dpIjyEvP+balCpo3g1dFVsu8lFsrLZckNrXkv+
JgPU79cl1ftOnacmMBxZAJInAr+JINjXVfzHyIavshUMu+dFZGvezpAInzodsSRQ
W2SqriLtSlsvmRpoqXiz8rjDVFP0WCNLQQIVNOjHY6dnBzzaua166Z9aUVIijKjV
eqWL4mKAiLbaGdVJlLG7qagu6QvqPTwSCi5lQj/J0VMG/PzLYOKQv25KWBaRfvuN
4W4IPmZBfF73ZI6YOoCmnWEcmIowXRMX1J3p+YTuZUbwuowE/7E6xXA4f2t6Q07h
liPEDr6n2KrJ94hOlfpc+CshIX9EwXBGF0Z6ahl+JY71XDJ1FtPdN0AnWOTIQOG/
tL8gCO2xdJNs/N15AkQ3AwEjeKTaokJdW9w4cUmniQIMWyDdlPY2u8StL4dZJk+7
MkSJYWbmPIbdm02L8uiHlbdBv5FhZW9BK2HKCk4N+SITM180NxUFOjBY81A2vm1Y
htC4ARsFzcyRUEuOh3TABHrcFPW7kpc9kUhbZTVK2O0GZihoCcPguvnCMCtF3IL1
I+2IxnntaYDi1VwP7dP6VBJDvD09wd1/Swlor0p6vERsjKmRiFZJ/PohCAXkMt5C
hqW3glAphHYEgrAkNQJ1/SQs+nztUeMYSbLnzYcUpZq0stDVmH7+/kIl9NLPViqo
Evc22JWGouD8S+UppsFtnU4OoLypSuJ1mryONLP0m+/kZts64e2dIflcJbeI5FnM
8yXuz7/ozS/s+aXj06fydiYnVs3cNV6p3kWSpn2wMVovDAhvKIymQksKOsnqmiWt
1HOYQ6IVi1W3kqoQ0RYfIl1RIL4YXvCk7Sl6ZjXODgSZg5vwEEoBspmpPJp1ZHcx
wbX+IcMXh2fQjLn+1j9PmkG2rxKzWNE5CI4fmaLLRxxGYHiDcUDtRCpdZe1FcJ7/
QOmWNZg6LLQ6CvkUy1Xbbjb20hlSw1KNCu/6FY64fY7tTvgVSH5xu5RJ3R/c/ILy
EOaKqViJnwIOUnP5QD7a8Qh+N4i4XbTbiBbMPKGEKEVmATJIgcFRjhloDX+QEoDq
EFQdw1pSAo1CHiQK6YT8D2OBlS8lWsXOoZWXNcNMdO+Ly9HklMmrVkBtk8SugoSW
etLcQyzJi1IdwG4qe7+8bxpUtCmuDM4omE4pU7cNcf89Mh98OWfYci7ni3m05nLl
9TAIRM84qORoKX8npELPwHMkVmFUqDQRZ03VWbEde2rYSti0YcpHHWWbuTHhiMKg
jpFLKnkvMiuNY15P5jU0cWU/eb8TsUu+Wvvg4dqRGiTTlu/sboVJfjvFOuleVAFA
u6vIr5O3DRM45EtDaq3TL66F0HY2rTeZlmM8Y+WYIoWJxvv2Ldl7Nevk0Drd7euQ
Wdh+oaYCwbAcAh64nYyj05R4CE62t7Y1tOvir0QiCOpnvuPeUicYhaS8Ii4+scox
7+s3eYxGpt2tFZdiqmKGfRGMwFpkfYj53odzeZ3xEL7qZMbci4sl73j/KAT1UP/j
wJPrYsoIvngwc7djMMZi8GB+zijNuF5NZ3gyNH9JJUb+MVunDA94lb1R+p6REtF2
3/8pmga7icvNLjJU4qoRhsEhNFEGnprLrw0PHW8iBoi82rpgGdwig3dVYjccNaBk
ilXxdiMdPvs4MtXyIodKXGEXlvCYIDrb5ZttIzghivxmmUdQ363vt+4IXuP0lCr9
zuu2or+n61ha+S+etpF3PsvnqKNrt2D+rcbmgrB9nmFUVGi4f/kcnLUqATTCIPDu
MA4lkhDM3y0uL+m3p2E34v/wq70YmUkq7KAp4quN77fXpQlZz1hvuNKDp+xmw6Vq
usJmFx0U6y6JzihqeWevsWsgM5McZzn2vUhkzOEaAQBmMslPOGnpZGiO5/Ia/8Sa
DHQCUxFqSrp4Pr896qcdZ3mn4t/gUjpIs/Mh7NILrVKEwwJtr5k/MjuRympI1nG4
KAr8q26zXu1dZPOSkcYrZZwaqhQW5iSAiHXBck7DQ8Y869djDmpdBBiYlHNJagSg
XOMK6uhcszZgtOHIOs9CJ17VSv67onL8Mg4DpnlbePGD/RnjO3fuFEG39qyvfv0T
0wh4JFwMC8dU8JSUWS2G7zrxODPkoKe77htJDcRuku7BjWMX3I72LuY5PyqorfjZ
J9i0d5CXgp5vHv9ovhLyr7ePcrN+rptW9JNqHpnQHJYYNtqnKjSTpcrB+83VhQAm
wjOvqRQcPyr/Ou+dWOLq05fU+4UE7+zyK4nJvLjLZ1bfop/1n5BPf0e+KBxfLDhR
KX96fvpLcKvD6Bz8moyUHtDq4Iu9uMTNOIwjXxSTj+F6AxRPC4Y/ksrtEAtS3hMD
JeJ6PhHM/b/Thw4ACS/XE3fgomQwCQ4P8HYi8CRNjD+jccVSAyONNi2A1uVJFIop
HegAP2VjadxBTwuVW0eDh+2mjFf1CtC/Os8cW2hUhLaHahp9QyNGT44hfM8B2SJq
QufEti8QuzLouWNGZ2H4cddBVWXnrxUZzbU2/89Zwkb98PzJrUE9tIP3u1inBppI
1j0kxouEUy9nl6EkkhI1a1XIuka94MT8XRxhMpLzC0GxAlScEh5t8lZuX3fyqGSD
IUleDU10goWvbfXyD69nPt191BYTsu5Y9aDsBJ0UL4GQ739j42G7M42IQfxGhAG5
1VIAiQad2UoCbVeLVpkRNuHZsdXcmcITnBxmus9/gTUeBSHguF8dWvcJMWg313lt
yK4h8QnT0bK69qcgKXiG04mGvXQ80/pJ48jtPzuMC3FM6P5LQuAcWdxexDjq3OjJ
cKX8MM5cQXujn85xhZqF4a6mmNV8zZ8D2F2YCtRKzJTBRiBPceQLnVME3Ngtrx6I
VGZ4Q3HheFJ38WMmP9MQtyG5xk4spbi5iRyLMl/7oAhSrc3ljpk+ky4ggoeR0xkh
BX7xNRioLYOGHhKPc/w4/zAOTM+cOOmDbF43zB3jMWHi/vwJeQb7qT+QmvWliFSN
oJAaOX6tUKyKwr0bEs0gldwikIdLPf5C9SUXHC4nRee0hnXTg+IrEwiyukyleeIp
glY3vpkYG4AXJXw0Gd5Xorh3Go1tiwiPh9VRHkyURLAghq0398aNioVzsUrrt/EC
nK+cVKDloGYjv6MG9JOvX7Bxbjfc4XrVDzseT2ul17mO8eFjQhq5/09kW9fQDovC
rZKNuHfqP/kV/GzRpHRjJe2cA4WkpjnLl6hlNtE3W88laCz5yPoduVklo3Neyo+T
sbNKvJpurLoAg/HIOpHqegf/pPvF9eZTtq769FDrk7U0BxsLmp1r2KEukxK49K+x
ZXwRw3F3KEyr9hcgc7I2G02slRKSuB/PYWMKy2PgiqXQZeSkKNeDB+4UahmCX5zz
jZPO8mMnCtZmWmC4SV6n8mrDXfg6NUN1af4Tk9iql6YocSIzjRtktZFB3sW8Qz+Y
BRepOQ/OCUga8PQNRq/IN8O1niLtlHOvdJB0204ojdq5EQhH1QmUxnUck3IKnAkI
JHnaSodjMfb7v2z7MNQNJJJq+0u5poASSR2MSMpOohKWMBzRdIXXHml2YRZYkzD8
JQdPreVy5TXOKn70BF5b8/Z8/aI9PlFXl/wAiB2oCNlCk4I40IUPWzioXwFHJWdD
x2HF7KfOJu4faGH7F4tZEx4ZvTGYJgyqR9doZkIFTW2h821/tsa2h1mY4tsMZ0+E
mVS045fS9OAL27WVdZ11E4yLwls5oeL7a9CY07GfZyBRSFghAFi7jWU0PaoiGug0
uc0/J0dE6ieEUr7M+KQh1p15ptHKuDEiibnjtt6osSbaMbLKyCBkKETdeDG++/un
+IPlvChJ7OYiZUhGVgJnsu2ErRYGzQyN3EgbEWH9yQJAnf/YLjCM3ldez72E6d8T
7E0yg+R4qjpJUDPi6kESOaMbB9RfSx2xcoZPstCYTSFHH+HmvkvnvSQEml9lTgam
ISAg6pDMKLOyZC9CTvE/aVq+5tds042Wav9du8KjMLKpC5Ft4YBLSLsQ0IgTgN45
bqaKVrOEPrKa0XBVrkAa8Si0ODQIFgPWIvcWZpjqLw50964alkDNkwAqdKrYuSJ5
e0NLYsnq1BuRUP/y9/jYw2g7OTNbIqCBxRD1O0fexy774bRBQvfe/b2DtlxzneUZ
MedRTuba7/Gda694HzabQSYuelOK0rldbNGRnFYyM9xUQU6SAbZKnpUcJNyCVhNn
ROjKC5wDStydkuENSDM3q1Mhd5wMPkNc7g2FnwsZL82O7nDQESNivcefXZMqahe4
uKz7Pw63RefSo0YpwXdkX5t6qdI0k5dUDUqau9aKMX0C/tq3hypvt45gak4gHr2s
OV6CdKkCNeC/oBaup0xN3CUmWqCOVfVCCpbFkjZNolNRfQx91UghGtxV3fnX1qph
pxTY9UergMECAIyRHm3IgAmOuFoF1p0FJ12hHnA5C9yui4AdLw8Hj8xW1fSQ5haV
8GngXLcIy8BkOugQosv5XYLgMJKBvwhBNsD625ACN5xbCeFx/ereSvyP3e2MXTVM
WWEUAItvLDnKo3Bi505ZkNIe1ZOE7yBUKioiiB8+BZ8hXDVBsytqdfB5y1IcdS57
0KNONVcAUPEYU2LE7RpCu0l4HFILFzhkKI/zGDbo9xVm1LlYFEAqusvqt+Xw4XSd
7VAg4XDV0kDvcoMI8t3ewnqc0WF2oiNguGDMVxLCW3RS4zV7wDNyjLGDZ8QnUkwY
hr85y4a1si0WZ1yqV4h7t7yWEMnDLBnUmqaQVQM/9KfrZ//szOmy7gfDDNWSXyj3
AtDDyrZhdmP2MN/Kvpqi8udFJ8rlxVwD5s1r8xDwgW90lZJu/qMZxPdJ+7qaKrHl
dvLH0P8PEqSLM47bq63AqpTOm25JNjBO4ixSo1Ors+LWFw6/glB3+pretoxpVkxp
T00R7k73qDAz5T+YJOc0xJm5qd1AgY2tpLW81boigBT/um4E1JOd7bCZ1lDekYOs
7tuDMlUiES7cpYEmybZEJQCqJsQOhqptrrrBXZ021RZHN6gqxw6ZQ0LuoC09/q7I
qY90KbDArLk58Lp/M5heJLAV4HltiCTOQ2JRjgB/xQFzd6RM4AJZPK7WLchaCj0z
nRln9yPFWXDyV5SOA6mP3WAyloJKBq6/X90ZCj0z/mPolGbGK/qZmnObvQ5IptHU
WdOb3Pi9ENkKSWhNtkLWBuAhIHuTq6+yZBWtpURYK/QYwFYIWSomFwx3jhH8HpgL
RTZ/tHjhLOPHam5f2gRcvSY/dsvMbTCcYRDlIOs65rfBqIubc7eY/3D6gwSuj9du
KZ6ybssxAJh4TaP3Wifbb2XTHwZ8OxsfuvM0593EZ7Py/Z1EATt02/WvaNJXrj4e
UmTDoCWyFXSj51ueiXbE5BSnN9n1bvMt5WzmzRon7R9uJL21mStD7y4Lc65eN/2I
9s743loiytD5A6WDo0grpICD2qpiwMaiTr0YWuht8lWjLn5pmCgwSLvWdlk8nwAZ
b7DnqUshxZi3NKoTopv0q7ckEQkBIZ5XyZSkiV3BM/YIGE40vlz9qli2ENoyM1/w
ZaktlyL7rv/KkPJe+czDRzjdsDMBU0NbFFYznTKvLhUjaHmW7lk6L9JiBwsllwDS
lL89dFs+Hngv14eebZVcPVAL/6uA1CbiueiYq+DhrsODMCTJgx+oTF3pu9MBakVP
Kz47qLXGRupUYFNAMNG5c2Tc8zBK7MmOYNx9bkTPwNzno409UpHpJiOkbJyPkSO8
fSafly+lkOK8fjhsk3uEtLLq8r+JXSQWmvCWWia5U4er/eNXcfCuIxz0aL0Wfkqs
id7CaB3wypba83jbEKGkBdnXKjTrAEGpCiWsvScrE5F09pIhI4gGIjrQ1eI5wkCU
jxBoRVuXCEhcSBgOpFHTCu6MneEQqTfnNPRbx13emWcY94zSDq87IRb0SEaqpctG
7pAbSFTpkQk+yiVPzLHGyzCKAmNHqnd1synfBBubVARgjphUEmvYEptLLdbj9VM1
DE2hlkL5CvhWWge3mipfXTBeOeOjotIisLOaxlFbQ0FFq1yz5ALQe9cTw9VUlrVT
loypYji0jhqU4E4Zk3uEEqTdZoyqcGjbVYE6W90LV1pvaXjbUFlV44fssaHn3LJh
DqZn9m7i+EftgHiMKeeYKlnsaw0B0z3/+vaZdh7hZDu5IJNi0OC5cM+Yt6mn0TUy
0TE/3IUAmTNnaFe4NoS0uQiZfeu4Tu2HmTq24IRcXsn9JgcG1SpRkmmb8Qn4oTCY
kLXBhc98axlsWxlaDrh5hsJbw2RWFGk/7q6n5CHHgH7e87TYVc2uy+eg5w2ps0Dw
VQSKQhsjLBJuS4gYPui9VPBdjbGolGbmCl+Yf9nL+Q+/GYXcfxp9Pp/EIjaD0z0m
YzlE3hzIqOas05YGuVewCPjjE1w4yay0W1SJZxmFo5ft4LFDSpNhdyk9RK/4AjBs
2alAwEhhKtTQCOcx40zUrYUlhKs6L0VaWd4Zq17fTu/EfNNaIfDi4ChL+j87npQc
vb+ZcFBJgjOxbYiO16gxWjDO9D9jE6pzNJ9CjHA5plQHdLKEnOea+y6rkNe6ZYgU
pDG18RnMrRyWDTYY/aKWJcS0cCXoWavoJb/AtupJWwee67BDCjbKQfkXTf2JpS+a
tP+48Ei2LQ3eh7r27lHZqLwCCgpTew67CS6756A7j7W7UkkAot8ByKSKK5qbWbr9
Ly8MEsBjQMVK1gSBL8VPVlWFosSZpwxeFb4XWmZAFW1+D9H3Bfmq8FCGujapMW+g
39OMCQNGgZSw28rc6AAS7Ck6k/HHqlGSyWP08aHqK8t4gKJirmvjVAKELTVJ2S1w
+PAwm489BpIUZuHjUaffGCTP/W15ogwsryXm8P1sQ6d0Lv8dxVfbCZyc5QMTAKGp
7EUUHrJ+sZIUtWHVXDuPAd8nLXubIv9TnxpfRIwd1KImLbUT68kL6RKykSURycqt
2HkXQv5ix9ivktmDCZPfDouN8vz6xJ24IBPDafgBdgXLNhcX3XJi3dS3doeHyYXn
afj2WjhC1B92N2Aujek44om6VFFxrfv9sItEOHBVxNAwUpKsDtOTwORqZ+AYz4Aq
zyuB2u8dAsZFjT0w2TxFCOwBsakgFvwA12zUEwa9qkGjPfYC01yUexmTdOOOPc7Z
zwaWymUQGm8wOZ0EydI5QBpGBuSPU/nz/PAbFLcb5hhsPK12xe9ePHduDnWU1NEm
HtQvPR4Ki/gjwheWeryBiMe9havfcrkl9i1MJuSH046BeF8nFo2hKQ6O+7OFUjqw
lwiw0PpN9YHLJn9Ijy+CCYn4Qa/akorPNrFkiGfoXe85e77XdHGiqCH6gm9gXkUH
IzRmd1Hh18+Kze2aEkFO6vx4zACYeoBmzkeCC2TpZkP7c3kdZ+Fjyb5jxjNVw0WU
W6SZPrP5EU7eiAWs5B4LINUpYbtQrugwGnyynSUYtJe9SuB2yLsAY9sVdKyUOvUD
GIytItaDZYn4lKSQIBmc7MSVszObqdztEBnPwig5/Jy9rFzaliPwURs4GT9myrnf
KKtdzLyAS2UbpvcTURETC/AnM9mwjh/boDkyFo3Z9kK43R+6vhCGfP7HJ2RmudAz
lWz1Xk33Q22YPDDkV3QNGXCIFITKgDFzPQnji/arnZJ9/9hDC5FM1YTFDi+EY0ag
1NpfjRQWSuVJDBikHvI0mhsrbWP7+ImUbr+sBoyKt9bMO4Zmexe0Gu5KYHnxvP2S
UwTJ5IYSaRAKv+e2TgLFcx88hm92ATo1A8kYk7KH1H8V1nwmkt8TZyvzYziu2yfP
oTJQM0607U6YBF1HEsJFBt3s4zfy+yTwStlXf6RWCjQ/hOdxVNtG0rTiohWBN5Rv
rNFaCFEk62KwZ08AeKS88J6Bvg1VTQcnsYZPDivKX2venAF0MNpJ3f0BAXAvkwhO
wwC/pgFDQN6o5i+ZHCdJSskNDk54CSjcHGTIXv9DjAREKM5I1py8q19STuwwJNRv
z5jah5XFTzqXVxOVijKGM6KtXuAIw9MTDMO/PZQlJm2J+WEE9ZAnlCtm1H8Quz+4
6qRSG0Z0PUjxLyREz80fhX2EIJ3oqlDEpV09rlbtc4noQREz6sdG++xpv/P5xLYu
7gWKkvxmBJnrIz35vvLAGXBhI7/8UCSQtlRuprT0pqENHItQN/mJ7kuDNUJ9Bpe3
sGqXHp5mfuT8DIZE/rTYgMylUqx/eU6iI5ZoTfpr4MJK38yPxknQbicKmXpNTWA/
+OisxB6lQsDvQKYc+TQO56pgX0Sc2KzY4vjRG8ijPDGCKiJSeFmCQweLC/hqn8Ra
QQcuynUknTfwEBSFbrDvzN2FHs6IvdiTFlp4d4wDYDSzE390diwW67USmODhq1zg
aFmiWll9bmq9jQRQl6D6P68CqHctYdzUNmPLz8B74cEka7EEwfmeFS7iAs0VvBvR
OpIDWfsEtuG9tNQEz58ie1QQmAyKzs8fokQEs2YYq8jIM06Ga+kr7wA94EEPfMMg
5OYZycpAp8ExHeNNaVwdlZK2fYmfWayBVW7KKQZCdvFkioDvJhyXaeHCGfoxqsDg
4ZiTkNZv7cHtyUnlt4rGnI1hN0i9S8AcvQHTWr12b1Pcjehd2MLVLl0xqqMjMQtZ
DnyK4ShVlnmU3dsa6/7Bf4Wpyk0n3rx+QP5Y2mp8+J6JxEpCxnnhDFWMA/P4wcx9
EVcB1zCUWEDNLyoqJunBwhEMTw431ZgCP/mfmiOGdpRR5eWe5Dp7BMmIENkAJ5MS
rkN4bmTxr9OXXfOYPQH8qxkNdpaKbkrsDSgDldPvztMPp8+wyM5ofwOMEksbFJ+m
Ht8OhNBmjg2W8/2Va+sp0grsfH78Yrsr8xiokWysEt4VXYKg7bZv/p4Lk5YzgGOG
09fUO2T7JiEa/cQheuEULO/xYeuPeY6TXPSq8fTqOjjgHzdCLnpdjrLoq54oDWWu
/BYsNabsPlM+LOv5k4tG/C1j5mDc5BK0bCKWr4Mb56ACrEjhFLg05yIi7RDYIwZ+
U7HWiG57U1Lz+l+Cpj0s9DaHL49pMNIdb81MwGfDW2R4b2Qy3mTHc1iyvTNWD/Fd
MsBFc/uOxbIidvzdMr9Kcf+KPZpBwGYmDlLFb1xcOYHpisGClTcLJqbGc7Hwkv91
Gqb8QCLB9c2MdVVUvRCYo5lmrcGUYomi4CzB0Qdw26s97EUZi8L1pViYt5ewkmBv
WeSE1ErRFdL9qn/qLl/nCRKYAAYFdc4rcV/aAj8l8KhYoOlnlg7GHizb52sdd42i
V2Imf9TjvIHZTBE680I6saZnY3xQdP2y17du45X2N6hpyl+RcsZDBRlyEtIUzvdv
z3qy12Y1mvh07cP9ynzqYUC6Cvr0Nd4vXyQf/nlJvzYfBNjclMwUJETDcqArjHbf
7FtSpGX03G342wmZyxffBBPgIvJ4E8jxHcs/d7EKixJQYtTxdENrSYRiRh/D0bd9
aMjDAx4zdcDnyKwd3K6LAGVOHTzx3F6gv8JznDA7dJU1HqKI3CDJ23Kdez6riGqt
/OVCnH/ixJ9DYspERZJ5rX8wp+smDl+0ZXVmvUhzvcXjThIqZ3vg4BSHToI5ircz
l/h+lQqbiErYS9w+/i/r+YPW+Uib5fZBm13LlzK9DJa/TINtqV7F24uyTqh6yf4n
7bu/N+9cvhVG/fiSO3+IiEx7MV4tmcsGcZOtue9SDyaO7T88HI3WrBiRr79QJ1tJ
tyDzvetuIz1y+nR2zM04PgVNvCCBiVIGQup1NMD8OV4ggejQmJZEeyfeCrPnMsxx
JQ2ejsOFXnuz/fsypXutN9cE7P5BYHj4iOqZt+0+Lj+DT1czSVD2R1Sa8M6664K5
9NwjOtKiPyPyhKeGSzJXuu/EOSj3Op7PBiAr1D2BHAvXkIqi+o22Sa/8xALEU1T3
+h27VJtYxuavEuH9KolqbqBS3CHRUptQLglTTfuAg8peDqczo8DVDD8aEAGpsuXK
RNv6gtM4SdSbl01Mc4i15Iggr2qt1YGPa1V5rDTlyJoD5cNoyqYwrhBHpRltlHOH
Sxs69rAA0SUN3OLEuCmjtMiPtcv2hN6vKC3PBgsSZfEAA5g7QLU+1NxE+n3Fq8yR
r5HM1wTAEb2hgBp/JszkbwF7JP6EylSQFz7sx0tTdgx2apJMwD5cUQr+t6V++m6X
+rhXPPgpUaxtXoMTz7vkFKEwevOcvRZCeyTOXCge4nqjCpfeywqU/9rb9ueeaxUE
Z3wLecLrJMaESeMp3tqb2HvvXobB+yQCdXC86IqhnPqkRCy7ib7Y2ugzNASxl4no
5E2xWCFH1PZPVVSGhEgN4xwDiQtbI8RqoOJZHZMtvGcsZEDvX3xZLpIqJ4waxyk4
pRXHeE9rd2o69bSqp/d+rFmGSA1I1uXTZcEGtRDf8+EQ4/VTHCpMPhQ8kMqeopKH
m/DI82Vr/uie7cLro/ihgSSVHgE/niQxBHmJOr+C+WmH/QlJ8IQegzbMEpfRNt7f
dxp0nx0yfH4OpK6WnGQSCkh9GNGr1g2jLSAQAygTyfJt8NLg0fIpJp8JBG48MLZW
d+cQIfcRHkIlN5BauUlQStaqmcbAv553Yv6i+nMdjhm09ae9gF2n6rSXHJYkhFmH
yQVPniBVVYHWB4BfEwPZq6ZbsGGLoZlTyXdV41TNriMgT7get+aQj6Wh7diDt8Vc
qpcoaEbjlaAp8BHUy6PptonHA7KjlkUSBFMhwNTHj75CqzfmNSD5XerQl5qxaB9/
TYl1nOColwHc7pVesJ5diw+wywhiwe19lGxqnAQ69HMtCxjxPgaoN5ZVqJRgbckg
VhRFRVOHT3PT171ZFV46qJzo8+PkggdyPW8ir3rvJp1DhLWXdidM5aUg8eGyu5U8
zX31IK7X6lNh6vsb6d89MaAotqtUgTiSUpsxEdFgnkGJiffUkWdvP3cGG1LlMNOY
z3V2gPED5xQxudh09OL885Z37xEHM498hvbKNq3kAHUJIXU7S7eh2FgsVBoqMlxM
qU4/mKIbww7MX/17OP4uyp/2pmanqUYkoo/4OdFmZQSMqWV6g3l3iKvy4Q0+5X+T
bHg54rET7Ml2PFzdPLw676/HRQ8y2g3yOlYHJ5FCNoeG5clcpI2ywwkrMiy0MvR8
eFi8QpkKrurl3hIP9SGvKIHD5kQVo3ROqi+Abye7ZhOobfsYh6gLGHkX3RkXq7Ih
0GO9pTynh0DXYDFNbtFL0GY3mUrrau83/cRkJE0vEJZnL9aAhcm7deGS3GzOlqeM
neoGcC0aKxp4IddXbKknMPkOyDbMC8KSE8eci+ixVyTUcXwjEbu3e2z/HHuqqA2d
X1lSA20kpyqkbJCU5g+ZVPtyRUjAQuZrd6FAl04EzNupTwMCA7NCqsiZ/MDKuwHh
rVqv30U6kdLRLXxWAqKV5wFhtstJxBJVotG0hrNEWZOql0RGVDazQ7bRfZtRORdR
rsYoplX0OcOUBDZU9bMPdBJFI+jy9+5UnxJKsMobhDDuEkBS0SupCMe93HVhORQX
3Io529WJN2RJw4IwmhBPSsDGw8BVVMGH1Qdke6R5+fv9ns3p2Lqz8g77cbA6ISDz
lYpmNUHMkezH2O+cLCvlQFDkTmA1WWyQjY67PJ5mlxMc3pFWDhrijcAFD6diyLdS
qrxeVN36L1HxXbwp9gwFRrax+AfAujTHkl5Wm9zJG26BKQF9Qvi8orgYlKDPetI5
yO8gi+Il8oSxyBWgX+5cdX51zZ/deO9hLHUHhc91CvUepWMv92j8RmBqp/2Wp7KB
fpdOndQCoz+gLShKmQENgd22mud0EniwEaOrV8EJqrENfJ6WyQXGaiw3sMVBW/cV
kstYak+8PFNYI4PMZD8Hq2ISeqJZYOeaQuqTZVNcy/r03955wLkM/77xQAxCAnWD
tHSMYJzw//ZuqxC9w65adEgZ+YbqtcJwYKVKPeXQXYCNxMrxbe33pdpZfXiQyR3c
YfYO608j7XYO7Ear0/vRAi3vUbUl0iGarWiI07IO79TY1XZvM1eWfeBS38QbThl6
wl023xvtKLigTjSa2N9Y7iDOE9SD9Jki0F7nlHoCfteplgygV7ZD37rxa9dCosNa
3KzPUYJemZfyosdMDPJdOMitxEim5CigF+3IBZIWmoHhJ8l85eqz2OieiFNJ7a1A
TP6pKGTVT0GUrQV1jY211XNCi/1kkR/82tFejk/UzL6gGn/dGShfJ6LQOR9r+3Ug
CXC4Ioj/eYQ0ToARKLsjtrLOi85MhxM7GkaTK1gMtTEk6XqMpEG3D02o2qnckwEI
93ihjNOrvIdb4rDM6xZvdem8EMar1avZJhChfW9Jp31TE4fq8Zo7/tj8EQLUxuYt
23X1Igk2A80ekthWoTyFNr68K9AEOUqyPqjVza5WJf8ZMpPa4bPAF4yPRu0399Vg
fajP6AgEGSdJilbBl6fFrEq09xBd31vwmOodOAxpFkoDA7bfIiV7vF07tN6j3ptT
YJXUhXNCVVB/IfUnseQmOmRnUYuCMCI7piAKZhrDMyaYSWaXIpE3Q9m5Cv6jNDCa
Eq0p+IBWX0E82ikEEiE2maoHdQpudallz7Sj87DaxhhLKWeLfC069nSrgWd3WdoD
/v2LiEc9zCvOfgi6KWuDksjQjmIo1O+Vg0BidT19+/g2y+8o8kcMHFYD0poK2aFd
il2WWQxFUYEb2OiYYWyzs3d7H/BCCXb7/UqRF/jASs/1cAbPk77vuo27NRVR5B+Q
e/q4066aQCNXQZiQzLk7/eDk5FlPkjyr5ZF8kGDfBqhjGfveVbOIwUhkUx7gukEj
FKKP54ezPcEtk/iNoZqpNOSiEdSMv1+T+LhEao/XQ2VaWE5Xm83Ockw0qb/yghGI
atSj8n1LU+ayhQ80briTubdwX1cVdQzBj0rDi7ixdnQAwBthmvxQk4aoWXYmddvD
SCvazLycMhPaE9HVp2xiCqA1ix8G4192fkq6VQpa2xUU4wGpEAgvBdArqjIKUMmM
wLLuZtV6+1uVF+l5E6rIs6XVpKjIYEq/Tqr3O8+MDfK4mO26QT+cDoSdRSlNZeLS
BYJ1FNIvlgrz+kg68CXAX4xjufMkLvz9X4PAagoPIW9ifbZyfxI7IBoMEnOLeR/w
9h7Ll2KrDBAHiXOCcdFPZfi3In/+AzISABdzY9QYIAAQV2Cy5f96Vcorljqj830i
RCWIvzp532oIVYP7ejo0g9PG9Ww692k62KbnJQI5QsS6nvAqbCkJe73qQDlFdTzy
Mtx/IzKKlEqFKBFpO6Ale8NNaoH6JzjA4K14+c7ACvuBugXFjJFbuopu/IHlqnCx
cJiRyh2IGIYQlJGvBoey/2bz+Rfam/Ct2PSsWu6AsB/65tIO83f9e3Lgz0tgf+co
q8QL52uTuji9aFqYJPXOEn9TOBAyLwXNPqBLv+xjTKQ0sSMRtUmEJs6hWBYf+VbG
V8ZjlySNdh7D2eAD1FgfJRb9UjEu5XAFpaPKR/5Mxc2CgS++ZeF+/I8mcFJe+J6/
GsJg0/7OsLvoYZhPwDBJuQRW9x6xWGohS3UmwXFKpEqlys6hWshTkG6SG6WOfnVt
i9uF7V3xJTOPSajnXpEQaS26cF6GG42Ojyy3c8nbKItGX7Aax6gy3iQHpmHMuZa8
bcijuGgVDWmtJtAihdlBaO9CcUrHIVLR6kADsq3645wc+kKymb8vnrvxN0PWa3gc
FZoPtI3RvbX5fN45DKyrdlNBP7KpGkxmXy4SJmp0ZQXVlYpJp0YtnNjAR8Vm3KFs
ZXxZjuj1oUzpZSfiAMJF3C7fJTBzhbKOsf+OJ7bjuWA3XFT/oEr8l4gl30/FfUrK
G+v/XeaA8+11JjXXM4Zc5OL+HmQJ1uRWj3oYvgQcp3gY649CP//MfWHtPTuctDUM
wvp9in82PFgyYU4H8kUAIBDpQOAvZdAR0aoxqWWAIFSgMse6OHvl3sZNKpDXXD3G
SH+Z3pUXt27irexajq3sly1gPn2SkS18W+cNPxflXSSFK6MHi8l0693yjFaqKz9t
/+uAQjdhRNgmtZI8gYHLYDixV+DtBQiQGfV/KULvNsFad4vUUESXGPlvW5uJzZWk
PrDDivJYlHVXDYv5wnu2d7NZk63WsrhoqEwm0PYg+Xio12JHZVb8Qka2i7igFNgH
UNJLDkDp0tM7Epw4zbrIQtlMOwnfl95itkXN0hC1x1DhrttCErJFJmLFydHRy6eQ
W92ksfHbsih3ehWnOsS/IaBgMlLq2Qfhr1mjUaIk0tYqVPe3FD7jiYo7MsTUQAUL
QCfkimb6IpbOiB/cgU3tOrNGDZ/HIcuBssfJqrFBqz68RV5915g84+N5ts9bcMiy
V1GmnEqSC9k6wOXrIoSnbTsmhyW7RQ2TwWCTHyuuBSRQqQVS4pXq7/5gd8gQDalc
9+ggu7CPyG0RreAW/3WCyi8HaMI85vH0qlTIB0GJz+hUw+IvtiDCiQHD+3l1GuI8
eFZBo6zmOe4O08c1YNtl6MlhLmTjGPnN7dy1j1Snu/M2ILBoix2pfh5TrnHo+sYI
aD/f7DrUgd8cRyYfkLqVMQQpRI4xVA+zGWeEmElY2Ew8JXfTOrxijQ7ubbcwvf9l
9WVLuv04aBYF77ECl9tx/kjQjBj4SgfSolzDfA5D+ZI7IE7vHv85ySf+rvKbmNXQ
QZHcIvdmtigkm/uxEHTjuivoaVCnfrK9QEeX6msv9H72hyrIRUC0tkEv2RTUSRjo
b00jqq6MxkqTb3W76iMc7PW6vgMCGdunFRoW7FgvwySwUvi/OQBS1DZ3xQwQaaAa
GAQOvZ1kHmyOiW39Qe9SukJCVTfYCesfXQArq/3EjZqX3W+i3U/P8IggBM9Ri/yV
tTMhrtfpbUBnm/0VXxx8IPZxI9hybqL6VgUm3aYhQY36awFK3PFZk72yYOKRJ808
AdB9urE59wt4+nvTfNDjdNqyD+z3Fhtpy3muHR1fwZPve3pAGYPiU0YUtAlABQVd
yreTKhsGjmjKrbNGS+1rmNSauSsfw79aZhd2Y4+gXpYgAQ1W1dPN2lxxQ3WShMo6
WcxlOvHRZXB2XDR4+8ap9W7+Gn31BjQwRqNOALOh2L18LjoTFY2XOD7MxWb6Cykg
n+MLAiy8Oxt2PruDuFPhAcqBi2UZ/I+gJk0wpfTLH17YiVWl+XW56pCmQdYwYDj2
abUFNOUZ7Q++rvmXJ0737n9BBJbOIUc0Rv9NML563N4HE7JcugEiVQc8N8YttvVs
WmGONvq4m4h0BBydBZacNxjpfpOVzgrzMJFTY4WRaSQDs7rrgJiProS+lD8uAbGT
K0prRFQIjBNlPwSrXJLtpXOzfE6sjagVDvKEKFCyLLyYIw0tLvxFwT04dXWl+OWI
A9sFVdbMmIHdEsbdhoAnvyj6E/dUeBQYcVl29CuLp1ssIRwgBP4AWNYNWkixgqeg
7KWrgT5TEKMZnhPQdUj2r8BeZYKJ+OzXHj6whR9PXA+nC/uTkrMIxrjzXI4UQdM7
U3QbaLk1AeyfG3Ca9JAoHkG2Eto7Da1bTGk+uiihVe21/IM8WTiOAhIYwzyRNh/k
5dBIyPBlIW8/CGfj4J2xAkW/z0kjKQlaXDY/e6UmY9+vanK8Ahb8YN9k35BjVd7s
kPXPh0oHsa0QqT4XNlQd/r2WrFwJwxqMcc4S7AuwdFNOant7VpJjpUJ4UwAZ9SCj
+oEms4ULzm4ChoWSOQxCFXCcyLe6Z8RSJOLdV4OUl7KvhG8YGYZ6YSf4AsWPKMJC
vxIGHuq5/N3N1L2/V8uuVJPdycDJkQPrUqP8xzT3WpzO1FvkBzte+hMsfjCNUYXX
Zw2ENFvZLqpovfS1JQSrcuqrVOZxaFi3tfIsuxzHUhYAle+uxZcy9HgtzatzNmj2
Z2JljpdECimLdBLtk3wFShueTs0f0yZ1mxZ7U/m0813ugbnn/xKMPCAxu58M2Lzm
bzlhXyX97s2jPDqY3vQTO44lEvQMldYWKlmJYPthrZRiETIgaaHOLJCYgEyAzrXQ
T9p0LLsEpIaq+vBOD4e5Y7+BDBc0+6KbWV/sAg8Rav74oiKC3dqcsUsJCljXYQFf
OOz9b9fCea8Fe20H+TpvbZddWV8s6FpvjP2U9xFmFEwn0rtZcCdiKA2xfH+NiYnK
4YFwu6CTAXwmUgmowhKCXkMlyO6DtgUq05HrIKOyfiZHdodm/Igyw5WM0A1aSl8V
+cgrM1DFXHpCUI+HDQLMEwNRW6/V8F/cxjSm9LHWCy/+pinXnR1IFBFrSVnJd7aZ
uyKVNwG/wnADEgznjLQ6sCuoqhZviJQVgu5C9XO0A6FDl4beynKtRXrDpUhyJSxt
pUZcyT+8q7q7C6tGnSTF1K0AVVLyMD/czrT9V4NROIdUQEIj5W9RUEKqREaOjU/z
RYGGdznC1UOdhGR2hDY7C0a96WE00TMfGY9PWsWpPvtauuV1Fd/dBULYxWisnci0
qBysWoC0gRs1r9eUt8tydeX6J75Eo1MLzjXZQ7SGXLmFk9Fv0udeiqUj0cdD9CdS
72hhyFnXwSMhxjdyXUdhqOn30rWncQDK1h9DPFN+3PBPbrfGPAy3Cb4HvZ/ZTJ3b
pNitPzyysqFGG6cuFPWpOVgISbrS7xlNfnwtQtsdz9arlAtnehJk4x2p02VCUcMK
5PPmFgvoWkb/OX22mWJv9+l3h338mkC2jU1TlO7dJYEl1xZcFE3Cowg4ztPZdVjQ
nh/vSErybehkvhq1ytzpShlPDhjqFiB/4OH5ZRQgExKMtqIfXQtCSAqiIHCrjQzc
AZDz5ZPbhLvwfcnPplCkUTnNK/b9QXb5ZUNXR+EdTGQe5iRONCiuPM7aHVNpQqH8
N1ihB0PPEhrKanuds9fBtJo7lYCGPIkNGTpUhsJ0fk5O4czY0abBFa4Iz/knK0FK
8Yf/xuQBMk6/k69S8+3NFHEotT/hzU8K/zHNXNoM0r/9HMq8bBMOk88ANoY74yQd
fiq4LY4cE1g5SLN5d41/bqro3ix/cook9Ws+GPuHNaR8I/enG6ktNgWGscwt7mgZ
2j16USS1KdXkhMStY7C7rEQmllzQfluqDdsqcaetOHCsvpCPRuMhTFwuBfwaCPgz
1zUgwZKJJ0nbqut34k5YmzYlTLpw1gYFY5RpqTyYxOgV+oLepK7Et31shFhaTXDB
xotdYGp9p1BhVLORF+SrBuWcDVLdqlUybio79XdxZxKFsRkttKP7zFDjC8xXiYCJ
yNw2KRisZIP9aGGEbR0IjNE9uf7CGYL+O3iseXxyQYupGVmpDUMXy5jHWidmSADM
kBXPdVd247gnLdikd2TgdgrEdkbS1HGml9xrA/9TT2uatnQr1hB94E2MdofpvhoY
prVEC+p1pEpbv09CiM3DiD+b/cOzVH7Tx4Lx05QulF8pQIlfvWqs5/djBUDzmR6s
d7/lDn2PNG/5HLF5pqPc9kbTpvjFjsYwmbyAnTRV9WOesYK9k/yDXZHKHhAHutjj
r8DdB+zVu5rb8hkQ9o7uZOP1o9ocKBDwAX2OP1517zrNvmc1yttMU3Ntj5SQrLwr
eGrSRCVXmpCfdbg5s+nR3kMRQlFkqt6k1lKvMv6nkdYNEOB/8bWYRSZ4x8dMVSGL
E0yrZTKyjrNZxJWvw6RgWT3VciXnvGYFIEPrK8y7YLPrcm/Hem7jtJBimCoHjy20
1/wwYQTIxlNI4gqw+duCDTlXMitEChe0sXTEer6weR82VZxDjqH5CUzT0Lwg2Cye
UDoY8zPkCGphaDX83eogEJstMWnvPKmMG795Ig+HWK20IYvaYngC/g6wy0bi2nLI
nK7vTTjxqx3jQnqU61jVr1SpeAe/oDMMun3LJzJSsauwxF151dP3PaZv/y3TAIsd
OOw9ua23OOQu2k1Up317Lqy/cBOWsuLTzdVAykwc5wDNgEfOKAtZY+mXe0MYytie
NXwfDnGV1NjwXjKAe9r9mFeQqwuy+YWpVfQ0N7JVabWXY7RoDnHCdQW8WLoKhzbX
+LhHNq37uw/w7fbNM0WXn4E3KMOCGPJU+jSKRBgUsYfI6hJXwvIXLtlvdLAE7bRZ
B8DA/J/KVhvrudm2sLs3IwhxvtVhAiaVAWKNRRagO9kXEQe5INTuAA7K+zvMClyN
Jgc86euLEyHNwUmslOx+GV6KkQgWsY8N3UgELbYo0N61gu/WyNHLzbJ046sVsxmv
0yV2N0mLB8EWpAOd7eoMFjPEn81jrbTAIU8eneM/v2TmD5IuXvqjXQkwcj9THu4y
OD2hZ4oyiW0gP6CnQdqR0w/+YeZbQ+IGPZhACErhSQp/OMO8zD6W+Dneu/fuSZze
BvzwbkTYCzSxtZU7LaMq3bP4qiezyxLkVFSlAm6aB4yTUja5zDsoVa8pkzvuCvFK
G0UrarL4vzB0HjMScKIfyK13KK9iokROlxw3bjO0WR22/AUKTooNxGKHyHwKgZ3k
xb9skJCItDyHKgWW48Mb2hTFTPfJSKf9+2jk7vfR6wpnbX3MQVmy3GVkuhvvWcry
0Q69k1meX7W9z6Dp6oUEoqcLc1tGDJS+CT8EZZv6suZPS6KZMWe62aRJeccbeKmL
82GcSXRGc8hD/KP5nJfoGVz60AxESOG2ZZuAbuFGENxOdRDMpMb+ugIkbjBbu8z6
wtD3FnpprXw7FatlSXnGRpog2lv0e7AwszATSonSMv5IUg/WBcWl0HwcSAinRzKP
O5x+UKZ47mIoTJAMqp7yOKPzIczbOC0oKwejmV/w23akawX4Yo7ksgL/a0xd1dRA
bevRSbumI6+TSJlVuRe6EUMSx+wK8cg2+zeCi4W1Jk8W+H/RRyNPiRH+91rCZJJG
Tx/zKbPULdkCYJVvBfS2joCwpmOzkj1+9uavgtEGzXCVl9ojc+8nSBP0FODTvAGb
uhTUl2Lb1DyyEQXL9iz/xF8mGjou0J55ZzpHQrAuEjHBAf1qVyoOfFsaVY6/2iHF
1ezhS87+KpzjHf62IuBumt5PRnWn3nKUwqsEtjj5biWU4hEAnU0tQ01Au8baS8PH
eafx8MSu0nb1vY0xOY1Mo2h7B0IkTOi7nfj6IG1jRP2YF0IeXHrfqzZkXVBIwX7Q
HmGcYD63aEtFPokeSvI8CDvsHVmhhDrvAdT5Th6vbafhK8EuxHZ0cE6h1Yv56h8j
S0xj6Ek3eq91WZBp68lroGa3fsCUyiDRvdkJSuW5egFBx3LamUfhpRad8+ck2eNm
gCjXyrEo6/UW0SRYKbXFemCJIZ7vAfUg77lMYt1GgOM5O8jwHbRK0LNtV/XelyLw
8AGnSCqcPWLMD18P8QtZjPZGRNtuurnPofowjQUlRqjxXFeOK0JsckNNCsyNghvJ
VWp77RoIbL9KdQEFTcqw8Oxu3hntmxbA/3xhfediwwuzxekM1EJds89GnXeHIyim
Zqx81USvaNlNyD1+ra2MEPJJqZ6RUvM4KtpxJ+ZgnXkLUAxHpLEFqGVTgLkdvUQg
ky3qRIAGAw8acpu46LT/UqkKvk+97wsGUnCJm+KUCyh3YADol8yLxtTz6SC/g86f
1goaf6qO1CUVtw60r79siHFX5GGLLYUOjP8+8nQgZ1LdYxercvjpXqdVuyMnyM9I
+7Y2t+IDxEcB/YL4OWD40TFG9md7l2dxj3W0VtE9eUTb+NXZl3UbXeUeQlJCbrPS
ijdjbrndvnU7ppJQPkqvqsF+sDpKhj/YikfOv7I4fPyMo88PmJ4S7kikTJYH7WhZ
obKbVWc8TxgsWvNQeJU+8JGRzEwVa+W8m6DDrwksFRwIIalP/rx4pELulxnVIkJM
qA8GYBfhfmEsWJ9pzvbn+/JD04DfyboXkrXUDYVHvJP2X6tfnXB9G7g2ie/3YABg
EFPozcrhUXP9gPNzczTzhZNAAEBE+Qx3TkKofx5bpdoeeqmImgcf8juovWEPdFuL
vuaBNEVPoyeMqxu9RUDQ5r/Fqkr5dEMW+NQMLc6hoCvorKuJsMEimOHp4LfvjZbn
iYvKzGymobGIy+ae872qJm0ZucUVYyXhEn9qbXJD6rOKvM/4mp8B7O2X/zjiM9xw
Wx1WTd7FgOtz7KKtKdL0tW1wwvtMiGr+K29yHcRK34Jr/WAYHhPx81de+W8zmGBe
24Re1Qr5NpyVG1a5WodOiJUm6vhrI6eGZFwVd9ztY7GrEz0kO3wIfhuU3jjqJTaq
1FwjLCsKsc1YTptHkGB7vlNgGNeWwAPjlM7X7TG5k+HBvyCByDARd0sJOCI2K9ue
ISbCFAqUeufCVI37xzCnR11Y5LUkVTdsQD8+TYj7toNPZDkTJXF/usRSghCegsOR
ysdhOrYxZnkllJzYjUtBXHwNEE+77xzUaEPJzh853IDSBd4h5JuHk/a6LLEL2F5s
5GEn7I0np+MA6KX2mHVOpp/rr7DARxDauehAs+F90oYCQatVZ+mPm0kCzUrxGkH8
zo8svzgT6lTR/6GkrJzitC+z7EqX6wIm1zN4f1lkcLFOPWNJfu5lfn2e6PAw8VWn
aej3iQ17PlF8NiDxhXw08VtLKLST+4LPgSmZ2fWRGdno3yk9JKFRQimOMFeaDDCm
CQ+lpxcuC156uJ/+Go6AFK3AkPRJ0gC634ZVMfkp9VYT9yoqeexOTtCDcSNRfAoR
ffd1byOXgAjc2jK5Woz3mCSQEehQO/1JwgGJq3Dcxhi0W/dnEbMWazlv30dDsaR4
0YgR2nokSOhnExggNZ5P7x8jUAKXTYonvWLxAAAnjvXky7cQcFimFj1DyEp0wRpI
VrlWxxLV1cTkvKYp6hu+EleH2pAiYQrI56A1G9aHTypfi3x0yBiJtsx0XB7vn5zI
cFp7AlH7N59b1KL24t9PepRB0X7alZqldEjcqJN4jz1WH7Plp3J67ke5Hq5AIZpc
Ldt1E6B7c4GXJqBUsvc1c5+jUQzVAbQ0SAZw8x8cuEkxG4J0c8bR9hwqFuWA6XKp
NMYytrlxdK85x5f4XdFiKv4BmyDdwav+ejwxELWxngZH7WVqpQ29XsFsYqpPjIT/
odmq9aM8c1m3edxB1lGCDNNWlU93ClooL6X41TE7knJl5lTLy/0T3bJTQgtywecd
4pErLKFWZEB+KarZqXvWuUXnW/h9d0dpHkW6qlPGEnTb+tu+CyFjrQqN01FRubC6
nIpTMHHLrB4eTOROD472ANdrQZcwYfwK49DFVWySNYUW0e+cXL62EEqsInDcIIoJ
P4xXpimY7NQSGZ66b+WejWXEpdXmeLwV0q2cxZmyJsNNNU4ruZeDG7hHQXEck4Aw
+jl8UX+XzvDOxtZvGdTUW4kLVLm35IeTO4+nUHFCbgg4CDK65dAlLnUOyet3hmfL
P8BVnz6ehlsH+i74uTTRawZhwCr78zAOwh9MOWpPblAmQ+M1Joyw4moziz/E3DFR
xm6ChmnP0pwqnFGDOGDGou5Y3W/5VTf5MtQwEUoih9CII2teSCU86X85CrkAhndI
oUfzzB75S6mRHfsrvEgM3RgzrvfsgXBCfWjZ8Tx1m3/L6dubktHn+8VRLJXCGXZI
P0tVQVevABZ5cU3WI6EJShs2Kj3cwXmqaUue9m3oEcB5UumecSttZremaQjyG7Wz
HE3ni4QlSKd/7KEVAkL2RZYYF3olXhBJIbIGHWgVk58FYqm30gUsYlNHO+sfqkVh
pM3vCRiuvy+u2tSlfYc9w0Qp7NU8Xc78xTyFjKSSgLYd0k0XftFP3/9Fsh7vhvI2
T5TYSuwOHV6eZXf5CRxPN9pTukGqXlZP6P+iU5qi7H9vhhpqQ9LXh5RMxqhbnMap
TdAk4OvfcbK8OacovM74MhxfJrnpyTWLxNDQw/1qH2aCXTJzYPqNrsEbLS7eCZSS
HtLGR1qXCtVkHpZi3RdJNBfbrDrTUE3JpQpSHV31gdHszWfG54YMa9UmDRJMIacn
IQxITMrQ08YKKuy+airfBydgBtRoZEf/meUBO2Rotwku7rUUC3LlXF1EpVM0m2pp
sWQj0Zn5k+l1VYM1wVdZiBXF0jmtNtloby8peCaIKk0URM1ULPuAvtNEdNSbM3f9
fNAyDCXEnzqYdpntS7XiMNWtLnbniuayy3xAsPRmZxMwSN9HVwxITW0GvA+AlpKP
I+AwlmyGDUDqrrvfy16SMVqi01DA5S2RPnsBE6DOEi9P2oy3gsgOMhNWbLkutMul
rBbYaCm7p1WvFRF09/9otP3ul+zmdjVnVkV04/U8+WdR0zIjSemOKs5yxiPx0RTv
gH237Cwk7eaxmXzNhy4gf+SD1r4Tsk06fdJSl6medqEb2H4eo3j+NwJcW06q8vnJ
8lHb5go91GDD9Pvzbyb72MRhTT3rBSGMY4erBuKK56S93rPsBpZpvkfkkO92n0ex
3YxJaKSDgXH5b7ylTJGgAmgtIte9LbkdJOCb5OcBwRNVRi46DStjDXKz0uPUnAq2
ljYWCPCAgeDR4pcDLLTKXMLRUADvJ6evPT3t0jmp29ZHxDS/eoypPSdRycNtH1ZZ
pifCVpNwDnFhrk8qLK8BpHHNyAEyIhO1C0KH8ONv7r8c7heQhctRCfIOqlz65TUq
3WRzPX68S+htJ+E1FS6SiMk6mnuOp5Eyc7iTwkjbGmYPXJ0XMWCmvCy8H8Avt7WP
MUKyGjho7QN5tSGto+Ime2n9gHSlUL9BiZgOUIUX/gai0f40mvaYaE1y7cIV5vF7
n1vGUstywRpnxwVpPKjkpaiXLu17TLYc7UIFv1VJWMzoUAt1JoXsuNyMmLNBP5mM
mvgpEuEvg63fWahriR3WL1k9uiYvRImOBVHy/YpwdHv1nP1kLA5utwtGXtUp4bUf
94Tt2gnHITvyMYU85wTeAxK8xcMXqRmBowd+uRNlyOq2W3tn83psJEmS1EnSTrJN
vbofGTWqdR9rrcug0ZRuXsrXfuqiADirS+UKkCZA1CUIjwBebCwEqVFpPIPsYSXo
yqS9OcZLcGDcc8+mgt+EN0SKtq4CeivlR8uGnhyUObL76ErFyxxq3uEgUoIdEKLb
Yb9bsDMbWXiMF53N81up22IjrUVDqodwB7L9IdLmxXKS8ZHnNPaCOXjJPLPpWU4J
Pcw865L4cxOPiMtLSG/zGw4K295Nm206ehaj5AuQ2Vm/9CMWH+lyaHDvcd99bY3s
8ZarIvzX6WO3YHBsDJo48jSdWDpDCZ+OzO4lbMZDUWdYUb7D/USZiltr4FRtAoYm
HglTAWjoPIsICFQv8/keU0Y9dEQO/enk2bL6TKf5MYT03L1DmmejmssGaYPFH44M
zFmNUShEjNNTKcIu0Z1doHEgDNySjMcXUY96i3rMYFIf2578Qs3/vY0uz772/rvR
2mJ0OqMHNv/99RZuEJR0L0oAFAidlZI4+sp5YlEWBeiYl4BZr+9pCP+f8F+Khx5B
7EH8El49SmZTgZR+G3wdDde8YSBFfycO/CmZRfzEk4qRdU2E/xNN4uLK/MdFVR9v
oGIs7mBG6Hd6AuBuvS0DlC/oW5eG4crSlAlDZ13/9J8iFdMJLROSO4LGp+lexd1Q
o4wtBjGcq7mKK93ESACYKgHKsGwdi8XN6StAPXI1SSUIs6hll75qDC6BobxahAIO
vCHLxlVrGKkTEfrNTBBhnNaqzmuEkpx8wgmfgVhKQtvS13BcrYH26hPrjxR9izgs
6PE10EvwB0f2ImtWuY1dKIxbl9lUJaXEp/VA3U7R1zHqMyNF7Y5NnQeagnO7yXLc
IQZ+ey5Se2SvJ1sC+X0ShTVm7Ew9CAeN7btmiXgt0mRDrj+MqM8xGoW5GYN+35gC
dHk18dIrztiPQz8DvvQxv7z9+Efskx8bDsnpgp543Y1rBcNrw8XIRJKgN2u2B0My
FWmxWAst7fL+YtLEyEfFmBQNu/ikfZN9kV4wY9kOtec36EF5krpnbV98LzGcTuJ0
yQnJS5vuASTM9h8RelEkqjSDwwd4OQstE4xhwWeE2T6dfl7Cyla33xkoTWwsRmB2
tsOiVolHpBTH4wR+15hE3+fVNaHQcXJll5wuGkkjCPyphnkF6QKnEE5PR2f87M5K
/N7jO2O884H/JWkemUwg+NrhbAbSZ0D+ZL1O61PYOnJWirY9Lv6hwy19kPMAMv1z
9M9z8y72baYqQeIZYSZT57DMN7m2DvMoL8imXKNhNEAEkP20Cv1wzKgTPBYhT6X2
1GD1lMNB2nj+sXMMEgaIFcOKuMxn64hzZcAjAvRfLxV5Pd9sFXDr6LfqB8xrxH5V
a4eYWVFrb0ygGe1nm2R8Rox5GRiX2kg4c4TDpZ0bLCILdN8ePE5ygPEt/hUIWBm8
1OPBL8s67IHO/shuiIEFtDK++r6aonBAHqYJfIsdEVtLs4Vypy5Q98DYynkcXxY0
1MuiIHc2JDhCAjmYpHKpSD7Q8SBebINOJWZi6/HIxwjTw+dPkAFdrcKVlbj9Yq0H
GYn1BO9FKInDYU4TEDOgJEYEeMmMAqSGcvxuEAPVoCfnbvY59WnbJ0wHBtXQT2aS
L1PY7t5hXm9Ev98Degs+lrPFD83LQZjSFuYcHu2vc62L85WTUPyuePQMeEVAxaQ6
84ZkqgevCrBVP4ebZ+G/03xc5XzUFtSubrFpJdiwvtetIJOpAfQB9BZlntLupzCq
84wtzcJeRjltUuA7Nw5aE4cvg1YTFvqGProJFrhD09l3f3vh2YVL3dwMZrJLx3By
uO5nuFU8qNUu2AFeBKcgHe+hnqTbRW2U7Ol+4PqlaAftDKP2oq9ZF9wbVU3MLRu+
Pp4xiS/OjBz9G3iHqIuM92gtBoYXWS00uoFro77mdbkKkO63IKqqsn5it1+WhOUp
vq9a+Gl/+fv/BahRazaRq5DyElkJUkRW1qEXuG30A8hw+Uo+xgBeYXrRe32AJy9Z
gHogBxrWbAGcQLOrersIAGR8VXODROFmkrINyqHdwu/AKuAif/HgJIBkx4GmTW0y
ZHCeozdCbM9/cYWHboI+6KG+iZEM8Jry79kkXF3FCxLdqTiRCo7NdgCj/6VdzLEy
LtqPB+4QbQQs75oKUNmL5NvHS4vou+z71MR4hL1xDcW1477NhkbflTS7AHJ2r66H
S7+cIwrGmwrbJKsqVsS29Rzoj0aNOhmyN9+86N4CsYY7k4yZJiGTDSHLPNGnSjLM
Shp2AOsnHYrXo9ry/Ty/8DDSlb07B7q3eZften/2aHw4pG4Nav3Md0QoddpF7vfM
ickTr3sFIB9Wr9wXupuIwGcz21G757m+BFZ3ziKerK5FBVzD8FF+Em1m8KLosRJt
1NYiGTpx2h8jTmMIm+bd+XA6sZ1YsvWD9kvLLWRMMnhNf1JaAgYZoK+0SuTs8iqK
aHaMDBuJNV6u+vW7+zyCrXbQT3hXV3ebj/XJn5yeJH+iNwHkm4+9hRI9h10sSPOF
uCb16tqR+L4kshBfRimFtMz40kpoH7M3BJ/ntGKHSwc9cQtDrLclvTA9XXHVdmRh
+u/ni69TEATxfoYp6GakJphv/lT9/xr77ybotiSRj60wZ0Oc4nlx0rVsqZNzNTca
sYc9aGPImwUqoB5MG88oYWKzJkFhFUZ1StsY2ZGV/XdYEai+V2wURw2UVBkcTBmW
/tAmNFvI1AqTRzZXV8edi1DlwkSa6RKhjAGIqy2b6uiqZ4CrFTPo1CxzpG+5rjBk
Z+xannrizS94t5AoWuaMXlxv55t9yBJvdzDML4eeMqoEqusGGi0yhv/0W2qR42fF
u16OhW59WCVyZ9/0hOlpHG951S0+rKOoRdTsfeLa5CPvEu/mxDeESgcxbgDI7jvr
5Z5jKzUzY4IDilm8Vx2LG/mE7zru0Qh57WZRbhwHq0axIQ6drGii9mQBaXxAq2LZ
IZKKCI+sD5nOekPuQGMMHKAIXtSlY8wC6KIHQwVJcMiLvRoQ7i6VYKUFVA4tDnVV
pGx9b6bQenRvNcHpf7c0V9OLT1o2skt8fG62Tunh0jHcNI8PRf2utgviqBcq2Jzp
HTYRk0S2b70ZSJB0CGUJwfYMrGamkBTmce/JIz75IOnBdZaXc5carP6ltbMPHq/E
ohQEy13+WzcKNDqPA5DcgrsJSR0kksVLTJKoLTeKqBQn8ODEIqIcr8OzZClbKDJL
4rTnz3AWofvD2lzGenCxfZd5khSl9bdLyJJQ3q7sqBj3YA74emEt1caHwpgs9tEQ
z3Ge6ShS7tYV4FSBFLSQYuH52K42BWE11TnZ6hyFYZMvgY5tsaMW+35X6x3hejrV
UtaO4GVsn6DiCsYn3gCWC4b820DmH3O0Tp73LcBbKjikO7S/dCgbx3I3aRv9GgS3
F3YOiD1hWUzAitaVm7711zieGpgCQZXHSnzHB0j06AgFwiRHCvZ18DzidtspqfTH
PCfFv+GsSm/dyhysXKPgYV+AvAYoA3N1FdRTTsHZG2VyJUhQwFq6aWhKomuAm2p2
24n61+gjioJIwnQmZkSckTXCst0Nv81osVY3qRPidZ896Eack6kL6Lb4UJic546p
2Vkw6JlqaJbknpsD6cZDl0+um8eVuwTo30Zlm6PCX2Eo8VAw7UKjV7hX1TDVk1+Y
/ztWovPrSSdH+VYZUXBrzNnW00lV8CR+5uL5j/RuFTro1zVX+2TZhcDCJMxEQSDr
6z3TptmzfjSrTDhvdn2Q8to0DC49HCRsVxydRutPNrPoqbmeYAunXecVcDS9jDJu
T3WC6jZaGqQMw7WRuhnNsCqhR91MBCh+Hs/YWolCBmfPkIz3MuUb4wMfDMTffw8G
sr1ozOf8YAVkk5wu4bBRv7RlAH3j2aG9T/fSRDitdYXmsduhhbKY8WkLS3OE/ri6
/m6IWrKytOGuipK+XkyddtzjATkY4EdVPPghCrvWKZXfSfxivSkLJ2amKn5sxmux
7LTMr6Q2r3n+7tO6/B8eZb4SIkxCesXIWw15O/nfaQHcm648oZqgdsRcovVVeauE
eGZu0ibo3YUNPAyTMpE9zzxFiYUe7jVzdUw/d8ZWlmLhlU6HgUf834Gg7l5mFdlr
vHbcFCEX8dXpDYDysnEgWLjWypyAJbcOWL13PVTZdQ7ds1P6jVDssWgrC0SZV8AK
3vXnsLoTpPaoVypwAkDc0FGRyf+i4DhsFzZusF7tgq0tnQCMq5ku4o9x+dG7ynR1
EEpLAqSyywmj8fIqhq8Yn1psxOT3HKko81XzCylTh7Z3ucCLOyU9D5v6UuTL3TbB
46C/bCWIvTxvgpHLIyCsrVKFwGgSbEUUb81MqebwvikzRBDJFFICl6QTfv8r0nts
3f1yk8KPYbYEhLZoPJXKINTjymgPO+PkOJH1uy+Tnn0Yyo8JCRfJRfZRomIcXcwd
za7DEU0yKBTIIICcQETk1sMkys829ZYniSc958g/TFqaihPbgzYLr70TIBj+8KKO
CDU9boPy9LXWVf/fXbn2RKZTJqDiY7TA9eM3Aa5q98d+2SZrH6ecO3PGU8ztGS3q
fC1YCFolXkgLejLsLbfPUQY0CKXSjmZb5nD7G3eucmZuTcpa2DiOYtIn4S3vTiZJ
W8esBbsJbZI6vdV+iXms2vd/16dFwMFNP234Z/Ku1kfW1AVuG9qWU4qnqysgTwyH
Ujqm7XYUNgx9d9vas9qwKr89YiNZW5x7ciwCx2MHV9zf3YH8+Ft7L0Me/a0wR2BD
9iQvG9G4KLl2JldkMpyheR8pWKiVLYQODL4S7eGCWnk7q37KPf0Y6eYKj9ahYJ+Y
B1yM3emfp9Bwo/M1uOF0wsy3o37DOsfdhuHMK/eaympE+z8NUV+gnqqAqGxdy40g
VEnAdW9oUQIAYHs+iTkUSfBfj7XjCTI8o3HBg2PvX/7CX487f2DovR0uTyKGkzXi
IkfNqwcBvEe+uDWQjdkKHU2U4bcmP06ApRX7SWXiIv35h2awN/IoyQRLcRZmNXUV
/XyML6bID8BikZ96q/tMZyALYo9L6LAvTa8BhpmdRRnFg3jqE/kotEKVWA+iyIbJ
ehLls1lT74vJP73F7ZcAaIEmqzM7hQwU+ifDzEqDE2HixNvdAB/rzN4zyXdjyT8b
YszmBO9NLqxAoDwgH8/C6cHHs/QHQ0krazgQqgkimLvCB2HOpA8bWsi3RfPsfjMY
R97sCB/YbI+OYwe+73ZFSEvB4M2A6w0PVErehADLPm4IjM42sbl+nyrH3yHTPhyT
2K4s27yNZUgVQeu2GVAG8CBL/Po0l4tPTRgRUvpCQDcnGeOXJfDPEK72CC+/V362
TJ5nVSRGGOkfEFp1vsW6PsJSJntvxEqN7R6TaD/rQi7f4BKlL9lhbAG2Fw328myZ
ebJoY2TNWNic4xpoRpO7ffvaTNPZtDOz6jVDP4mJMskI1JSCNHhFjLVazWBvxO1E
G/9rWpIF2S5Z4awZLaJDh/KGcV1viYC78ktO+Om5U3ZML+mGCZuixw60BY6kJHNG
xV/qXi9D8xjPSVXRXxORDYFh8u0A9i2wSAoSTxesEjX00CHD7oI9kFO1LSCFF1Ct
gfs9Ebf3bIJzyYEv1YVdQcITT9caVyvorYjZY3Aur2mYQww4LGAxl+8xSV3dzW9b
aHe0Q+9bayQYoaGBuhZsuBFECC2A9CEB7oOEezJShOX7JN7rvIHTrcWc5Pz2ixXf
794u5chdfxsTBp+BWnRpGFGlQOSGRYe8gU/cIFC02L+jP6gKzSLUn97WEE2Cjb/o
bjRyddRiSKS6ZPFdV4x99lQ6KkTotclz5Ad5QB3eTDdtpgt/cnfy6TC6lELHO0HP
RdjovmlRobkpgx93nVFtHQ7LhANdi6VsguHNJ2McOxnJTKMKhwckADwvHt9gVrb2
XTl1N9kGjKoGy2dD39FF3QOY6SSe1xPLU0zOuLp5JVv7n/5VaKk8PURq2Pw0KgEz
WLPN39TJn9lw+xx7ZVZTi2yo50YNoe7NKAkkIdDAoak6NzZkyd1OvijrM0xgfYNb
CcbtHaNuikxq6W5Nw80wQIjaRDjNF6kSPKgcvB/7MsIdP05CTTLLFMQ4VTqB60qW
mo1y2WQJikvKtfFSy7BHM/FmCNtP99K0x0sy/oZN6qDxPjiavT+WPG9Xjbt7Cm02
xG9FUnN8Cy3xkek/H471W6WKmJ3ZFuYrpHdV2sU/q7CcuZ+QzN5xD0Dms6EBdI44
/KXvuU9fqTGU04s+XZhPWkL8s7Vnd/qF5DcKXDujSf6vA6Qn/QgQWG+EJpfbSUfh
VHW0N03s7IT7HZFkfoOjzRppfBUhNofl2CwHTd/CY04KEaRfb9NGeu/1nngbG0Su
5pte9n7mA2ifwa+AzUAOWjqHVQAzGnWKPpWy4HByaZIcEcuuy8NT/QoEAQI3Wvvh
JktgthuxrEuNfNKVuA7jeGen5k8mqqCk/zhG5J8r1h9oDDBir5BmIVYrfVhRr3l2
hmgdXq1CKaF5Skhy50SudqOIfiJXbeWsaPF5MQJWFDKBueJknDVxztsUERpKI1U7
K5WflF0J7sjbLuXfetFGMaLSQYUmOlyyMwFJmha64M9247725G7/6eVeXKFm41bi
h4PiK1kaDoSKC2hYeqKfDcfvie27XD6hY8kljj0RJF1XR41Q02+5awHcDPMtzzYU
dpquMeK+rvOvy92RtHj4Qyvngl7SXV025gzqP0hpwYBU8W8sqZU4vx29vG5yiFzl
1T7RLSXp2g0oLSjpcbtk732zsey90+7taSQhXyOKolDfsOggHnD3UMeiJXLgU3n5
Eq7lpufB+Kqm/Zm/NFm+Bjgq03QZ8nYAgGmITd+0kSfgjWjwUqnmMhFX00h9WtLb
OKBqfsLukKp4ezvaCTLz+X92hJNZ1HquPYRT18DlYQ0A7I0g+QH6v3rKwnkvUU/7
WcEWH+P5EAKmoQKVDwgOcFeyeGqkpcB/hVXUIBdZOLt+zAbboXgwne6ng9r2R1WS
5tnvMVeMsjsB8oXZyu/plS9PqXldcRk1muKJzOqdPFL18/8e8CqJH+I1ikfzpRcB
SbQ0YJ3bOpvIXuHtm5kz+ISR92ZsvAnfShCgpyjwSq/c+IusquzVblhce+xt290l
nCZ+q3S4gEMZlMEgBpTa+DloATcK+mnaNz3HURf+PnkGDyw7XYoaE8vV06sjQ+n4
FsEkZSCYypW6znVBR9vdvQB/isKpBXTJpHckaC0nL4fIxMAl3TVkKlh9HlTak+jM
3zC8+eGR86g0pA2p3FD9UdnaiRZilMRBaee2Kyn4EJtpjCuDk2ja3vQh1wMyGaW4
nuHbfzGGAgCC8Th0UDIRLkkJBzJCeW8IwyoNB37sy4WsjFPixDJp9YQqbeZBmwG2
4c/7nT5yXz77wTt4j3VXg82LEGdkdD8FCMXFMh0c70FNOUuMdwDDrr57QNIiE8b/
MsLHDeyE1DUKmMP2UsJhky0IQRIlaVNllX0QX9FnvG0VGWBeOzWXGR/X2ncAXhSo
WEnyDilQ8V+9YcROm2U0KSoqw9/Km70PCbl/JrC0oPl7Yj+9Ycwr4GdiPxb3TrpA
XKP0vxrk/bhqjlrP0OwNCEyTvZ1Q5epjKdxfgkf7r38KLbto0NYwkFXAH68YIjWC
Q+GmXt0K4ojafuka++lp1T4ADdNtHavL4Zps5yuLEQF+5tYHgfB4lVuH1/ewOV1Q
IfElmGPBsD2zJ1kCT0oHWZeQoF75ZTGNarrYFXAZSUpOpjNASa5F2G3NSIiYrYTz
R8ZDOCDYTjTuDTb4JtLzulEQTEzXPFI2PDZ10w3DzAOK4xrkRgSvpT3SW2zZM89h
0Q75tpZ2uTarWMkAwZkuGAwIVz+ectKOitb9JgqX8H3OGYFEcw4f4clp+FyXcQMX
dSDHv6QxSxhm6aYqLBZXs+98FocJqpvKTBkJGwr3VDnmAkw0r0HaYMsfD/xRtcVr
i/be2BEWTHx6weNmaMACNYlai96WRKBzRCkGv+O6OueLgdh7O3e1/+xof1+21txZ
v6xgzEcMQSwOpTJl5JZwshqrmzeoYULe1kbYX77DvUF+M35lkLRk1zjAQQsDL4Q2
sEhw5Tnxdv9HPFOH25Xaiw3orQ9kHg2rciK+q7UliF6Uxp7+9+3onfp2HG0dwHF0
5oUUB9Oh7LdZKW530uSFaQaZlKHzDh/Yvq3nNaE5JN5Nwfmph2sZ10whcoeikqU3
ugUPnzQ2J3jMT4KNJV/8DgIzb6px5x+Vvzw2uut7KS4hUIaQvsTgoqdOLgrCR2FB
/JFHgZbPf3cOEvaueES6kiGOPuxzOqO6JjAboEOhnAlTSFBex8fJ5KjH4PHyvEdu
SYYsJiI9DjkUu7KOOcdNflN6CKmW66Z2r60JXwCnO7uvkW4avBjONSSMS1B+IA1I
R8ib1aZLn+NetgtThzfp3PtSvgCN0aMt/C40REQvejD9ZMWdjKogL3aXYFIBHoWE
e+dk0UcpaFDpic7IHp4UqZJ/yA+RNYFRx4C2AaP7SaxjuCt5cB5Od8M7vQIXttpv
n3CBzmvkD6NhrXRRHUbkcs6MlIipUzEkTlThsSpwTePB42iES9KjY1CxBVXa6Coz
r5/hnhxea/ZC3gL9athzUHZ/GMITVgTBGt0wbXn5bu10qSpf9gwoNr6RRMlG7diD
qI7F7o0mQLOHo4kGNoRl7a6xPMtLYxccbKXJ7unyMBzu/jkFBkUD9wfD6ygocYU7
1J7dkrjALAf/8BIBj6LBF1soa7F+aOfzmJLhx5FhBC/i5aU9KfhJlBe96N41KvkS
K2tn3OhRYzWeJ1O2A5eVkBvzMDb8VZCByMFSnyV4Y73XW0KnTCpn1ZHVDv2Fovbp
R56dnfr8llU89VRxHjRtFki5KKfom8Jar1kiqWLoZWjTAUkIq2jIfMjOTHXbApIi
3qwi3E2hx3F1/1vo5eFqFlVnWcJYwjI2ApE6eqSKClIaOEoFvD6KvTbgTuRtQ3N4
csqp52qknxYEjqLhRGRc/SCzW41of4bejz/rXQ5GituKlQrxdbNiPbLiEDju6Q0x
7vzsEJ7Sfx+pRxcADnwe2/hjVVcACGoMKINXVE1A5MiVmdPlTC0eDMojKJfH7eJz
SOzGIqMpTUZuFcGjocpMh4a7/MhEBjUUuxrksnx9/ev0rgLfcRsviaal9HzObgPW
hgcZZnZq1DJzKu0Yb3G1SxQmzDbKSpu8mlMuCgqNQWDOpPmU5f4gbcRa0L/BN23G
+6SFUPvhTUyO7k7ekoGj59/4+9HM/VAh5ULzHOiCj18GJtg/POdhBCCAkFQXBRUb
1ZHe1eMa9V6tGu5p04JZWmTPQZwDSdN/nSNdX+Ojcm3u6i2Qb+DSEax0A2Wdx8IY
KCBEgeDoAQF1Ed3f4T5z7+07PSs9jmt7B5a4T+Vx9BcUszKCzDTfJIJz0sNasDWD
RGTuvKHW44PNj4O0IkyPETIUQ/dczZf11ZiVnnNaN3AlWny/1iPiA7FUXhYTRjAg
BU+KKdH3E+dW5pdfm3/7/mpUJLrEQgTyp06593IbwzzGfZMcf1mYAd5bM/WaZ7a+
GNMcay/ctfRDN4A6s0Reakr1/CPu9H/xFBR8lB4IdRiYcL/+jzL706QMvbNnXdw0
P6GkwXgRee/UGRQUFXpO1VG9f3KnNo5F1G1gkA8zDjkFl5hBTjEXv+m79xVbFxwq
np0aMjAXZOxsORP2GrZqmveK8qLkLlUdtIgNJ0K2GCchgL/r5eCkoAywQn6wMbXS
JpIXLTAGOtmH6AfyVHEEYYPKjKcYE/AQ32PNu0bNnbp2gsEtv6BUtCoR9NJdRPcG
4tCnG1V7pIljCWezAzApiDTzqpD5MxTaM2uayG3twCHfIlUWaZevlRU0KCGup77i
nUv6zbyfgCV16zIHr3mgl7Lv+52FjF1If2P8db/0GY76gWOCGKzYO3aflEraGxKv
yTJyvVYwJbx1NmGEqOubsPEcRb74lLeVw3gQGBT5M/i/Z5cIivndmU5GpJjrTWYM
A8E23FCQZ+YxrtBmeYFniW10JMlEZwDtlw99PjQLiM6JxIyFLH5Igt2FGpRpseDv
n5qZ0Npw4sUOi9fNhRcHVoShYITugu3Eo6qqn2GUKgaEfDe+a/a0w0GhhuQOXjVu
HrNS7iG+yIG9uDob+4cCMJokOlwLVrf8D+fx+KpHyJQs0i5DXPF/cW7TJK1VgWLr
WHsu6fZkBcxGtDSx4CIr/2kJDhM+ScSP5xCcEvbTYMFLFKr8UbVvZeg/t41Xoqad
v3m0cjZRoIdsn5l6OsTfOK/iCBlI2H5AzbMZ+m9FDb7Dz0LUMC4ufHE4NlMBuRy9
Ypo/XG8wrydzDUgYfBwRtKpNnxvWrMKKCteQ2eX0+I7nx3SrtPFzD90EqnJiG6UL
cDJkN2t4W238ljS/byzjWw+TPvLBg6f1zl12nv8/GFaW7s1BKD6q6Q/puLy0WpFD
ckR/AZ2ndLR4J19pHNua3vhAn/vKR9jXY/cLkTPLxxJ5fU7B8HYMOQa3Y+g40oI6
v7NdIxg2ERF1NtTS1qz2/arbT6Qj8PQ2HDfP9gaklTODuKQwlTFhyl+sidGU82cP
JIp9kU7Cms9mPuga6DL+1+XD4cWCl5S6bGPBKc3wnbRhICZNwgvFHUJaEVG6RqZd
SuLBqheg4xOr587gpRqPIve0d4gswP0pRSFDekUxtjmqDQ1PUq8BKFuqfcV1Qw0Z
/p6zFik/hP830KwYyRhAF/0CRcwP9/Oinz+GWOYGPxvEAC5t40oG97R+FBVPTQbI
W401DyYxN9/cfH689gYq3aA5iDLeYtZ79IW0UBHcnuxV0OqJ9z/nrhETdigyV93I
DQcDfbT77dRaGT2nIYBtEujyNYuknYBQdyNiLUZuVWR47rcdKykoMdcd509VG9W7
5G58nEBVOr6IHSRrUhqAFblh1HpdQAKRR/vy6PqBmAT9xzcl3j+Mu+1IX4H47lxA
aUIG7nG1Bzj5wtbI/5tXWbAfh1ugTQWqwAqmX46rSNU6bCi3+fgKb2f6fQCMN7mM
A01FEyMZ9WsVfNqUFsihaUEzA8bfx2Y6X79Jz7hKA54BNMUq6BGwBsjUSKmH60Zw
14/m1fEmbUEDV2GwxOeow4aUDMVkDAunnSaFS52QSPAcs49TK4m3jlgpMlrSRkc/
yrs47RajLfYuI3yPcrAqe1+sygHUP7+uPoN+JwgVaw8j/uWp5dN/tqZGSAuURFIk
jIXlmLJB+MueaTCD2UnobRo/TcCn9UyOmMVrR8+c1ukRyAMeLT8bflt5RDlj4zVv
nW4Kno/Lky88CMk1y+6Twg==
`protect end_protected
