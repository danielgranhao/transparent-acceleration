-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
R/YCSGX5xjOfyBtERhm4yH1/Uf3dQ2j75c2Jg6gPIxBQwk31cYPSh8SRmxm57RGUxhShx/EdhNFR
mJdmQru3r0Rn/7244O60U64gxuflS2hQ2Lo3GMRJDUZ4Ds23kI4L2KoC50c9g+icGf/8Ruv8//Rs
f10C31ahbJZqi6CL/KpcIaANljJlz2Io+FIw+HkZ8HwMy426h9t+1zD6TaIMv/PXbWsg/hw8ENtp
xUpQ83qBtpMu17nWSY6BM+ocCdAU7LQt90wP3pdc/vNZou9l+hPx4yyghO+AxBYVnpGisQc1bi7m
ZjK7lgaGejPjFP3zd5+wPuqvk604xMBsIMiL8A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13248)
`protect data_block
LcGRj3NTmHu/ZyJ2fzquaSYf/gATtmNn9R/SgzOARD+iNhe4dBKs2pfttfv4OV1nk0X0QX79f4bd
pLokTY/gnLwpymAYkl+J1u7wvAZrvmFbe90+GnEivq5ybLMZqXu6I94EJJdJ25zn41ZDNVn4iRR/
qs+OurMCQswanmyVk2geUk+lSPEun6r0X/pEpn3aNnA2PF3c5kTxgwJZ375RzERmmsS98iD55hGy
VvCeNeliWAF55/eweKb75wHfeL9fabYxxf6QAXbOIcAmzzC4PPm67AljKFricWoW8PamlVT28s4x
pvehMaB0IJI6v3q1djOII5FBWwwFAnPZIXSX10dpcAYtVQ1amlGrA2fZfRl0ja7N5jSILVns0OaN
mvlEPYtAQEd/nQ2P3GiNjGwWRtZB3inHgwfvLonvVRfNOSEWk1C8V2rM3ostjMku/Y9vvoyW39XM
HKqmTuTV7xwuMVDlSr+NO63anOMNh51ImNiWvOs6MS+Gr7PcDyWCnM10IV7MnE1PdVZ9rkZW8NRC
rHbmQUEEziRnZpt/BqRBzd17d4HGnECuyOG6o7YXlyhYMoK7HwMQTaMCK/HmwIP5q7yAHR2CkM1C
fhUT8XQkZfSSt/H5KoPMnBMfvFzeT0SIBUsUn4SU5P0AwxrsFtTGL02r0u1pi1iufgdUsmo2YlrX
t/DePixYxPBEdwN361st1yq5l5IP/3wCNLqMDwCzCjnVWTisFXJjb5sWH9I4jvP/MBDv2zMcvpNu
NVHtd62GosEEozdloDqi0IsOeDAtYm+6D6vSiRWArOIcf1ETGIvQJgZj06JlQ/ZGBlUBT9NLoaD2
iiYoqZ+m6fR7ruD6Q5SPfe5qcyFcycOzWehYIuWpt46KGb7a55WDhLiwG5gn9k1ivz1g9/Pzz9eo
2k69rg0DpOq5qXgoc10Ax39nGF/4YZK5PdLbIfqLMAfxaYOenimQaX01x8lN7qeAmDPvDhsTbjtP
+ATrZBGvboCI6OTLCX8iiPPgpfSibuGfnvZMpV7M1hPxcOEZbhESAJxnHM8wkzxXV5bC87iw5SUY
YtyvyCNcNQ+RUJbT8nJZCQ3LCgK/bjRLLGg2qSNUuU/7ovux+9r+ADm18s4Iw8fH2MhYPZtJ3QXI
tIf1hO2uuCEytFCPgdVqRksjwzwTGXOwPJwtY0L+PbFxdA8zd1AlprprN3whj8SXEsnT+afLs2VM
2UkirHl2YzSPDABvyTtcXkMB228zn+pxaF27x+BGq94dZlFjP8BydO82ursFkqB0Ncott+lEm7C0
b+RHBSsU5m+cTYhUQKpjCeFVpy44PXV7IuUGutBEovZFMgFblZEH25x6wXx4bYMuQ/kqcdtl5i1z
pzZCu0ntqpSwdJUjaxu+YcT8n99JbRnoR7pcPlop4scnEs5O4wQ4jFiI59NqiB77H3AudahJLNOv
5E/8h8zl8d/GWuFFbIg78JhX0aBopQmwxbfurN4Q4x80LxuGunlhK3O4VDvcAfdFp8qVSMxvfRnx
/3ZO0QzeYRyqY461aF09/4BRvKn7E+2CXhaJwCrhVH61UQafP+zgaWl31L9W7vXiXs9WS9ImoOfa
Vj0Lhn3GKgGQ65xV0863cEjNBmsgUbRTnEUeL2tYu1jRC/qDWJ/oYyh1TnHhDS5dqY0zQxDbQIwb
1Qy/IAv1jaC/KF3yPDM9E4Ix0EzEo5DJth+yDoVZl8yyULtLgPexZI6eqnvlgWFM+N+QNbR6kACY
1Mj/tTsAfBg4iKsmg6KNVFW05c1mNqFgZwATpNQce+S8toxQaBrxcV1Oa3aXpecVIFdGWU7UKI/9
M9KhZa1DUQfS5KU3ZcudfrvFceiGizMgCPbaaMa8777QsfNajA5Ccpn8SN6B/NpinEG8J2Niobqq
YV7CxuCbAwcpl6xA5bgXty9iatzFz5XRa01v58WiDBsRz4p4mKlxhwRpzb3slDxVg9tqkZfQXttO
GbbWScHTSnFjtBdbbCgvuRIdFjoLLZ346NhOs0rkXVxwXZ1AsGNPZGUWd6BHxlTIq8Yzg79rr2k7
Cy3uisB+mzO00AZSHqqlY9yxArsFY/P5kb66M+/owwvZyGFmUkq36ZhtXf6vi08Z9Fm8kKkaxjF0
kg2RWv445Mliw9AAS+h39rwl3YxV+KUkN5XYaH3SGC1UQVeDOOLb1CSg7qCzcvsdFMUrWErmi3pm
yXLaUeP2ZsC1Ni1D9haYbHFnKh+gAoVAblWwZkJz+fCiH3JXxrfpXJ4aD32oDsvM1EL6qp7ptHy8
sI/M9cPElsd1Qxl8dbRoqoGvHndoqwyLqAiVhR/sz8eLLkMXmMhAxQYX6vOhdtTnF97a1OSb8iHk
JgMh2WaAjMQp0emlIzxmLJya0y+UnXE5wxdnKl0tG8THEt0F+5B3T/IffLPWiGD2z44e13aJjyo8
4CwUzbm+NZxB4Vxw1D02UAfTx6VPW8W1ARsboDC1spwxGdW0yHClv7/w2UqFfkB6sxfg/K3QYmoG
Ud7mBUAMYjXH6YH8a6I5z4GqD1/0GFwh4vj2UT1f/N9cG1pbXS2Rf9o/iDAgEhL66z/ZhcI7qaDN
1sdwfChKaz8ny3tQD4BKMoeonej1k0Dc5LgAQRlrdw0MRk1YmWUfjNrv0SmxCRgA3QjLOf/6xRo5
XLvhHPjj1hpONBQB0Cyi8soVNMCGpsa552AjhZbn+6hiLpS5L5/Jtn34ZE9keMsL3hVo/G+wN5HY
qdrDekr17kyW9ojaQD4unX5DAmz33o6ysx2VEIhvj1vMaU8fXzxFL43yKZflEEq94ULndvMhg7V9
Vt7wwZ8zIQbYRLmFzzarb3eZ7ANylz3GS7+CKoSZ+oESDdkEHFqnMAESJ1FcNxwfZS3ibnAIRunb
k1UKltyJiX0PwiGrmhCGiPDq4ug2iwgx2ISnADvXeCumpt5vHYng5z8LOA5WFQPIy20DVHd1ZUC4
NopOM//iVtgNVleohxfdByWaU8EDA6J5l5seZ4bzYfnrCzGdviQM0FlU5ONNRg9spaG8cMf3GSCM
dAk6NyrMCtcCYiLZw+Czx1SZ4M2AvILlWXHLhct1dkRpr45MHBTlqGlUJVEJRthcJnTXPtn8/rz3
2XlyDMZ2+tXDH4fAoplvc3S1IXVK5t7+VKzo4YqLXvjeKQJ7kcV/syXWuOiHlswIKAdmTfSEin1e
3gSKt9jsCuIA94fWIF7GuQT2d4P4ye2pUnRzKm/1scMGiAhUBsEXfSHjJ6AHR6GGHt6vx5OUq8p/
ZeHWyj5G78LOV9ZL1OxpGGN7ntHOBqo84fZTvq2iqTamJdx8koNdm1Baor+hQLNBDioptNWdi/Qt
lPF1VcizzGQaP7rbOcRdKlJSLNij233rgA9wE+BnDTOZpGfLF9tW5yeR+flO2ZjBazs/eyfgY8ay
PKn9pGQqM/AzPVvNnRv8zHr9rloDfnRrVcDghT9XuBkSFh/+FuN/WWdRbD8aGYGBqFBu9VmkQRdK
U2iemAKZJ4Qzmegkxi1aPYDIjJ2pa91VTbQxr5rQnN3Hl8V2nCzBa8ImYJaHLAW5JP3WhgbYjzQw
dJlqTY5kkZv7jPO6U8PZIcq8xzy71tXrfmVAVRELVdIugIBb11kBe79E8FIvHkGS6wL/p14PnD+9
ZlQNxHKj5bX4JnU+m3xdrqP3v+ijpCbVH39X9Tg98LheEGoLu2AFrD/GQkyf7wSrGbDvilErlc3W
uGtJ22K4nlagAtTPRRGSZ+ETXzhI3lFk/k1qMGK2kYEr9wNaT0qapAYx35HRRoRceLGw1ZUi1DkW
GPxOpi+ghzPQsRaFBf5l/Jr8jbU4hE3KIlyQmurMx96qh0dPEmP9jnOisM4kJ4GZzcXiYiSePtbx
BkvyZJh1lo5JEBdKVxCzHQtFvqq7cdtlTbmbi0MJbB8bVqh8BhhSthkY+SmAciVwtm8eZdBvbFlc
te8EQWKj0nFWb9kmLHcP1vmvMpYpvHS9/gFhY62V5pOcdLXaytCTYrHpy5caQtvmVHyaZ8EMbENM
B40aT9x3dYt6R8i5a1xR3T3dGbVMTM2RntmDk9cpM7SvK+i8DD58LgOQDhkzm3wDZkcXMPbWCB87
2kbrtdksUYztBv/ZIXYBkQoah1Qn30PR/V2MSgt78E2Bsz7OWOU8wUcH57yaoQdkpG5L9w/JjR19
MbVaHtI/YmfwQFDeXy1gIJa4O3mP+vySsy1yGxkmUmMlZXMDcG4yXZzlCS4A6IYMviiBhMMc/tIa
rByuSvq2NySzm/ftqJNXyCIO/BZyWTY9xyzwfwDQT3EM/kBpney6kGGvcM6B5K/falFBnazpI9t6
H9kfqEvrCcMG/Kb1pO83TaF/gJFhtB0ZVC7u+l3efuXGvDa2xDBBzq582+dEWujV+/vHlK7EiSE1
0SKi54431eqbgNidwXG5bOFY9i2p4DZHVhDEeQelIbCI64kTFX0SG9y+Tsk1eKssXJOZEoT8Izd4
g/ZjbrLz9fO/d6SRUMRF9r4+QW1QCyR7cZKuBrRAew9q50Q+fs7xV1BVuH/DabF3Wa5bKwfVkNdO
kcO+t8wGaIA/6tPOKpDQlY7SD9mnylKsBEI6Nzhi8UNRHLPxwe+n4K9iNwUO/cE9NZgQSq1XA+Y+
L/hJk8EAOxqP1lSxM5EnLY/2WXn5GMASdJrdH1wQdjWg9Eb9kPv+vEEKJxK7UWlmIwK4zpqzGTSd
d4rrge6YY4M3YkUK3VEuNioRodo6+hfjVZO4E15tB53SWpnTnJ6ec8NLJ5eGyJO30foDnTlVw2u8
Lz9xEw2lfgEkvjaeyAxw2eXj+UqILiceSvW25uG3xAetd8VMhsMfjC5U79fcVByDx6tPdhsUCq3A
q5ifZYOsCg4dr5N9pElqrmXNQorrBezH/Ag+3e3fbn6RHmFby672V+owWIBcYWi1rGUXMb81tCaT
iRFrtH257DVyqFf2OeNXSQ3+W4gjg09TMLL2kSH0o/cLcmYL4tWDxb32i/Xuzh39oXisSpEaFqbs
WEqkgxSzGu1k8BMDWmFcvhqmt2KNM0wNOI3EfBziTZOkdAd78KFLw2DvpXU6uunEPy7T6NcqccsO
CE9GWJz3eKLUzMdrJ+p72r9cihNdO00IwmO0Lhg3iA9y8THp0rzkW4WMnlUlKzDW2+g7Z17EJvgt
a7TMHDG65aLIVayyStDdHbPx9E++MwOsXqTD/QYwDst37+yjSLk+nONJeZFIkEKscj8bbrrC+/Zm
PQ7ms+FKbWe0qHKZuEJ3FZByaU0fORs7IZQz5aSl0ruglBCNJRFEiCLGG6cS5uT9sLjrwcgpxsPT
jFp80unvW1CIWgFKikTd8wQB9rHpUBjJK/CDzY4lzR+knKnWKbilFpYmj7aACQKSTzk2Buw2dd92
1qHTadDLo0HwpcrPpHRSdhR23/zd/wHAW+SwhXAHahDfAjgAF2NZhsWfswIxNQXqO3Ebfl+L9ee0
B8WwkjzX/fBGnxG852hIB1YGoR5t+/9ARdlCKGHCp8FKndFSL102UGIU7FbVtv+jWIDMbRW4Ulw3
v4fD8IubpDarQCPYU9fIodQ4/wQcYBDkxikcGWKtLssRpqwKYpMMeDIBpS4JxX0lVPHDHA6gZxHq
hf4AeYS26t44xxzvv+tXT9MBzvd/maPUThzLLiSSboC7LsLOwLGtsezDm/vgxsFd5kPBL5tiVfYw
JDKKmEbDDrVz60BzSG+GgtF3x6h1UnYqDIDtQrpQuvUVdMcY0JmDkIm+2LtSjRtlbJcafOEitwyv
N9VNff+MoubCDEFTeFHOSEY3gUIFckLwpEU64zunFWcyO8ND8DWye2KxNs9W/PIkw8PVjjFfSGa5
L13y+myYKJLRK98Xy/AonP0ufUObQR4dAoWpczsQ4ey5uS6M/qcUYtJxjLUwIDloTKQDOSG22/8e
sPIlqfd2kDCDV79IWYbMwHICsDVBKe2oa3gbUI3VFBO9UuDpNnbrF60BJDokhvfJyb1dIO1ypo+n
0CK3e4TGWDYLe65LpyxXq5TboFbyZjhUXH4vO/2rtn+jQsBhCC2WQ73akjJlMQIzvos0DH6/uGtA
5OFpe0usfDQX/gG7f3MESI/91MWbBDDg3nKG2DSOHGgNEaFdHy2RPugXRd0CFOTXkYGu3QnL5G9r
NoxXJgAMf4HyjOD8Y5eRCEyhrE4QFcJiJn6lhr1JXU5nU20YsuuhsMi9M2ARjhaEPJzzuVRzYvO4
WnvFKX9aaOW5rCunDVRONxJGJ/AMZ8oJB513dXrhJiPVdm8XE3pZe74chUzhNBlxkMCPx+lsix8l
k9nPZjUMj/Y3zEKzb8hnSvJVPagEzdmoxcEvQ0V5EAWVYZUg6s/rzFT6wLdVVsdh+Apx0F1cnz93
cj+bzrsIl1gW/ghx71/z67MpMNQMSXwhkJmTqpobd5EFJA13VyTRiiv/iVxvZDxSRzLEm2g8uHRv
4NAZb8qvg9wdu/SLVr/dr1kW4Fei9U/Vc8dFupgGwO5pV8JXHqqhHc7V8GdWmaXrao3S9hRbOMQT
L32J2LZJHjfmHxdt+cBNIGycsoN5XpAEvV1yc7mTHNDSXNEVG/VJQ4nQPofejCZKuSfqGO3HK2nh
EkxR+XqQGyeJgDkrShAoUqPpl8nsYg5+CqLR+Em7rU6M9k8/L53CYjbPJF4x2+G/ENn/kLtrsP47
oejVACO57pxFjMxR7UihfVyxKlMEp8U6FLWL92sUVd5R+v/msv/zDTNFqnJl48CgSTf4tqwCDjQq
m2Tyd1qmS5Nf50uCCW/EHIoO6OV47vHTiTOUazjlLl7nd5ETgXzu+DkBLr/NTizYvYDoKWRKpSxd
pDk8cUnhqSSX1weFLwnmkAtaSN0ULrOYpvx96HTlb4wyGGbPjD39FIDXnRMm44FBObdAp6kYR5L9
0k4+DUwpWizL+sTbUVN46Md2fxsqvceiN0IgDZ2IyI3Dlu+tb2++z90IhetxQtdrrQ5FPdoqiiRu
AGcX/lMh12TKObnZghaVS1qSFiEkHPzHScLzVFo1mqWar/ZYjyvASbPEjU9VCkwNFzJZvwcGzhH5
/LwXY+/Ki4VDn4+oEgSlZHDc1OnA2/j+6W/wZa1UWWYufzIp1E4FV5RL/+qWmkAvRBtf4AXzAe0L
NyqxcH5VvgvLQLGK4NLuBrQ0Kcy99eL7jsgThJnv8W975Jh+SFyhA4WTQE4DAMS37m+NX/9lCvJ5
RReE8Ky4wnm2b1bm+ByQyV3aURazQcRiZoK7G79YCY+qCdM/6gi3ru0E2WPzehWozvPK0HlqHAOb
OyMg5mRsSOBXdyFj5r8ECku8yoNpGWXHusv1pbvPwIC8FSBbErClELCbEcxmlQ7pUoxS2DfAR/qM
1hsMjvklS7udRpQ0LjyTilQnj9uVrDee2OBpUeVR+zKdYiz+gBOxRC2n1/aOwY82iHC/jxFcrvVf
1Gv+jlW9+9Xfa8s9sopajd9UeifnGq1HkriMnnO9tRQF/+DSaE1M10UZBkDNGREo8VyDROOGm8Zd
wd0Bgu6A+J11kHoo3O843RL8Cee6nZmVTk6lzQg+rsryu4QM7vFTN6mg84Lkx+g/6nCVg8G0Xi55
GuZnh9DwKkzK0s0Nb+Mq9+kpLe6YjE8c/DDSptoWe5Gkr9yZxwGHanlyjDFOTbEBkpbF9kQIV3Sb
ZU3/K9UEe8UbKvhmj4fwBMZkm3t1wA1hC/TH38jyySB8XmKC6UvTVc+w735/Mrl/HmR7mpVnttME
BhOWF7055gBjiDt0BhKnccLTZQtESMh+enOQDVfZKlV9JkDVdjMI86R9q3aUwJvSRxmNNYKjVuhs
qtq2oKr0q+5eEBx10OG+S59XQpknwjGHLsM0dT1v4V2tH+utdeCIjwapuKbbB5kZu9YzXF0Cg7Y5
AtXxd1iOkuDGy8iBb5vJCokfzcryyyxCttO3Oq2Dyao3ho/xQd6VsojfKfFsXn+07O/oIV+whJFm
E9TPyTX4leDS3qK7X13LOe5U56f6TpaBzxn+LDsyI6e69AGZvkRjkRVEfMUgKL3u8C8vxfHjuomI
d+n0DTfXIstV9wGx202NItBWrjTqkFwZOuYRJQ18MxUCDOrNucU09XjGoMYvBgFUHI10W80nBTQ8
pcVJHNhsgvtkumGcFFFcMEeU5WO9nWPR8jWKRU7T+eCep+t06GLD2xJpf72ZqFVxNLwEOKn7XdRs
MH6G3Nc6sHeI3YSmUi6eqsTFidv1cQpbdPtrbSVyg6XU8Ua1spfSOoytXXU5vYH8ERoa3XhGKP+l
rr8XUJNAQTMA8qCbykP2yFnVBQWvY7KD93gswCRbDzjXtr9HDTc14Pc8QZA45t29UNbt8T8coHYJ
+OICuYEoU3Q8oP7zjykfEn8pDorAwopkaMYp2othIcElJZok+R62NghU6PfXzJ4CatI2IqUTEvuY
8Ccn6dXffeOaPgOcbsBAj2h9a48e/mGx1FKPBmD65IOZtzaOlnvyM6obeOKcJ+rpZpKhIZ3A71UF
h0QbT1cwLwl6u7yWGIOzOzJjILMT8k6U2GYXt9my0hnrbMgdO3ose9n9iSDgfZIOUCIq2fcff3JP
baZkZVCUhhCqkgrz6upnTT4vgt9r2XGPTc0sbd/nT7lZNA5nKG7WJ4qTBRoNLOqgf0gdoQ8HFiTN
fkMbesLqo2JVFW3ZYlJvG2jnKpZ+Abx79xFv4CHgfxuGxvasR1M/PKe0spJVc+yke/ot5Qwdg9wt
RybkgHQaiksqrG62De/KlfNcZqyMmyGY307ui4MaamHi2hvniSLQgj8rx97V8qzdrPNMncvByLFZ
YC/GKBM4blIpltsXotIMyO2hSFOUcQihN5LygXohMAzCvPyITrkslGgg3r838xcf99tXQ/iZRafN
9SIFTldQln/VfpBG60S8I6dAww6VdQKxapXZTDYkiQkaUX+qZ735Ia4bBGetMO7d8ZTZRx/EFbMW
P1ol6oOVW7SUn+f3iYRjNUXeHW+DLKzZrLGRxcoZ17StSHS1dz3ADaEDa9qjKwQz4vP4aGDyPfHl
zaxzvyEKikTNQApVe6RDPiEj1LdKO+cVp2vp84pAHinQ7p6TB8xUSSlUMvYZqD1sHl3kYcefVS2F
zzYm64/+8cqMquRBHkVLbqox9F26aACpyyKaIWRwVZ1IauXPbmeTtzPgC769raIItG129skQouT4
xf9iIrMAdJijylx9gpETrGMswlSkhL8WwYSFtNjF/+99VXiuIl1DBTG540NYNKN3f+rqVgSOvpwj
JMbNM7j2p/A0d2tusYTn0lfW+IuPlCIZGb4CbcxhGEI7UOSz1TiXTvHJbX+jSgo2gB+ECgMZoW/t
GzlL5sfg0f6DG0CpCFjstNBVMgrmcAg5gfFyWF0sdVC9maYhcQCgFsDy5RxwkQW69BHj+xx9l4RM
7QciKg2MrkrsJGShi3QEaYQmsVlCi/yhyy+RfmKsnPADWYRuZLFLRk/z2AJN7bK/AlOrCp12AYjR
GhXusvMHEOXYLfVR5w05tddGZzXtMVFcjEs576+UV615bQtZwe+jZPrDvwuoLXhLBSZWMCpVH5BR
04p/rdZkoX5VwV+gC9OJZi/ioaBNG15tDOxNlHbuctSjii1RXXMv1XmhPF7LDtmDmb98v0/GR2c2
nX6TSsGopFtoK5tKwoBPaDNhbM10wLyHlhb5SekwhBEy/A+XNSlj2ym5T3/lAx/25nFA1T77VQgW
4Is64ZkFtUcseDPyFxwj8TVoxvEq63XpbVtyalYqo3zRUYaiBm5sOyh1m7xD/fR5HIgr9C3WodVo
1QtVjcAv0YwnjPuKceq7PUFrhXZCDL1LLRSjLFMgKhWI6ucNgPo7TlMaLPc7YpBaf+Abi+DsfazO
uCSipa8K7al9HiS5zZVv7ZGfbv7TMtAVzMdCJCKKGSKliRyn2ArS0a9x5Vm2OtkH3Qg0CsiV5azK
dxVsDLH+esGqgYOLeUeZxGOps4cdIsbXzd8WGmPEwtPr0SlzKor0AtPZDnY0jbNrs0hGkA1WXph4
+egRIX5P+K02YZ0jq3u/5ORdGzHB7fGfVFviYZ/h7gMbD7OC5vdXlXPC7SodqcSYCnGIcAZn4Xk2
3hAdADE7DSNdEFpg62gaKoOibjGAZo4ll/h1B4s3VqGPJw0WVPjO1n6bT5ce0PafcZ8aCZZIEGw9
act/sIG3wF3G56jKihkrmrvRwoDtbKARV0bQV9UH3OUKhKZNnSC/O+BbXCCgyYuoFGZ8yHWjkCG4
3fQl5AUmCcGfIMbMPLlSKdbshOEsSyfcFgEiEYsCKWidJc80BFswnADFRKK05Z6zIV/ZjLW+7fhQ
qgTvOTJqtm7l1/BpqyMKvK30YKKXZeeABiCeJaHwVIsSv8R0Ed6GMgeoaMWfKJKpEeqMCAPkudGm
95Y/fr2mwhVV/cKKfD8w/RrziKYKRIYKsgU/nrkZaF0S+MX2W2ksvWkQYhy0Av3T9lEYr9eJW5Tt
omlItpTPiEuJCUXKvoEugRTx47dDwXOJZtpiv/kaS/cLei38Bi0Tx+S2x56jCA4qDexySeaR4k6i
asUM6fEOLtDU2Ho5KH8gNFfrQvwoN5nlzUxv+nPOTlXiDolFw8aytGyK4jjrmA8Yqh47yjhEMYXj
3Olx1fPcSjF0XWvG1ClTpKoTaFB8nH/75K+66jdsNN4n971bbISgFutI5Ri9/3/46iBuQkisXtUo
d+O/4PzD7PBdZi1LHSkknZhkxdgLwonXEaPUv9D9m4WmI//HlWNM4etJhfo77pJOUNx0PDvHJ3ug
nCtzciIdif2GRqztp0/4E03vzzSgdUYZl9hvuNS0+/H1f3ynW9CyuUJVA13oK4/PBpnOTyv/qlyI
hS93J+P/CDe61m1OH/FzFe8VqQT1QbzKQE77iA4/WzEuBTGb9cK40oyDGoJp0z43WIYrxjeUgGe0
KhGKyrAK2+2fDPfcdmjHXxKIYg69SqrnildlTBbwSYTcxHW7PSL694whg0ChaOqbNp0ZUtf6JOQu
M3q1uSOxUxzl4Sx6x5Lh1MGkvslzsJyEDilftIdKOJPzmOVLRaYXc5fbNZ/fJ77NLjmAaGCyqtQy
Wx5pyU/Q0XPl0pIdV8kJzFyN/45amAI6v119otMUjyUtdsRVLM2RoVhAODbirpm9Go8VsbavV1h8
6Id9/WoWK3Wr6gSW94tgQ0JmHhUZUOcIGRzSao3SUJ/ApEajY0iVNE9NR0hq4cDoQ2iI1DKJgWcP
AFm4XHQwwcy6BMBTnpW8MPXxkHnS1XRlXOxEcmwBAwiJhuPEzyrLF4Ma04rfTVTdYAZ1N37977eb
NHYnHya9gVll3hsGAoOhcFp9xc2R11dpkQJAJNOU2PVwG17R9/y9T1cIM8X2eeLcpWC9Rgjh0Yf9
LtaAF3Hvpv2lrwSPnpYREx46dMNbp3ZNLxgDEbRbo4tWu/bK+o/xrV7srnfxCE7ohNiIdvu9GDZL
dwde/suG96LKFW2Np6bm/HhbbD4ukz7E0ChKtcPjoTFxxuFHowRC21Y6jacIDNxgWRlPRPGbQa3/
34D6OuSS3yO8RpUj8cB3snSRs9pmEJF1NfOE752gutHP+16Ql3rMA6tIAxpfgicm/AK61v0rP9Bk
CdfQQzWXrWqH5ygDdtZj0A7aBDChOMhGEJ77UdsMLETm/NBifpwx/5ZCFInK8pMLic3Kt3kdI55C
QxmWVR0ZWTnlGKMCPz3zT8cv6KlS0hD7RCSU51E4B3ns+4XJrB9OabBFKCRMm6X3ffgheCqFMVAc
C3UptjPB3TzBXlxmFCDcIAx+4BNS2JDsifJEqBEBDYbSeOo/Y3pCrSJ5oakpetCO9ZvJDOjRT+7X
GzIyLkXAM963okOGR7YHcoZOqbICJro0dczkoQeMpb8M8k88hjd0MoU7VuIi3s7j8i1yxj/yMIbF
oAeGxmmpaEvD+cLrENfKaOYUz896aTS4D3lcRKn6MqOK6+ywAgGIIqxwpBTb+sgz7Mp+WCD84/Wt
6DnZgLtSPHQ/zLEPzIomgGkfUrCKAXdjvXbXWzreo2oRQXnmJFwaT6R+gOlyQdW+z8WTui7lz2vn
3RNlibza0dvOHgu+rIuJdRp6yjXydn5o7MmNcetxgX8FZwcBd+JmN8tItgwNiDHyn2ijNNMhOUCk
JcJiBGQ7vGlqIjN9eepw+cErc4Xg56mwExwhWQ6tX2vXYI/+UNi6jjyooAkF2BgXbeU0gKaS8oYy
yRiDC/eZdZt2yGiXFM02JchugtfbVidxEGsXzS4vLlvyO7NJiyCQ5ue9vAOBhz2sJ3/3ryuTc/V/
D2R8jNt57F6fY3gcTYOEbFkRRKQK65fX5Bl5O//7iIVbsedOiMcM/XJIaG0YM5GfK06SEW9uqFNJ
VgY3HqqXZQSdilorMSimb422di+gM0wzgh1IIU03u6vyPW5DCYjYtAwpyqa15YudJJPw0PuButfb
J2XtLvPM2ZNjqmUgA5n2pF6x6JevtNbvgPlPpsfPzhV/70QAumnDGWnZXsN/x8/bGNXKz9VbLJEa
fUhcB4wINa5o3iqBWnt0eXG+bglwDRMwsJaLYLWxqorOWQLs8/0EXrF3lvI0DgwkPn0jWyPl8sd7
bKBgV9KzJI7OVKz5dUhn//1pEnyMQqfqPHtV0FGpS5leBqTlo0Q8wul0+w3v8tLHM5RIVP9d1PK6
c62KrVoC4G9MP//gP2OB5IHpDu2as2FIRzVBbgZsI9UnwWOApb2dBEfNd/cGHYHPa6Tu3JljzwAW
TGRzakstfKMnQJVHuqs+nQwmNU4jfLcQRaDR6TwXv1Zd/U35qWxC146ghDXtWN4LqemWui5LFu08
Wwjs67XYflHqTWQ28fCg7cI8nnx7mF+CWKQ0x09j+z14J+9jMgW5YWyb5tiLaKk+uCxLRBRt8tEF
flQ66LgNzoriJzAL8t+20nkxCjAzOUtISQ44lUKAij2Z+Lm+dFWzHetTYXCZBWasTgPUJNe7ikw8
62u0aQYXh1D9CX33oVSj3yYOSZjV6dGLS82Ca6EmUnu3Vp45YrmIz/szFk7h0Uehdh1VPZnYDUPQ
9D/5YbU2T3PTOhC4KVUtuQh91YnyexSLlQX9OQyzLzPkpQISa7CF4MNrzra5EvJrnuY5yaplE0AD
jRHf9HxDfotk/53Fruxoa1XaXXTqrdMhcoCnMcJ9o7FFfAgobx4MnIIQAEjwHE/D3eE9zi8TDnEh
zRsNialPpr9fESY6D4/2pAZV+vUyfwmQcJkS7cSc91On819c4w33X3jwlVCJs7Is58prBRbuIQJN
n8v3iV76F+jizBfOkdVEJrY5Cn/TYq0e5+i+m7ikh45i0Reqc2jKlktGpIciNTK74jwo13uZkLU5
XiFrQmkRihoXgox92VTQ8ILp2k1sLLEgpbumenl3fnphD5+cDnmqlV1Vxu7FwEeqj4uYOXKZV+dy
hsSnOCPu9jZUy0ob3/5ymFu6hhaVC4IwJFPKPYAPfkbQLN9FKRAiOouZm6xkiBdTatNW+wi8Onbx
7Jca0Dc7sEmW5zadefBjgJkTPB9oTxAJUQLCxTuuo8CA78CidpxfFq3C9HcbyerD1HnhQuOPvpkY
dngT1TOGGMPmax4wLiw4/veGaj8YA59dt8+PVcBC9uMOEfpUOnpTSSKo8DvMPGt1H1rN4v1FKUya
KzQFt571pxFjTNa+b5FHk38aiZGhxxssT/GGs36p6pxXYwSHvm+qg6CkI02ljylINunD9An5x9sT
L6mNCZ7Yr74Q5365qBtJ+XRPEx64Op3Gi3nRcnYiUyvQGuyg23ieYM9h2dDbo74Spe+MUyL60V7k
hi0CiZ4qrLsCiavP7cOdnvjKA2T7qFC8E/f6BWk/OTvblxh+tIdwZTaxDY8OdORrL+6YMpraY5lT
cnTNX1M5D8un1mZvMw66WtvvE4lyq05ZgDQlQqSgVw4HjgQYWr/DVKnJnA0CeLBqIlK+/h6GtjJO
BYL5UtCaGuJevp31ZXoZCV07TNceveJcOALGe4xN71hEUSAUH+7w3zMgzH5zcZflv5u0IR06zPA4
EY0wO8CTyVzda7JjRr66KmFcw+WCX6yvECD7pJXrmYr9gYXXFAlB4EqdZSPUgqh45Y1LfYTQLSE7
b+viB30/D5LVUabzWNAPHkynskUbVPhy3VIt/rsyH3+FMjus9Zq/eaShMlvkWENMxXcQ7AQq0dWB
wO0W7P0i8JoDrDx6PjZxJC7bP5+FwYliOhhyRMRAczN2U5qxJuYSP0O3OzBDeAkwOLUom5q/rE5C
221o9bzTydzySbxnyi89k10ltb8meE8E8OkqrLkU+w1xif85P2wKkgU4xo5pKOtVD9wKQbkXfTRO
9Ytr+K0jRtagb1C5Cn4O+GSvmtUVpNkXebyeSezfnzKGHNLLetwvWzpSY+BYSEpii48sCKJCJf61
AcH4CowHBcCi4GcLgl0DGyzDpY0fhOY9oAd8QffWTPwru7x7kTGemtFGA0TyPZVWe+9vdBhGmud8
qPqO2zUvaWrnfVQiam5D/yTz04SqF2qpIZZ7HzYuz5aPx4NBkmbelGiA7RsXvcgeHgl5uZbGK7qZ
DfDNSrYlJiitxEyQTcA8zoJePE5qMGVAr+pmhyxgm11nxCdbmvcB6nyQa+OOKY6Zgr6fb+/N1fQn
48yT0mfd/YoBMWsXtcRECVhOvkbs1AR4Jb37AgIC1nb7SUDVFBgZpHDW5GZu3kevsJ83G51x+jpH
WAfXQiINMaxuDO76msFkSE6qahqlrJUNGACCfgPYZm0Q9E4RbN3SbfqsfgjaGrYP0QahQnnyE+My
Abbff8oIRiJ5TDI/VRyGrVJ3QaTzYZIM9PS2EpHNgussAWRzc7FcfCDeBiz04Hk9q74QgWyC1CXw
arusRQkzDw/5g26c41Xk2MVFAckBtRftLtnL/Bj/TweGcScPYuh390mGrAQSKkWJOKQiHK0xWkf6
eRFOEypX9E3JndyEpDn1o3A10fisJYid05Ja3EKXQCJ1J8h0rH0t2w5E2Oz9YGyXxiMu/+J8SHFZ
0nPBzaKYtKuSbpBxkYIzmrXo5smxFHGzPbSW0fd3IeG+Me9w9Jo9N43B5AsTRQW4cZ1gszTke6Vl
gq8EyDeYZg2SYEZVFoHvYUwBtl7DhWsZrs5b8AuHegsohTPIGBtzs4l8m3HFnuMnw12+4K1PW7v0
SsnVRIq1cF9q8o67xrwep9PmLo0YsatzucET9aUMOPv0N4cWj5AGoJ+/osm5ACAGAVtRFH8Vio/K
d4KYO6qgCNaqDXQoR/DvkHqma2T6IrpQEmYWd4vOL3ZM4RnidRrBs/8xcdnaXcV6sIF2O4XsxnaF
FOwV8WB82/MG6lNyEqnVySklpkz9NFBpUgSRX9NKHSle4titZpToz0pzpvR9V2yHNsPCO8fzruLR
LeNsIrkY/Gw7u42BpOzg9wLVo0DHe9ZquXoEuZpS6mz9NGDVUkGKzZKlH+If/2UukYivERNs+QJj
2iGjsEF/VllTsN7Pi5AbuNc0xGpPy3eJj5lZHb8sXcSLH5gUwpSgaJF8rUI6AA+QCrZgZ5TxK7Wf
S3Cg4Fj2t/eYbeKGoQKiPstKu9CLZCnesS4me/2ceWtiDRUV7rX5lAeGemf8gesHjgdvNt+C5Q5E
pqt4EgB4iP2DwjLD1aacAjed1nTv5kuERz6dnM/tmNjlhGKc8NnWNOc3T/gkMW8Ab2kJUESLPYvM
FPYdp1jbpiuraDRplyrIYp72lnEF5/bV73Fnp687whHaDCrS2jO+N9v9Pnu+eqr3z0Ry2e95Htn3
3PnJEFxO0MwIW/pL3kTIIEKE5Jc/WSqKdSetGkUFTGLwcrBNg+DILdgSawov7WWiQb1KiLM5w5x/
/0wO+ZoQU1LDHNXObpDKVQoHjM9gClWW5GZMz9Mc29R2ezNbNLRYc3GTk2Q1UsC8A8YL5PREjuCr
5rz/Mjv9zhmw+7EkyvfNKemIdrwLn5hdiC2fAnKjRvnrMgyMqcPtJVX2cudTabJlottr6ph9NBWN
8LlcFuXieOHdMUFEEZddlI4YDBLvN/JdMqa4/Xe9A8NJHH237aEbMlTJGiI+uPyVgcGDypZ6UQ0I
MHId+HBhm0eqEjrIHhUPdzOIhSRNd1KeyJptHEklDctEZahqGgnLa9Ytuq0m6x+YK4fwUJ7Pst15
0mMchX/Z5lyikRVjEuhHE2scHppw0DRdzaGZy2ImLP6atLqCbn2z88+Y+SPD0NESTpFYrVX7My84
pkuMuL6xFs92zOE9Nwj36BFrVq0uuFr8j8RMQJpmU+8GyOAP9kXYyeYVjwNhZmqsyu+DZMwnCLac
y6GOX5sJbQkunLYxSOQ+k3f5AjTZLrH8t1sSbqH9vjbOrOGSe2t7jSFm3Mx1g6PF6/mmWWc65gRU
2lvlsgngBGMFpeRHZ1omhpa44YRy3FyMEtQmW7fl7rI/kYcwajuWB9+n5B9Dq+wSlzgCf1lEauf0
eJyFAd0cy89HRCJ+zsXecnhWOazq+jIJd71hCPd5bADwfR9FACEnkUzYOLyOg1mKjqbi77uOehi3
4p5mvdgqU5tTeD5us05ZEa24XcsXSQdnsGnx39MOggDQlSWbC/sHbLe2HsBscN88DII2RRU5OX6j
qZxZjGv4j8YjZdbVvBp/hnea0sZzFQ9jP6Ikme5M4mKuu9qbKhX2zH9qX4lsXULqUcmnH+B8VA8P
aDmECo5tOKCRQGrzNPGb1g2dswhkAamLylnnAB9ePghh9bdjA6njAnas1YrzYjDVgAcMJpaJdB5l
0QgUWuZAG7Goc/Ou0HoZr1updurXbzZKJhUU6bUW4gES5d8AzG1stcz/bDiupAk6INPnotDoSaLm
OIA695q2baq/Oayo0d4TXVgNx+jLwJ1WwYc5Ox0k9PU70l5yyB7ebBUhEbQcaNeFqUZSH2lVPPMv
ksHDjtE7s+lDDogZXdiywYfgDqOU5iNTzlz6PXuoXwszE95FF0yxsx+OYxmynHRsgLMVk6xROtrk
gz0XStPmsESoJWBZlmuG+B+FoXgFLKMVIDG0F4BsRYbxKBSfnuZdUYfKbmhz/oPkj2Mev3+HgAXH
CXRNTfWxO3of/nz+CTUdIP2Zaribi9f3mMH/tFPKgitcUFTbBtqYHL45kOjDvGpKyi8Z/ajG0nas
tvTXbhRUnEppeTzNWL91qyE/xhFahi9mgboM+JMgVj7QZgK821gnjmJkDSf77SovEcO1aygXagGP
WYBh6pv755dNg/A/OCxPIq0MPuZYhYfY8Y7A335gvC5LfUSGN95etPz8tXLjhyEmBIKkqcuqJz8H
aB4d8ZsfAFZ1cyIJf2E9N/nBmoq0gFOvpmQ7dhKvc5A+4sS4i7js1QC3X2YLpcd+n68yWGs7cy7j
11r4O6p3RGuq3yt9sveeY0IQsfLh4jraRk5LQQ+v+3WU21IVtug/5dv8yoiJH2ulKJoNquLLenpO
2pYdEocn6t4RFhupKJkwAmS8TlKfFyxOHkvX3q/AioBwx+UGVuzWIDqmfOzOGHUByN9vwFL+tOxl
femfBcBu3dkWeeLx7OF3M7wJ6Geiq2noSKRyB7a7gCYQwKBSIdjya53zYDvuVhscCMRMdTPTYaag
ufGoApnskA6qRtNawr1DwMmyOZMZhgbq
`protect end_protected
