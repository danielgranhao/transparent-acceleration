-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
KM45viPywkgpbKxO2GmHzXGlUIZWtREB9gbMgK/syscfqgxMDcQ+yFtiU4usz0Qi
WzErzyIys93CNWyxbajNmnRcd6kcR2P0b49KWAGla1022ym0feyEREfa4zH1SBQ9
OTaBs1vSX82Fr70suY3QAGtQYRiQfjmTTKyOIL9gsiDCMv4g50iEEQ==
--pragma protect end_key_block
--pragma protect digest_block
6YTNE43CxTVCqLAiaC/nVM6qRpg=
--pragma protect end_digest_block
--pragma protect data_block
J/bhwBZXfqlLWZ5g3mC9dmC1wkij4X7AkGJbEjYC0Mj/vonapl5Wx5t2O6MlLBLq
ZB6WelQdI7rmdTqAsblE3tdNIce36y3fn0+BKhL6vVifOdrmmuCe2uOjknMPYnSQ
DPhr3kqf/vMRw8xWo+7qFDmqlfhMqBdBLEx65OEsMaEtKyKRz0YuL2JQ15i61BNj
oYBzdxrBd9ZOxagM4H3AA9J3qK47TD6LBPpKI28scNuW4OsIQU09r7AYvhhgJpBT
1Q380wJfMI8jfSrwrpa3+gQ0QIoKSQJCiMf48BIPxAFsasJZJfOWhaAFKu7KEG9e
YDuJqNt1RRJwrd77zIsYHk6euDqufg+n9AxgVNyqeL3V+8Erw9CJjQp87UTyjkXX
nrAcQVxiNJDAR+qEXknplFaFxdWQb4PIPNp2BLt+zPRc9VQRamS6m/NrAC7e6P/b
sX1VdG8nZR5X+9a82hUaTg6KTfX1LGZPNAY1Ctzngb8Y296p3v7igoyVeQbrJZzm
0DU8ahWtltp1xMccepTEGBjecZrQwdCVdOpaCvtX344SWcjS9otw2Ve65w/LKFF2
aX0jBFjT/TomWrCXIC42E3zWvu1hhNh/nHwp6CQa3p4ikBduzzuZc5UxlEqgM+XJ
87tX3p2gcsBg57JtMKObd0Hd56m+UF13ZljUszPuPN5oYgtKnoqEfIqGyHvlXSXV
Pa7Hfywrq0iiIqb2TG7JC4cxMX+tqy8jGbSh9bJcB4/7EVWhu0aJncuhumEOUatw
NE19ufkMedgkcFmQZCDdTDMYeLBYaaq+N8XrT9f0oAzA1db0QuHleAYWswOpVzRZ
JtCEtZ2M6O+wJO23Fs1TsfhT7ywrh/Nzl59He15AxMhzU9qBgx+/O70alzrjdC1i
EbueZmiONa5pkHb6RaG5ZrdaZ6DPupznuZFaa0Z7arHoklPdqC2QMgesR4H/D+RN
I+L+RVs9xpu9dQi8gJoxiTu8DT+OsFMtfm2UGfGj81Ew3B01yBzm8PPXL4iOwATt
OCoRZB56sAE5G8jktjWd02Y1Si2/gbZqGHhoIC23uDMZv3LoG1Et9KEjCAU6kKfM
POkWD0fOhHx59bQK85rulxn6aDa+f70x6uFV+VXDQqq8Iwe9nLsRgVQbcUH6TFkx
5+VT4V37JpXEiP6h6dE14DONsM+Z0vow9Qoj3R7j6WJI+1XfKYGdIi+tNqlZDw6g
qCj38O7L9IMFToAAwxQPWJVVlUVMQxsxxWaC/xarSR8TdM9rDuYbf1rrYPJUgQR+
h45oRnoMobz3Edw72Qtjlmjbvr6LIcuXSgwPR+HrOMdSyDo/EyBqqVdKEk+wjJOK
vRgTKqx1bVID8a1b30qb9enYsmtktMKIUd0KwA3OVFh63IhKhe+FQI5IzphhOjgl
+UEhwKNrjewwqhyQKB7zDrJ5n1bylIU1VMbBL7dir9XQZJAjUqKvS6sYrv0rexoH
XnepYNfPPjhkr9NuODHlu8uG8p6hAK7VmgYW7vsn22n5TORC30HNMg80HbEsuqZc
LuCZXIA2wcu5DXDFj0tLKAHaMaaZ1jV+xT9luqbfhp74gmpPKhzAHcDA9Y5+KUUh
TGVxHDFBmw3534MflW0wvQ6Nu8rBvCsjA/FiY90kQysKTp6Zem4q2ySIZItI+oOk
nMIahin4bnAuyeYhlcIKTeDo68B1WhMyRkkefrvFQxGBzcdq6wU3qJtMZS5PD5w4
Qp6jdHoj3ebZVFVQOKIBFPKFHp8WNBdeeKpWmY+syVjWunFo/rL7KtcUy1z4iXBT
0aQANFc0pernEJMaEhPwNv1S5m8xxW2fPWCjx4a6UJbr+U93YaBpSQ8kBuBfZbd5
DZdRPlMA+q1NchB+9CFCLgNzl9uHwwOFXK/4mbex9dgA8IBWHcnuvyVJSFrKX722
O2AwaMjJhyd6HJD/ApPsD+4BgIEIPxQfjrzx2RYSuf3hOHH5NPMs/ELZEK/G0ZRl
pmC1Ul4KjplqPllbbryCom0H0f2swwtjp6rdAbehbBHJNpkhW9Z9PYKhklC9xivJ
542Ccy3JT3OvPPiirqMdXJ5uXxjebUZspUqaOFKGNpXcu/3FbwUnuPGuUb6l4/oz
KD9p46gOepZXYYvuRY/zbbCF2Zr3febvvYWKro8LaErCetdxYpsjkcLbHlWjKhYC
wL2v7JwsF3PJb/8Ku7V2Im/zqT7uS1EuEy/GV6ghEtAkngdImbMzzjG0kTTjcUDO
VZAHd8rQEG7tATS53+Ewd09REwjWBcBFLo9uakdTuGkkovzrZrxdgvvxErzLKFTg
jZdBn37oBZjklkuArVjVkkBbvyccODQeQ+RukHo1VF3/7xOgBozabAzCWMwXzJOP
At5BosZdyBTUdOifDua+yROXFs5iyChPsCV8VVLqIodsk2kNo66NlZkqpu35qJEM
8Qd9auKOAVTneOEoaf/gldqijX3B5EcAYooDKTEOqyyYdN3xsipcxxmCXv0h/C1l
x8LNcoTcK68VtVYSdMp6FzLVt1TSNEjIRRqOl9oFqNXF9Cy9Hem4DcF6lYHAEIBH
3wNtEDgnkfBfsMmdiDBeOhEppv8DXZNZo9eSp99MdQ9BTAn/bmi/LUNpoPpn2Ugg
fJl0opAMyY0M4XqlaZmtaKKtw86TvDoq8YiaUesyMKXzidx7NgIhEB2TLp1YqU8T
OXYXGNnO0qzpjVQJWhh9ZosieFR7Bltqr0/ZhdXdOcAvg7ucsq4B62E5AgimYWCu
YpHQFKPreG2nY0dGZlcpd4y7ojbkh1CHTcZX15LXecV6Ecn5bv0LQnHD5O2Em0ti
Ocq9VuMcr6dFGkIT71i88owf7j72IAfWpiK5cDY7/gHCvZRv42lx6fTysKnhWik7
MtfrtctgNYty2fW4dZjjKFuxc4ZdZ+1B8+aNqwLRT+0XeA17K1+SsoTlGAExJUUx
uVRCojdHxkckdWwkKRTOY+fKYktuZjw3ErmR8gMrUibJn5CH0Db0H6gFHYW/9ZFo
i59QwB/ODerFd4sl4O/evtQZnZwwIRUSUmwicT2Hz5JMmizz7uXNzS8f+T733dWm
Jw4m7By8UKmwayd3AJxjqBh+gTTMm9nTfKhAmGdYRTvOvzwvbmw5raLpBGrXOeWZ
PtI3D2rfy4kIRxpQK5b5R+mR9AbnZBygp5OfqfFMaFHWx9fomXNf870YaVk0OZ7a
rqKFPw/DOm2d4DILQG/M8NmUr6EubH77540lDK9PFbc21NYH31voBfAnapjCMVKb
fD4sgvllaZ60EVt3Om6u2ssW7LojdoBtQWks4lfgHiDy4uqbSwvr+ePWbAjN87Pu
jz4+4rAWg5ucY5Rt+le8i2bgugs5HAdCfDjovzWzqEwEshDUd4ZTedMhx6qrNx5M
dToWGPcwBILjSHxyfyZ5kTt4CqdxIgr/32dG5JxqVufsGFiyMntV9RceiS6u2E2C
vTnPtgYA49RlWmmY0UskP9Mvm3zUFskED8FXT601fyUx/z0K4+IdzxhzPQkrl1Fn
hJtBbWOgeMq+HmcHzBejozMQNBNbg6LtxtuAt3SKAPUfRzp+x0TrEx7zSh6VqAnR
iAme/m/XjqeNAdy9uFGi6R62sPex0lK/Z4Z5nfO821k0HVNtLQ8famy4QRdQf/mD
HvrRP8xbn+u40Getgaw4y4jn27GlfzFPQgROMaC8xA5eaB/DHiFMcpeY7JQY3yWa
0f5A1/eTwL4rRJQ0RJe+b86/AX/6erq3elPMv2gk7m7SFqes0rac/phyWMWYk12F
FYJC6HCLSH8AvfTc5U4ZYlNdMN+uRJBuMr8C4RajPn0jDNgDahWUrLl4DtD5lxsj
U/Nh2CSQaQjLZReCphoElSTVZpHirTjqr+M5uM2sUJhtbjzgbj/IPo8E/AR5oaql
mv/gpAnZW5dEoA+Lm+Lhf5iX6aoHJIRtAxGhTFoTd0O8O2smJyPpv8zVFFMty7vB
YK6Ue5ugg8FeiU/R+TojTAC1PeQaJS0jzvnM/qd0myDvQY8ZSn28hA8w4cjmKqSb
aebFh0NU7cj4odcUGzRg88qe0bQ77G2OddhziXMr8/zm8qsoaBjM5X35cqdtkizC
QZ/GpIrpLAi0H0k9hK31TpZYeDyrCJV7SAaN3QP18SkouZQ9oiZWEEHoUBsfc2PN
t07mVLN24mgpuTWHLkN9uTODto+kvbPKBFXQRwXXGvD2PBnLWgQ3AaU2FhUoWWhp
cmCIRh3IfdrF2bbzkk32wrsnA2p/TgBNoEncromLpdvp4tl3f8wbrNVIQO5/Fi5t
CPApQW22PmuKmPxmh2bcyQUd4d65d2KY3U5XmnwJAqMTNCIj6kFAFTH+BdNSlHpa
kdDEHd2BG8PnhqBKdBHHQGwEsGkrVXknNz8Va4Do0Q7VxGRnrZ04VjWeeAufCKxH
yODOU1Ks8GjKcc5BD1a3JpZOjb+hUPElGdnJWPsGbG7oNI7UMk+vKQwmjQyVOs2V
wV8Aavm+m+4T5Lp5WhMyc9C9I2gaJtB5Nd6029/iMw+uovEaBpsO+5kzZHWwuuQj
M4At1lfO4SiRxCcn9wk5Av+n9j4or1v4rDQhswsqyn/bvORzsf6mxqSpIhXzei8f
v2RYAqi/zseiN1M5QIF5TLPOhViinmupPyr7qDanysy5OMSDJVkB3wK6fgQLaV+C
8ci0p6YUPdeIU5oNYXjSDrbCOTl3HXoj7/vZrGOaykQ/zrb0NbttcS0ycN1FWkrj
9XsDS96wyA0NELbl3/U3okYrfpJ4u0lKc/qi5QshmljnOiB7BlvSEjuTJOWHWs4g
TcqOyi0P7mvOo7yLiJce0HnEWx1aILDHBTns0F8aAu5bqx9rpRYbw5at0zWyvT3z
zzfXnj4182UPoeyY+q6MSj1KHUMFxJ7yZ4t2/7RPuvmTfs9ABzl3USEKAlFoSHZw
hFWQ3rCMwbZ45DKjBLo12rvnfMAS4bVD0KQqodcMuC1inRb4LfCsPC+Sv9/X5jJt
EqcFCIR8GRy9z7eyTg2/vgmZRqBWg/H7Hz7M1Z5aoSkgU48nTQSo/2ufQ413/bqG
eNgkcS0oue2o4E9hHxMMWitb+FvAvpaY7Zo1G9K3d48XjmwXWjnqU6hv9JzWww1C
+iTM+DO4i1I9Zi7R0Jz1FzCa6j922qUSxTsT67fry+bZXCt0JFc0oWEVU6lk2DaJ
7mo8Nmn9CHrCRMcKmpclKfmSBCJUzlcL7wFiyptaHIHu5uZuH3F+jmphXIH8u02O
KME6i3AFr+8+FnRb6Z4JRtjXe52LtjTHNO+PGJaYX8Sw1P6BxyqpEcoOXq3nokKi
cKtyxoBNOmfgZjC04mNDJcNK0oGaOM8Lkmnx/+wQhi68kQPpmL3Zy+uQqC3HZ1Pu
bA5AeREIVCRvrpWmGG35yzyhlHqwvFutWcxoufUC716SxV5uYslMqPTE346RM16i
UMk3FkKx1Tjzci4eRPtRGAzYKjbPHN+tr00+o2fZ9czRUrfstVPECzv4hxGqTOeS
WrqpdplmADYTD6SNPQuZFS+m4wQDIGCdGRqzRY8enklfZqR8iq+mOqjcZjnv9r6a
7InMmgYrZirc0x6haGe/AYxzJq7r65x5TXJQeK1iCPHSlshAciX1Y2dETicTPEuR
QuAzDuYO4xEuK8vt56albnmzo6L+V7vBYqEXYdSZw9lcs0xjj63JpBpg1zTVpjyT
jeOZk67Sngd7wJCDoTF/X+QIcuv6tVQHNO61C5j/oiv1uAAIV4rgr8e5EooZLfI2
N+7FILJYuE53lwScBj7b1zE992g9kIXypSbD7rfRxr7ymKd5dserB8OhWzdkbY3K
naSUN1lrCsfL7xpxmD2fNCbToYo7xfHb2cWoWLU/+YYMCjXBL+zoBtlqCrUKOnGv
9V/FI5j6tWinep3cvZBUGxvR8ZyeX32m/iPPOjKvf7/G3/A3ifNG46bh5h1FVqN1
6RKBd/rx5lkl68/wwbKRIKLObpAig7F5YmibC1k+Hfw9KR7KKo6BOpu4Jp3wHIuc
eiRos6DtWK2Ux+l5aVPm52LaV6JI1ZYqlVCIVEZo4qAr3KVf5TpUjGsrSRHhjHA4
uaVB1UBgFdd1CfYast7RIPJJ3ArXgr562MkP/5YOgS/D6DMg0Q6I4E7NVgC1JR7Y
WRk57AL8BKzW+s7mY7aLou/a8dhsYz3cQ5KhraQSZK+TWAlaZH6YiFoCu0RCtOY6
O7ov9Z4Gua7KUUp625VTW0yu7bpjp3j/nErBMms28TqtkE5Wrz+6Eqn9I8IyTBar
BvIIOUmq2JFsbJmSRXSA1sn/aLiAFakPcIm+V2VMYJFicpoqQkPPvFnyzppPo1E6
0N6LP+68jrp2Os6TdtMj6uKB38W8U3jtSz2p4TJpOqSRVUY13Xt3O8I9ddZMXL8P
0uQ5TJQzBJgNEDFBnFwVcgD8axW055vDMwZ+AmUh4OoW/1fRWj6ZVVwS936BKnWD
Z/Oz9LXyPaDIvVocSekt0EkhVbyZ0Ju3cH4Un7FBks1dmM2MZbp40RlmJaChWm17
9i2i3ez6YJVp/P+erCkAe1GdxKW6JWVtruzhz/fKH+oXV4+2XNvAkiL212+c9JvY
w+sHXsbOlM1x+nbAebwJtdKl25CV1G9joPF/AtF06hpIq3f6dZOK79+n48QcxA2U
+u9sVf+5up2CUena+uEn8bB5I7Idrl7D9IWLRh8WhVoFvhWWw99/oi1ZPN5j9+3b
Rae/ddIYcy7dHWrco+WBPmGJFePqVTlxWGCfv+I9MoOcF9aKBY/B6zygRm2ad5xy
c3zFLp8Js4mViWH5bqHdssUzqJRcrWEhiX1KOgGIXuc5P5rA45iq9c9RE/EzpaV2
Zt2YO0BnbZY4je6UBEs8UGZasE0a7aT3y2XQurBS1QMr+gBTTsNoAGB3YJt5vA+7
5rbTYEDqA/QdZMauGBDzlHxRAJ+aY48/ADE6FTmpWEPjgWLTiJX4bVk5hQcgNTcS
mvHPCw32rqQSkw0ZfQ+VvXAnA/vgzzwCLTpxrsFdJXBp/xmnvDoTMvpBAYHc2aQd
07K4+lOxKPzt6vfKu6qdno59tg2ybN6y12Nwxjs+e7Am3mPh9I4pa4+w80XvnN+Y
8RScxxR7PY74wUT6X48lWlZCuPTVK++JHXcbnEn1KeaM4B7Mts7cyNlrLdoIPCzO
zsTnjVENkcCvLO0d3maVYHNeNS8uVJ/eWh9hWjKUeiNGcJ03I1xyqM1IzjPEULPL
xR7DspcmsMkN3+Ru0XrAE9pmqcQvhQa8fSyD7Y9S0hjIp8jdICEfpQmPK3CejUYW
njnOxQMtq/29yN2wIvBgY7q97X/EYpB7GkG9K4AuPZIv4QM7jOC7yOxMecvX6sqP
fBHdgM114YVPenNKK2XJOsVtbH+Ylka+8F039vxHoz+DMNA7YV7XMNMVku/f0gXX
RqDvSQ66QvXH2nBan/auIB8SvWOvMX+IConQXJ0v8ReKMGRpqXViOZXjsRu5V7k5
htg5DciN31H0KqLTzxJKuixu1R5JwqrIWrxbqVqafcYJdy63/ZFfvw0qZRJI7FB1
Ggwq6u+MhXzXztpyDJAggbd/qH3GeisJ/8YbHjv5cChAoJtvsQwuCX0K8OxLq8RD
vpZw5BNFc7m4XqdeE6J5exBXfBzlCImK2ynELpuffjyVt5VaYzLBoLkoDpaQF3H0
Zwcfy9d5YM1Me8Le8SMPvrvlpo1IURru6TxD2l44LKp2DClcCTmNQ/CMJgwsPOze
6qqgMzJpFPBHzV69vj+VvTGudvoti1CWhD9AO8V4jdzGWzh7k9ve0+6gn7V/iY6N
pVstDiMZfZDm4tGrS8X2DjdmOKqu6RuIWb1dm4oiZWnEuoni28vnmbno+Jy0AaRS
bOirrcQPWzTp1am7+cHdHmonl2DuF0z7u64YHgACffXguAZby0v8h5x/wEdSh/77
1JBevEvSfZAtLvSoKv5prTMbyEX3dTm1DOxf6kzWDdsgnJun8keoPIBj2jp89dE1
uirvYfSyrhF9EMl85Xa/4qDyGbw3xgTmk1skoZeObmvKrS17FJkCzUL6w+9UBnsq
+meSDxJqywQVodiTJMl6nN1Zyxfhmx5Zoy19//e8cfm+cPxs6zQG88zeZhANk4F8
PE1mEjW4Bz0099FRD8TSpswb6e/y00ZWxddzpSkUfCsqaDV0xapKFGR+PRe9FoT8
j9iTajPkB1o7bglUXbhY6AZWvTixcXzrbDFeZP06dwRofHUgisE6LiNI2KBWfUOr
BsOzZi3Dd4KoEyCK0NA9/55iqtW+J60uUkLMrDjJoO52YFOD9nDQDXdUxHoQ5ZZs
g4txUY+whWZQwCSoJaKXWM67CGgHGu+NIjbh24Lwt8lvynCRqePAhuSOtnQWREXr
UxXbTePIbq7fYHbtks4YAYe199MOxIfknwyTe5MqzS/+ESZEQDHMtbcw3Ls5mexq
VDWsQosVGMg0dWsEsuysoRGdVPhtzz3HS9PmdI5oldh4XqrAhVKlHcgmjOmWCRk9
xME4ku6nuDk2DqRyyfGwadB3i7L6hJxajcGv1BD2mEkM/tV7jFxnDP6wgw/CIF4k
OxqaXjihyHA5G/6desqRkyMkGb4DNHuQfXp6LpfndAzvx4GS1kpVlhFB2FStimoH
lfqT6nMe+uE7QsBJHhH1h6weCUetMz8UC0MJ8fmzrlHh/trZmib1IYh9mLYkvrpT
+lBzRiOf8IehmLIHbVd0SAdv4VUasQOrZykSNUGryCQuITh/L9fq9+IseQV2uBiz
RFy0hnnS+dCWeemX8T5h8NpuWRcIjUiq1N3KfIcvE138QevCz7m7skY/Mz9HefEJ
EUOWsFtxAS3OGqEGrnVmMa3+TfPYxro2hhTM+HbFr1mVyv/oTlyoc1LLsVEIchbp
C2fyqZdcsXNT0F/HJM7F9F+mL/3m3JdeeeY8ojwY0aiZNgYf1p9w2I1EYbDowDmX
vD3EHI4MCHle7tMiqf8NB8wqbz5YGATXcV3mgH/1hAtma9d8Ypko8OK+5QbJXrkc
ocPCnaB8FbSzf0Nc5tgqxqnEU1SVN1RCiIPXXHujilI3Q1UoIT49WSdBimXQj9WN
1/iIOd0CRxyAcfatPVczd06G5hc9tDLYVofwXZX9B4CLBE0Bfko15nHNIfWPKwx8
CVla5XlmzPVCWijPq0GJCvSsdWACLtWBURt+XNjSAfOVTneAv1j4OmHm5vPeFlMb
n39aWDbfS/shGf43JbO5zzHcfbwusuqRzbNrNdqfmfU7GI2/AsYaBO+4FB5tKMdo
kBSmm7XOyQo3y+v0Wgg8/TxMxdzqiP+IL+A9VlTfSGa2ybHBc2ef4Hzq+WuMA0Y+
5BWqcZAOFSr/yejwdXR8lryjY6G3AkjKxUwVnLiKKofd9HvCH+eXppzn9M2XOaLZ
RIedzP5drawlfKSjjcvISkDzqXDM9etZVDPGXpDjdz5Oxs7D+pkBlTQMXI/ylJnJ
3B0fRw/AY+34EJh630n+/iLihS4SILmSn/cTxcgJSuefRZJxmQEmdUNtoA6YF+qz
v74+a1odsWyMH9PKGod3mKm76PKkgaanHzqM++s0XfWQL9LerG+aTa/Sdg3g4kZq
aP5p3kHRYPw3fd9Xg7p4tkXkdl37fnV7wczyAkqeky2+xFAretyuFCPV0YLzxDrh
lDbTGt+AgwoMI7FEH7rHpUtzeF8M4hnFUUqxNoGSIPvZhdvoK9C2ryCz8o+i3zYb
lDrI6FlGe5AdBrVnK91W22ioz15mHGUaroOsKvOYxQcVVpUE/49YOIADiYcpFzLP
Xvz6H0Vc3wsOm1bTAP0z6kIzS3toXlPs40I+2p99Ox+92tU30sVWheazWs+DUQh6
VidlJUnVWpa6KaX0MZ1PAO/5yQvp47HuF/uC75c+b4sJGYrX4uIilTB78jfNadNa
C8LLnHjnLK4XbO5gs4Mc1X+R+zg/jlip5KEvpbcOgVPovOiwe1OfyibuBCzrzwTy
p/0Nke8r5SpzCz7qC5wZvrSIbKPHtoyX36LYAR+WEc+8aujwL5Jm+cLJE5o+M3yZ
diG2OiomF6khGzvrsMMpGdpdBAH/6/XFnHD1tM+iIT57dD6tR+0HU2UDz3oA9hDZ
D957ONq3h7OzRMYduFO4Ct4T2VROIfefPOCw8nKW6/oOF30tkDHwQMQzCWDiV4Wx
7zbWHO2nyjjvGo6m3XD60ZvLR0Y+6VRseTIWpxkRmT6MS6VC1a19j4CFZz0jGxKt
L9rDTKKZpRD/wGvqrzhpCl0cJ/xaL6OrP3K0+e7j25kfVqVsxN1syy5zg6fPCO7m
dW5VsEPsAShyLCVkjCcMTXymgSqxNXaLceNBJfOHCULTjKcH/25m5yplU3uLjWwV
K+pUap8Yl+vud7KeXJNOyriirV+1GIsKSg4JIO2Y3fpQlL7Kd4KyjObgrdEG4wSB
u3cn+pWWZ48Gt+ujyeL+Lg==
--pragma protect end_data_block
--pragma protect digest_block
9FnTHYvzBJkGqz2dBCcFlIb2bDI=
--pragma protect end_digest_block
--pragma protect end_protected
