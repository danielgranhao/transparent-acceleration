-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
GprAMlbfvwkdCCWyXFwU8JwXxnoRXJHlOyGBT/YcXiB4wgIYwPRE9ErCEdwobDif
zyYYYhkVhwMYvAWQIs6zN2rnZwYKPGKf1Rwoa62K13wNacYX+vopMNs41LVwyLJA
KBt1Ec/ZkXtg98LnniG02HDunJuK2cSCX6GzLzuMdzDv3LgDCqrbMw==
--pragma protect end_key_block
--pragma protect digest_block
I4NEIjWlhXzalzIb4Uhoc9zIvz8=
--pragma protect end_digest_block
--pragma protect data_block
3x3q2nZzG3lOepZEu8hv1VHLWd0sMu79E4pbCVY10VUkujFnOIxAkAmuCyA6zHEf
NZI5nl7/kLeRZm7Pw4CEktw/qZileB44rKhokseQTYG5RwaW5DiakIam2JdGTuzx
lKJ4gHYNHFTqvNOq0pU9sWRFtGNSwFF0wDJcntgcmghAd8lavLG50CE7DyU2iNzI
1bOF2NfccBtdp8lYOu0S7LLM+91wY4O7QRowVBCzOdDsCdiDgC7M/TWus7Kq5Cqc
3Cr2xw0a0ee/iCvtZHkXvG59HR3t3l+QcYUp3RVnwpHbZF7wtVWGgwi8w57+P8rJ
DK4AJK87FSOG6xkIF6dj44bWDK2fGxcHSy5qEzxBIe7K+LaWRlrkfo+958G8gFX7
oxcVuSFKUUC/pS20zYtsqpqJxRZINHf7l/B6IIwd6QyrQCA7FgYfMRJlrok6lerU
tWfLWLCy18g0TiYUaxp/5UwMEP9ogwxgos0gF+nCv9cIp0Fd8kLcs0EoOkIkNQT4
Bx7G2HVD+iMiRVdkzlrG4G3pmMGrACErd671z3rJ8q7WgAaJ/2g/FZPwUnGgH+z8
juuQmSs1+/8s4bw/kzEFe+jffYL72JwLc8SJj/UpICDmM1NkWZ80Dy3+9IhZXuLn
91IXL0fdlWZKkaGjklDWWxRtcEhdbrpGLqfWsp8Th0Q6UIwG18E0OaxuiG+2bS8E
KsGN0PTDhzflvyEz8e/jR5z8xPzXGlQPjwhU7QPYtjMQpkB85PJOYIsyDFh+1nCw
y9XUKebgWEZiIyt9AVKAMXuRZ5eYSjaYIkaanoiEtJjVhEeSfzDH8BzQivC9OdVm
rdLI1DP0tUjyN4DzxJ9Ir9Yj4dDCO3hsqczdWxZDZYYg5CMvomiLOLLDrOBVCKS0
mnjZVevLU0cDoCQd+cMLZ2XcNWPEfmpURkXVue2DNbgTpFaZD2nSZpu1xusZ7VoL
gkfQN4QsXtH4j5S85MB5+uWmaB9WkHW49dy9Ul0Z0bsn6IhoJZk7pIgn36tY2umb
h5TcjSqu5eaP3Pp1EGjYucPzG0c2Tj6z3x8KpDpdMyriQRZMszFtE1DbLMZaxuaI
mKkYM7tC+ImriLJHJw7iczqWkXZyAFTKm6x3ra7au2DRo+Aa2MpgY90DZ3wJ0d8k
6f9k7TJjUgtYbggniOo1BuOgQzu45rViOk33FbFstL3c5ieN8JANUOfKZD9fbQOI
a9JOu6TBgkWHZTid5AWqiWZy+TPW/4kn8x+0o1QJRKtlRSAJrza8qz1/Cw17pJDx
SvOD2sHEqxFZ2prBnosYoevy1CJl+qo9g1ANfywaW1DFr4SlSnmCIH0mQgIx9O5F
/zvC3HYmDpovy0zvCCC812yJi4anHjOqhaRF1MQJvzK0RS+7ftRI60voth2ea4oT
M7R7nr/RCEWouJWl/mJALQCoO9v3mYpNrzjESmpyMMyGEMHhFIb4e96yQEwW6tfS
mCoyZSp+CzlFFSWrSyZgDpndVoFfI8E3FuU/wbhCFspXLUWcd9+9nh1jXsa5Qw+g
TYfSfvI62weElJmFKbCy3CCgCY3R/ArwTRgbCLdL8bCyowaC3NuTYbkvV0D2P5/W
LCmHfKH5niMGHJ1e43oNHZOO3s6uH4uF9jnsJnHWroEx5KmMoBT+g+PX54k1VbtE
DBzA1cCEg0utDDohcYQmOIWf84X1Cb4xsxO7rvf6qGVaJsJMQ15I7nnVdsifQUiG
Y3Ko4eTtHvaXucbbrazaL7fLGWsOx+oyuENlgSPYkHQlK/30/13vfK+TpRWK3Dnr
WJt8SseF67u//zRRNnp829PLbJHo2KMN775AGYDF0bZ5R0HZg9KUPtu5bvZBOfVD
cZSRjdwsun09lKWiAj4KS6/vz02cCE+yrTV0R8hi+8JPzAGdTcn9CDiYy9otSdO5
ncM2WmPdOkOKam3j5/6ZJ+cSUUZEs2wcKvAhf+weU4oAGIKF2Ui/D/8YObUALhFU
btGkE/BFHEUX8FXKrL+NU3K3+B7U/5Nk5XaO94Gx8eUUS+ZH0Lb/G6+XglbyN+G4
JYVLUAmPxAgBBzxlbUarQhVqJ5S1Lt/eaBgZ3eM65A7P5uH2wuBNuLnwiap20bHw
xc11hXisYXRgkXCd99RbUZvkdR3mkrGLsGZ/BVo8jqOkbnWqPBPn2IUa/t9mwtST
Jy97K+jrn3Mz8VLnUDsEJ1seXGEgHv9nh+r22gyJ0qHL4S1SD3cZDQrBApfRc8/w
6ggS5UUysUU2KNIgV2x4HK6UZKAdUM8dq9ukUosyOYlNe6gufQXCNYoYCp4lSsA2
GSFWq3s/PNl+xiVnqRZHKlfgUYweXL7JQA6+IFyGXSmCNQn6LJCbqGYtVWrtjh9x
HZj/KNBl4sfbdyqNYinoLIJPc+WNbjnWfBSv1dV3ZFRQX8nMQhZ8UV9TwAYjibQm
UGvXEZfKtMxiu/pBzeP1alDl3dS5ZlX0JvfqmgrpNJz4n3iXrIM2F+hew/NLWdE3
MBXXpzQjv3YRGx2rdV6YCUBWtISdARLBvcjU9g2Dh1ggNM5SwMDhGEavovLbVcaa
9rpfV7oAHYWJrFMpJ1mQIXWcf9xb9882sZ1zImAaqu4l/o3hckHEdefZkfx3yVVW
UcfFmvham2+J4N1jHm053kuAlqYQGJbe3HpSbjD88a57MQGJUwBsx1RpMSls7XxZ
HlBYjPJQrcBHq11LktoLkyr1NEkTE5b5fzC76rH2l27GVs41dwNSfQ6T+wrGsgL5
AxKfbZ+b9cDXzrAlcpEjP5AoCuX9ci93wtCeEG+apqxCOFDZDdSs8G8MefDPEpR9
3r8S7IDHJFKOv4PceCFERzmnK6Nx/w4t4V5LV+tZ0jFJfr4k3chPbPQrz4Y8EJI2
6o7aaLVrTqwnAnZTLFiNS1irHi3JuXMYg9SRuSfylwdZBf8pAz5QCBDb9eBMektl
WX+EasJxQRtzjw9sm+dWTJX9QN0609TljJDCbOZYGN+AAmkOkiOdKA885kyrpflW
uG/WuFFOy9Ug9EEa7Km+RqeqFTUrpkCIwcmhGuA8rj72eTtJQsKx3WVLre2D5dYR
HiJjmNQnPwkTBAkYUrTQDOOkBruFuhI7ixMDn+gPtxMYpHBMT3LZHNmUCqVDPK3K
OIphD45vOpUPRmPsXlMAu/hPlVE14YAWd6dH3r41ILLE31CxJVMVXZN5AAKWshXM
Lrzi7CjHrPpDUq8M7nYPBv4OJxWs1EKX2cgWtxW1/rAEQlOQhueNgV4RGDrciYlH
ARN3s+b/EAfPNolxDUeWidpbh/ERXn+5D0sB4J9+twqXylmRC/mVweSnEfzVFAlq
ALdpi+n+ADBlDV8VLxniLNx5VdhwI+FxcvQkAsHACminDmglRlraV40SE6E8Qn3R
w+C4dKASTrqWSxSs2E1eYyfCkWyWNfYn5CUshZGeUdVw3xRThJt/eZJrMraW3IpU
RFQ+8YLVb+gAEW/us5jh/558bXbz6LGcmCfUFNnAd+OKXyg8y+7sEKtVumkjcQOb
szgL0IAU4caZVSSa8uqhLMru0b++LolzhcYGBbYpTq36+FSC/XrU8eShxfsRLjyv
tJ6H3Hx7UPFd1/hp1ooYq2rTthC2o0Ix93cJ7LMR+zN6XvZuZ6bT2jRidve5ZDN5
yvHxloqr5317TN7t7AUNLridjnVNZ7vC0Vw9lPZZah8VXY3xYTc4Jj1e/sJn/v2I
BUanDEgubLXr3r9wQsy59OfcfRwncc7uWI8rR2+GL5M0Jdk/4Gu7H+HdufSqqeGO
4/oxi+VAdrrjvmOXUlhSvyPUcQHFZeyufG8KqcsFgd9aNY4wbzji/ZLrGMsCGt1t
uHmbJi2BHIu9E/Pk1piRd6VbMASDkipLRaHZi0kba92aLuHk7CGUmCnCvgB0sXrX
WV0MF6ipeRmiNBMx0Zka3uDP6hUOhmDXWn3/7Z3bulUu8cxS0LNb8XJqcKXxJ6v3
ZbMRWbsWXTfVClKEfRWvNT8S+N9xU5KgevSx9InKPPY5hvi3tC3/mIYZYdaU5VND
yfCGQkaDlRr4TdcYbCwIv30MxPut28jk97f9y607v4cJ0qolqsGfrt2+6oONA9y5
DfK4wtox/nyY23KouDMSYuM7Vqu6NFf0H7BslOk1fB1B0Ax7Zs0qV8fPvgcJZndY
MTffLbYJv+UHhdoJZ6MBpW+AikvSfAlTeEmxbuNydOUXV5a49mAh6WFr+CLTWNfk
YiPC9n6CCUW93xYrnzqBqablRY5zc7h4Ll9LsWf4g2nPlmqrkFdkMOePG0AH8ia0
duo0JTAMhifyb0xyUWabLg4QB6PocggwVCJJYk0N0EnWSTJzLqJbWWg2eRyjgMJX
zyeHHRAd8nJf3pCQP4K9jNNT770svg+TERnt3KXA3GKF7yd+jQetAcGGTTJg3yrX
Jl+Sl2A6Y+49YXl/O1LMXtEHU2ITkqvEFNdbEOXm3PMNo4syCVjTXs8/RPwkuTB+
rhGdykhK47PYZDGprtNP5F27MzO2DOWE5h+3ORsauZkuVSReOv5ig3RC092bz/CH
4XCAJ0G7tqBDlgWbFgVfxTrkkh3wn1hg2FvpwbQmCSqWgNTa3pZ3QdlD967mcnhs
c5JYrRLiLCyM4YxEx/6J08fbzhPYP7lvLghDrSsFwA+z/DaVFcV40Ghgd9nEGpS4
bdfsznkzblD4D9HqAmef1N8drFn+FVHqqUaruWva7EJ39CpoqwVf+lomnvUZlSTG
pP9rAqtKkmEVUrRAGXSEjGRkM1tC00BEhvasp+wPJyaY2mDlwTkBNdAHW51dPsm1
Tkp4essnzt0R5z813WPJ9mVsKDPWkxc7JAIL1xS1xo4EWPGi/Ps94e/QXgPLIIrP
JRoHEKN4tWYfa/yXFpquBqO9rpXl4KwNxjhm6C9uebheUbHj6qOqU+HqAGLjcltQ
HpsSqMxlABeycuHoBBjqLeN/TRiGL3BVd9XIzY3KUmHWmM3iyuQWguwJUz0ORZ7j
gPWmqvyvIgW8axMO1N82W5h1rZhr1ag5gV/JCvNANE15JuiU1hYaMeFSAaUSRwEa
OKi7NANXz70DTzHppo/5+HGIitI9WOmxLZjLrbu2ZrAPF+Zvo5LtezDRWtPBxO98
Y6tI1rwubajVJ1g1UbTJ5QlW9EQWmh1h8JUNTqPfCC0DVV2XpEzAKrgvSZlpUQYV
q3fVzNamxWusBsmiHk+F+tJYIQQIOt3qMWkRBDV1lptepuZd6SWPsD988lP3sNYn
0s/S2RSwXbdzpwu8KZzfKibe3hyu/us0lXkcIaKTTr8NXlnbhuqNsZx/LDiZaI+e
JdStUnSCrPVBl98nOOKXf+DQYjctgVbhcJn3xhwXfGv9B7qBN5b+8fHSoW/NI7kA
flXS8EpMQUzV44a7+GcJS9rOT6jMqdUAKQ46qLygx7R/hV/9V/zZANOFHDoHA98k
G1br1HZy3L/xwWyUG48NBucoFZUWB2SlDtoLJ6T51YnTt7lxxVk8sUeGVlhhs9RF
nX7rHeq0dzBil1Xa4udLzgE+VIjwRJwPY6g2a1RrpQ3/2PLBZuIyxZ1U49ezlvyZ
iSHkHH4qONs3V2/hqsw2Dglun9YgUwSjta5HRe9kukMImh67tbsyrPbgmnYdoKwq
C5n3J8FPKCdy717ceuAAQuGU0aptA8AGKAEtnhIDiqELRypnCNG2qAyKKleF0Mvz
J/i17v1M+ZUwIaeEImMBkMEtBXcELpZv1NspEC6bAOaN1K49rNjDm+sxYypbLyyC
a4vaTjwesdAM3E42hDKzQKkosmSHvs71RhfNHrXhTCwl5XVNW16uoNORYcE+B2c5
0fXGs56TubFk77+MPgGfWsg82vAA1dHaRizBMHtDbtWoVDJv1qzTvP1MbBLt+fOF
vUfhGdkUFLF1VQZOrq8DYgcalkQcztEMgEopyEc3uIkE0kL4EWfhvSwH3bz2PC2Z
XNv8L4Sqs+HkFc1qeaxWtulh0Vi51VdzhqA+zeI5MlhE7r9ANfMMAWkE3LzTxrkT
P40YL0elInpopWXYVDIm6fl9GFjlCK2myvNjG2Cp9FLmcsFrXqhnLwq0/uuvaBa/
8nafALEKN+L91O6e1Nusp+AyoK/lKwG6Z/Kdjuk19VUnR8jUFsGf4gINPfYe6ujM
Kwep2K2MT1FRKTUpGGFBVyAtB4+5l6xaJ2XnOl+PEFxWyF7PLI+Js8hr2TMTNWdM
7ZVZ5tt2DknXcL9mLt5HluXCMZtY6qZxNy6AgxzztixzgTqf8zoC7xTSCLA1H3NK
VS0HI36QgfsqKPzlLTsu/0LUXuQID89P3a+OnOAolgyx0txTZnDln7G7lBelnnw/
rLKPwsXoGp7ukvNoAfaXTGWwtYr8lKSQufX4Sk5dwY909GvVOYIzFqz6xlUg+Sw3
1geLiEodrJjiQDNG/u5ictPnnCZdbPQK8m64QFZQu8oXmRRVVLK4YHY/lH2irVzB
tyMGpvnui1Pg3dasDrl3S7q20BC24M//sjHKdFyWBPw4o8d8+juB7y9ekvj/Rk8T
4SiKM0kbavPHgiVs6fYmJIC7MfUTBKXO5fvCJGcl1c2ZEmtoJlI7nImN1B7a7c8f
lgJ2iJJs/xvk/gDaxyVSFOrAbxFV4RIkSKeNpGwitAnqmMQ0VIpYvka9D7QAsOJi
Izhx7ScJ1y6RNADGD+StF4MUDdcMRUMoOsEfgWQsG6H997gFz8W6I63WHrHWBMfw
xjeE0F9BkCRQYoejiEpdr3MuUwayc98A2Plj61nItzhwCS2vtwBDUV4vAVO6revE
qYlykA4+RTVx4+uRoVd0dxnezGufauFR2YMV9sic9MktX/lF9TXwq5OWlwc8tbHR
d9+DjBmyrXMAjNxUnYWeCyUH6hA7atdBiov3uJVavSNvyTKt1yAiZ48AwB5xDTZ6
D2RfBaWn4mn6cplm+kndgYt0+rvZBBOvzmt4WwNkbT9IZDMyLYOtbHnY7zX31/+t
L3+CueSg+/B+M6K33VXd5EfEgDDXg5bMa+Sru1RANYMJt0iF9r/SG9CV00f0DrxA
vVXLOXTql6A1H2EZIvy2sLHld+ruMqXExioRKTVUXaDW1Z5tnwddKwVEoUfn+Wx3
w+aIIFJ9wD2jjMI3IvsfEG6N33L9KSf74sEAZxG2dnkTSrOg3BfVmrOqgDpL51CT
9+3/UoY2i0EvAVbOdSto+Fm7ABpV8H6VtLJedokn4Dg1CBUe6RDzz6BsuzxgeIxY
m8IcL50WYmWBGhS5t8gBeE9cU8J9k1L/DM984uvU8hcrhYPfpWuj1I9+iZAYgJm9
k2pKyvQGa/y2vFiuQ+QyeNeA173cTuLi2I8ZzW+gdDnAnwWSsu0d1vV2MtnteSbQ
LOg8XQA+wj9UzvDm34jylO5DBnE1dfl99XVONaCJJUBJm0jvXzHZ678gWKsMS7Yb
GLFYjEEpyqkXlDaYiM7lCnGYDv9HoHcgQxtRrnOVKb9Jh8yPLHBPFiRaz239YI/2
ee8kURN4l0DNBmEol2Q7SdwxQyRnkuUB9N5d4dRsRyWrWUBvsWaEQ5HogkKmthuJ
6S+o+uFauFv4rOC1kRabQ81o4DLP0z4fzYjkEriFArQSKwYGkwaRcPnKPrE+JpLN
DousAMWOKAGWg2ZGwkUeD5aBFFa+fElWq9mXfBhGZH8rUNUwYIdzM4UE/FSSEFql
Vam44hW89G00+AQG6MZfJOaUYXSEGLpfRBI0pAL7WcGXfrF6g6Shf7X4qwC3QLvo
H72K28Tan3QHZ8hk5z4Tnq9uq2MzHb3a9x/x8stq3oehIMZIW7w65wX4j6Cr5UGG
uqJ46obbJlxW/f0wBrBKEVIBaeXxZxWlHek0JiJsUchw/12y9yt1gtmwghx01Nfo
8QK2RkrDuzVFQOk2YSdieZsnI5W3HuiEELnu2QrWnsb/5wsRS3/IAQ5zJ1bzIy8q
/5e/1agSNns9fR4i2DA5phxlvZ5soIq9uIdmT2gxT8uwT9JQqHNb8vUK0omqa+pf
mbx9QVNNjl6wnjWUcnhGLu7BHEntDF+mVh1bmClWeH9BXy6OeRGdG+zuyFgsEvtO
BvbR2EBGwtOCY082bXsM9eH27i/KcOvD3O0sqF6yDSYADAwT8xuf6laaCoEtsNMh
26mZjhxCN4iCqayEdpAgWgR+Gxk4agVpd1TgAvBjOkEpfqZzJmPbhO3rH8w4BBlt
LUKD7UaFQdJ/wdr+XggcUToV0pCfC2J++CTD91ilBB8XxFgsCduqpLAMhGSAeUDg
yrs8PDKLteacKQn5/7c2F9Qlf5wN9d+3hMY3SHQeaglKLT4YoPj5w1qsD5UNSJGL
YixWRDuo4kRCZVGWnB2S7HWcoFEqe2YznL6hbueozSf1Y09Gq5LVGEbG7SGoc0ZE
0MflVdi3fDTL4uSubU95TbUMOpCTPIZvlTsmCmLJ9UbMPepbhFAI9V6qxw3jifsE
CWri1DbgB/O07GG9KxdtodlYtRTyro4V3c8T8Bwp30gVb8DAkYFSoMQO3kUDn1Hm
Nh83bGxcjib6nrGTDnHKyZLkTIOiFDNdrDnxfhZRV4in7AdzXTjWW7RXjyXmLwlI
rpCozXfGtdqec/GgdN6z4ZFwDVEVjpQW1yiVS9gUJkOHfgmRNEbnylW1NPev9T61
SD+OHtXBha/694I8yhgrM5WeaNC9dzc3aqAq9I4R94BIPjz5bNWwE0QGveNtD13c
93MWbXK8tJL8tw9pyBsisewULuKPUpJcPI2ixM6CAI2O0C9xh/oFLcQ18fICg/DX
d50U2TewTz3cPfYImSrkIaZsznyRmVIBSsvHUWZRmv0+jmftfj/Kje+AxTxiwfZ9
cuMJfe6oCzgrhcI4L0BUPFUCcufXQGqtb7m9R+0yoLlwBXq656ofqzEoB7/ScAVt
oWON547XYZ+9hYptP89RUU1am1DItbG4RAMsyXqsGbM5ThySAM5rg68EbCMrZUBd
eVcuS1khwkCOyqU6/UHpdJxurZH4afkpgE3xI5dBHcXEwD2cf0+y0GYP35m3elhC
mKFrpE0y3Jmh8h20ulrk2CdQuSSPbExPRyz9prlsMZsAtFOjKLPO0JhrPtQZ6H7g
/RolGHIlQlhKHnscSCAeQavBZ8NPWXj7h9C8gHP3TChqoBZgEQiPXpePnIX9pJbg
zHjhOiPQ0dik5zk6lJiHBSKQ8TiJDW5GLZOzO+dmV3RXDqHnm4keM6853NyjNVB3
4f9jkxKmZkVEJcS1tYozPu8OAMjJiQUJzfeNfoXAsQCX3/Z6G4UTeAAmmaAIS04G
IVppQBTfspP6weLoyn5T4QkCll0ll0FVptzsSZaMLF6+9j3K9OTnHUKH0MCrJBxg
MU3ADRpd+hEAQNveuRZohOgGnojmNPslHS8fUH1duHZWppx5UE8xolApqQidhPdN
Tz9HkLYArt5ccsJPNb3y1TK9QI3soEKfbubXCqZ1WNJJX2AdPkVegZc3ypMwnTh+
09i/cr/Tk+Js4VVkK2Iyvd2xd+RKcjSbhiy0Ul87MC78D05coxW4tDt1OlZXigoC
528Sa5WnYyqUn+vUl7lxEg3PGSKWUs5Zd5SQBjMcFkAiiF6/NZ2FI4LSmK50N0FA
a/8ve2Wl3gGrmsHTO0/QnONviXXJgczA/B0Eb7ONroXYLg+juq+32E98Dc9NDpBY
tpIz3iPNy3QR4zw34C/hcBWUkDVDkXMfEETD2U+lExALjAzRiNpKa6nfN0CDSbb2
UF9pZujShFHl9VhlkZe4o1XQFCTAsWZ/OdlywEwxFltEpg6m0IFzM22oG57B3Huw
ofdQRDkM+4GqEH34FVjxazKXdETw7VK8g5pAzKV4nlqhF68Lggtn4tFR3E6hZkRx
Y0VevzTaHUfJ13zz3h9oMUwUI9Zh8a+Ds8zR6yM9JqONl++TXXI1wNkj5j25E3YM
Sj9T4F7qMoXTVDimrDM8n/3DL2HtyMbf+HIoLh1brqEEZhzMd4L25WK8c8Ndw83z
ub885YkDU/1HulUApEa28gy7IdLfppsX8yglVoU+LKIVbjrAotuHyeXZFCYbj5nc
FKujWUpVbPhklah27JSCcrNqCwuHXWkGncOZgDeRbj1CumLDtyeyAi7Xlrnt9ikr
IU3Zk66Y4BcJu0Ss337MyqQRV7ed50Gz79bfTM/wKkp2DkTA/s3dv5grPUgAp7uP
wH+iGDJoVD0DnSvUmFZoGxEamyGfI+nBP6cki0GchaXZI8PDIKYHHd9v01EbxZfS
RA4Ca/sJCxxCdpDYsR5+cGtbnIICI9J/RNIojG4O+C+I/jh6soIW5RyIzMG176X+
muWTTb89zqNW+HL8HukZXRlnlV2z1CFEdlxmCoqsEOX2l8jUVfuiVD3FNvNGNmIg
3jyP8hI2TVeuENun8TWIVlIwpabB14Ar2lBC/MY4QKCDn5fQIg2tA6piP/nj8GvZ
1VBj5utyWz6/TQX2UlqTL33gxesDYoN2aFt78Nk9JTzIaMgIrgpEPRgE5tx28d4k
8aLwKxyxxspGimOSJlQkLoovNOG8rK8phs1fN4utrGZ7qDWbGOPI7/PVABpxeCyO
a7In9GqaYdq/W7Ph2qOK5jMLLC9DtE/VtvwTqAgtlMKE1I9Yooc6sc/S7d7O2o8H
o7coalePH8ubHbnpUjSpk7So97gHSxi97aqaf/R9e76yTPzWIus3pdUZk861CMxk
YH0xBvCRUEB6xCetaswhB0Ayl04qk9lIzew44DPVyxJYEUXphDSctfIZAHsSKeJ5
HYf49vpWJ8wbCPYAAluh6Z8XGCxggeyKsrOsn3UVJIEpDAGwuuYVAPxLL7K7RE+6
ubiZ5TqvssPoPP6fynfn8WZ3OXN3Ez1SsDzTPuNq4TJ5n6BdJEbMgSXLXNYksp1I
1qybVrDIHawxzkJOhHakA+MCTpfrLdM9Mim/n/HvPw/wLrGqqdVZz6RLL0AfbKOI
Pq4yPesLll0KM9Xgj0r4WcrBBF2evdxYpYGR8vy/ndQWt9dNUJ27eEIRHecFe+0a
iWgM8hEDlNypb5PFKspyVMK9eMg1B+YbxBW2RSlqHiVv18z3/XQqTrEoJMTjdk/h
sDAn6EJKLHKhw3lvqi15Nb83G5c2ffStka0eUfwCvNhgXD83vhHL06ZukhivGM+b
1V1Eg1McTfQ14Var8KqstgsKfuvA3TfSW0RLqNVfVUmUqRzd8xZsaAgToWbcOiL0
W/OZ92wDzWgGxq/I1UH6bOo4a2e4+weVffOE5RLMF4oRsntfGiT9vfco21zLIVFX
1IStk+4yASihwBSZ29aZV2VoFnQbzow/ip1/mYjB1Ib6nnBRU8oI8MG1411CimGM
cLLYROlJGwngYh3WTZ2CTEIJnk1alkAp8TbUmPTnS8w0YSJf9XBLQVxSXVf1FEEf
9GKEHqBtOTpgLZXzpStrMScXj2iNwP+EpGVjrikESos95oUMLa26Kdl8s2MAl1vD
UUr7gqutAl03+4vAFOtAxTsH/14oLTFwFqZ3ghI9R8j9/ugn3qeMUbNmQ9xVZUWM
EoFCm4MWM2NVpuzG2joyznN8zlAeARmpi8/Zounm4OGyu4vDnr4fkJyNHXodYyKT
05GLJX8zUcIYkRRNcXSCctwIpZLtpE0JGx9dzNwGSe8+D/C9HY6qkFvJhu0tt9Ae
obtmmdE/6j/ZbJIb0G632uKPhyGzD9QPwqjFEuFkWacaKvluaUNBA0p4NJwgmFQy
AVfXjEdz+CA/AefsEZqhlb+J8eon8O65NiCvinYWhYYiOejKJpTyS9IDaIks1GXp
TUrylQhNemzG5QL/9ncbVLjEEtTwX+cPM3UXNClV4UpPyUUIRR1Tluhsy7Wna24v
UFos4yTg/uet+dsNsQY3bzFQ5QJMvjdzG2/qyw5kRn+SEni3Bn7s4SHfhFZeoKNp
DxLpqjx2/aMK84CStwjgw/ZbhwNlDZe4nALl28LhLyho6ONmoft6ffnrZhFJZYLN
WHPEZIktxyIVL3az7VXsvTFWAVVaWllyP1sjVpsxsCMWU7O23pGa2L8KS9rqAjoo
zjb2sH9EPTRz1fmlEyylriJrCrBpODCjDcJ+MC+dUIRnsmQfv5paEGOKzghlM1xp
MDMY3ojLC1Glt7cw2RLzWDNiL0SgfWJEdnyl7UHYBgNh3hfQdaHkA9BkrFMSzL34
vZoZC1QtEoONJj5Bd8MfFQY8q+ijBsV8FnjsvAegBOlC22vOfeqrlB+RzMBNEcZz
kFIaPhAmIsoudwL2WndYEVdRib00ntOVt59zGT1GEAEVI2STbIlYKq/p+kK1bPph
SFXFKq2h21kVskm+OGKXadgs81DlPWyfP2oOoJShmb8ZpNFhtVeElRUiTCJllwv3
OL3PrXhOx46zNVJFLJ11Wby4MOaCXUdlOWIHE0ZhfKbOdee+DqxYZiDjC8cQ/M4Z
wrBgswqk+Im5K/TAgrEHBLMWu5ulu/uTulg5ENU7vfQs46lL5zYXEcxqiCzCQsaX
7btlTjYbJLt/iKzNdpRJfNa3emrSnT/D0jpXyTEBWOrvNdeLxRIN8cuRephfIZuP
KLHFCyt2sK3++vbrktiCxkeAwuQMeQAobeQ65XfXbJy52rlOYD0lOU2NOeGGCc4V
ibKTJP5h1SNjtgtzrjhma6JZFnfvcdFigi8l0VIA2tQVZQ6XPMAOE09q+c6uQdiC
INHc86tJ8W9DqTyJikhIPHcIYRcVgHyop4hNSViTVBoyeOqQCohe7/4h9ntwCDFv
ek4W8Z3X+arx1n/tIfJoCzmpDnAH16Y9SX/Vk2mLXGLsjXTvUEIis/bg9WOuXXqA
wCsHfqJ+bR1DQjOejMiTkM/MskT1N72Tq1Rlh/YPbXyHbU4cWSIoTYB+EL6d7ED2
qSoFhWW/EimMzeOkwuy6GCbigHiiGkx8x2xw0bSfv7JVWA9ehMKX0DbqYTf7PNnp
l38Jia62JBCrrvK9k+0wUcX7R+eA/jWfLtcC0yC73FmhaJqZcPGrm1rJlFk5Qcb0
uDZhjMKKUYh3LB8RCvP9D10VC6wmsxZ+xsDuVsiPHmH4FApD+ZZP1yMzpEMLXYvf
ndN5MGBjUbqq3sUVO5PDhtFpT6RMQAeItLReSAn5DrmyqzvEYbdmbrf1QHWlDcGZ
/i9eq8U+ZgY3OzpQwVkf2FtHliQ9AsBboJeyvYjAW/TxU1iAh1Yy1/4WGALqMIGf
L1WyS8aiCrQQQ28a4CIzSHTEtAX90LPJaQX25c4vvWWDGSM0GKyN7FM6TW1ctQYo
GwjcZq90+7yiBQ3ZbApFmLjb5jrizuUr86Y7O16uMhmFSGOxAktDy/GxQ3VmDd/8
YjgNEQviS49jKWgzLxZXooggEzxKJm4UlVswy9xGZq9AmgeQyGXfvjUu7dY/EyKo
8O0j5gVnfuyQkX6tiYuM5ELGJPpLwDJ8yiiLzcBnEnvMuv4Vi9j3Bd/iOOiDHjPE
HhNggTrFgcP6DC/WyHFsVrqCDioLlRT7X+zLmjKCwn9ziA9/Guu5DmreT6eXk0qu
8/w9LHyJGlWHuUD2Kj98I38AbKF5PR/u2yYUgQsHV86vjTVlAOqrcv4O6dQhb1UH
MhSwF2s9BVcf/COeivwzcvkKbAh+WEqvIUi+BOG6OwOttDcByCR2VTSvJzsOpda5
ZphcA81/GRa9fNTltxLf6HOZPttbQABY7xVvDdJJ4djQ2ICtkHtUUi051PxK2/xN
gf3srn5Q73BrcOjz8HSt20Y1G+jRFA9UweuyH9AwbPrpgV+cgXG5n3+terK4VB3V
tXxffbRrLjmR1/DnrBDGpnPPGjrdmeKZVBxF418i+D30KV0h8vxd6vtZoqqpMGg6
y8d6densFKgCEPepUB83bbP0NJhnAgxrhUig20b52Umu5DobD8hnFkK8gBQ1if3L
f/wZICdqeWIDjryHr6ljOMYD93crvM3WysWsXsT7vVU2WO07T4VSbbMszQIxH770
Y96tHJn4yGdDi/pYHcwBN/ke/G0bEfjavcIS7CMGJzIYT28EHUMvDezgV+7cXbN9
EYAjWa7KV6a6IH+g2EAyYEB6QyMc+efn0JKsi7DbU35aOfP8DJDPCadjZ1hhZVsA
8tOBrhuDtbZCBg76Okff/hx52/W8i5UziogtuaXgqYuL4CvV3sNYxL4avpTyNLRI
rb+ElJbu/YbfXK0OXy4b5whNztQlbxxyPKtnXu7camCwT39JK5aesBhOqFTVj4J0
mnvoFIeTkTgh7emsvuNFi9JK2cWvGc0AZrfAEBig15g9pVMVhyEb42vs347X0VCV
enHhdVAN00YTWvAXA2s9V5tcJvKuULGMW6d8Bsj3obA8zziL1HjROxEMzmaWV7Xw
UgRz9c1zc0/LxVTX6ZpgusHxUfXeMCVdAKN0kE36OJ+d+jurCG59OkSApXOS3r4/
gwmhDIBaCtU1aFpMO3w/OhiuXVHylnu0XCCWgX+ikWc+rcT5lQByrWN6ICKrPPbX
ilBIj6ZvRHuA8A2SGkjvhEPHys7F1iJXYf7zda3/rRAmnVFMQepmXQcTmO2oyTc0
UCMyS38r8xTuxU3UA4l8odUou0gAKZ6aWPmVeqeWY3mnPeAOOI+rIF7Y7djF/+Gp
Jbxrw2NLXPT8xp8joLIxQVWvoFn/FzYeUMZAv4cTm8clkO0ITKPa9u4bk/lxL4NM
Qp6N5bjGosy4x3l8s7Zs4saeamC9FAWAvGBG8wVnbHWqAcIoaljOgylG5csORXn/
9umiofIeCJ/xtsZ2bsPxNluxASErXonhbhoFjwboVbxlfwypL5MTtnf71kGih3GO
k+rMzEybj6GVP33U3MH/5UKQbi+vUdrPDTcTAJKC32RFo53uYjs+FFDDAFOQ6FGK
5dCEWa2mBxpqXrvq+gv1EtqCXlUosOm6NnRmU+3a2K6XTIG5JQv0wLoeQbQ3Jb4y
pIueGgXYqNAJpjcI4igGswEJhMBZwFN4aCuBxUOCfhvwMU/2ZFa/ZS4FWUyxoz0F
te6wWUMRdU0tim8rNX2JS8j6P/UsbCnNwwLfz5OSzMFUvp41alOezZSPnsBVX1nP
Oy84BZPDaHQtsdAe7z0Vl/5XKpPEilBdYAau5sEOD9D7CW0MohIhmJZv2aRNJ7TI
/xe364fWq+jx3SmDW8oAgTpDOfc63sHsMiOqCOdQCCPgOmKWVSTAbqL6MhLEdXuT
P5ZpWCD/j6xx8CkuyaoZQQpm9ox3DOuQslcJDnNWa9V85L46bp0Hvm3D5dqdw5Yp
FrAvjB/Jtp0C2tHnG4Xkz6QLH92kNjqODp6mlIV1FpulhEAAN4bCAX2tS27CbcZy
8rgDekys7RbX4ehzclKoAd2kaFMcukYTEQh1UUDnazrf2uPTki2uChzzyuW4Cwy5
CtKwRp8gURWsl70+rcf95TaCe/lAG7KWhNQozCPWNbQmhK0qJ1Ck9HsK7sFHqprj
O3K6pGjCDGAr8XMiQejvtWanzaD6wGmnJT8qxN7zdMdTVJqMkKQJS/x9/p+vjuAS
w4zl1rNYLZ6kdBMK5VhpyzxZro5m3QtCX9a+GmI0lM4zewrdu7++IZ27raN8527j
mRQ+62EF0XGnSFuxqIaLk2h4hr4u2yEQa+uw9K/ZsF4tKINjWk71w/t5zGUi7rLS
M89txCbRVfsIMbYGraavEC2W6y6mzIF3rYv9/qYofPt+N7iwmRp02S0r0pqRXDHK
yNGuh3Ix8RM68W1q0SQAR+b+NJZpUw4ZSI8P1m01ar/qVe0n/dV2Yd07M7Mf7GcJ
pgvJXCUQlyrkc4+sLkgidLTUP9tSODFKJEf4Bmyr3+hice9JiEvTSyg63YLB6aUM
WQj35NFSLRXD4JjOvUbY5jq975CRYTYRqmi3/yWhcDHXM0bvtRY/EQCiV9YxTpWl
z9lPj7bx+oM6wbgeBjLZYgcDEeEvauizaPUh/AJocR7lOnRwNQ3nfhkpyO1nWqim
7ZUiVGHhVVHjaKWmHTKssAGumk8vDJ64V+eF5FQgbN6L6wo/0RuWeOc1n/LcwcZ0
G8SkimPS/HS0qyYFkgLmPdgzSqc6p7Y9fjF5a7Rupgoa7k47yjLzA8RnUSnlNVNN
B5Lg+NExklvvrgqCspUOKNxISYqHjmlyGZAtCoVZJWtRy91CHEWHsAUrp0lYEx5V
D+8iNueraNLLqCIvF0ZTX/gd3N/HC0fH/TWFiLLNJyr4uWh8szCvHSz+uGGYtvex
Hyq0xNWiGYSK0RNy4LAmEjz0/W/s19NRR/U9crsEHKHAAeJDPEaQpKXggQws5+r6
0wB8k2Fth5Z/TYzbctZ48Cd8qP3i39KzpUDSLmtXjdLffuHPejf1KcbO59//Aq4X
/g8VBSlSYJmVifQqjZihZGnW9+gbzkn4iryjvkmpyUNnt9YW5E9475Id0mzvvAwa
tRtg3encQgGX4RtZFX1gLQc5EGhZNjCobjF8fk1PRCngMDN134119hyaOnOVCTi3
gx3VQZRpY0J/i9ZyjE23cfRa1XzvE2xFgPQXDSx6rmQURYvvPEbCJNcK8gfYUk2j
i7T+x05OS2mFusvehGsgQHxGDszE4aYUqQTJ9hYOyHjh2doOOepH4EdKPuEDfTM2
81yBHdrcdNnIHI51+dfJmKeyIrOgfIJQln6sJhAZat7aKparCix2zJgI3AyafAro
eZiMtbHFU9yCian+NhGi/puRF38svThi7ENpL3SUjRY7kEq5g8T+F+UCRo/Ep71F
iHxawpWXtIPbIRTtk8AxFEaVeuFFabAza7uCTU5nLyl5acyfi2k1LLYzxlsWHmlZ
upUoEDNcSuuXTZa42x7BEYXE/EuRvzW8vUhcGKvL4enIVBIaeJ7fwlKjfMdqbiDR
MoK0jsmoXSb98UjGblcVISEM0zUuP71Jn5L9Ga0o9zZNr9JF3ms3e5EkZXNw5OmV
k8Vm+EkJOSRIjTRTaGJ0P6oeqmPgPiIa3r3ksK72/XOxQTW89LGJuhEtBuShiGO9
wfhArPhRgrAAbDRlEj0CavCbgW4qBJ/stLzV3g+TyWgDrOAxARy47nEJTfAki41r
tdriZuVPAUeD5n4b31j9C7eoQPYP/6+dg3cGFy9q1zJkVvCGx5CFxYb8bNrlnJoC
oyo0uD+8kUvcXW3Z8DAqiA4x+INYjrta6xWL0PvvgF3668uK2TAe5j/zvYBL1PRO
WPei3zKZ/ZUBfvPLyifN2L7mFyFQl97sB/2fJqn3tTVRQwu2XMW9N7gl8SWGLUQt
n57TsJcURZ2F1jFO+y8pkzlIm+GR9TjP+JAELBFSbfsZQYc7SvEUajbgd093Yjl8
jPixoXW4yXLUMYc7xhOXE2BopEUOXuSor7PldjMgRNgtPW3GNiuY1CqEwzS/cAuO
ECrDFQbpmO4Gsb1jV9XPtdSOWZOfDvfokTdWWlsjF5SvBAHV/25yQq3PpTbLRDH/
bQh1JEEG0FMITkBMnfoOM/TcBiCXXK2cVEEn1fU13AP2lVH14dz1Kxh+PQrS+uUI
+wNkJFiSX0F+i9kMBQMsKomfZ6++l+eojT5oudjBDFQpR+IrKU4nuIjnGknWhsg1
jJC1Y3k0LQL0OJwKyjaztL+0dk/AS+ykmqGW4LyPfmJ4y4ZivkznPgclJFXNIBjd
LvBgRkLlknQV9JtdlIiJjYuwCxPkxuIsEtHuf6gLyH8+BpRcUY8wWzJ/h9OZn342
yNnB+6ZHJhLMz+3ZW1FXLQLzPfL0i+i/kEbs8Rd9No9YwfoKcTKhw3fyIM4awxbY
qmHiZmE+Kk425PN5i3pqom+Gn7KJr0RzjnfJ0qy7XSKMFHVNHzMSw+iAjGvN7pq1
sUO4F0iKhuGxwKVfZgz3Yyrah+jSwKCIYQ7R6SGuG3XEaQYrYDNib9q2zm4sdKcH
wCvy7rYLVNygwmYGiCjBeN2MRt6jrGWqIgQ4F/9KMMqCkbG4oxv8TZzIyUeUn13A
2rfBt2PRO9lSsQ+rMCfeKXREST7kyY4Bn4Vj993DwceVvUMsCkBbQHQrQVtbaqYD
SFUIpbUPpv/pOEU2Bb1Mt9KaAwtiVzr+XJ5p3z++YggqImWQ5vOB1mlFEHJC0vyr
N7pHLS7ae9l5YK/1Us/UdmBOabA8XDpfUDRY2BXTOtcwuoDqCh7yF157gtUIOtdj
jMUwN8kFeiOwG2rad6du1cfhx0AWta+WWYju5tYDeMMrmqGggnQT6X2Gj57x6Hlk
Zx9UvyiktpVdtCO2urvls2zgqNuHRhKVSpKZexyRvi6T/STirSVx1ei2j901kbYO
LDo3XFciwNbIGukf4rtAsOvRPfcuJPXr1lE2bIs2MbTkIqhwC1iGvar1u2xndDBX
bt7O6mZAvidMXQgfIv/fhJwusJxPhxaEAyhfO9kihNdxrSr1Sds1KIrWnwn9TKuD
4Ok5nxIsU1cLRMrjr8RxZFJiiWX0WHX+/uVGHc/CpQMJi/8PeCweqiy4dwSykHe/
HiSx+bBE9YWEyZ4k16857A24bZvc0ESKC2cnPxFN1501M3JfGCelcMhP3a9+B+p6
/K5jdo529qexpzNefYM/nhsWOquK6rCG9Lq52wgvXW9vOtkikafuv/npGY+nm1Mv
981Mbnge4/U7eX9tlc49fhST6qLJmQIf/htsxilkWIREe47Vo+BKrzy/F/+t8aLp
CAiLEofXSZyBfYvvQGbO6FKTW+7LT8WGHWuRVnDC8G9HRIKNToCP3gJ64VEvjQaR
a2eaCiv+hR2P75xZZzAgTlOnrIWUrrhLm2sdoxiVYXaMmK2PLuHfMDfxmIXwq3cf
kG6Jaj8YF+rCjw36hpKnbfhikDwHrZaCeaUY97RYisUiojmL/kQFv4nCKYXpaVjL
/Jh5WUPlN/Rb7Rk/QYDHR3inCp6c1WFp18fUg+IkRKEoq+qgGOPQ/4GAJb09AgkW
U2U6L2D7pKHadQn1qirZkIhwo3o6sLJziftWmsuD9GmtGmuCyOVploYW1USs1JEx
HyjwcnI/g0VUGHWIbVGke3nf1vM4TQqiLaR4ZRg7JR/r6sQ0cmdeQAGqFl2+KpCg
LxrkH/IBb4Zw/TYsHKtsv1TOpEY78mfPjokgupM1mJXE+r1nVhlQa5POjlrG3Dj4
9566lfYNizcmQsUoCkR5ZDx6mTHN4/d+vecFLMsejXDMLOOYhL+f7eFCTQd58aw5
cZQVPOyBkodgwycj9lToVcpcHddilEf1AMlL2TwIE3TVleZ2n7/7VWAVrNdZNx4H
xpPNCUmTsNj9M7EXK/+n9zAwFy0J/ZsuT2T4H7VP+NT+HcDN6Ipr48jXXPaIpuQZ
IGlzjrxkNUu3HgfgYmfvKMyKDkiv9NfkeS4GA9UB1/bGsXIXeN19CdeRiwyWpMpi
d4zvKEcX8PwuDQDm7LxB74MCghTm76qEJYTMrLNB65hIeocn9saq+DWKrpS0nraZ
diGRTahYd1ek+HKg4eNEURnKKqesSw7kYmWZZJqIl5CnNnrrzTXa/vA9q+ZLFuc0
4K66oQCtfSeMMkoi2drfcVncgmkA4nyhm2KbtoZPSpro2QXZr0bNHpD+hCHfMTHT
sX17hIfnzC+Yq9tS9/M7gU98MEfJMjpgw1VwpIQ9BiJUnzbz8FJo1O67+84KR+5G
nGWfxBJcrHkuuZOCwmI7O2I3AZml7EjgZG6TxmGPK2mMzDrC8R1MHS9vcbQ/Llry
YBXgZLp6Tdb0xGDZoYb5S3v4Ke41ZGieU/FImEZNqgQHNLsG5+uyo/NhGku2u+GV
++rFFsTg2dT2SoeuURk7/fKZI1njzUPfxWejl7FU8X0OCvOA1lOSxKzs67je25KB
wOODWYCOn0i+FVhucSUt1F9iV9iT/s+fJpGyboAMfg7SzxP3JLVkc9aKX5KOFCUj
pX3pzYF33Xbev8yi0ttwKDGOZlSV4+MxXcA7v/sbrDbXu1vAL7ewX6Wqyr2uIRtz
uo6r2zzHBcQUot2pUSWzvWfTEr6o+J/ozLNPmGT/meGvZaTAL94f+ZGSzzINdcB3
fWAYUjEDbgkFmpwuFgVuSekalqLkiTJ0ol3AeQAQvVK6yPDgdVGo2rgSDcw024yA
iIGprsbjTAGU1/BhPzcIB59JnnlqiNFJEv8EvuqbsisR1JuJKF87FHUDZejf4ulx
NztPOsceGrIQY66MxJCOp8YbuFz0HVYBEaUvv/cZfPxWozvJMp1YATd5Ne3KaJaO
VZ3sAIKjqASuMFaQLBkmHsb1RB2/984DaOilsH8gQj5NOrKR+dr/rGqQjLz2AKe9
St8A3Rpyb4AmhTDM4PmGMK0vy5DYn500Cm3FubvWMT8Nyl5KymkhJGc52AW7LdLd
KMdcD4vC1ljOATme0hE3DeufBnI9HeNi0OJOHW/OgkQg2YOsaAwNT9sfUPQ4wGwS
ejRCQomQiOsEsUzPGPqjReuW4B4xXf1uSwNujC+DJV6HuuA+DcTpidEswKWhhBO3
I2Sm3WFVswtFIe4koi1miJOcIrN5p/dUAOGbXymDCITRwXkn1W7Qy4po1KtVRbHH
WoxKY+8cISh7BACU/fjvAR41o2MooD79+ql3RK362iuNOPSADsH4FlY2EgZ/qUln
2dM/O3Ujj4MH28+pAYd1YkMFqYmXv098JZdcfrstf3D3c0yfFtjW5EDOx4WSmtgf
E+8fYOYqaCMN7pC2aFxRct2ecIQ9hUHORLzyW6uXujg5oXHw7j/8GkfOx4hnjoA8
hVq2mAdyKrLb3e0DL1SkCJgUlSsnRDNWXGzN2OYhKfEk7ngFSlerKSzAUIZnVTwX
BYacrtGkaTtQ1AUZUMRFvBCF4uA01h6yXovFGo3fVcY1rajcb0xL+m+YoNsavonN
0Qtg2xQ+U0qoDuirFfg3tzEaaGIzr70Cpn+hKl9v42cyeLkBeA8eIjO8MFNfa0n0
M6ryPCA0jxKBHczQN7DQqTw4sdnN7MZNVxLu+GL0p6PZTTOV7DZ4ggNpIyTaCxQx
CuUKIBupMLGsOk5RQCTCj6934cMNmYsiT5dzn/Gw5adbx6rew2b5cg5HkFZJDvnz
8NVaszwx79ELb0UgsVPvMXtsZI3aSMiovJ+sJQBm5HMIcxTRp2gwxmeEpd6UJq0d
/LoWfu+eU08MIdzBnPPKg4YOaQgHDMeEnSAuMHMTmc0sZ/evi6yARhhsJjDP62mt
qTma2EftHpA//Edv9KPOwej44xxGetFxWClgIKIZi2PCLghCYMEICvRgQKh8mzQ+
mxmVndX3gqAnjjlqwZvLDG9VtOtRxKDYl0jfkgCV30VTv/m0F/GR6bQYTeq1b/KL
FDjCZFit/JNMwvEKjsaSt/vG0fkJ+T0OHZml76oFZW4NaAXW7T5Qi70VbHrha0mF
+nJxcQcVDqTyPyQvfc+R8Yd3ygmzKpnt4ckw55JjVEgXBWhA0M+LHLTHuixBqsba
ui0Y4gwx5ukUJnePoQe1Y0uepXGrR34ukn2mPbHcrs8V4FVjbJGznWdurnSVbx0V
7aWJSNU4sW1AtxArFkbatCmq4mXr3r2z8Zq+fpQN+VyzscrkN6t9ntvQ+V1aY63y
rtdZFuVwYdMOTs3FWsel5XXnwv1HPArpX/tigHhWYszhJl21WlnG5B09Ovc6MpAG
tsz8eh66bMwMi8k5qk+CfB+BX/VFu9PW6gaYtPoCHNkqZn8X9ho71lBF+j5VhvNK
oYJVIKoFV7y54ywA3OmzIfFaYkFaAs6xcxkOsfq+LM7sQ45SrlZ5S8iLqOJbqoA0
bn6w8GWPWE6vAT5Hgk0BTT0W1afEweEnFJy7FEPcy510UdckYbS9xiTg1owFFm/F
1ubtpnXPOxR8mPr1xlGyXbFsaMF/04feYwVge/v9JnsQPV0Egu8JKnyQxbTGM+Qo
KEYxWiGENLXj+HbSQJun+y0XFZIwQClIMvPGLKh66U5ecKA3kbABuFm6CMruQh3+
F71g5JUxVN6GM1VI1BSHYTxBeFMNzv6A6+UzfEYNOt9FIGjNYUmI4Li3rQvhLms0
pJ8aoyCh6n6Ww6HWh0Whq0YtshrA/4zITliUH8/sJ5dVBXXWATV+5LfcqoH4vdxS
cwUA+9wfDWI7cAyHRsneTepPzo4hrTqknWAsG1ldzoqIgf6RXhhIEaaPtZ3kKI77
DGZMxxFjqqyiRJelagUj+mixaByaqzQD5tmDVV0os8dJyg5Xl55GIw7nU4drz8Jw
aSksqX/w5ys8hD19gBNSM065X1UbT3tjPI/kg6kRot1eSpzo0zP0qlMHmgTBnTyQ
Mk9FyS1780GaaNqQPh/uRaWs6emcf4YlsfU0CZ98wHLReY9F5ynzV6B+GVc+D7FS
kR4BcxN4j/Pi1jQdDNWbTBUr3bBSsn7Utb9R9Xvid1OtKYIyMF02nsipsSZnsvo3
ZLJ3P7z/k7LnJqPNcPa3Iau21pHKHLSkNb5HR1VsiTHmjCNuhPPISlID3s59QAiV
ievsliHkY6DqIDWtYAUebjIrjxKR7x6zavNIbzDd+BgLU497PIOAG8jBHutbhg7i
zCkiDeGkmCwIpVZdhsDHrRdduYe6lDwsni/nkMQjj2aVoA7uSmPkETuZ9HNwR05E
OCrJJpBkLc8gNjU+A4y3GhiaB40Uz+Ga4zcKUi4hPzH/2LQbIGgt4LX0v8Q6UTy0
vmIzCdbGDbSJR6pXqiZoPdoSUeu4Vd1PVnelb6CSOEhqIHKYQRBUOvAzm7wgvbxa
SPJLKM/hl6anOW9VT9nvVuS7cd56a29NuBa5vd2zRkQ/DyR2E/upvA7PJyhDYu5W
1iaNOlaCeot69OeHDQDCBDkvjyLIIILKTNYcAHqUnnG1i/zL+lT3MNAwrvUcAL3Q
gtmvvgcBgwTN32SMi5qvIBCCcylBXTpgzmFen+NT+W+dpGltjB8L4jAraJIda0CI
0h6vcVZfKc3tK6X7/wkbb7FSPJjv8uYD18i/W3GKy16JlanugaSmQoBosphM/eMo
E9ltOvgx/bv8B433dF4CfKP0FelJ1tI3uRajN87GOaqxhXPQVgAmBfiMxhmv9uge
SCVrYBUR7dQqnINy/qqK2jVDDX6hrDzDf7Fsvt/8AWGPHE4gAkuB6g95u8mDvYpJ
Wryj2RhdeSXn55Uqk5FHIOCELhYUZghEb0KjX5xQ1dFP82jzBykgru0FcLV4fFv4
Ux4XNgeFLcPlMfs/GMlVrCXzm0Y0S/N7/NA7DKShlmxTfbi1Gbt1C/5n6EJEuj/T
LRg7giN/+QxKmHO8j754yCMJSscRgOvKp48AiQ+TTx56JI2qrbFsUN8mAg9hVzH6
i5dX6XtwLXUKvByY/INuLzsMeItgsCQKFWivLNlEVg2KZwVZnC0P3DJf9zgq/Wwz
02e91LBxxlA70cUeq9qIYlwrmJTYSHgg8JrGCC3wrQ7kNvPTjbtDLHlNaUMqLOOG
Rgyw270uH29kgrqT7UiieKsTLkMCYo2ccdWEQAyYPOxE/jej+L4ncVDN1TJwTVzb
CrcyxS11fakWGmATUevsU27xYPFnNuhOLDsjSoT39LQrRNwk8A/Y91FE9SAFTKLH
SsApxQlsOLmllLleDbYJb/eBdrPr1jfh6E0RJdAI+wBqW0c9xkhluZ4tT/UdCjPF
4ehLmEPgqvPX7L0s0KQ+178WKAGYWuZh0k0Zk6n5iCNLEyqt3XeBjDf/PySgEuq4
pz7GY9vfHqKzOYveRV9JlwzL+HCROSQXGiRDalmfmTzCvGTubEWLyaCHn1Gebvaj
pYDxF67TqbjynQKtDjKTIy5tHnAF/BPNSMt6vp34NjTF1nqc5bJOUeShCpVRGd2B
Wz733B9YpakLf+I45xxl51/Muv8lixjlw7SUbz0UtGyzc4Yqr9BIIMHRi/BStnee
ueHDanwMQL3yc3DWgTe4NuHvlQYbDqUhF0npKEjJ0yTOWYIzF/lyb19uZXf/SRdo
8KswQqQKCgYT/FzOrSwwAXNpRArTGI4bYlQ/EJMHTpY+x2UF0h+OnmcwKl0Q9XIg
UiB+u5Q0I8m223YrhVsErnapy+QVMkcAHuqg/SAf65p23otCwzOslAFo9u5FlbEi
ONLfGxcdjcEEA3zIVV/ymki9lT8at3GWSzLbBVqk/R2Oq2g9EC10G6QH/WK7hTMZ
v7YVI5Yhl3pIJg/hAait4KDPsJ9cqqfmG5XZtNZ2xLLJW6KWsG4ArsGgC1dXJVYT
XxHT4gWNRW8aBOKZZG8fhY1DgwVfdTUo8HSyRljpPPiB6kE9Lw4sUDZpZnGgoq7V
6Hm/24rnRUgc6PGiW2kiJXUGtIHmiZPt3t6Qci30a0GG5td+1YWj2p+S5ynIB1Nx
U7sHUI+y1PA4/FusrlDmvaD38HOuFZnf5+hHEoShOcRWDyi11N9PCoFqdAkXCKng
mIvavpZUVx6HKH6pSwgdshoR+fl12INgZb8dM5cG6Ahkt5VoFHAQ0MFiAt9xxgZG
eZd/W2qkv8hzwa6mxBXTovCE5PGFTLfq3g8vCsBP7lk47O1793IFXih3BGkRLxNW
JQ5mEToMfnPAPk71F338VDcOdNQk6BjaYFHL4n+NyabJSXfxh1sEiWWpO5SQb3eA
4me8+UUkC3kIcM7dS6opJxbHX0xFfmkn+TzcQJm4nyszw3m+GwymumHhmPZN2Z89
IcORAyvlBrRhDquo+rgKTkykF1d//3w+BQ0YAWfxnwdNOGP1ba70dZPnfqQOrrSY
4gW1V2z0tCNokWZK315lSHjhHeZnrVLkdrUuCJAxHEzFjU5Vejnph6L38E3kIFjm
F748nNWcV2f7E9LvEhO6AQ6oPTXOnA+55U1BWkouUvHd8ZkmhqIVldpAByBk525+
l2FBfipkSM8XRmh6tk4De/aNcGkXaZ9T8lSbZjAFXWsNni6Gx+7lAGpKokFteGZe
ycb93OQmC+XMqNXyk6uWl7cPVoRkqhNVngtSDsZ6WGaOahpbjmyA0izuh02e4GB/
lCCu77p2GZG3l9peSwqkn47ZuRe7aOYVwTuc0usqF75djLUOgxlBVRHtyIuXMpnW
Q/O4zUDI0Is1ZEo9Q7Xi+YUPHiIJMYn43W9MwxVpd8o2N1EdmOn3vDRsFCT2JDU8
+vL5OzQjHZEw2Kiy/6Oh5V90UmbkYXzgZQmX8oLNfXiDX/87W9sNOSZcVeLRQ/cr
0Hj7oEy7VKfA0sujUZ7pHVl4XjllYpMt+XixWVdIYV+yQKFeYtv+eZGaj4rRFNXT
S/DBA7KpQ5u22c9CEJVZ0fe8k5BfbkLdgf1bfBTJ7WnJCSNqrPIV1Yok7rHyPZQi
ZmU0oztLuQahKzEo/ysfLJfes6S8ShBzyUrzvAXacWpixhgvlGCzbqTuhMa76tuf
HqFkVtQK/v4rq3uf+SKZzqxTB0Mdcs8R/zOPQGT8TWTIrIoDltEmfmuavmLhTRSs
DUL+uF/PFA5QVc/4Bfs2hfwO1QN3DYV/+LdAeKCbY+pvpVY06/ltzNkJC16xpLek
qF0zzBmsk4TgUqkXCXUdDjgfAXJvnS+mF9LTOct/nElxgMCpiSAGzBlRKynfPatr
sAq/cGOLzw45pUrJiBUzF7mWr4ilrNclhnJdJ6wjmJziTfDFeZcPSV+ZmFSYSsRY
yhYZSPlow6gesHwCiUwcm+FVcQpA/zb8mACPaA4O8R51wXqOgNH22U1ZEmzfMetP
Yzm3+e7I2umtABxIjOcYDvwC5gDkEGW3Xu7G38SukSye83lQ95gDeEfMiUJjnxFN
hv6x+hNXs+g3F4BoaZx6oIG0QKrMRkX9ivRth97JP+BpHT5Y0wslPx0f3kZXHdOk
QbT23eyExJ0vze/cH8zMxyFa71Pp5t1uZbzx+KV3WF5r0MUf3aWzGYNd61w/cUNl
YnUnriGLce8r7b2292Mdjz11NcU/YBz2pYJqpt95RjJhKg5dgpmjlV2AW57eq0O4
R3njNclKye0r5b8Kimqyvp827+dtlTRrW7UV6L9e8er33ciqheG6XYAMfNip7fro
bnpUKs5rFv41qVp156BNHuJXUfPPHIOFULQc1eo3YYoB/EWMeMSd3eiBZ3QwgMwL
QyUiXvH6XzTUDHhpIu0B2R0Y6AqPK1e31l6B6awqB8WZSjbdvrRL0FjFdo9dyv+o
fRnpkuViRtVVvkp/BZNtUC4B0w5txvr6sUpBqp/SPxM9tYTrb2eXteuxBmzks3UI
91QcxFuJwcdx8Qk3Um+DdMUyM3e7UXRFLTtoxORSeHHePCykN6DTybgEJs9ZnTEU
JHoQFwIbdt5YpAqcWI226SkCAThzn5+V9K5MaLVR618lDpTUouo93NdieXVLJ+1P
nZu+IVywT4H6SubCwWnzoZwwz6+NxH5eyYlfLqtobUcWhsl0F0zRI/xbDBZQj+0+
n4qhFcBP2zPQ/rfZWbCAEHieMBW2W6XQMGDLvww5pFfHSkA0VeyxkwdijDLzBWY5
9lCmLN6IfTABMkRQY8vysqLYXmcD3bA5JeX15Tic7ZEZxqQ2pOeGNteVjnFWOvJC
n69LxfspmtCJwTq/+c2Zq/XQmFw5dmpGaSdYFIVO/gV+E4cmMcIGtQTaym/a4F1k
1uNN/o6Sc3JbmdqwbzU/LZTveJ5Hdmov2BHSkBJ/nZAhzvKeiUnRMfAhviJvz94w
ylFGf6IChyaSLXYxkfnUqqKuY50LpCrc+Rzn4fx9kPHcM5dkXgUneNR9PkuC0UP5
VMczcNimVgglD5+C9ujOsWs6H3WyCO3XLnBNiAyC+KmUjVSD3vR+/xQllnEQGyAZ
34THhmK18d8yn3muiT3NNvmMzlnU6XB4taxqC84OO17HEtiOprA3YXR1hFq8o8wC
0/AL5nPT9u3bbsLGQ2yiKKZE6b61pQNCLSrfWPig2g+zeRVw10DylZ1mHP+xNVVI
vbgWIDCvyYmIkO6EkgfjJgWalSe2TgRBmrL9lavhfU6u/DlJa3glyn8utfGq1Y7A
Q0uD1dPAmQwBH0xYMYDdfa7wG3UerbCKwwgvfY+GARR4Mnd9ojK21upoFELqCqjM
iO4D5N2Qq8/dvwCq5EJoQpRnsET3Zhi7EUvMiuHU53qp+GQrZTKhpf8uzo91zU6w
1pORpSaUF69oxeJlKrfDOdBh/8qF5q8fEyKmdELLBP86L3LMBl2NiehTFHg133dc
/kraffnZssWMp7vN/mI9YVqe47rI8bq24y3cbnHY6fbYQPY/Ba0zvuVuPOJgfNDs
eRIKRGLzOgu2iWZ5x6xNHysJe8D9SD8uSV1k9gZUHG8ZrsCh6WRE/o6LRx4g5p+L
gjCx5ClS32Ja1HMLfXYwHIUEY2GdwHNeO3yE3SC+jfSloLwmN/PzuuxVcQy6ru/j
EGeeLAxxg8UKyxtC2qU55UD2QftkZsmNMDrA8XV4qZ4nqG4t8/m8dS+jNWdRNDgD
jvuRcoX/bKgL2FFBJOn7reTlxZT1cV+kkekplgljdiKPVUchbn5YI6N1aExJaX2j
W+TKx5Ssf9Fm//O4OT9h7PONQAwoW8W04IohPKGNasP5T8WssS3bIxsXTlceyvpL
R0LXSt0LFd0XZKIkBNST2ugWcHMxt0ma4BhnD3byt33QYaAp7+7L2sFimWx5qOXZ
YUAdeC1X6JuQUcixsZQpJ+P+JHy7M8T/ycbeWfa9PDfbesNso/vmF1kbsl75kg9S
2oh+qomlEMjUD0l0jyPa7GZFybTg95SjZ2HGIdCxsXdHZlMDa12Cp/y34FkaWqUU
erchjVOkJisDIMbVdugVPh9mvFYqF1OIXMpaDONr80JcbC4G9tEeO4+bhueHR8nP
w0zTj3co2qP55v/eGIaV/eQqPAGB89amdl/j1zCNiq34CUjq2GxJNS3FYlt1Pabn
cX96Bm+xVsGUXPzKPigjLzMdF6LSlCVPjh6qZYA3aPL/NlWVRfXwYeQVy0jHIMXo
GYrKo8qVsuvfw1kMo7wDd1VNCbfa2ZoKQeGT0bPbvKvvy2I3IA/MxTq+PZT+Dtfe
Q1wGSuxAXSuNPzr5Dq1fDkd0o5YzbcdF34KbF5WskGL+6g3VkUBt+yeHEoGziYqi
/9hmrIUrVZP1ssxYe6kIMPq2i+auZwkNASiGT6FgXRu9R7BTHbxcwGOnzkZLsExf
2adYw05MS66l7OxH5XpldWHppH8ElMiwCoZZTfdpAWsfk5/LzwbPJyUFA3dSHo/A
xrrljuQeG9kt52T7UDI/0uyqNBa++rjaUAdEzPAGG5O1JaxDcZ5TNIRemwombP4F
huMBL9GdDecn4nNviMlLefCTQKHoPUZuy5bCcNI9aSOa2dsJtueBT+gVpTcovXZ0
z59Fx47r7fGWzCo8YX3Mqq58w0Gy+bm2vg4fBf9x3ynYXyJmitP8WMpnOa3D1QJ9
C+IPVoMKQWXbgESf/OpUxd6MJmbpiCpu/gh8ZDh4sSFrUefe63OhlvlepKugRWEu
f+8oBVSoiPZQPAzwU06+V66kvUcAFAeVHQtbdG2etEUnWTs53tOsNLnDADfCvn8R
Eix9qJeX3ik0C9AS3bctGXxYWQDa5lGFsVRN0IGsjXDA6P3rOqnfjJD8N626/azj
bPohnb6eeRgKCDBO7FGO0r+xCMcGJasVxuaBOB2+8wof9O/ghwivb/UnipP9L20Z
4eMeau1rBfDP2O0wR+IyxwseEtV7nyoG9yyFh2H6CUtqdhYgVIOR62PCXX+ZIBv1
944wWXjk7XkBW8eKKbWoeew0UnMuKIrgQ9oV3YB555EaGkzAZE62wqLS0xU5Int8
z1Vni80vzbrDpN06/2wnOWBPE69lC6Itwmh1krfEZrlo1PGQQrzcDrzRs/P+m2SO
AaSboMtuXN5jNCWXsThggtf18pVnp1WhEuDAQBTDGo8EZjY4W/KB23BmqcK2pEY5
bQgwi7X9Im+hUu5VT0V8jPMrKHkxFq96g1IeqfN9fYu0wPXFK/Mj2TNt7D/sYc1w
L52LxpQsZvxBbkyGKJr5GXklnK73BvYD31rq9mFot1oE5Eyj+ayg6rMrkhSA5+to
D9pTBoRvnQqWdGVaZdeK81v/7CG9V+3h2aAOcZ8L7lV4tImG4ZRLyg9dr8Qsq61z
W6yi24QxIihyTM66rnx6EOTlXD0JiAYUQmWjJ1CN/NLZt9J825GLna2v+Q/Jn+uo
toETeO5J2DFa/gldCYQflPDTcoma5zYJ/JHLA4dHqiUdzPoh4aomTzudb85/HXZZ
wSyFu7WP+UT/Uq93+e+lt9RIOL4FIgP3rXRY5x75wGOrp03rZBzyx5yoN+9/2zYl
n+wu3eZr3PAeGogyW6RLjVK0XgjidJJcCONQNtzvHd+JONzYvhLqXpF3G7rB1x0r
DBSsIblHLnpzGj86xu6WrdF/2yX94dw7B/s5Bdj3o6ouHTL35vm/I1GogKTq5J2a
vmhi6xxkECGtpq52uhY50lh7grqwg/MAj+uNm2TULkKUFy8vu7znhDU9mIPe4pg5
RCBKnIBOgaCCl4XnEdVqj6TWheIv3I3djYHwAleNWwRf9ARV/oyPR/j9C9700f5I
0l6ufeeO+H1bERe8X56RtM1nqLBJMjVhrAXRrkKN2T1FDVVgNvJLNMyREqlZDAPP
NWnAz6aIFwlR1E936DvNQ4aScwkUcnyKJFr360jkDt4n5V4aQALiGR0fLKzJZwEN
qh4nsXLEYVvCYyPnXsK3LM9utVsSHlTTRPg2LL7Jk3EIEwXqEsVxVvZZ/gdHn+Jx
C1kJjuO6SaCelf/ZvbEw0iuf24JLEVwVApfSbZPKNenBAFSVMRe3xl+Zh7mn9ODd
/pdikg5cbycYzQ2/ibHCZF92VkVvqKuNzamI8Jw9v41aF+yByYGvKat996sruyJs
xTfz3UG/qKGWD36S1VJPEstI+lvOA5+x/pTgj+U03+i60r2a3c7rCCU/uzV/bwRg
JiwGeKXivYfwK0JxetOExKixRD7cAcBEemrNCBAUkq4WsGmQKpCX7eoB4A/eD6Ee
SJititVQGFevvodo4ad9Rl5pL1YG7CCn/0qx/XuO/awFVrlKJb8ot3vczvYn7CC0
Dvc0HXzgjoRAmDlw6v7hp4xSMI23myaZKl/HMSH28SqYrTvyKDOjPPkQF06xpzuP
LO6PTGyC/HAVljg9KcGrt18whccetwTJoTsd9e6+V5Bu6OxgenZ3gHMHYLvLz8Vt
SKNBRh6KMhdoEAtF2pY7A3qjOIczZQR90Rq6RXkpfwIpvzYwylqvVwMPL1l0tzgP
R+BT2nwWBD5ChHpYgveMPPqa2tJhQ2q+i7hlbxHWfdRP5F1X4Fvl2G4ncIuDekNk
UqqwGgZ6hD5v4ATv4CL2+o6HyJd6VcBKuk6kuayTR31a7z6C50w4W9Q2ofWFjArS
w0vFNi41tXqFaqnI+6/HltatUTwQvZ7U/fdENLY8EFXbJW/Srms/faBb4iTA2uvC
DiC/U4mNSueFhu9g5pAFedMwdd2NI2UCoUoWSmFZnkd5aGQ+15nJIFiqNevxaYUK
jvgqNjO/7XyK/kPPYy9bWo1x8gySxY/whzWfK/J/h37Wt6xvX6d2/2hKtQcjcwfQ
Y4WzvVSZbUfILSA28/E8xrnSGAM8XXDaDVEFaAqLeErz4xf0JTQoWhGtXfNblZKB
4WsH/exclLJU4glNWc97G/cwTUyOdm2ilZ6y14hGWcmyU5f9kVU53qbYzuH/M8eq
NwEU9JjbR8bU5Bit73KJD14UbfJgAaX4qYhYo3sIygUkK24/X6kC0bP9vRB+nog9
uC7oMqr+Xxcyw6p/86pkyl+ZvaLaFLIe8zMDBgxLTwyGjLprI4PnTiP+3v3o3yi2
72FEaWKvNWC2I0XPNhSr40EL7X9MYcSF09gDIkJHjFu4BCoTy67qUA2E37D1SL2k
dSnud6GdnuNqwjyFiKSAfFORXRH+iYXTry4+/lIrhGXbSRPJM4iRKmTKwdudx7jk
lPViw47Fy1E85dw297pf896svhBiZ5N9eWoAV0Uircbylhn/uJkoyNvwAGoF4KVU
2GNQg+vN3YX8JlXzyLAAAg+TAVtfXtdZ8DdyX0JmwWDoU+mjeR/hjyHruCrCDC/5
73YS7CUcn5BBEA1dl7VWvKr/PcMNeN5U7szxxUCOcxew+FR1Ca66ZSQnyJR2H67K
BS82Z5TXjl8plxkNbb070qxW4/dVjsDp9WKOBOivpaUtkM7GkV2Fpjw/HM0JtzS/
RYr6d+HU4ZFDkfTEJ1PbX06LmE/77hDBsnqVrOrr0bbvwPwyB148kZjjtixfwDLt
hNjSXXrZukvJJUI/kxFYhESbcduG3kx+tivHX9usutTPgP+MjyZF4SGJUsKdYxge
OsXUt1xcJ0yY33LNLIFyn0DUF6ZAvVzMEWFsrzLEG+QIsfDA+pZSnOvt1GdSSTw+
MpY95c//RhyDtb10Z/0Rcy/7S1p1bkSEu6HEpDeCGEcPqmhptgxocLffzA7v0B18
aPfKefyA5MxqcuxvuN5mlOJ8OybvNRaX2RnuRHBWgvvXuwTOIhK/17rH3Nu4hpZB
7899skCT1q9ySL+PbWrZIAzri8Up64tIv5XJqIKlEC+ieDBNY3dEt7b9dLr5tvX+
BtA7rd0zSzfeAA4A2AMMljIycOZMs06yFUSRzlmUngnJKXiyQZeSMOPMot2feJaC
zrWIkKl4g/iHt2OjgQf6CJ2WQUG4t+hC3MsvBJLYpReq8JgzHp0/aahXjru9NngV
LqHuz/NDFlbJ22uTajQovqXQQ8hz7x4dVEhEuRL0TqDbGzgmdt0CmTK3lI5qEvFA
R6lZLNUzBJoI0YZWnIHfb+9Ihv5F1a+po9uY3ZMeqZ3zhFyCS5lYFJkrkKy2Az2g
JiCVS310Fad6hpV8hFQGYYZqEaK7yue6CfLhDGtv7TOKz5yWa1BZ2dokeTclDmmL
YB6tczuHidtQdxRwKKvO+gQVFzP8mSbhKveZrb3oeOuL++roQYs9tdHWUbQmgnLv
6aUZ/FgvFV5LIVLkskTRlBS+ySeG6txePl5ihAMqsToBAPGQCRI3YR0cV+Q0+14E
KMMt7uWk3of+Lg8Ndrb9RRwGW12/t4XfJFtm4GKXYBPZSC1yciuB4HC1dnQpnB6a
NQ5x17+eT099KHdLeRsk3P+Q6A4o17U94LrfdWoQmnB3ODKBKKbvwj3h9Rlc9izH
rjMg/Bytzm2oXZ3j6ueN82wrYI7TIICIvtU1kMXA+Y/gQtEyD7X+r5E13i/kwq25
hvQtvVSOa+SUTt4azAZBZxn4U7LaMCOXfIyVUduLmtYVCyyJD9R1gwdUGU1iZuVw
7RzkbIz8s4mLLKQfDnq353egudpVYxyQlZKEX+vCJ0T9/SQGvZ1Hu5cCJ1QtoOQB
0gebc8VAIRvdBQLNvbhvW8sK+JISDi75g0IFLsjI4STvsTzWsLFjuCBsiTGkYEir
oXFo4MHiL4gsNi2iJmwK6IP13HlspYCfBFmNITEw+RZTnvbiDOMddkFofXlDhwMq
NU2CrGhWcdhYjZZyvGp5xCdaKQ23qafNMwAifTp3DvLPC+9h7eXyAtrRdPeMohPP
JzFYDS2oNf0QqwYjGlC4PAAKp7xKPVeu3Ms3NgxQnJspb3aynisxQqLK2XdzQxMk
VF9fyMN9YOhSI+ng9EwOsuOWYYAs1U0gPdeRtl+XqFaj0YpRsNIX031qdzhzqvyi
nb5aBXS8/sQIg5rWeV1xlL+042Q3woQYij5IHZPOo0Q/NCE9mYPvO61VzagtPufV
x0L721T1QKhePcWZF36smK1MmmTXjNqFcTazXaBGsP1j6n5VWgbEU4YsvG761zuX
aR/62vdqDYFHsMzUrJuvuBSv4BzJzCf3SVeFZjkr4vzEc+ZgAtc7P6tSDlVzMQIA
1Sg1qr3Y2x24mPVEXazWsfMGLrUQHW0h1ksds6JGcljFe2O15Yis2c9Hy/zrkpyP
IVs44NOj8g4OonCOf+BBkArbOke7RznFnhsyvquD3RXQeD11n4/4PYTzC+2YPtoD
V5lI8XQjiWgyu6p15jInhS2qSsX0i6lJ8KyxQh8QkhZp0oc6m59+H9sWoJsmgA9B
MiRb2Z3bzNnUocyuHWMjEhzV6mdhI1Cwwr77eluligWYZqnX//2Eyft16H3T1jRZ
cEwJKBwcrJ0bSr+kOrzFXG2sm7XcFmFGpIbxEy0lC+P0SnmiQKDrgtLeJF2xa8UA
BwEFdZfn0YhFeT8cTMhBVNlQKka4MJZoZExHEKt72tzUfyyRXrFtH4PhE3dNZ6jY
2iyWsL4Pm72epPjscjpXxmymeRJTb0gkN2ExJN0qk1y/dQKsW5BVaNe2Hv5bVjx8
iHX5QS9b5URuLqgHyA1L+m1Wgf++K9esZmcT85IcWMf3qw9wnN2+DP8h9UoD+YpJ
4WyHuYSOw+xuia0OWWrotcZrsKFF/JpjWFOXWpXdkYI6k93reFuxy8nRmIsbnhaB
g5S+RfWbU/NsmyXHRC1O+NPJdsyqL0JnoDf4BlhdO48z4s2NnC4OKADhXY6Bzhk+
ZEFimsZqq9z0sNJBcv/mpj6Q6Y15GqHZdpzthNA1VQpFYduSXQ4Kz9k48dYKfSs/
gMAnHLRpo74kl+WwbC22VqbGgG8PkvakuJQRFENC+AoMs04fjjjs/C7kOrpfk/J9
gQULb/+j01CbtEgZRr4mAwsWS+6KDotQApoB5Rhk/E8GscZQBKCcjsRqeMoDTBp9
TcVpapyjo5GNqGE4eqpoO7hqXIOYwzA85bCoo/NR/zD3KWQNcKNCSxZHLGCueQL6
qqbCSCrTy8/g6k/4yn8y5PBL7H15jXHssjuC3MKliAx6BdiM7i+gDauPE3x5dac3
01MULoyGuVjEw+Zvmc11I/cZGha7iCUPXd0x/7eMrTFzr3fFJKfwNizk/SgcXihp
WbAvYSstwJOvp87s8BRpLckHzMbO6RAd9RRt6ckAVOu5NL7U8DFLfb/V7uyJIS74
ICRc8iyyyY6lVizsGEp1ctSK1GRANpwPTmhou/kant17qiomIBN8fLMbjvjphHHs
H5NfSo6e6YvQGSoDyU5riAtanKUDSa+3F3UI6e0h+6PS+uYeYcY1Nfj4PTvCwbTo
YEJq/YPHdnmtsy7VOhAxgwykmHQ6fCbDoZslMCrT7uLicdfshQCH45jKk0APab0Z
XMHRD8N1b20J4ld0p/Q4pQs9jDlzyL11hc0GD6BN/RB0K8cjYqX9sSElsi2L12uh
cJUUzJEjv2UUtYwGwVgGpy6EcgNoSvryAq29BK7G0nP8dFz0ZElPWkzP5vy4w3CT
5D5G4Ak7hPKbVR7sXrz/u08D3UD9Q+38+QOlOWNUgFY6cQLjJrMcnxTmtykSkFmS
QeZUbL7NZjD/d3Ko84PvpQdzvAhLT+I3cjuV6Tzhd4TbvoCT+IdHX/eTBok0O3WY
kjBuj5UpDXatQVtKUnSrQ175+GNyYVrwJ/Mki7UISt8c0Re8IaJq+3SjIR8Mwbvz
LZE0dDaT98tyCGqpUw354OtXJtIFSiFtmwgVqpYYgxhSkQ7gNgYrbCxYqrXxYj+0
EbtVrWu4jnNmITNFVZR6w0ZYP4rCxsywAHjPEYkUpWhxJ2fjYDGPjGW5eVCDGYOP
Bda8qNGtA9QaPFMr4Q5UntfB6U+qiXSobYyeH7rn6zd8WJMRhwel5OYifOUTu0+D
84UImcq2ICeZUaRaVLtKHp+8rvQUTp0+OQXb+WjqkM3c5c5n1ganUh/BSvGz1Wz8
2YwUNNh5JSsCeQDasbf3qSI9s2iKztV6d/S80xTg2HxJ37CWyKGlxmbXlh4k3mZf
RpztI7ti3tH5TSysl3IRcPyoTUG5bxepvPUpx+e7A138oMW8whvHFrlL0dU3R8Ml
BP6WzjB4zmd/3ts26mn84EMMmHXSOxXlWvuoVaUV7oY8ZfsZDEe3rqMxqMZoWkkQ
IZz9xU7w0Jdo8vTzq45VVBBth7cjCm6rtCiXapRqRTnIxnHmJkHlM4t+wI35YNtN
dOS4y3Xg3dAy5N4dfFMBLoSYD4kyO3mESFBmpYCwP227TBrQUSdgbfU1Zeh2+KD0
Dm77uSpkbNwdb01e8lrkoR4VmXSl7M4ZwoqyQxwTIia/gFCjtOrXbHEZR2pY2RnR
Acds+eg+jtiznaYrhXO90fVekmO/VK9bgE2FH5xkRfb5a+OkNe1Y4XLs5yC96w3S
fFxCapTEHfabLM8zDVu4Nr8tzmJERbledAK79+uDXvWof5gqfwZzN9I5PbVS3+g0
fZBEPBG6KRIFIj7IiKXFBONi/IipZKprow/gwg7W4wHoeDdtZq8++tfkpiqfb3uV
uRi6F+6ndJhOt8XYd18EAZKAQlPE6SlPnXcOpu7yptZE5Eaod0lGBminZ9v2kPdr
TygXmPyAJH++AstK07MHdorIal+lsrDvfqWBQdxSb8b+Op31YO5sZPtfytJFChVj
NJIWimbsDtoIwg6tujbvAQg0Z5rYXwLzAPeUplgqd1TBt/scmCLAnqrhv6lrKDC8
u+vzo9E/XoKdQPgf02pDy1UAJ5eFpZtQGLitRbTlxQBXmYpj6bpWDwT1+Kl6g1sw
bAaiW+H4cVj+kmqu7/gfLxyJEJys0dEucPrj1FOPQLRJtPH3XSwJcvFf1L3m0rov
8nwk1Hfqs7/7hhJ+cLKIepI59zD9JN6CIy0jNs/F1122dfov/tN/teQDGMmHRUtM
8ya1IlykiYr5h2LFr/1oY+y9uBxf0qQFBrtewGC5ZBYjLgcYYM9evm9mDjvqLlo3
siTVn3U8z3Gno7IorveGsvW5WgWCUBZOeTjelGy2HcbeIyZ3mI1NKZ7KBrzkwd0J
RscSywolxemApD0abuvcqC+K0r3cOsckUUJT1xiDq9PPfNTJx0PeScMdd2O3EJEI
e5tfU9X1nG3SBCl1Da4fJoXu33u2cD6cvK5o/uHNQzxoB8OSn6K8Uqsjo9QP+h1t
5K/qUduPzJOVHSjHE+WE9w7+7GmkqXFFxAi9ff+ZXh84xDJOc/fJW6XFK8GKdmsg
PqJl+zAwhyUIGCuiNUVWn/Kg9acvYBEpDMxqIpW2t9w9IVkl9pAbQPE2XioT5q0b
AcO8aw0Qe8pN9FJge2sFVfKcS4wreHAKnV4z8LCSiZY3At8ytD9zK9hNPkcZNLhj
rGR2KqT3qhO3QdhKNQIy3V0JtJuWk/u9jxoyEu5gMOtAg/5HmxZ2lM7m49bFqEsy
WliACk2ewwxrG37735hqa/1QXalHBhK1cvgJqrun6v1aA2WBAxhXHMVQ+74qusyQ
HiOTWyrHnObuADBl4Wm1qlCxtzJmsaef9uJgy7FHlokftNNpikMQqn6IQpl0bnGZ
49w+3caxZwu0rTrKOUVuMAVYN1A1kztpVLyrCTRh/RFhrPdcHqAYYpV4XEzqemsG
Phcq896gXZsojLoZkKIFQhEv2OaaIcSkn8hGoki+f62opsnILdKSMmCqWIJVpGTc
WLiMDrEUkOURv5CTXvDz/pJ/i7pW3aXjjappy3HbG/VNsCgYKR22wR4oTuynM6/E
AN3BBk6YhXJUgjkPhwv3OdSS3r2385XWZHKvwyFNKZ+H9ml7itztFqp4V8X+GHjq
aCjKAHf2+ZH+APF7p3qGn7/79LjhUn63aQKy2q1dB44M5AXroQ0i33Cj+a88F02/
ubQsBf+/v6vG8w9JbFSEkkqqng2FnHc4C+Dm6MuXUHRnCgZOj/ROLkt1xBABKKnt
2TTDnxBy9KC6lIFpSzk5/QVeJoxtj9kHrQihLDi2vnE10BhAiwj/oeG/eROLzAsK
az+EfJfOp0v/Wl4Ml98L920NAmgzkq/LAWBQZQsMeMhaMArCPXWCpsaWbhaHyuYg
vbLYvzqXLp4gkTESrYOrLHRRkZ4wIbcCn9l50nAch4g+wCsVSiq5OlEKAqwzAH0R
4aZ1wdoPTcqtg984XfcjhyshfFVW3GgN+zAc8TwkClXqZ80uQOswYnpEOfIHdsq6
JjCBvbf7gRs9lisTIrwPIDjRfhl9qw37Al/gjGCXaG4bCjHju5PbmIR+UhTKiv3S
Kn04wVCe03/6TTMupvZ/O3pwDP5zn9g7wvrpHxJy7nOqMnbE7UU3XpekEVUKfAWZ
pS2XWVFRiiMpNwzG/rF2OhGUwhuIBzC3d76V1oYz+QzUzPld9wuGkm+FFziiZB1W
8F6EO+pFhhQ7wxQVhHTYJc/AreO3txDGClArRAudbjkeQUwQ7Jy4I1FZirPlFb6L
isIF+3xSls6E6f7zK/XY/6JYqzW3ZRZuBWa58K8/IXcEurwxbDbqSSKzxRuk4nT/
a6kkYFMOuMpDCzYdjNAV6vEvR7NAKQMyDAX7F9Ft2eF6Q8MNKAPnW9R/sy1qVbNw
WoCaqDq0eoDnJTAtdVVQoWn7kPQinRYlELACFSJoSAc/RSKq/v4nTf9IhZcW/qtc
ppuJmiW70G5bfNwY3XqmxajxA/zKOjOZhvo2kVU1QDxCegEuSt45/RFOADNZxGgA
eE6XauUFxw/6Te4BirzuIGG1CV7BS0hX0g3maUwi+JaHtM4erYlu06W9SuZGNrrp
IgVmHE8PYBayqCO6hSIpdc5g7HGThEpA5KqGJz/LBA3VX/I6qX6QM1FR/HCV3oaP
U/y3JvwnSDx8Ct2NPtYms0ZKFkW/VEODk7565U+/7ORoBtSz/NDUmrfoD9a+/HdB
ozLNOOirtDnaR3cuzIHF3Mg+CgGkQQ3INhWSVOuY/WSVtVZaJm7OOMPAqo8YsGRB
zUWURA6LgAGqslpz6JedOGA5c+Dp6wbpR76rhAY+WuxXDoVrY9l0v+e4+EYHX7Sn
eOy3BSaQKezuHzxxEw9jao/blShqCxuFDhmXmaCNSK4A5+XYgHgDZtNnC59ekrw6
QLUJBEqPYDVGGhO8ESDelR6KW2VNi2fL6iys7aIMwfDooVom9oTMT8JiJv+q8kin
F1hFxf/pITa5hNUbeJ65mA6QRg7cRJjd7ilAFJcR4yMlZK3KvQzqvbKkFWwygwsS
Ivjm/cjLCq/kY33UdWt78fzjonOvdvZ9adKFQel69xv0RRcfYWwoPDxzmDHXVQ5q
gdR3Zb7r5TdpiySoi54ZUmXub4LgA+TWUb5+UNsxMSyI8fr0x9JcYdlL8PJBAU2P
pHeg38xtFKklPBQbTs29K/JvmMY4OSJ8MEDXn4fOcsHTj2nvlexPn8MgPbN1e05c
GOOf4gvZREGkdx7J3uS1biV7xNA+gEA6eCtJ+Qddjt0iRxNTsip8pU3CBbYbzLCy
KW02Jns5uMiiWZ1ecwaZvonx1xrwFXeJS7t/60ZDA1SPQGt0+cjJZizzJPsvMCDr
cT1G7qBdXfzVFY6oXLd6a2rBLu0DQ64AYruTIAd3k4kpcgHq3T+P1mAlnrt4puPN
3rRMt2kNzD5CoFWqQhY+6AodTOBf93WznK8+LHSh6yf6Ec2606hsOAXA9f/+mYLO
9voRajHGJMNue3s2zZPJyhKssGSMXPKSwpuYUpT86YRQntPo3ZIrc2ckZybFOMwC
RHfwnWQyDv+wds8MZFMpL9lP1iAB0xAPOLW/7m4BqpFJB65TIY8PsTebhlB6xz5L
P5jQo1c9KV1j3JH0VdPWOQcVl0a8W2irnq8GoVh00hW90g1cWvgPfSM1dxEAJjj1
rCpbo6CQKQ/FzwmM/IO3J3KVXI7wMEpogC1+dCqf08+O1a8ZXyswqAY5NWW6eS9A
TtQFV54bIa6fbrl7OgFZ4HvUn1Vc4kakc69PJvYxS3KnQO7vv9cRKROGRe7xKfGl
xP8ugX5x4Bs9LVn5Lj1a2U+bp4vLeah2yn+Szba09oe765LZFee2xg3QX1xsquCJ
PDhgmthoXZwWHQU81fgS7gEKGy0bwlAgGWWr97ydF4sVj2PsLlraDfbS1sHv8CYP
nrfBw9VejgRrUzL+llvdXRegPFnLa4LuXzJy0Z2mlvRGotUGPAhIlCv/M22/TS+I
fVXryOth+Bg/9eYW9541eBNpQzwXXEushY8knh7E23F0DaOof7Zw6zziiE4j8de/
u/AbEO6RqkB1VdayhwfIlZBQLUWZwfQawRVW51vvbutgSrDOvzNw6DKwz7WnKytg
H0c7W3W5RW8Sw6Cjrd26uX55WZNq3c2/exdX3d/wvsJT0EFp1Q/RyWl5t2jkVKp4
+BIhrKC7cKKYUyoEgJER7Vz2m17LJ6z3FDdoz/zziYAuEGS45hpB+W4s2tQuKE2K
MnldpmGr+V01/t7yQJ9kWXGXesmzDSVDm6slHqmySj9fwZ9xIFCI/McbGB88+11L
EXeDU8A0D6G3+X8d00nQFTy1DTjv+XOFC+niy55fTth/QFFGN1Id8Uuf/jQgcan7
LRL4lNA/Ut1CoHdlu7EkGjzzZrjxhKgexxSvm2RImLDW3bxSrVBEl3/0/YtV9dCi
6PA0mv0zF2/KBhZYMisqLCxkYgOsAZM3aFsXIZ9mVy2jQ71ASg3Y+DhydJMBejMg
Ug/Vpb59YUM01zCfwEXP6kOBdJ4O+8DbwwogBU0CqNvOfzZlijBgsI4rtz0+WIb/
SyQX3GaZwS3zpASxoqLc9leoMMRX3QnVgAyj9NN3PIeJwety3O9VaM/LM9HRCd7e
CubZOTQHeApFQ2eAZlP9jnQL0OOvE1Ka2ESst715qFtQXTZr1JMnsJXIcdbto+H/
3klq/8qBuArXeR9TJXgPsDdATVZ3lUUL+qzSbmb4wMFhQ1lRv9wndE82ao+fM9KM
xqPw0nIDMiiEepXSpk0DEClT68eV6odZNFhtkzIyPI0qtPzlpnAtiCGHiRzave7S
Ow55nTNsuj4WMFLkj1qwrmRLGH2NYrC8UL8kKntNyTYi/2mxWXZcL761zf0t7urp
jWMfGm4OLhZ7FFyRynb79ikvL0tyeLtNBhW4ER5k7rT93BDu2hCm0IN/BRH4hOBR
DaLxL+zBvxN3cukIklWaTw10AQF2F9RB13D7plBbP4AA6SnblAhwq18iep+5jE9U
B9iQ7x7Pbd3OE1P1SsrLkC9rGjFoHIx0x9bQunCeXIhKCyN7HpkCky3msSK6QQFi
yNDh5qbiVsmQwB+1r1Nu+L+pwLDOIeLvc23FzLO9c3diraIs2zX9MOJADNRZRn0o
elB8dpbywqPVX+9GOmSCpLhwtmnOAJQ/cITJv418+VWvI4Jp3hmAYd9AYN2WlS3/
RowyyTsQ3u77WQKASrKv30UXdwKNcidLyuoU0wpcNBBHPFu/nHZ68UPEjm2HV0X6
0B2cGaYFrrM7lwOfl3nySULustWTAD2/8XmveLh+39lcmmuWulFFGoIZ+gJErtE+
k+fnGbSfbRG3LF6LutCdZmRDGNfpCyyZv9q8QDskkhaDHhUBgwO1r5611ftSIW1K
sPD8AEjRrFsUukIYJR4IrvHRlTpefnja3Tc7aFvt+lGaDPrgQNPd4UBlN7clpi0I
ytkfLAQzm1UYfcSKVYvVj2nU2h/xgScNf0bTU9a++ZfIul8Wa6dxOQXVMoTMVrj8
1tpsJE7XzzRWPfJTbteZByzHBezVuxY1TWgAs1JWa0CX9SgbsgV6pvpfv2bzw1V8
LGS9zpLpPLgsDgn6yNgjLWoe+YkDw6QmvTxQbTdxkQiA/BJTGPlFGYXwUqrfp6Xd
ZPjBdXHPamERDk2GhyZOlw8dtM+LZnNfhvdCZ3v1yROWzd7V7IYFhtl+sejCvuJJ
biWUiuiGUZ4qbXI9rebi2BB7kQivk/ryc5x5/XTkfmQ3B+thk5pHC327G/5QJwp5
0pBc4BTQY+nfAL4ccGCEm1UVKf600lEh+ZR2D0NepIMNWJFGr2XW2c4/1TeIg3eN
wXq2n/P8KnbmO8+Q/ekE9mVCNW0fRGNPYA4BDUHxGhLRoDONNOBK0GkGwvrA3uxZ
9Fao3ESmm7v8DEGEPQSGH5GRqr066GKnG8y/GO8o4KBmfcPIexfAmygG1cfwooq0
3peKmnZ7UWFGd6ENbr7kbFVYZOv64uehKQHWRiuniqIPlYwcuxeNldizHk1XHLZm
/YmbW5Elqnk1n88kgJszzztHXHxxNI2ELGmcsETrHkaHKIWp7E7/mr1RcePx3sJr
3bJKhdPzxKdsrHk374H3e4v9fp0vUnCidtrknSYA466qUnqow10LHcpPV8KCY6gV
cSWZcIpH9ryTgjsR3C8BMKTxRgRh0+5XAOo3Z1aXfaixDT0w7yxvgZWMH2lpSoYC
gIus74LpbwqVYAHU+j8LwNDDUeJ9/gd3N1YY1F1Vwloab38OIPJh5J5aEqrBTGqz
e7BxUajrOvaeieBpnQ1WslbjO3UTug1r2ACLiYaZ8ugGJGHld5nsvEPBmUPkYIBk
XmAKf+BOhChyVFZmAIMEXiLQpGP0HoFfC2KmcOXjW1uLHJOkOtHzP5jo7E5YpbBJ
TE/QLgabPHeSOdfZAek0/tQcC8OLOnNfwRyYpuvBnXjGW/pxHEIgIRf7HMXYUIzE
qWbviiJyA7sQGW8rItkmMykI2KOjKjNvVb8pd7Ca0UJHtmSSZH2sjeY2ml1EIrgR
qlO0Pf09Be+7YKFLCy538adQTE6tMtyLhxog1MozgCPjCfftOlztgyw6+jXka7bS
Pm2hfgN4pYZEv4bBnrooP+9+Z6jTQxgCroegtMj2K39+U9FpUrgvsOCTDQiWr/Gq
MhF8L0GqftH1LeOa3r9HaisxgqcvMn5HpjTyYlBqcPB2CwJDm49+iC1YuNlpqGNu
CfMjrRHbxtqpDHmn0t5gfxrQTvNNlhfk+A/pR4ml2JhcIP6qugv6zCI4BXet3KSi
6JPcF6MtoJVQSNAk0e9WVl3cyIpbYe6GRkl5pQxo6cv2AI6oEqlY55dmx+CjWxr3
T+cPi6sFJ9OpmlZrK+vDhY6eRM/5RGuFLc8mPR7QLmSd9cKRa+knEaRS7enc7BX0
1se8WgcZ5pzRwTN1if5ZEijZqr6lFRUrPEYzZ9oNpFDvWLSeodR8XF3z1+rvokf7
p8Ig8s7SNv7ruEcWQ6Yx3ydG5v5IKCKc0hUxTCunYOgP57l9RpwwuirPFHBAiJAA
Xb0R30+hU5Zo+UnosbPzJxhOjSPA42SHxFD09EqcQJwBAqkvHGUQCLtR8nRXEdKr
SkIHObfSp2Tg55lnSYH41AgN6HPxM9RFNpxs0nOf6Pc3xf5alN96Xu/kfhlW3NZR
PIVm04myA2cyoCnJxoKgwtl1aeT2i3CdKTtwr92PpwoCk9kPOTblt35rMb3RJ0RU
2N5Q0nV+JeQQZh9nhvVbL21RQo7eSCDFw9Mqamnrh8rnn+Lw3MV2EfrBrqMsbTSt
Dn8EQbJMXmmXkS4fULwkvoobcdFc+uVio0swzcdteYmO9az3mG8YqlPGWex3IyzD
KdS7ZoCb+kcvy1F9RxVwBHAV8gNwvwFhEC0/kefgd3V+3Bw6EwnyXUxNTq4+aFHW
u9dQIhhVccKcX6zJw++QWPjFDz+0x5lCny6kGC0UuBLmUfzMYy3pfT8sHIGIffif
sMQa9j1APL4s3AqRxrgyVuckWVsbyaF3yaKTFDBpS+3xUYFDx4b/yExPatzKmu6e
wdWku0iDmstuLfsyk7t+QBbIr4EE1fU/N+iXF/ZAIE6oLkiMtlJqlidQZtHPDTq4
XAnXm9GFsUodr71UIO+pnI571esIE/JpsreIX2QW8grt9cSuQlSyDIi9g/o34rdi
5rD6UbxGar8SB+7HqGn7oyS6niuFUYk4pq+7lYGIbfvMoLpSEDhuWRSB7+O2SM69
IjrBBUsYN4A3ZSTjA1obFnYpNJBswShGcEslY+3npC0jq4FGaM6tfTtZSGwm2FRn
FnJhk9dQTF3uWn0GmPGdeTjqtcIcjoC9Lz6A3z5QKgE5wI+urscu0eB/zT6sXBb6
PCwT+3qg5N6ogzmZg9W6ql0lMOszQhtuHAUbN4lS/IPlI+dP5wD9kyNkKY/Blr2O
+n7lAk7VOuv1zAhMBoGFCBbQUa3YqZa1yHdkE9E410E+a6i+azbZrgGs/snQYQ1e
IjAN5tUZKKqiKlizis9lhD5qlq/qZa3b3HJyF9llFXYx4v5f+ZhAj89QLNIoqYfa
FWC/6Dmm9xGUYiwx3VtB8c+C7bc3Xq/ldrFYcduy36lJBubGPXt1Y/pg/xBoA56H
UznO4E2gv1aY9AMAH36/x/UwCMWA20Sdek8uPVer99mM6N770Alw34RsQ3Qqq6rP
slMmkxAA9i6v1cNeVmLj3ORaxSny15s71LqGC2oYNB44mJQO5TGGG7bJl5A69JuU
Exs6Q/TSAW5yepU6uT5yZ+hAChMs0cSvY6bEJrRoHbmtMkIEZlqj3SY2+NiCkBst
pOAv8RNbYE2+pzD7XbnVlGCIZwaurmxFz7EEeSnEo1OAgyNMM7CbRi5I99Tj8bXY
0CgeBj9hKREHlxEFnFwBQDbuuvkV16W0WyTmepBK17i+4hIDEdMejmMT1oLiDZMU
35H7P5OOpDOK81rt+eJSMJvYr24Yu8s5ZTuNmopiN7WlDWN49LWW5FXuOn/lcscM
Q0cZVPtmax+GZDHlkOthjGmUCQ5C0H6G7wx5nD+jvH3BQuK1k95yhm9A/oIwNd6p
We9PgRdNptGfIZVf8PrHFHw5OHYiBK5qvjFlKAIVUi95Kup4ZoIL9GmDVY25w65a
/sD9fJTqkLGzIH8wC5anhiquHjX7+2SjwFpB7M2lwpIWaxqbnrIaBbeMcSuC+t01
dwtNvAI8W+6y+ZdYZQrVYYZBSEA5maagGK9VJe5Ks8k9mp59Li721YITRz8l1RVZ
Qa0wWI9SwdAcNvLlTmLd0i0f6EPouzCZj/DsoG2tsP9q8pd8ev87Op5tQ6hGZTgS
jbu793p9Wk21F2Up+Fjd/LplrQWk6kbFur7WN0nEJz3TrPt/HGfwyyJC0rETw3Qw
2gDtirZhGR63DnKAZyIMWG6qfYesJxk+wHbYB+o+DAfPPm7BXtAoc5jmgmFSr4H0
TXxWqdSAQ0yiE3v6uX+iDjxCCpyJx/+G0lbJojhNTKX2cAQ/lEfoL9U4HFwYg43U
Mz4LwGYEczCZ0Ny+2OLmq1OKR0rR9IugcsTqUU1QNGWiXa80K+HV2dBBdlAuta5Y
XOuXBM1/DyNutWHwsnfgTVQ/gJhW4lKs9v8nuNoeNzYsiFgiyatpetZIkH+GbSF9
ZazFNrmbGSSOHGFeCBOhfHN3t3Wq5IRBhdCdhtFcqf3uub2cOfr4dT+NiDf0aTJW
o7ORYv7bjQ11kLrLJfaxeQihQxWl0Hcb4PSXzVDuI9CmixemD0gKXeeOA5b/i00I
cwAyJBPKS9JTLKhagrEC0PYcgK0UvTcyYvKa+TJhF5uXjzOATzdHnwsECmSe9yFm
vH7kfXtRmvnoQzlhHMSQxRZkmpJq4u8ppMO1+pOFu9vYXbWUmW8itA/wtslMrcca
F8hKRZDExOoWfefBQ3duRBE4sFKuXIkWSt1PMxlyHzzwx8/JQSQuSAN6YNZxYuvP
f4W/niQxpx8TkwIGv3JvfR4Nyzvtpzsb++KY8+w/wDMRdhbLRuHScIXLdwT2ntpU
CvdPcfo/L8IjEERbxsitH7NoM0127fQAD1cFTfHs8n9DcP6WuioEa8ytDK6uEfCZ
MylE2PFxTQodfvwIQ2YQ6j+iGyKC5fdNUFS5ido46SQvkMEB6mykB8CtvycaEHkl
f0Nacge54GNBu8EKmFFgQYAvUBifxhDQBWr24Z1U0JIgmDXK6ChYRd5zsKl3uv9p
VBMjtTKGV2ey53hREkEL6kcIq3uquhQkyZ0+Ku23OFW09hNCix4rR4aLV1WAVzBU
H4o++SCK914n3B1yChzO5BdtwOgsSOgWprGdM+sinwNJu/Ng6Dl1YZN87TtJYBu6
J3ikeUVKf7sTvDsV6iPNemVwQ0w+OZGulGDVBx5TMhVCHf0KqEmQ54fgIHYZ4Tot
woXQ/X+WKN/wWggyqFIwoHU9uslsQx/U30UivLI02vV3pGdyvEkDoKg6gu6IYOuh
9XTJQ7h+Nx8Ny4hwOOC/ezDBKYn7c+TfvyRtzDMIf6XbrTubpuMrnL4weaq7Iqly
O5jmezNW0CU/gMTtjdIe40nCFRDOFg+gAeLkj7VxPu50/5ByXzmFsYwnscUxZekL
KzjqqMbko+2UzkwpeO3FfS1XiuvtFaPkvVS3f2TGFE9MQ7jeb5pbXeeOMfDpb4p+
G6y7Gt3/I+RuOgtiFLN00hdvxdjovuAYJe8aFdYhwZVfhR0lFr8gyDKuRmgzHmD/
dAgyCtaJjRpD4tSEzR15KAQidDL6xUA7xkUS6HAJXIMtxRsYvaL1ds2UR66WQmQW
D+k4qdzcWBVW1p34wV2l7aD8O69A++RNAuOBwks+h4SSx3e2HpjwlkvY4ZvgqlXx
vV5UT6i+Z/qMI8k5mr6uejN1p/rSZaiPxCReImtDr1y6GyWZ4NIVe6LQSEXsXMRG
VsOzgg4o8MzOWzKLl+iAMfeCfcU9CubKVHWOKlv84gXKmo5UXenxe+k22GqcyYL2
kuPg/8E2q72PJJRpo3kfxluOqvo44CCsxiRluaEGgVCNoh0CE8EgXPjuY54WFUYh
dtfhv+r4R/MYIA+GgtOROLp0dnelH9MKV5hbg3hspSesFzrQIxYeFytxZn88i8Kj
hKRJuD9TFXUMpJP/iqax9IeVydO9OVw+w5LdxPsjBerVKLvIHIR2207eJCT961W7
ta+ztKwdSe5bspuy6//VU2mTx6uAWCigYikoMfK2Bbh0JmzopwMDA51cTj0paVIV
kNUBJcrETsaqXxunxNEbDLrljQgegk1J6nHMD87jIO03R0os9ja0U3mOuhHKr7ag
fDEbwdujp328foZnbtwOdqkaM1GIi54vFAgxY+UyqQuci9n3Wyr27KnVO3LCVaGW
gHx7gdGA6XArS5agwGS5pBvcG8CzyyV/PxNkSTH2aHcO16FfjriFiBIh243BCMQZ
msROYz4jJF7suQhTfO7XXuhomihXMoS3EufMfIMJlfsKTkKAsaxCe+1ZgRGGH1EQ
n8VjDmLrp6y3M5fX7RAfrTdsUubSs7ZiHDmYKBr9uwnOYz4PUm3MZ6le+nBY2bvP
ptLN+qbkmL+/nliMEYW7WywzSQB9bGdJlXOMOjykqfiThURioxrejObjOTiICOei
HuA6s8JFmA0/yudw1pkl6sNpVHIccTXcPhjZitWGt0QZfhksWMgPEcXReQIuUmvM
7zcRRZ5vHW6wBtsI2KOpZNous+HpX3OkO78EKtecG8OT1+mJKdjxqIYLHi4GxRdP
VYVI6Y12wEP2CRr35h7HmNIlCokD9g/gzw3IvzVb9cbP1Zvgc9hEdiODeEWlLoJN
BvJljKP2Yjz4ZilsJZQ59WNJq9yqIY1+n/adEwYMJnAJ/9gc6UxYZjNy5aCsFXy6
y5b5m/3hjsUjSBpXNJTnhHRJS8fW5tCGHBS6Cua3907NAqC7fkEi5jkF6LUXb1mD
4CeJPPzBBlQIThZCfL9/Sf/bi1ofFRYXgpo9hms7fqrZH++Q9zfMkOxV56Poexv+
cP9GO1eHiNN7lR408FlmKzaTtBZYOtAjq0sMB1qSBw9JWtCaR7LKk/AvpaWXBxSB
MJum3F3lHG6zzv3bAs8y79hBxN0aePPO5BVMlwrECOUPjSMlcMrzbp78LAzvOwxs
b+sWC1ivhpe7/7LqIo5YZSePZmZC2bYJ7WvMXVreF+eDAxA2GumXVpvmT1WY3JJi
E3pb978kXhnJS3MsP2/tEpWrVywta6RzBiAuFSO3K/hICKpMqtRMxXOHovnkK1ra
yJZCRtorg8WnD68pKb/ej+2GTdhzNymBx/UQKJWpLwzG8VRozAacV4U2ig+jXdIo
jY1eXlA+YItFLxVZ/B1MkeVZZVTQW9nFCkvU3C3ne/XOmhxJnHMOCAXTuOeaXW7R
OlcUZsyZ+F7MvJjbBFRkN4ZQJiYl95vpFt230NE5TL65REzWobNV6DDcq04+Nmy4
GiDS4GG2LpNd+8fQqGmVV1ULa646fP+2dCcmLpSY/EWBW8dfHA3X6dJu1ea0lWiT
Rm1cryyaKfirVI1wLFYQtiJq3r9UJMJr3wq4D6uQHRHP6V8MxicN2S775tCTPYQU
eA95ZLu7c14MYcWdi3e6/LSBpRVbopaT0XY7sebIbu4j2piVXBypoo+W4t3i8qzZ
/1Iy1Zg9ObCSxh4aCxytYWdUc+UAgqNk+iwLJPOier80lsRjS1eIjoY97qDL13qr
Vnj3ml58lhunoDXdCmWcFBSER+ouA/dysd5olZRiapxt2Sf4nVuVlkUVu65C7ZQu
xUFrmhRnhFoHx4pYMimrxrgEyV/T/zWz4af/gNQ9fhosdrINlQWbk32WqLs82toW
1ozay7jFAnwhJ/eM5nod0Wutk2s/p7UzkDWRU0fkYD9mzLQMABF17dpVghX36u/o
bgLKGqhI+Ni46KzqRdJkUG0CDcjsPQ+nCDMcqRCsRoHuoxidVKhRLpdZBs+xfDg+
6vtmV9EiiqIlVFjR8Q9fX5lA+U2tI3BoK7zpxvTMuBQE8/t7QMwJAVGSBtxTfRAz
+sKWGsrrmqNAcd3ddpKZz6sbSncbi1fW3L1VZelxBpIDkKL26bj9nkNYLzs6yJnj
KAsL1h5zQrwumknRTsL9IlWj8l2Lzn71zyfxJz77Bi791+6/YeBBHmE+Ic1OkHLb
JzzXcDsk0SfVpqgRwR4kCHDuLeOT0yXVaO314aHBXt+fCrE425nM6FyL1CSgKP4x
Cq5nqM4c9H+3nPe9G69Oor4pZ4g9IiZl+ONG0CAb3IYCw/dCezLUIAH3oT9QR+cc
CRxPVsEZTGCERHcNxl4i7zncMC9++J3O346/K7+z5wFhkSsSXliXo8X4dcqAbiFm
u6YRvtEsStzqYohEDYH/O2pmF9/JT8czPh6SbOkqhlXgf2e+KYkKPLtBIFZOHu50
0O6xu+cOjxucXQi/TAKoPRGRvewtQSzHI6RNpPrv/6yhJy2U9c+nZz6h/tHbRXw4
NJFBLoCfgemOvByMYyeisGXMeYNBnwQGEnyZF8atUlxmPhzurPWhRZxR0bGAtLVw
5e1rl22uGEEorhR2Jl6YezYGHldi/XfEwut6fTHthCBZLSg9xqKTW39GXEkMCyNO
E2e8LJe0+nbNdHA0WE6ur3BnDnVcJbd8azCy1Tw3sCYEniAk3ehY1IpGwpeDkMlJ
D85Yr6jetK2HZPVabTps0Xc4ABI5DqW10cRk9CJ22YSdsP0G8+O/bhhdr5+9Oz4O
4BfREtKxUZrPGD7VpHSlgvPvQtZ+vUOqy+Lp7vqI60wYeAdI/AF9v49DtoiMZVl5
BWMqKZePLtr9NkGKdJYIJlXe1Z0f8LsD8EhLFTQ+gKN13aGmmxTaNpeytxxWdd+d
j+OsAnWpVJugW1fGa36TMsE8qYsybRc4SFyykOPfH+VcyMDCr4IV15RKY0nYUNwz
AeOg1AgWSRVhwLnXkiCr2fgyDerLU/zwL2qfcQy+LutyjamHddXV5Sh/RPqfTl64
66k4Ik3tAcq9JdyFi4Fuoer+VI0DU9FUNJKhJIXusDGr72KCzOM1jF/RCDXMkGOr
ct/0qQ0UJUXH1aOmVVEey0czTQL+3axuc1vQAGGhxzUTLB30ByLWZ1p3+xvhU1q0
EOH7HwOquTYCx8qpLAtALIAL3qHjQULzD4FlgV4GC776V1bwLYyurYJbyWYlh8BQ
Nc+l4USvO483hG75ijnAKc3wivZKbU/bcAIkXNVaZuIf6LZXGJ5s9L9480WduQfT
4T8wu2sR0UfH8DRReMEIM8Ufsc1MJEn2sRN4I8xiNiVlevvXXEFu50exxsCxjzLW
PrpT/+gYTKD0s+c3KGlnHVRU58580UqAYMozuQHyUY048+Wekizhe00z895bHfaS
iL27toix1cQG0/N9rWcH8EMYjtASknJrv/wjLb5JZyWpNFR/QL4IA6IRxdo/+lka
q4zd3dlZuQy3H1e1idYlH+OBNZbgY8rqh49a7HkNOpcn9fx7VDMcwvSyYR5yb7IN
HqkK9B4BGKff3engcpS9xepH7Auy4hG83AsvhJgA8arlJ4bV0DhCeEP4SDQAiUdb
cZ+3P0bbpxGkOJbQQgsuxmOhSGJs15fRxKQ0bVGC0fYIYQrPVN5JZQI+tZB1gcZD
dhpZ3bmSgY8fMxGR+k+YJ+kFIlgpKaE1Pe96RVSGzRzLELZVwkHRiqL0yGlfaeY/
ui84joxLyBXD3h85JRqtCw2WFSGsjb4/rcH0YHKh+K93I9eYiBvja2JEzTp5Ihdq
wenGKuDADhdIBbp98z/GrBNpYRH05op7+0Rjaa6Vv7xeBPe1NDrvjLYNIdBR2BLU
Mb+rpTlgsCp+MSietSp6dw0kYpt8jkoQwHM4mJS6nBKPvWBt+x5xVVLr4Z73Jwak
D1Z4zTja79mr9uKwMdsIoIInXzX4turwDxdSc//CXwklih/chERdJcG216F09W70
JG5heTkVbQ3LqebQcRxgt2VRg4WSJzFdJOvFbPqLgVDP778bQI1PkPS9dXmHCPkc
KAegIG5EXh5qYI0AgBwrW/fK+Ywe93qCZ42KG+gjrcJ1vuNFpsOpr5+kFExLbJZK
ceAIpZhb3JftceDNKCE9ehc4jtnjo3xvORKm0tStHNv117hIUHTT6MEDwOknmpzs
OFp7q+4Bf9PQNnQTJr5T/zqGeKD7IY8JaH0SQo7cYedghYAOfsUNZyJxlKzCXzZS
aMvObfIxOiNX81Ihx/DvGuNtbmYORX0fX2r6kQUW7iZNYesbXFj3OBHfo81WvsxV
npXKlIdbUWEnhxMCVKa4QF3yZinyALisogkupRL6bV0AxuMX3o6V5Yhj4kG6+ifi
0ZE2NF+Fu7MTC4eDFMr0paFRBY1K5waWAOVyuWVV1rFaqgCAp5A9qUb7Jl5u8uSK
TiVR6bn8LQGLn70Zs5HsEH0xWyGfFK1fjrjv5CfV+KDEIzU/+od1EL36OOr7n+Bi
WrvVY9agnAR5DHskVpirns+TyLzLKfH69HOaFcIxgvvKyxKMX5SpiLXYcz2l3kY/
WrzBUQEBmdv4AzJXn2zD0kMBWhG/rpybDtKLUPG7wFvB3iRzVZEokBkeEErlt9Kx
tXOkvQQf4yC3cpgwPM7uOBDzs84Q8w+Qg85QsdYLXi9E4airfnKpyV4ZoXDPjaSf
KMnn7ziXSbOrXsdiz64t4ReUhsOOybGavtdJluQxfQL3fNj7IclSomEH/nypwTgi
73Sg+U5Mb5SM/lR4jwsCCgjELomtkTVmBcKqwG5Xv1j4numYuwPf2V+ynZpSWjvL
W+Om8GeySeXk1t4vamc09MBZFPQG/UG2mnaYtTRgLxIo6VVXhFL3g6mftYddkrzN
XVHGZhl8YzQulyR9g9OXzcvZulTB5pDZ4PgwQxhHc7rz9/lHBpdY8mnfNDGqrWKI
uUPw4dyvwkX7zv++tFAfq7p+z4Xwt7vJF93dmuw+N1yixC36MRisXEDPQlNik4NP
UML4zFLqvLkSwXVBBYjwXYVCbrayvK0xvtQ30o7KY+A4jwmMyHU4fIsnW+64PGIW
hHXbjLAswncRercoIvQ7TnHcCb1IGZmMiR66Nv9XIe+6n4nwsc7scFfz8y+VixpW
6CtNzSLHwtDv0NWH7/OR7G6RkizCpyb+5Dp79Jy3Cl147yP0XgEXFLu+yUFDYpvw
U2+Zfa/RbgdvkrxVtjuPSrP29OGjSXGRi+MtbJdL4W60R6FEcnxpo4nqUJzKz9Y5
ZqDDhV12vXmkThJHzC77HAsHIOJnG125QcFwS1g+PNfXZ8JLRyCGEqkFRTVJqHTQ
9mE9CFFECDjoMfYYhaRKnxP2d10QXHJ4wck3rJPDXRzpgWO8mzUdIopo4uHKWqHV
qibdCg+bVwKlYmBHBKl86A6MgusWOklG07vDh6yl9hj7SiuwOU6jE2NgqYBw3lmj
KsYS3KMCfLoBs5MVpgMSkrDnT76NL6ZRzSo+ANM8N6n6kDAZtmFTHeg5KGK1y+/n
1moPJpTCR01VxzUVpK6UlrhUQYea9TFRGAMRJdDo74vQyNKI+A9oqcrMgVxXjsXR
cez5BkkYuDLeTvH55kVb6FdPWuHGZQF3fweI1+0xpGO6KljH1fjFUArVVMcjt6Yq
MmV7/+WsjD+GuaDlwpZ6VDmcM/ERO0rN3BeaddO+aGNoHDW86WYAPQ25v3vlmxvS
13xSNOtyyUyYVBlqiA4IfqWk5QR9rFBY4nXqp3Ws5zeHztcsUc7g8uAgiKFEQToJ
SoLGZDpaoC3gM70OyVw67lf0p99fvFzTuhoon6WFeddhkH+8KFPY7adqQDyefYw2
lCztV1Od3qGuE4IE/t2iZhaSr/NjgAe/W2nyYUThhDY7Ksq4QKSq/PNgkECyxFw5
UEV/Dxfn+UopaUZ9Bq+7WN7+ainPqvt6FNpvt+lKHj+mKfToNx5L2NWu7qG90bCO
5Fs7sGe/ODz3NX1KTDebNsrblDmHT7D7Qcy3XuewLnBWnpUL84CuAe7PiM5rSMxL
BIZ6sQi7oeLcYlU/bU6ZsZ556vbqiKM1csnBuqKQPK0WPWBPBoT0ulk8jThuQdca
AQ5m1DF8d7qXZ5J/WxhS3+fkFMnqv7+lVsg1Ao6uedfbe9eCwJ6mpLR/CYqHr2y1
KdI0tfdyBNPGxLwHxQQfIZ0PPzF39LLJAFX3abK84CEYA4VHVkMg0xwNYxHTjWzq
46n40AC9l7UgxG0RlZabZWfkeuNJ4ocg4oqd0lnj8pcE566nnSRsrGEpAWuVk1J2
ybmJirD5dFoP0Ek9B1VL3YveqiXM/1ZaGelmzZVBjMxa/Qelfd7Mf8hI8BO3Cawo
aF07f/6wd3lBIalvcZ/wLtSAxTI4SINoKtumzcgO0nCxjO1aC1aLqUL/jMyuNBi6
ZMB/833818AYQXnLXW4S8apkmqkgIgnuRPtyOIeh5vGO5aq2rcUJrIttPGGL16d3
P7kX6gduBYIAueGtlEsNmLdWRTAGr2aSoYz49Dr8ybV+gz4rKvtnBg1/iqoEXAeZ
ky/sKocMBFc9w5dopkE7ZJduvbVeRYhtYBKeCcDGpfKMO/V2vsG4Z1nmr6Hm3JwN
aKhipp9PBV4OW0ie29/q3xbThC3YJ29VYSNb6DCKWAUngkjLia7HGEjyQ9PtXLyW
H0K2MIYY+fa0f8AqViUESO4qHuUcy4Jc33lp192Boweg9z9mMMuS/MInXZD0a19Z
EOds/YqnO+4GpYpLyzK6RmJiyoYcLP4G+oLBNhNKd21AATclaAYlqDA6/ix2rpX1
H/U+A+pRLZcRwJR5AxgL8dSQYyf6SJHmkzQ9XywglCZGj8yOuT1zP78cz6GWOJg6
7nqo3X+MLMguSZrgGjSHir3tvZwtlGfRLGvjL9Wo4/vW3LU/xKvOqq37M5YQ5ygv
ASu0JG5jqui7OTPYRybgsUUoTNsPGxG959BkFmwNz68kuZAQTd3cLIVeWnMyM9SW
dxouAaOsJNoewQHDMctXv6c310Nc9ylGPNz7wZTsqNRIHg1v9QwuMBO2yU31qyaJ
tUJhXHKRiEod+UNJvQXd+xamCfCzdgKcrxRXSQhj98dmLDdNzr4N1HUTsml0ZDHZ
JaE7koczHiD5ie4KWbrFI0UAVYKwWSaARfW7XTjrnmS5bVZA1h++1YMcEYjK/L+R
C90pzcUI9dOd+mKMEFUgvMS6pyRYZfO4xfRjTuRRhFUIXwZWzlfqZuU+BU3fuOnx
LhRuIc9+eBHXqlyJl+NBb1yJFpRbtVOpaU26eYRfnuD7uzb3m00FGxJf/5PmQyTl
kGp4ppSlwr8vf6wj9bOycLQabRJqFujHVVw6ItQPIi/5CjYv9U+eTM4vGlO5Ftso
rr4QqV/GqjzljsJrmBFCH/AmMKItUHlA/yCNr+5mL0grokz3+3SrPv/YTzDlypgN
aoILr1CeZOqiCNHBG91H3BbcmwYmHYxh0NoZEm2BGNrsRi4CAZ9yGqhm60mgxFNf
rgLu+mjIvK1jAoV7CV0C+NcFHsZLop+uTnCZyRF6Bze36rYXbrcGuSNWN9hxrrhV
53lR2vvCeQP423M0w/V3sMKk6byoxV5N2XU3r6Z0xq8cBpRtRl25LIET3g5/BwEd
0Kl15oWFD86SdnN1z/Mus5yhnX4imWKAwa7JnDnQbM340uvGRZMk/lgGf+arA5dw
3U9IPOL8K5YJtAXHHaql0k60LXZWdPpZ5H6/xoYLzpJ71yT9Ko07DoK3AotexHtb
xeJSJzOoFomQM+YUhLihGgARMVGEk7ohv8A3qCLDHRXxlcsnrXGu/MaSjvGM56Dj
6yrt0Xnvs5SuPeKTDttAnsvzeosbz+/lyb92UFcT6PszRnHixtdHwI2VKhrxxvsw
HXvXcVd1yilxeXSC0RP6+YCLORZp4x6ePix4+wJWl483EB5CBz463J8BQGOEzThn
Vx7bqv9wAMX46qBuw8DTYQqORRfX4J+zbVrJj1GfNwsAyO8kuYg3jWOrVmpL81Ff
Skort7mW9tfKEbmnRNcE2ueELL7HswqHX2S+BmH0ft2k366urFGseZOs1BUSPm14
X4pB926K+iK7YwV5iEnKdR9Om2WiwSBhq4qSZji9mhSqjqOshnffNeNEDhtyeIoO
5WVig9Vn/z1ctTWG2V8X6oSDh6rLecFKUbmI2cP1glMZpiqQWGYp4uvJKs5Iggom
LvWWvyINmZRKVDQPHp9Z2eaY8zz4V4BHi5LG5TlAgsT9mhsDGbzAoFwBOMG8inIX
fcowO7drxVaxDB8YkHJezgY6YEqvoykiK4E/mdUSCkEYmohS1tcjuIrxMxjufTi2
6gPFOXdC7e7RULoBo+cNyK5PIXGmNPm34spyS+FCyEC/3oUp8QDlPN+y97cLd+8+
bZYXxZ6j8Ci8HS1ySJxjJ+hHcbYeRaikbCTjsc2PCqsnT5bwIPSybrAUt6Fq70iD
VJA9mNggWj+SHrI9VFK99Yv7J+Uflis6CDTJ/Fhl0z5Z6moJX3upcbSGLunwNaU5
K89iYJVVpD0W9C76+PUQlg40S9s7cCNJEHV/HDVm0WykVxPHcvNjzqCY0f3pEZZx
ebr6RXPlgVfdfdTGwa9xshZNIaAe2+87FjbA0bpKnf3GITV+wp0Y68rhsC3M3Dv9
V+WPVlTmHb8CpqT0CVzidq5Go0+HNWWR55YJUGPsRo0aIudMgeqMLuopBghVf6rg
7vHw9JNTHHq+7S9MHiCId74lOre9nP9rO4ZDkPcaESDD/WRvS2SfqLHI3+UG3ya4
RYhC74vc2TXoVDhVC9jO9HgIjAHuAei7CKAhxeG6RyND21WDlJq8LNrUzIx/ddgD
61pd0yhn8XVcbJXGZT3IaCNp+QnmA1km2hhVIWJsICMEWplDecQOK3sM22lZdzyZ
Cd3j6+mJLmKnyJJ3yj72/NE5eJDkIhCKjhdEkafvPdOxQ/OAI745nEnj+98Kunlu
mxkCp9K2dWGb9XGFn8tFpyEaoW0H0sRsayi8/61khkxJLInWtzjgExAfUV7HtJco
j6keujw5Is3mTrdPIynE6grmEIuvNzmPDsv/RbdGb0X+OX7YHu9m0wXYhmfroeAV
JeChyqz4wfB0xiZDUPxkO2e4h5PRzKZ67M8+q42PmYpxeq9PYLi/A2ljyMspFx80
87cT0dqELUO0T7VRg967NeKpKump5jOEZt4tAj4MhEz25k31eM78YUAVMsHIB4O6
cFWwNjw7FJH46kOhtCdCVydia9LPqWciLok4Y+Gey3o/r6uP+atJv8we7dbA8yhD
dYhdi3oUh7zvQEzTo+TjceMWCq0BcbkAVomwCTWva1pWNPDGmvPQf44XRJXD23R5
QxVF5jt6JJ1ZDjnpvRT4vQ7FyW3F90AP2V8t1PgoGZ4C8dGBx9oq5Oz9zfbZnHvL
aFVo795t55emOi5zaRA9uqedkv8bmkajqYwa7eDq4CLC33bMAEuXeOk0T8XS3OqV
3Hm9qjSqgJxL+WfM+1zoKfK/lklUZTfsddXdPowRzdMetw8QoNLTpjSueKyrEguo
92OlpxhD6Ix2gaU0c+xPnPEVh8hNvCMIEMwROxewQqXlgQyv28UYgbG8QU12DNr6
RFQ0ew2RGuD3qkFUfQFhD6sfT5tqsdNycPvuVm6xGErqb2LQFjVdCokf+Tr5TCsm
tvh4/PbUXVyGOK4yhr8k5ckxVQQ8L9Nt+tdXfIUL/5KsYuaSJgWhkqq1gS/7jAq7
/NbQ4J4sEKME1Rkr34UCmbpLyFA22Bn4ZSIwmTVGXZwKOPqh453P7R8dF8Q7/UEx
KRHcxCqKjZMC+bEGhuRKNprQS8qclI1Lb7iUk59tp05sQKl37/lLsRjDM/M5tLDo
LfJZqNgCDpkG7XRazWNaLvDrUvJtnvMYD35gpgQx4B4ZyV1vWJIlYZ9TVdY56JmC
3HV4M4gksFSERR8pFfPv/PlPhU6/ECbJQQkKYsaIahQtcbNpBVvIyNBfqijT86wc
5PeiUczGSUI1Slg9sxNoE6sctKyowHI6ds+5tfFUVXo+nI8d0bQD+/ihP3QN2kVn
HBTYPlw2iouCIrpODWZj53orV+hzc2UVgYch3k346sAssnoVPtX0+K5kyFzLEOx5
ZPseIJcHDNXhF30n8TXDg82ijfsPX2OfgcjbP4KSPk5bxW5OLODNRSHLWOO+a0/u
fFSUzJX/CpvFmMaEDJ0aWn9yFw8w50dxqPWoDlsl3mCLEEvFiMNEU4a0/QKdJt0/
+ApDgrjJyHEVD0Gub7CQ5g19pxizj6Taps4iyzrNFFojLN31Ez++dPjZgcuoFnYM
R44exWZGjawFhqs56QqR59i8bQGFzJcoJM7xOoiIVPPJX3hfVMGlgP7TRc4P/yhD
PDcyt2GCPLqHorKS+FA5N4xnG3eR+CuzVGy6f4HVhOXGtQJRAtOuD6BHLQSQ5eoF
iXs742c8Z6jmeL985oS03H1O1Tj/YDKVJEHk3wikN4lkEHjkO7oJfH9Hn4Ql2+Uv
BFz5eWXOET6UfrhRIAHW0xp+Y9EhTqPx3EwUmALQXNci4iIki/3V2JrQZR8WU+JY
xE56f3MYSdCV1xeWIsJpH70zMF11ihcMhW9Lggu9pHzNN03SzKGIEJiV/hnEPmz2
HWjZFc/hWuykU3cSGJucQBhCMGnaJJrsif4uQgatNT4vcbL+PaQ0VX/rFjzxiFZr
OBfQWxHfxOfxHURrMlWN6sbIoDFt7ATszN3VUHYzwXhQZVaCq1PSj5l8ShwXQtRZ
gsht/+BavyDM1BDHitEFZibJpx3gePrZrMaXrV2UfsKrV8jSDzgERWh81mi8xo4j
Tu6GrnevnkAzrVGnXzJy/7dLTxQxpCyxvpLYYDxIxUE5mZ6N3B9EOAtTpLqS767g
a0o0Qkll2KQfdHQB6jDigldNqTmcc2gCBYHLsmxKHdgB8Nyl3Qbykag6XKG8Kl72
Um3dGYr3sBjlKr8MMtYVZtT7oACe62+k2qdKS1e00rV+bDpiSNl/Fn8MuX3b22Sw
teKi/lKTtbbz7WW70nvw4LUo4Jvd04DQxwd6uYnGjlNB/Huxv+pZuMyTOE+WOCyC
frudtbBQfMhlT1F8i4ko0cK/0YMfmhYEevfs6UB+5Lzo5WuETUANiFiYEG14VY88
Z45chYUhT4H2Y91axAgggeEEz8G2Jz5Eou2kjdiTaYUdUZX5J7k8MFZVv8bXvloI
i6XamZDFcPNh9GzVS68s53Gi9mM+spK7c/uoRmI6KqkTZp1haw4B/e4Nl7M6/08c
WGYN/8B+aRFmEX7vWsOsr6IWkAoGIg/NxGZ8tiRi8Kk6i49tEp4ke8i1tdv0Hk0L
M0Ej7MXzJVzX6161Q6LRD01841e+CzVkxg9s9HFlTYVm7SrPkYmZ45U0+DuUmnyN
XwCOCGWVgOkNoljIqg0fVvyg2e+/iZlThAagW0DtrcqboctUV8FfdErIv5DQ+p+w
KfcuOSxZ7UOjXcWMrmgKiiwN1zyzOOdnwBNjuS3UMJcTV90j5Kdc3y+jP46r4h4T
JUKrtvhul00zaJvf3n5btQb4HFmAjCa9z4EIbJmeRmY9PvgdrbFZOrWc9xmaaAf/
X2fcJaKqzNE5uVMOcZDdiBY0rtivL8xJ/H67inmEmVeZ4Q5DMubGlAjUei27Y91R
X97myyHzYnMhnY1Ub4mmKF2QSLzMqR2FtDAMmNEd4pQdcOj5o0zEqusPe4D6vPol
y+LsW5I9J4OvacR5femgbeMQoseantED7zg+UvZKb8nh2ETLckmzKfORP3qxLCH5
bGli0JZdlaZvdYwaFUtAoKyig5nWRRM6VggMI+vZhtTQJIrP1OwFGS9oHejLYaq5
o3W3yVQnJ6CS8UYjHhtFZOfNXnLfgALk2icbnYU1q7+PJvPSnJBc10ToJ6xPiYrM
msL4SphrDPCESqLMOVC++TYFF0+mt4HqvAHrfWFBCmgz/+zHeTJ48ECWQxVJDDI8
n3ITvSevyur4IqVGNaYiwyTLUnnbM2ebpEWzB3KYoaq4w+O3oo0tUDJFNVJDYwgM
hvp1fTkirdCU9iVTD0l0a+EiyUZ1itCJjaHT2iqpNCMBKIlGHAMMwwR9YD0eySjA
Tjuov+bmaijOrjsxVrGW7PAF3Y2C0X7LPzcMnz0xaW/C+BoBg7QEooJWpo4UXylg
EHFXeLSTRYttpfSCY+HCLYi5c4pKcNl+DuB1xuKOxmYYJHGYFKXnlk6j3Wn7Ge7F
Z4xBtaxgRFPG+/8kgOZxQctLPOIq7NXgYlKxQua5ShmTOFy/6HdGWIPRci6K4kEw
skxsm0w3pJ6GNQ2HTJxY3sNx/tUApW81MJHNjFgFSXvfb8ZYgMUGFYesQc1Ah7rz
ySwDOAq82JwyrkJVG+hGKjnikFjAZ/yfIFYshdtG61YfVwo75j/ggXSIzgwd2sZo
OQz9QNFgANgJC36OvrYuWfowVlS5JCQ82+jLOz50WCw0rcK49+mR4D/GHeBkxvkV
jBhoiZL7mm2fRVHnmlvgoFiWzyadCVHtzjB12iladxi5+iNNkeE40yJDNhvRAbJn
HxOW/ZWt57eFfmfSB5G7ZHdZBTpd/hOFN4xPLHD//X4RTDd6fzBfEjJEeyFYp+vd
ub0Y43GO0ch/lQslnTz8g3DjePXn36+go4Don+M0bU6FTjadjDgmhvcsqxJJqNxK
sGBl6HR/Yob3sUc0oTQ4WfTSHL1hJ04S0g/8p+UIx7fxQx9WFbTKvEEGJlZh3bKD
OVycAvwhn3nb8bzn0Vk/kUkM4dh9eFtgx+mY8IensDasvDgxdJbWcAdKtkRmVOwj
A5hIgMD3AC0kcQillSVzUpm2lF2xgdFURR000fZo7meXYv/VGNW+qTEwyM3gz8W5
mMiUMOsN+oohcxkrvZRCW4WDaaTxcO6hGJvK/3G/4QIt617JPMmZx9rePLx3ZrcL
pEm/h9gHPVDdDWjJs//dIAVQzTaYRgPFcdz4qK1wIO9acLQR+zpbl4RCxOM9WMLt
y5bNe3hCNgBwDzWuZSww+9m9vNzoFrdBtF3dbYHl3zKF6K5lmyy4MPqQ2pKwNHju
Gjsr6k3PuRcY9P2VLSmF1BVlfwv8m4G461gLyMBnu523IPnCQbMHm6ebVaC17T3+
WdXdCvd3gIGtIduLuh8uCnUY22EqCfu/e8JJCWx+FE5Ru7cppYDKQiftP6/Y7by+
wA3EWuLnWg/hupfAI7J9X19aFXpF9wFFjR9k/K/gJGL2ZLPJVaSzK7vEcI/LwdMM
yTYvjq8Xdl6cKNMH5FBGL7EnOdNk40jSLkmQGcTIR394CHtdjlmyy7GcAp+1I9TV
2599h+swski11nf9GbnlN6/LzAL7v4+s8AXKNuXSWhjo1rpRsx51euQhUzW5xpSH
yIxmr3B2w4aLj5WOYI71+qeaV/1Lbg89Ogt/rIK3UQo6N4SS8Ps5qEkUjJuqb3h5
wXul2U4RvSs4gQ2qh5xccrXpBhCbCGxc3GnbTSWilIHQg20Y4x6A3EqKnqd2Tsxg
/YFb0TNOySlCZeD9hKkzHvubx8J8H3Vh9qC2fibgwZas4CtyXcL5PMs+L85R+s24
IotkbiZ59DmDTodsMlsb9IdbsYWTNYHEFNsdmEoI0A/f+Q1vaI/7BDXzMzn1Pz+/
lgYkWJ1cFcVh2E+Lefswb8ARI6PY9WlqdB/Np4XbvnD6dWFH+WrAjqfjJPMCFn8t
4ii8o5nYBZOxvXckektZUYVUyixSnhTfMU1ezNXxzUmdlpZZY8eQSs3Z8Iqfix+E
OgaPy03vjInTjZVjkz/xUViLzBjLIMBvOF0mJQoEEVN2bk90SAeI5VF613KB7YLx
2VU/g6iKJk0WH5TTgtnbUydE1bpEnePsdBNdP7Phbsr/FNubhOO8KZUhF7cAH43R
zuG8l8GiP1CAJvGjncpj3pAaaAUgDd2YFQfh1jQxmC5L50xXV6NuelmQTe4+SwhV
IWfv4Ngulupe3sRrOgmFliVn0pun8LVEwC8ZLUBLeY+SMpp7id48PPb5ztUj22vM
kKaWfe5vcX6mS+Maa6CSRxiZtJCNeKDa9DEJMN8perPP9Jct0i40kL7XO1/3sUw4
wlKvMDEqdntMlMKniTOtKnuD0WpGIqCuDO21wm0LRj4Q2EkNJFMleXe21O/9sDay
GuvdpsWmvSUWuMb17QOoQOXWQ4RgLA/xyOHnWrQeutKA4i48o0yronxpu9ExB2yb
0RuSsN3W6rjG81ZHVqpWxXiFy5G2liFYwONH2m9RO/zvapL/w4AK+OIvkgSIe60/
6N/qNk2UPZQwfJnSPTldkhh7IUS9+x/ovzu4pGm7V3oWDJRFfqLTsrYmXlFoIW+y
DMxsi3lMdTRCkriqtTJJiQTwx1fRx4fJ3IUhhJNw7UMeCF0wXYlt6IMgbHc5xuFo
dB/SCQyKjP+R3AJBZDm0xoFNyTL80dymQyydM06AIauOtwWwqSQvwt2iMPoJT4rA
YephCLypyH10lFTR50AXnHz1/mcQmtdnUE+yjbtMOp363ES15VsExeqgv83IpDnT
v5TTwq1uyziLRSxZjnP6E1RQKo1SKIffvyeWfSB2Avt1MAeP623FumBs7HUmovJs
5vT+RFlfYooF0hz1ZoenNJDHTZGv/i3cDhqlyOJ9Vw5r7031UDzxGjP1w/rXAdlw
UWFDqETz0jk78rc46N6lHSA4oH5YqtlG7CoJoGcfDUL3ao1D9yS8ukfhLCm/0OYD
OM8hvQOPZpmhng5qz1VVoyhwzZszrAgMsR2YGaaeuf0IL4SPVB0ZzluxY36JfsTL
N7/8BrvXKQZdep61OUGqmnyfglyGVru/1tL5JAK/4tzPb5Z9QuOR3walbc3JFtr3
pI00BVXD9rBstYqbIoMET4L5XVod4Il/E0kub+l4SPpjpUBGhEhhkkYTi38PiMxG
mCzxHlp6QkP8KdGcf0VHuXpSmymuLpMmzEDSdat0rtldeK0pNLtkKHPwrUKX9SqX
T01npFz+zdt4p6N2RyUYjAvdHMMc06fTNVWlezJovhe3HeX+6d4NX9TgYMVKHTZ/
gukX5iTk2fL8oexONweRpG/Tann4co2C8XtuFv0WF6u9BuJo9Aer03lK0q+u14D4
ra7RqD4XvcZVNRZbjkMhmCQ26uhq/s7qGElrqSgfInsfW4jrc7OVimu+pIV67AAm
cV46YFQ/KWXf5zOXsdI3RHyXXVnl7KIXdxRnkWI4v9phh0ELCHnu6Xr+na/MAqUu
SGXXtGqVYh7ZGd5f2zkGieMZirQr0YolPY2ekQyyrjgvijLNK/Ubny3obc7i7N7f
JSXjxgYEAEjW2S5P3Jdl7t6fSzDXV4FzBYUuwJc/UC7umRSxA/lO9/LtqnUiyfbY
fkMfXoTLGBQxAPofdlZd5tXA156E7w+YIhUuOJXtbCr1ENb0X6gBaeSfYpx1vpbW
KNkYFh2sBEhQfItoqdirOR+qHT7uIrnlrRbeFymfmfzIUkyVV7nOal0PyV3o+LXb
Y5ySGFQFu1++k9TbdYyRr5C6jdbiViOVEEakfscLjTLxwIy3twpnKYvsUoqQNB1O
W25ImCqg20BUPODelVqVgQHbJTe7Spfp+7wLhRK7gpDlskkYTClFuIC6r2dvobB4
dg2dwmcF1JABPJQAeZDUi8RAsDebYw6Bn6B8C5lXE85V7+sMUddRvs1Z2pOYLMh9
iE4D8rER0KhG5H0j1gRbooXFmqeadRf3+2etkt2Z/kwAOEhhSGoBXOZSfiIX/PLq
Ch6PLbg4cExRzwRsb2exkDt/msTTRJ0cLohg84NQysAqvSNy97wu9y964vy6aHTC
RJ0DYDMBGH9N0m5++t3Htfy5QM5DX/4xWH5r8lHP8wzmkdj8SyI43m7D4SIxzHW4
/CSBtbUl8dLzHjJRMX2/lQUJkiLSFpphYA1NprwnywrDcb+73CaDNhdhdtnOugvx
hFSFzVr8Y3gZBjbt0R+OB0J1Sm2+vZReBaO0yis1wojK1h9c1lavtNGIygYXkYm8
VNjwEeNh9r8/TlUhZRAJ137IzfkIVm1U9/I+GNccjyeGPyA574tb9dj8/ZJT6frB
FaQFK+zgxR5JlRhoA3qQyZlt3Mc1qA8PG5iA300oPtqYrp/dVniJhwZ33sZD2HlV
FioUOryYIPu626v0H2+ZaRipsL79bwULq50rNPnol5uAna+IydVSdpdRl+6euxPu
Kt9nfFoyrExhe/53wX6KQpdvDVknIgaSO4BBMQyOClxyZd1HrD2h1InGHOzlB/q2
lqNsc9ibXSgJzC8XalMFzColGrKMXIqRV47AzfqLyH9g9wxa/XTqHObGBz6f42Ke
iONDNviDszPBVOcE4aX7/BUQXtG6ia3gMVy56s5Qd/URepbUtLA5ld/T6fib87J+
ZTAtT8YouH0cidx7DoQ7JIlQNnmt1BtM3bEYJSOUO1/oxsibDo9ILvXv9IJKdYlf
CvE02k4UH10EbMvGefSUL3hMJeKzbBAUu5Du27VIquTN8amPfeoemdqx3VdKDmJv
2CRA63HWmuwKAHlPM8TY664m3fdOathalsJmMx7jXntOQBXkg3+G5bwllImd4nwp
7CElNp1toGq6AYX5avdQBqTEwjMb2dqL1/Q9c7+Ag8u2fY6qJkKQAcDJKtHQybGt
yT2APjQXvsXtUqRQa/2qUj9GH8JQElTptk0b3Yy6K0dv959PB70UK7eG/EJg8fSo
bhX2vJVSEJ+C1WWM+xFjdb46wJosaz3cq4SMak5H1Y+6V2VFJ/Fj9O5vcDUtmKOI
BUvOMnfYdZCmc5EQbTqEuQNPRO1/br6VUYYywpTjkZ7Qpq1eDtRsn7RvTn3t3dJT
Yjzv6vT8rOK/y/ERaAsxfnMYLn35o6gt2gveTg0Iga1YIYFDwG4pZMpBMdJ3MhJi
jDzsXEsW7bRliTxX87YDo1JxZmqkAPBYReqpWcxezYoYHri36tDKvT+Jadt3TCjN
0sj63WO593R6LhSREWvLTVjkpE2bEOBud4Wi1Cu+nunk32ZE+8lRrS/IJ1SZ8ORW
wfg9l33GAKBIjei8NibJihy1B3YZULSqBSO92Gk3XC8tKig8VMda9cbTmxT4lfas
IxQOFYYb7gBgI8bVoRwiUMq3UGX6UQMHtB2Ruc1dPfFJRDRRrUxqZpN4YCMyUZG4
+zUsbEjaZaBA201POoJB/j6r6TM5DOcPuG1lO/mR3U8VPa5NWrTHvMCvwzWii+Si
MsF5eL4ijrKloAeRDty8gNp8yZSMf+mwcvlZc0v1dd+n9orjL74hf4SllmHOEoJJ
LFWZLJ3p/jnFGJauTInXpuiIQtTweZtAPaI1PQJiNuhp6sAda+ZYH7nfcW57EohY
riH/XeyVW49ew4uT9W8NB6STknvQqo4MXHuHrnEn/W7sH+vO1y62o4YivDau589l
yCBY05w4Oc/60NIocP0HL+tdhsNs4QvL1phpMkUq8ycskCxhejNCIsq7UMsRWrUa
svymlVwHszTJRujrfoSUi3WqvLJiwZGHD/AUA4lDl7WS2vAtQ7b+RpXFlR/vShY5
RHdt7Dg3FP+pJAF1mjqIe6bgvw5IGNQEIEhz7pvBsfPccmoIVM+xBl20mhQWCYJq
kDjwGayvH+XQxsgVvoMjuTtiAuleeVUX5z0bkDzGPqqej83ktLXp6pTP/epxsvaR
j/jV3zkgxEsE4SOa/Zhw+6kZuWfq7aO74T6f9RH6mX99+LT8euLr6wUDyYjpBLy1
hkVHCife2q6mZMsnKVZFwaeofgPZWyBA9cJ3Rx/cp109G9yXDLCzhiAZjVGhD7bz
cxklm9Cjf/PUvNDxJzqjlbJ9uqPmsNTsPiEsPYSibLiXb5+mwIU12juQVZbOUNZm
M8uyTEmeW1hcHATc+xqoC9kI5hcb3kUOUiLw4qpESEuNepXGgy5WwkWxXvCQ563d
roUSXJdWEPMQxmCmOYKjhuvhFYAb4qKRxtnJd3TAdIA0mbHQSSw8GeIlgxmptOBd
7Ho6jc5kWmcfxBbRnQSEgttXE/RSaQI/44Oc28jAtV9RpAqMygzoykTqmCyxvmmD
o6dO6WKtfG2M8v2F+bylefVEuOONJSXPMBebPwAvp7hCEhQVft/nX8HAe819CKJn
gDSk8aOmr0AUrFJhKprxfKWpyPDRch6Q7O1KYexb8VAZNTTCPnIo0bWd/g6mSCRE
M1SHvfzHwCCWfGx5SOmhhNiunjP70zGMjr/Bf9Ciflb6mnmMC4P24a9V4OqKydwx
NwhYeXWYqLs5DgvY79sYJGn5sdVQWThKtJ9qb8zqJzcPkECyGLvdn+JFcrhVaRh9
FR3doE2T9FvC7YtdKRYxnVEHNWD2WB00w+TzblW2D6gC2OhFhYhIYGxOJdSDAH7q
TvxlzngWo9rLcFyLkjZbl4iXag1CVdX473TmlevcPZkLaiHsvBG8VVSvGd2b4g1u
T7BLhrZR3Ag2jmoK+SyjCuuXeXWVO0Q5pJQnlJsfrt+w8yJWNrWnxlbFqCLJt9MQ
VgM1qKfEFVQ8fsd0qOlNOF9WlMzLAtemW1JhSWjbMH/EgjS33OxVrntXgtj0QQfn
qhU/2rmCmuGnnha5nDg3wpOm6PSPlPCtQUvA/qPrMwkzrKfosWLTAbKs+AniOOeF
1YZeO6vvmsJhP8ANNC6141AcowiL/tZjTP1NvcRuKybQeWxN2NfCwBAMeFstOEJf
C3fCBEbzFu1PhICxKAvpnprSmv/FbmuEaTEzVYyfcjwth6dUZXcNuKK20LKs5eVF
dFmLFTOS4AxOTQ9l5h+/Dg26DKHpAnqyU3XBTApipzRuxqpqzk38VpVWWJAH7+go
G6Qhl/arlNpC8JKqs4myIbrmV+mrO8pvsUJxoglXHgfjQUJMy4M8OX9xJNPrMs+p
x+KzuzxX7aDYnc5otmEr7uw4PwTFnH8M1I2455kzYg/OJKI0RPii8woxza+J5j3Q
cDgNqEItIQvnp1f0m3rMMxtF3UlVdlAGm162ypa0jvKJfL1YdUja5PL5usvKruwm
yXtz8/Ds46iaANA5nz7xcMzNKIB9mEQH7wlNLdHLHObdMy0iGMqBxhM41abslywM
1PFPsy2t+UkzwVuXrzWLzc4xTFBvXgLk6u3UJAHb/NZJfh7aLJc1rqfQxERPAH1v
iYrrf1wiNgZSM3GAEIAbG6pNjOGCxw5RAVCtF9+Pucm2wIQlrFcPs8jyWp2F6Pb3
P8WR4rAmmTWZHbr3oNc6hsbxUY+yFJXPhVNMr5oClSx9zsOKYopDNVRt1PC+cwnS
uvLQarbBxK480+ACIWt0M/Rh4GZipixs65S+rzz7/X8UKyVrHWy2Px6ielI5BkzJ
yCCJ15kDZWRd49Mz3L7Tz8ZPexqnmvT20i4EuMvZosoPCmg4W3Wewt7RM87skzVR
TDMghz+vOB27ZGPIZGx1zRqQnPmHLLu9S/xEMwvv0dfnsO4ukWnoMLJvgnHfT/X9
KE5hPcWKUjq12IbvPK5KQ1x64AGzSckbyo9ILJK1yD9PDTmZQzlNlzajM6xGWHhu
dqWQ3g/Ou9f9FgW6ufolUfa06IZDRsPJ76iqKAmLx6FYtcEQoBqRzTN5zjCyHWLt
9wNcbAYIVSBXZAOldav99e7jZ8y1tmorHvGeLAMqyuCPtDuJmQ/4GWirekMhCG7a
+2mE/KZo+qg96X9G/thsWa7//ETDEQLqM84eqilEBAN9Lkyqy7MGLdiwGvn8XQAD
4ro7ImKYxKZ7CD5wRX9ie93QWCaG5LXza4kZS2esCBHE0rGpmDUaQPXR5lUpz1fy
rkoWdki6Woj26wuV+6DsZYfL/ksSLaCZDkGtg2Q6nB1g6RcppVbnld81wQKOP2U2
MFKfvf/8GajcbGwgtcJtE8g8EiLxzHriP3oB2NsMPUan0RA2xrzcJyKpFYjqb88B
41fcaTARwY6dizLBVF1WbKjpAzbeVk4pcQdr1JKB14QosHIuH3nrZ9vGWTy0qPIf
KJadt6+kjYSsprT4T/YOP3bqtDQ9XFykZl9II514ea68DFFGSELVa+dLML+Hlr3q
OoTjLuKbLRUfIy7tawpU9u0XYcFBjdrT64s4x/S+7HWtKTQywfh6i9ASsGa94I1d
miq3Thc6Bskj+Zl2NhLrv8Wu6PnfokC7pM7jKZ81lnkZAE6rFkm+rA9bThatdtot
jqZSBHSWaAaOwTbtXxzNaq8Awd7qfUIhMsA4T4YiZKp6j2AkyiLIG63BroBvGB9i
TNMp1Ve7xYRhIXxe+SHqAgprGiL8RUhRHUG2jfS7QCpDU0AIy4kwfPTV0j5sq0l/
kwiWBWDhQcQjMDOwZy9baRdajc9Wcz5P8wB2d9Y6xELFIzIJy9y1xer7A5vONoow
FRmx/q9lECyWzNbICEBbYTezaNARGbFzPFy13zeLAPSPXhq/Pzat4GzsqF4+j+6A
74/McKtU3vQ647013qHi95Eks8iHHU7aQhUo2e7y+BAv18TzQgNJ9C4ZN1ONNhJL
HURjVxzRewOKQr0L19kxk2zJMKFe0fBUhmnPWZSvM7nxWvT83QlNYUdjzBNG+v2F
IJXJKvtbfQPTwq4BRqJ7HacpYlepsmgFNU/cTA5wTvn0l05qD3vXo8G4r/Aoh10N
FcqWf5DmYHPWZxKcjJhiCoBPrAxBq67pvieQ7c4fWawqdJAgAA0EwsxfJsyO6I5N
qDZGUxBhuflOdsBjNj/W/7U/8ghpeboVj0irdYABzElOntW9gtyz6M6KG8gHBNiU
9+Pq6F8slzun9ZM976njw3mnx/iepyyesx8CG2OvWFyhiGtQtFHpHQJDkz37jNRX
IOoTO7voLH03Qs3TMhf/4X1QpNewpwCxMU/wWb3A3MlzVTZ+6ee39/Gder8HdCk8
W/kI0sVU/gaMal5e9Hc2QHXt3GcVWsVICORa7k2VkH2GXLgNh5TEQa6FevPI6SV2
ZzVFHzZ8MS3L6rwpHlw0IlxQBO9AK/IQusb9BFsewddSzZoQrBpTUKEYp4rnig8v
VtEiAlw6ByRV0CEgzrF3yqtCaotrCBMtmW08ZUA0Rzm6CdmvyjvDnJMIIRABuwwo
Whd0WSZ56AbjdapjMKd2KEhIq/8yOPkQpVc4WeCz9AkEIrw+ofX9b1RIR7vIf1Aj
+pRPmGqaQvGpLwR1MC7KW6t2FaE9qFGqY4+0NRoQWe2SPq6scTTYY65n4fFybqoa
8E0DvnHxQ9nzN14NV8zJjfhpTdtiQtSuRxuQgBy6dvNunararQyTpmzXkouogxoK
oYxMJUlJgYPkyfciWg7ENnVrXLG2s3JY+yGhu1cPE7aXH0UtGz84a2XurczHmpD7
Ps3m/JxQJf+51xgtW+z78/vYQ3zWPkHd+Fo/wdoh08szOPEFXToAel9Q/l4WCj4c
Rx5y5lBIlxfGek9DJQ1uDCkJswPfIlm3z/HuWc23nVu7hv+AQnS0gME+US01eHgO
gc9K0domGucChCl7Ao8qYmyH8FByht0UXG/dJXOhr6V1WJSKSHfTKJ09umw9gPTu
RKuGpR1Qt5Gs30SpgcAsUG0Yp0V7Pz7/ZwBOJ8QJ7muwxWCAUhGXudIWew9LRpOd
s1WFXmyK9XiC3SBWgmNHWCeNyHcPbnuAi1LYhCKVy3Qw8OxyV1oVGc9S9/u1vPB/
7umURdVCGX9Xutn2DHt6Sl59jc5Glglgk4oHauC8tg9xQtmbFn1I5HMHSdqG1aOr
sDBcCefS3XBQjckgJsnz4Dr2HAU8lYMXP4Ggnd5ycugekAwcUvtTrL+BBjfpIwC2
aBzCjTJTyTw3cTAs5V1HtKm30lYej11ZwXN0HUewEz7XnJqbidk9ftsuAafg++JH
LL7nm8qEifbphEV3HQ54XR0hgn6OSDlsfcHTVXo5RcMoad4n+aipxh/IXlk6Ltu7
+cRrHzeFJvz8oQtiSz8WzGoHgwuasF1BiHnpeotkpbg11nGEGWHdGvO3iYz4dFWo
kK/v76OzAX4tGeDq87RrXQfkxyACTvb0g70IucQsDUPrnGLG0q1SneNYC3hNcUZM
fb7tfP+fQxoe3LfP/opfyc0wxn2z582ItzLUiJvlHDy8qTi3sc3cv0YMnKVEijum
5pa67qCPD2/r0iwmqp4Ce7cOG5YnjJDwEne20r6jsQ4E3xVz3BX/UBk/d2bLzyYs
wI1GASLXwkI0BHfP0Rz0na6QJz9w8WUhU5kVanvFZQSAmQRUHWlCnR7pRLsBOrmw
+61s+K2VsrqcrHzL/pZ8d+wijIQog30V6HOeERueHKHsDE7+ad4oU3sBxbFhSpTC
PuzHyLh/hZk7SvT4xCoy21zhIHWQIAAzkgMvuC5w3D/MUgPaH5uXF8CK63fX/6BR
X73SB1b1SGDU1seHkorHGSgPdQpV2tc84H0GJgb6ugHbCjXaYIs+iNJPI6Emn978
N118Q2n/jttbviiESZoos6/eNswFlYWYazm1VcgVV52vXtWEecziOXZjcQxZS8OX
qj1y2vWd6IpzLSUBmYAwfNZeiQd9FhnAtdVFD9STeQeY8XkFLhgHXp195QuFJ2hO
F/oAPQTPuGSVuG2YowZw8eSNgNFOKN2aB0HH5cagNZfOxi69c9b652gBfZBd73ty
7+BaQKTNhxNWrv77pp3Q4lsyAQJVtCQP6xzECpiR1WwAOMfyfPwvmr2DmBfjSI9v
4O9YeSK6goB99rUmgN7SLYiymIKjc4MS3dXp5zqwH0qjH6aA0sHjwjUhGs5mmuYS
syHnVCjJV5Ce5fOO6cDjmaIXYWI0F/iA857fg2f9MdzW65+KdOS/RTZXCYarS0g+
IExY6165AadWJ71PfwwUGmJaerYJOi2FNNeTK2y7PmEbZLJsNcvwB3/zcuh39JL4
7msLUxd0IImjJQ9jc5dq/ZIrYHL2ZqW6f4A1uLu/qRPCj3slkV3TLsKDKCfv+zx0
Coz8TVwouvAGQ1H+W5NBHlb00Osg6Kp0gqfNLqQgK/i+WvON+ZaKk+9O9HxuDIZc
dlx5Hg0Hp/69IaZ7BOah8czx+S9diTXhjDg+8HSX84x8fRZlBoWMkIDfFGfw2+u/
vRVJUBIHGlj1kES06H3CqiIA3vrsB34K3zgzImfFpxXwUsw+qgq4dWRH/1p46MqO
oU9utBuoamhRMFCy1or+FgtE8wxc3gINC/k7d/kJMvTtU9L7QT6oIudUoxmNg0pC
OM6TXleelTIseG+Z7bfVoJvN7W7719771gmh11m3x06MxUY9rvZxd8t3JA/CJezr
DYNKQTFgWij2+WvM22ZUv10tvGpPKDTNuWe4KPR/34any6ID4rUcN18fcQhmVBRT
MQb1x2bwxb5LdSTk2XaXvpi5C5lyf6am0KPBOGLAWgWiIvcdcMsGBnrK+nl1bOQm
pJMar/rvGFUz0PJcceWramr4K4sHO593Tia3YbPe73ddAni8lCdOZTZYtELAQ6pT
4n4g0Ao37zjoD87JBiWtE97vPBAiHb34LJ3UuOr+MeDTj3BTD78rQQiwfLqy4egG
bEJxm4XvnxLJyRmPITIC2xIrraw8EFyIo0uN1mXxXC9mhzowAIwYq7qSlwobWS7Y
HM72YoP1w/KPdWxESxvjP8oXBtvBnqZlN27UqEMte04HZAvOs6C5kG1y9UzdAYtl
BKrcRPIV4CIjg7q5va9AEiLqOM0H9cScoCY+jvQmY9lv7wjM4yB0NvKVdKsmj4zw
UYvmpILClS9IWTzxSeUnytdazjDguRt5d2rRAPiqdUShAGPFvcbl3K+8PSaxsHaw
IdvAPXNii3VSsFfMO5zbraEXGVDbecZNAS6hpa9IFqbJIy1frbqJTLYdfsEtfneb
/gzk5t/PhZb8ah5mgfO1rc6nKZTR5nUD0Oui5so8WNQoW6HRgytjhfLb3HVk6Vgm
SELs4NypWrdoKa0RkBdv5pI2qM/8TkF3GFL6tRFXEVlzLurjTIp8GhcyMj+FNPgz
d778LR9zUvzELkKiHh1js2hyD9k/Q5cZp91/6mbz639Y2zMpwR+2gDtlo5wSwHTV
6avYYdA6+O7ZuBj0FsSC6xmROMJhmMiJeZAjSCxc0KHMZTA9eTpAbPrI/i8p2kWc
LAc93ksy9unruyZgCIaJVdV7Ik/KUgQmAJEl3LQuCwqMByhBE59lCOaESEbuCz7M
RkdxC98p+ppdhI0mEBaM0N9aWC1NkO+b/s8euF6xeWOPyNoFt6KRZHVJ95oJWxU5
QoLPiJHBLMS9LbGJOAVXRfD4TUugW4BQvSnFeZF6D3ir65Uej6AijVoBsNKZ4ep7
8xi4rmX+PWa1sZCGF2dMu7dYsgkb4myBfMxJ8P6txYIsShndo6vC011izgVf9tJh
uWPgtVbez83vuIqCGyc84TawPlfkYDasI0wwLGWM6mL9Kgy4DNzXemte1AfE/rJ/
5Tq65XX7lIhyO5V3Mc3Q8YGtfJYkmmT0J1HDMBdlTpIACbu0qtAa76I/6A/TBEX8
WPOyPJrN1thpwp6sbunGaEEea93L4jdVIaTRAXzr8QMUEbtewkHv1BB7d/y3mPxL
F7ed6s9DLfXNEZSWDZJLCuya1Qo/QYez4Cq7Sc9sMvmzX5dZrPRNQINPlyTKpbHv
cf79CRjTlHtlbREd3qOEhakYvtAeRGKj/sjjMp8m8bMVKWH2VgJWkn8NUkkCSKMD
774y4FODhT0tl+YN8geYxfcvVlrzmSa5RFxwa8kKpqcQ1e9EySnMs7s6EA6lP0IC
+rOsM+guL4q7LkhPl1wW4KfAz/NrIoIlicsSmnEavg30h4N0Xk0/HArHshoNgyM/
nUOuRQbOUw8H3hgL+vHFc1TpdREZufV+q9+kCd4gF3R8MEmSCSLPKtXxEETUQSll
kbnvhlWF85rBJzqg0fjbJUUPKyB0LzJt7KzBFDzLUy9XV0BMdP7pOdNFrtQyUO7g
+SeZi/NT7nDWrq3V0UGX3GIFWlwebEXSLBXK994oR7gM7yX0sRVUFaBT6JQ9vHU0
Ym+Dcr0YGnF+NcaavxCWy4XH+kTIaF8cBByeQRN3NZS+sEOrKtf/YoJValrAWRIL
jbEWjow84T4JyF5G9j9uS3SvMTRUrvEWw/yik0gIuj1jFuvhYp/3IPsakly1KZ0/
xLrKpeBU5X+9lI1Sdjr951nWimz15MJsL9wOQbCURvIzbmHPh/FJalcbrwPyJs7U
6EzR47xSnUZxc6ek9KmD+tYUix8q4TaiiwEwDSNfU0x71vlvtD0fr3hbmCeTt4t9
O6BRoOSiPfPhM9BKaqc3sBwY10R3IDDTZRVVDUCxJMFTtpngOnGuLNna8qYBk2XM
9VBh5qwO+caLVqAKxEvkeFBPGrAfyas20ptMEsqF17jVpZwpg5jPEhxOrfKrav1j
UbQ+weYknwOK5nSyvFjpfJGgBJFaSxgvle1LMxC4OkBtneqOgq8hilvURnxnIcdk
MKONlixa3tIq0MTuV68G4vBWRp33cSTq3g7UXci5vME5wL6nfSEvmhS5rdVQ/Ykd
pl6GIn+C3DUpmJmNAexteSFI0445U7I/a4knJJOd/VmAYxfQBfG4axxfNkbnnn5M
y8BiVL3GjrL37X/i2odkMb41zAZuduYgCsAyJMcZPajVkjmHNuMrVoXfundZTziU
KV4O1mYYFmUV5Yo6AmTtU0OlwFFc2j8kofaBDWiOyWOnI+Fqo/wNdPRqXkDIMwch
X7cle7CcKv+NwBEwUEIqUBehbuuUZMUfLYIF0OQPbQ4xVdYjYAF8GmEwvpZGkzFx
hxtw2m+vkWwpGuvYR653Iw0IXtTkD9zNutFGHmEBiBx+7NyHar9wMxBBK8hp28p4
u9AR0ZxJUSIdJcljibTJqIVyqKBfnFwbSRCqK3ForVOpl1LR6eWAoMVr5/SxHP1l
sL7qVe7lmsldvjEWNSm0J8oQI2v2pLG/C1dnOzZmpb1Fvp7lOMH51UtzDwGwdRgC
gaDdVcSRT15Sr7/HMofgIpBjTaQiC5puVDlLXH7bXTVtSWQCcU68Yx+K/0BdzMMX
fyeYm6zc/oLFhrIFZFnNy24I5K2TVQfPB7v4HK/lON8i5FS779FbY77xMLDwVQVB
w/+WeFBp/3+vq2ktOX0SU6tub5QHT+fn2LiaXWSSAhGrVcJ4E1kGCIXlI7amI9rr
TmECxkfMQ2kE961dzqCwzlICV9fdoZo1gfejszsQwzOW29ZEK46ugoPaOjXdH5HD
QHI92Bjh6aABbrztuSkK3bombzQzhs1OnWhZ8Sljph+EeR+46ekHy9vtEwhxC/kP
DgaNGoh/sRpYKxdrYFgu0sKENgWVXBz9Z41+j6g11DJ+q2WMN/QV4HKiFY1nf9tO
PEgi2OwjzwrnH/o4DD7BPM1Exrpxrv7RSobk7Z1l8ZkrH99l9QaGXDA7Afz0rvfP
FeVv6hYSbYxY4UfwG/OfvyJGdSBm/2LU3uiTzU2Sv+Krh7WBSvgCXJ0pOAIIu5Ii
JB/NdYmYGzRmX+sb3GLNsa3/EYfxvu/vo7AoaVCrg7zvS2fi7QdIrm0S23HF2cg3
XrY50iBCb+8elkCocWEnYqKDFCaOfH9o4l9Sd1uEQli0pLQifK92Lyp5I/O0OytK
LA3YCYBDDiSsMEb2VDIDTMrenuW6+YHcKW57qZVZs/7D3FJIxYwJm4eECwoOvBTN
btmjqD1EmhIGhd+2CiDmokB26NPU7tJftq77KpIoAcuqBb/m411uk4pl/MWHARgY
9VoXXzaxXdrU4lBIWtixUzJet9nec/YKEPU6FcyJOz/Tveg5kLHWOOGWu2uZzBpS
BICanW4LSMbngknOBEovfot0XzOTJ5+DVTcUvYAq8AjIqjghM/bnIFKlz7sTNnlw
zT4JgHrA/EJ78e2lFECOUkAwyyPqSKURXFAWOE5V1bpRA8DZXqHtjjEg9bfTJV7d
+HKQldSgLfyqZmo+WTbFlcFw5dkrXftNcYjoEIFHlGK5/x0yS5UAblsPilSTOiVw
6Y/OONfJdt7cCi+TWlXUfbX3a+3WRRnw/fvfyel+SObPzCSGpKcNSG+uutIVIAR7
MKV3ucD7L3s25QUmOJwFcaGtkns94OayE3acmV02V9R6eE47qeYIytWIlKvLnQGb
/o97u9TEl0HCZ/yLkllyw/Y6TiVHSVAHmuqFzUSOrh1cqvbGJLU8F0XCvxeeK0Hz
fg4bctwbc6m96oSgeevAhW4wk0/EGnyTAyDiG44zUrE8UdIYoewGAGBKs9+Nmn/q
w+2C6Ofiz0TmlpttWGK1xDo2InolvvYMI0Tw8bWjWhyNQU+AllBFWPh5B7mMUzzV
mMxmULxtlyza+IkCTMQ+FMgjIqRZW76tFj05mQb67hB71JWKPH9+YWsCx/Dl7sMQ
qvsSWfE4wLHzIgymV3LkZxtHztyPzfrI8cvq1MEl+B7W0UqIXBwvBautVoqNCCcw
5lca4fU6MmXx20tNGjiyJu7Eh2v0UATIX+NQOkVcFj7/OsVzf5etc8omd1fOShuY
Ju7A5sbvSmP+whEGdymIXHSIvgh1NDicP0+0yk//D6h5ACdNIGvoG9kqbF+T34xb
cTvGVrH5sfGnWK+1RqhEg24hBmQR7bgnyze8CyVxtlsPowRGS/4s25HBBaQJkHRj
y72vN/6jnDDeB4Poy+ptf4Vk1QwrcVjozi8VtzR7uS3KNm9V5DwaK9UDNZOFPh7k
Ai6JOcp+ZZ2XPXaSumU4W9ATL0i7j1jqCGzESU/Isyeqcy0RZj92jn93o4rQ5VIE
nh9XC9Em/DTJ44D05pAv21MmXJ2T/TWw0UcUaaknWyttYrgMkFtAX9SeJzr1BBJh
ukNVmh59WKSJNB7KqJz1sHYZUY+JiQNFiHWHO0Wt1h3BiIs1qubwX5SvScbaAjJb
mCPyBhJ7+KP0tFQ6PJ982rDzjonrp8j4R9FIdkPuhiB1VfWPzrgQJ9P0mooC0BsQ
CDEX5gaS0bxMQuw3rBiHp3PwVwZi+Xw6xYDIrghzcqvBJikNrSAYflJD3+aKJ411
gr0A+B5FckLuhc8H6YeIChkf9Wzdu1wvMpo23wa+PypwrSmx3QSWnvMz+prXTlgV
kpLgDBD21OeAVsWZMz8JKyBK+4qmVNmJO2YS5l0STTsJ6BhpwVx6cjWJiW6/xN2t
B8DxuHpyagwleTrg19lfPxjOKe/1zUfMZLa0HL2KZPZ9vU/8mN1tiNy6vf6y0OT2
U5xMK3KFDRbOX+kaxecbC/2cpN8va8H8JMp1dYGj3Zes2NjvSEJldYTSpkVOvnBx
1AjpOV0fesTI/9cWChQUvv7BdVA+Bg57s6+aAPof/TbtAU1VrX/9l7nAv7CZL7a2
Cj8pGAq4e6asHg2sYHE6hhlTMhtk498mz9m1/p8hcuu1EFPPrqtOMmmEZFIKsduu
fCBFMKEasd1poirGB+0l9Dr2ClxHsZz0SdR/WkpYlv2XVJYSAmPTePG/DO43Etf+
vxV4gN7UEtDKuWTLyERm683cBnRUcC87a06grETHji/kGgPPDT8eBs+LYIt8AEMS
H9FpByFBERWSDvGoV984bOezkR3W0ZtO30Q7nbC7EBDolRmY0RZJWNwxfXpS0tut
Vy018UUoXdTZh0Ql2flYOWF20yypdsQdsPY/n+vNyXZZvS3MgL2M40Hrwb8HRx6a
joR0GGfmycG2mVfGuxjkW7otgRrOyLoe+PPjdODSbCzG7QyEy0D5JL89Of6Amk7u
HE/cpW5WeE2UlZOfXXO/09W3U8oojRV1oDrrGMhy3EQUx/gPKRS0nKLJjhNWIXsO
2z9CRVnPs0KuibPqK39HTpiWxOFVAA1Lb59xa1LggftffQxKPUvHyp75HFByCIbn
+VOw7NuIsiiTCEhR2ghe+DhBiflRLFBsBfWVPWz8GV7fGVRdnBybajsVN8KdI3x4
Ga13AmtEUEfrqP+7K5xxy5FlMsVU77IATJ5Ypgs3G6S2ozTIdbsgZxAbXoaUewIj
o3gAtNky1ImTimtaQ8pK3Uhcgv4IkYEkZfH1V4PUUjvVexQfpVMvjgcyoIX9EoVg
57HTvfy7IwNSgxnxeEnovlcgItXlfbx/cP/YjCgSY47THUTMXhGUY5j21Fj2CPvb
T0oKG3Ju1Bs/c70Uqg6284PaIf3wDmGCJs8JB1V0CQsIMntaK5kRsH9mmh5+8Bzy
E1QSDuHDiRJ0LuYNgWiZHNx633hLI+fuG5WJfRiGl4ZOLLgD+wys/13sBC0GnOlH
yECchnFHMFPvt8JhAaoV/k4baoWX5UuKpgUhAB/N7EC81THDy7TpxhXNBVNttZCA
QRORMe+2XpHHyUEz2995hcO+6i97egFk9JGczFCdB1GfhA9XirJP6QEW5CsG3B3d
mBF2/EoEqyneaEsyFPtOde32hC/2Y4cRCLIPmiMyTx08ZfBM6Ik0VKcFdNb65VLc
FsRWrHCuOyjauRZ3WfUnBhVqqWsswoZBU+jhQLRUuPjsIUq/ygfWpWiaVRxq48Hl
ujq12pKEynngqA4p2X5BVGj8WUEK8kEi88ZZ6uCJPjCrsKLxC4Fm65BY4VKIr+kW
tvr/qZImo6V3EwnSUXZnu036BdLh8e+IO5/jsrrrrjlJxq/lVt2eLhP2x/hUhiFm
Dckqka5TVdsuIb5Sn6eidd9GgI+e8ChKnTBAudTK13xfGG6iu2dV0L0dOkc6pIjr
WYbh+NCxh81zJO68/SMj5pr5SGD+0Lje8dPy78k+KRD9k5pG74pEdsFYSOt18AEI
NPeOt709035noWkqD+JUqDK40Y8Ofr8BUAjYiClRwyr86B6C7t364f8GMtsLDjSD
YBEf8uwOdEKkUTEe2OZ0F437nlQz1AVuz/h2Odsmz2NSSu1wxomkmQA5kuxCuzqK
RHBhxGN9MSl2sIswa5nVZzKv0h2VKj6P4vIdIFWrQRmj5uvlcEaeheeiW48y+oT0
yJvELHW9BVVlNlgLVZVq9eQ0qZ1RhU72QRZClcDq8ZytGpf0X9NtmF5ZNLrCPVL3
UjWh2IWg467uPqauxKn4MgKCa5EekKUV7j7dcV5sRS0ga4Zkgyc7VGAIEcE5iyTa
mEvVCfbhAOgZ9bLUcnE0r40TqOXYZ2lGbbM4eiTzIclTNG8thHuANvZ84Xxl/VCy
6UMy2IDAID5ldZV/UHgcNiE8vebLzvZ6zJKPSJFdBpIycGbZvfGE9jKL7zGWFfZQ
1l/TRRa/rfujVXLrGt4eDDuryqg3dN3qWYXFwegJoKn6yC+fudxAiqL6sIihAKXG
Hy0nYsQ5p0w2Er4V3cIDR/yi5rOo9wWesdYfWzwrCeKrtwSkkL38YL6XHPvwHi/T
Q/ShlOBc5ksW/XcrNTfMA23hcEb2vNcztkorxPphc9Zy8HD4c3kjSU2UQrmrDqo5
sn/HT9U1zaXP+EcUFv0do4VJHZJWWAb8Na3xDRVwtmChDRrlHUVU1S7qbCHn7Jp5
Y2qQxBi8Gv46NZ8hDEzlLetEXgYJLe+AEOp0QbyA/BFirzQ4weLTPSBnPAACB3zv
kPAq8GbQhsjmVDoCmik/Pi4PvvLXULxUJcwrVSpcro6ho7LwIgUUR95IghNLBvsI
33IXz6JUD6drH376hVDqwbo2c99y2ic2HspofrDG+IChORpZlLqGdDNTtp2aZDEe
La9eY9pT+Xe5JRCHx2hVkkdRsEqreiX3/py2TyU0gIF1kDvwO6T1iM0mdvtU4cTl
uRQncff04hXjtnOJWDEB3TrvMKjocAVgRWsuVgopY1G3NveFkfOUzjSWdalxoN5Y
ztTouPbzuegrE3kaL0WRVB6rl4QLhDItNsHY+MRQ0EINDl7aWtgbGxi0n083atti
OuKxeNzDYMOr35pAA8uscLxrMmjxRc628b1lGlWIp1FKjl5nbjBEa8gftmyCRGT8
G0b3Wj6/SDn3OQ72AdSw4fREY5eusPyxrRYbS4b52YwGxHj9Sf5stfN7sX5j4PL+
N1IU+mru7NfmArrfVCdwo9av1mU8qj8CGwP7rWRmWAoKwLnPEQUZWxyGWuAr3XQV
vx1WbvUIj2YYSr23/BITjzdBWDBAvSfUlDFYjWySK7Bz00WQTixw4nsIRhDk0dun
tI+onGDAs0+UQASWOv+ETm2W9sE3MfY5tvyAYdyhsTx/Qhv0dKmQZ96mFzqqL44X
y0DlY24Qg4njdzQRaOppp8Fs7X/ABW5ha6POHoiNYSARX8wn0oKziMzz3m4k9qm7
Oyes7oU59vSbW02eBgxH9sNJiQqQeu5OTeFpyr4q6aLRtpkmAQGUPieLpkW9WfaN
ZYjPQcegClg1xiqZIwVjultRktEcNvpHv8Ii7pZs/kmLDxB2V0VtI75zgXcVr4I1
mU4ON5YbYuSA5gZybmvCDSOa5BEuUzsmaLBLoRC4RDopmyOBeN8JPLoi4QAUd1DY
b60g8V2nzJ1laCBScJMrCKHP8aCEEirXU793FvfB5XdS9NFIFABYj7IQH2E3k0cy
VHfPB7eT6pk/YI9U37Hc/MMwDjmqeoZxZVZTH7Cd0XKynmD8KU8TelAl0hy1QoYR
FNu7yr2io8Zjm9qR+KhOTtPny+jowQIxh74Ag31OpcLhOHsmQRFmSuWHsZ3XJuRx
Mw/2Ak9XBwT4x4VSBI+cBvcR0N5+yJdaKY3dijt2wCbL09mVRamyp/M3fwpf/BBh
h24fqfIAF8w3tOg6sryYYOeyhmYQjvjlrgkyzAaYt7nB6ZwvIKXxNVZgDwQWvQIr
mut4DB56iADX8SGkTAfcnIvTrdSKOTSjlC0fimZYg/e0k5/cdKaE19pE3taNYTOE
NPMyaildOwhWI6IM3zY79uPDSKEG3Fx056nV9ouEhsaBiP94lsBpmtROnjwB0Znw
3ihy4BpTvXa5j6nJTwNugiky1bRd4xOdUqB7VSevdBTrBjswh5wBR4MVsBkfkXs0
ZOSxVqsuPX6fADBJ5avJgMLU3bi8UWvrWsL5P94BxElmXqseYPHgGG25sjYjtav0
4J87og8GJJjg+F7KJCwxTggo8Q4/2n0MNLzdXnAAQpx1V4vjUTvT5KQUsiwWsqXS
KYI3bXfSuxCbnxdIaBGplLQ12NdPCRF86Ya6uBhZJ3ffBSStLx7U6FQfy68YwO5B
uRqxmENAqh/Q9Go43cbeNq4UmEZtvTX9vMM9etuUctBWQjlDkeKCkQemsZK/8/8Y
XCbi4pzUL3gRyNnAKm8xAehAPYTwHfAwH3naknPtrz4TZnPAk1EDEtYTHjvtLJb/
PVUos1nVnl+8MlgatewF+mCvyiuPVV9DwSuDTOvkGol3HTCw7noSPopExbzWMyJO
jgjc5QuTyqYJMjPHUy/3ZXb4pXwFPuPkmWMGxsFkZNRqCoWSUllg9DQwixsn5uEn
hF73RFOz27pmCxEps+S3vrplLtB+iaDXzUXwMHkzXJ9Wzxr1ONxNHJg4MqbHvTkJ
G9WihX0pdv8Y/bArF+b9eh+HQG9dEQb7Z2Vc3wMJCeyqJA85dWWc2/FUu4We256C
TeToF0DLgPpnC+X5ny1RkccLQp+jBZbq9oiZQJgSO82x+NFzj1Vi+uonEMtZ6pz6
ofr+d1zk3n4PnpPK707ZXh66zysV3bCw46UVxKmbt1T98DDLa6SjKD/rH4CrQZoK
onj7KZHsTkq7aRXkUnKRo9LAV3UjPQxM/KmjZk8vjonb5iBouMBzntwmTiBsGiEk
vkgBP2JFQqEkElupOyqHV367hzXJ0yxx4ZqVDWa0S+kfmGh67YvhUvpW5DU89ZQw
sH7gZXM8PPYONr8Jv/NIa7hJY8yxUWW32l6mKM+UX+VjYLwzRDfsikHNHpctZ67V
VmbhPptHP8Wjkid1MMEWnIuseuKVQLEgaYIVbXWsk5tW53Ru73MyvzDsu5Gp+UqG
SE/21oPKSQ79103z5fKWGtcNdwnvc6wIxcGiW7bMN2tugftHXW8mDgsZnF2tLC60
5WtnwpBrC0F1HgHlxCW5a0HNSjJvGNYXmjTyOf+FZ+rTipuUqtYmIjwH83MXEzu7
LKf0dVqG/bgCE+Fv9tA18LC6LKhBo0HRzcQyPsH9O/5ASOym+zBBMVUjwItSXCTE
JGJTeyIQDawAR1TQCpu2Z8doAr1/mDi7vTMzrhPi+JNDjHghync10ByvBcccdYUO
KmoI8t9Tlw9bbBfHgBP+7I8oVgp6p3YyFe3e/q668P7cEb15aEBiOhRE9pXzzt2m
fjjHaZGLuzJaQgKLG0hDmAkG/1WsQ+u5FWQoYSsCL+Np+WKU3EVDCJmFBBYqpmuN
icA0h6wbWUvQTvM65aWw0Qw4ASHaZAd6ODCGY3PJgfEUyktlcAIDHbbiAKpFV5eZ
JLrb31m3j+RXJFQLfkQhTp/SahkaPzRH1tcON4YJX3XFBJtitJmHISZkZkJxYyFW
F59AOIOWEuda5CjcVEkJIIo/HXIHwGoPQYZ7+hjnxKUT0GqIiMmcIPBF05WFiDk7
ugzBPb6Ee6u6V7qawz5PqPhTblNIK7L7zblv2vOrqRSx9V5BjPtajct3J7jHGBcI
xeXT4lmTYOo6SDrinMDq8w+GCVSR3r0ZAV3OhmQ6PTthHeFfLABCYSEX8/yRNz3/
z4OkqDpE14xINuQ39Sd2VI4a/eAy670Jg9nedqwKEdp+UYrKH9cXpqnxzRKLuOha
VUSFEcOQlp67JCS7sohp3mNeMUpZLtJJF7sJfi2kIOJ09SGiJrIu/hcbmSE+LMls
tzTWbQCotuV8lD3tux0YQzl23oWmuHSgQhoPhw3wbyxhosn7TS4q5p65gH7EfC+M
Dx54cVC4s2OhDRk+3VwaeeDpQ1BEwmv+OO9waNYZv1sjYKqLuoEuag+Qpf9vAmaw
U4LCys2zrl2uLf0+4I18dPDP6fATFYvWy/Tq0r+t/EZlXGmA3THDaGUqPfHtnL+u
cfJW8vCx0/b10pokOtYcPr/YAYMFS0EStJgEPHjf3tC5BXBXki/CqHIVIP4h7BS0
+OQ7jweYyDaLSjpyZlUMqDqhQIY4IZ0Ck5SL2rqCcreC0aVMaz89xeX23viuR8FT
L3Dvbk0FLJ0bAP+BEl1jGAudsqWkxudbxLNN89TosVyZjedDKawb52s5x7F4EYEL
+XbyfMPNUEeE5mbhtnyk1BeIb1mn5v64EFXmhajDdwoQbNHx89plvJCyk9X1MWuf
PpDc2IagezG5e68fGMd4FVYL2D7NvdJWk6nDSoa30iCHc4btpD1ggV/zVqHfKbHw
IeBU+0vLFs4vuf/ZNlxGTrkbqGQy28mjocmt9hNGZXyqpkXTE3WPCqkk038YNW2G
6mhL8Vt04qbWrUYPaySDyzGH5t61uhnp6+iGFhx+LjZ+Cz8CEW87KGJgsQBmpLsm
bPIyBWEMlYd4ZoN2w3IW4KJ3KCsKzKjGMiQBGNHOZRWtDlj1EOdoZ/1Co0tc5560
Euzg0FFHbUFaIkdxtwOANJG2Gkj/SyttqFDul8j8eJXRYaoVOzhELTwdTNuFIwn0
RND7Xy1RU9GKKq4gjfOKEDt+SkB//PxVXrlYWJEHiPyIoGYSUlaGBzxyryOOCcPs
2ILpajDt2ARKJfSD4yo1YakALx5yfLXh5hSpL0YguBxKf8GgkMyJxj9eavGjheTS
ANRM4YChK2ugSJzpG1CwEjQ0JlML+JPa2uBGJ9bE7rMk74SEAeo2nk4SjQlHJlRD
i3XPsauz9B2hm1hs/BzeOb53vCWdOi9f9IkU33UvcJnne97KmECF+IR1kqFv2DSf
40o/L/bbYQlfa1NQbzTbN+2MDho6Tt3g5ZLi1rbmw0lqqWpFWrcJb64kaFL6zhem
Ku88QMfpl7CLj1gNb8Dm0MFhvoFbJvGbuhXSDBUgZkzXSx8o/4ZBF3THeG03A3C6
tiLp3SgH2z5kYV/+XSOareNRIZgsyLze5ezW4otiX8en/9IHyMmjasIyqRX0eTt4
tbwzCj+M+V2xZzD4P0D6oZnaK33Dp1Q0t8hhBdiPxFDXdkt+n1fcjP/m/o39LfaO
cX1cbMjVFgpHrsRxp7Xyx0F5ldUUNgGV31YAErFoEekshP1rhsO+xi4WpuscEC/M
yZsM4Declq7rm/KdxZm+150tt3UsCqiVsFoOIThIhQWYzFcBbJMW0aabAipmMKvb
OuKUg9VZJfMWrd586BAUvfRjcI5K1PCSwxjO1bsFr9VD3ZCv/3MOy8JwNvdllwex
kzexBpQhL/L9uAj5Q66IWc3fgPGbegz/z8FHXLMvziwcYuLWazwTLh+/QwNg93MC
bp7HhEaknki3DvFirS2V3GbYkjaFby3z2+Hq+OVkPjwfDDmhapb51Pq/x728T60o
HWCphl3cjAek6zGdiP1jaf9n/cXkkDNVknT16E59xiuI5945Dj6GzOb+2PKpQtEh
VCTcdaBseMkbJ9n5EvF6Dax3sr1FNQYnYdy8R/m/rtL+MwLS2MJIlM47q/KW5RLk
3iomjKCMiaOwanl1BESZZDxB4KtGOI2J+t1oyiW6+GpG4vrw8P3pwB9TDJThNR09
LTpxnPwhlGySl4iCdFcUAqoWBRCauqdyWRCWHI2hC7SWD4ueryXDpqe+KDcyilCG
2k990B1a0QH8nLrKSkKY4DKiVO8TythKdD3hSG4W1zZG+TVilVNl1LW1CveEgW+7
DeIwaM8oservW3JQPenPoK6a37ofYGfqnZF5nm3zooymR4xn07h4bKYw5/6m1h3i
xHPeo4+nuenbMYi54j+0Ol5tOoZ19i3X9XlNQKcwiRVIC5bDB0roN2M7bv1MxEK/
N1DJge6HFtAP1Ki9f3p3gU7mTEurTfxXQFk0Zaf2jqQlu6x8DnOBz6KqEu99xBou
Tvlb4xgIcOO6Bj5w4s0ImylfiYYkUN1OvYBeRdyO2jPKAdvk5wT30jw3JAWvyinf
rnvHBceCmBOanX8PfUK1uglSQJQi9U9aen9WPiiPCl4fPj8kVCR30McVX/8Z9Rfz
tKAZyl6jwRN+Df9RN35RC3jyztaVRwyd9JXgTjzrcf3sHxLRMH64vXfbvxNEcE1X
6HjFvIRWrMV0sAVkF+EDrRUog8kUVWBsHqn6WutZFHEwif7TdiBG1KZMufZUKPU5
SYtl320VhXze+IxOIPekoX507G57PjSTkCg7FWS4TiCyIHg2rqoJ/pk4D4mLcw4H
q1X8JrmqZn5UtYScHQCzMqW1BEYb5f4VKcnhMo6ZuFrIfrjmnkasks+RNvONmone
WI423VhzUBEEk4NLmDN/2H3gzo7Xd8lmHGR4Z22YQokmllMwsvO+lw5WOndWPdNc
kmJ38Cy3uCQuz6dfAp57e/75mpWwpoootJNv6PD13qGIrdUMQyHvlCqaOCTGOLY/
KVa3adfc2zfetiFEHJBU73B1eYmUIW09hrrFH8bpK/MhqtchzrUVahxIICB1bCQJ
Qdh4dSSapniLGM3Gw8bzjUlpN+41yGmdRy9yLi+Z4zfQZVJPMBeGBAuyYg9eK+Td
YtGqqAbXpvVcmUxmRCfRJSAJJIfn5z4xIGG3qapkIG1WQTrmd2/5s6jdPi5tUhJB
mbqvqesEuxKlb4XLY5gE35xwvuzGCjaz/2c3ph7PPtcukw1njCTpb7PrXcHQrXv6
QTV8QRCMo8rfYi8t53NKzsjSJ5vWpSHeNltM4BobQ81S0R6Wr5GZu7yrSjoCW9YP
sRwe34XgGbNScRpqWy0Vx7WkjjzEUhqfDG67wnE5W82z4M7Yi19982T2UY1Elmyx
5apfBhgoLuU4h32p3/Q3IGT6MGA2sUs7a8cHk3avm1J/FIz/h64qeYm0mAdP5n8q
ZmToqQ2pl0xbMOmkwv9MNW+8HXvTbG6ea0Wi1dKHn6OUCyy7ucfHqYys9eGg9xOm
lE+qK3Wbe2lz5tZCzXBlcDZ2+AeU/GIcz+LZVdzrrAf+ufC/DzLkNj+MvenhbLou
ME5qweag2zqjvRGSsAa/LitUMQp32no5DHlYn/crRek+470xoSM7v50i95cQ87//
e2seUrTj6DoYxP4FLur96BFemIF0/SBIiNYGyPtmmVxgsLOyJZPvgo3jfQ/G1QMA
GUZbSuE/78qR5AyTzA1kgjD6NjzfoziRmyfQIDQO1l/0xOLwTa/vEPItE0TXFS1D
02/RIQ5SopuC/qyB642vpqe8nsP+i7OMJOuE3kvMEz0rqdxTWrQkLgCkEhl/bN6R
DdVQ9bYuUEySWoSfjCsF7vX17cJ5ck8USBN1uPct67n08nqwlZ/Slr/x5B/kKDGp
o/cVU6BpUayV/+FM8TdRrz1tO41/1R7ou/9k/LzPw5OPDAXtwFHRFWC+TGov/Vd8
dsFmxhMh2u4H4r015L0ZuBzidwD4l0nEOb4F++v+LV6OBhl55cZ+JXun/LnvkJDk
ZUaLBYBPpGwrAJzBH5A0Fkve1ECtLKYbv0p/p10ZUMlaDJPiGMzkR8GcpJcAOoVn
14lji75RsNPybrK0KhcBpKloeX66AAbgmmKWzjliwMyNE4aXZLtS2zBgBU26zx6J
KpJvyIMEWcGmaX8Y+XfTYAV8gb/72Ljakii55zI1Nz7uXFDzzxJGwBdAJ9bsxqOu
g5GEeDuz32wrs3lS1CQ8yadQNU5ArIyXSqp1bpLr3+Wb4ZmxF10fDeQq+Tuz48hN
TbuQKXf/qQtv7zVigTa4Gog1WkfwjeVq1UbU4bH8F21bh0PH4jcVs+bhOrgO/GOt
h232BcP+/KgtaaEASw2kyRrwoXSdH8ns6Ikoucz5dF89Hz00EjdtyIHJL5g3QamG
Y+uD818lYTIWKVVDauOh4JOJocmI1kt4Dkfm/UBJ35IcSLMMH9EHA7xaKNwp6UNk
R3ifa01aHws1yHgjSr2fznkVyfQK7lYzvuFXvsBmmJgs+BqGC3+A7luRI4qRaBVd
V4XzWmSC+N54tEu1JXzTnxrYiHd58505iDV4BgFXfRRNZoi9eTCK4z8hhwbO9JEM
jIInoiP1KzGYUhoEtFRy/2qyhu2DS14Rpa9YbTXbE36Q5902hhTk9mCh3YmpzW4D
5yKYJCNZOPn+fxoP8LD7BQJ21g9+eVik9Hu2O9J6fnQ0O0Zb9nIxJC5ZUWNPo90F
Z3ayWo7S/zqjy+ROx7M3ojjFPvFod2U1N6lqssr3lK+zjaoRMbehB704wAga7Gi/
joQZ/Fzf/cB8c3ND/iAex9DcTL53UDnwcVvewZUKtIBri/KVBFUArMT13DuIUU81
5KEbmt0GAU96q0JtyaV5Uu+RVWHlsxlfNiSwBPs+wcI4POmrU7P5AEjPKRNM84Qm
IqC2bCZ+/MtC5Ac8JJFczD85btGN2w2+wvOdDDI9yhP8Y+M9CgAO9py7Av/+7LPW
xNBwW2WwmAjZMgjSsH2VbDxWxf5xGGQEzAGR3FmeFYeymlBpVzeY72+XrFGqZmty
7M0G9yuTAsXn3ZSkDYuoPvNESl+/nmdR78KjwYEzH8ck4HonLsvt/94enOIFXY/s
G6dkYfkPYSeCvyrCzky/TDHRBmRkzbGCuN/qqOkbLYRLwUP471XNUlhw49V4Qp9Z
edxnpdHsyGIRmmnUVMAzxKgcPke7jJLB93MRnpT/5ppFnmCR6tW7fFeERQ4h4hpb
Yf5IpyTewqy/QPaKng/AYwm9QJgMqEJU+ClcH2xykv06rTm9HCuauTso6ISHR0C8
dM+Iv3n294sUcjdpbcIBfWB0IGDo0ZgSw4t35iZYyKV3KUeaNM5wAIs0QKn0ol9n
EMn8hYnzw3cvpf5NRkA1wtACPNE+nJLvsBk9F8NIF7Ujt0DApdBi6qXbsuUJCKSG
4Gp+160BRstB2MYnFZVmaAnPFHQ70uOW2+9EcdI0YfloHLEJMZGz9uIqjZeQmu1y
OkQ1lTzLOZekyp4HnRO/alxArPIKvHPaaF78RyAtOZb84qcJC9ayvvlBN7A6Ge46
e4nQGL6tNCuxcL6FfuoKNcHkcCYp63MtewQzLw8t+B/T7kXopc3Ei8dMdDYHqO7v
HH5aQhUjmwdoMUWFYX0BB7w0lZnFjlWt0lLN1doUK5Ncne7QEEdG8LheguKLVsWS
RVKlKHCTKid/ET1FIVup/Z0Y7cYrTrzZks7MS6JD3Z3xwmkbDJeVqXKTbp7n+kTC
HUDnKzJBoV3wB+3dK04U+yQjRWmcGdj9P5Ej0X1TfkWhZCMHOwQF91erF2UKpzzR
S21BxBnzh0Wn3uNxbvsmnCOBNaNGCciE3odZEA6BgcaEotTifM+Hb5CrvsKOYWvX
VsMASPrWRYeEN8mRmNx284Udx+vsmkQ/6ZcJMXLjw6JdXOpw4QH3jcAIBRS5ldmA
JpxJC3A5tdvFVpB9PdXDqlTTqgDJEXL8YdOlMtB0PconLH+PyjgtsUXapVpCy2tU
OGaxsWSBcAAP8hpTJgpZwRmwHAcKJ+Jg6XqKsU0kYSXjlqZeaK2Ql/HOpfz9KMS4
IaUpM1oHZN7kgRdzh4WTGztMjfAmk22eD1ucTWs15iWLWemRFAF/v8EuN/jT9Wst
9hmV1vNU/xqWHCdx/fh62lqC906sOr/77n15Wgpxj4iZ+EZfpXiWLcnTKnwIR3yv
ObYGsim760+q38p0jjLG56UBKj6B9lLPAFL4WZVqOCi7AhbzDEDCMSSEGMMikZEk
iV0nnd21zisn/P2Al+sYpTln1TXB0qn3Fi3U4llna7SYAHBGzVHewfizXNlC50ZM
DjNzKxtcC1r6P6/IHXUknVtdQuk0gEIyPtaFTtK84T2uqRWn1kIv21JYJIPGx6z/
hW5faiMoIj1ZbkNOhpKlBWUzPMMBEoszx8E2CBEQGv/YPzpYiJA/LmjYBMseUveB
xPqMcK7yUNSBKfJlYeGBt4nYgG6g5IIyXA6vlVp3DEumfIE/D2jBf2BUp0qQYfuw
hCT1Zux8NN9hHkMbhf3l+KCDtx0/wNJP+xnEqvEJi4hfjQj0aNsXvoQXgqLt7FgC
bvVPc/Ss50H5y0ZB/KArFNxIHy8Q3YxAxe6BCB0ySwhWb6UPQtbORYlj8ZZTncrQ
iRWKeEwEQTDyybC7Tg1nNBl0egfwB/5vLkc5YUw5E+za5ElYQJERfinQYmrnuDJY
arD+Qxt4hI/RVqfm8VSmmA118nQpxkM7auo0PJFJU+RAsqbNfhEw+D/dGvuOITuv
4GgpBwAeEaPgQdwTBJBSf4rf8tJ4Q6l1+hDvymPuRV0H103Gzsv/01lpAi5sph2R
8judDNjBgNZ7CNu9pT80l9Bny24kNczz7JfpRyeCSL43Ylev/cz1JV7W1JwBWhVZ
pmHd/Nz/gUl2YGnl9QYjeXy9yTTAlMUrLjMgtbyKL8X+GVUfEB4rOlijbDTwcoWf
hj7r+8YJxngZF1F/qAQBCijC0SW+c4Kqf0HhZX4cy6NVcdTWzcHOy1oXkgRP/m5T
FJJ+badquO8trsCEbZLNSP8HYCq27/B+gpof72GyjjOK3CoYvA+w4haNXXB1d9BC
zzPOBt7nVS4LZBmzTc9PjGGDBJGTF7JCYXErfh1bblhRSRxvNvW1hkaBbLgOEw4g
joKUz0d8o875YUyEnh0Llvq8VQuCQO0UbM0hX84v8QcQB7Mv5y+dCYCO7TcOtpzu
E4A6eqklAVzHsDPV4rdBUdd+aLTeHkB0SwMS4xMlAWkd9TPRtyxaT+HQX7Xp5kPk
CMladHJ9164Rq2qC74IDaL8BXEhL6ACyaVB/ujzqnirsJ+mJ/GHtrVy6m/MzeLo2
YxVt3pJm6zXUBTUcqY8UtGLq+0MZ0ClHW2dH3n7VC0qiDh0tAjhsTvLQLa9EH/GF
UrdpTj58raG377hLe5VRydQUcpDvkx3rJ0+oY0+vGc/PTxB5TThUEfq/GS2hgJdC
sEDFZecA1dPP5p9GssQzhPjdfDLwRXO/iZtM3tXliRBVVaUtwojKE7cps2qVBXvU
N/063NHCBdjsieuLLVvVvnOwOpnvI5AgXeUEu9n9Ha5R6hgt9yCdpzB41KKW1BK/
OEgGpkGT0jMo+VPawlVzBLU80NPicGSqoNYhkGrNjmjUt9BWnYZbk8qqAzIkdQUJ
fLjxcTd0XkW4j/4h4/q+Vbj6m5bINYobEOjh6KaMKq0htQiNxH3d5zzHvj9H9I25
x9ZNoufYX7S9sRupGYS09NC9YI/r39kY+Uxla4XODAGCxJ3LD0MVkRKtxvX9yfLx
dc7DSO4JqQqP+8FrqGXXW/8yI6HlKjRHT4tt1rj7ZP7M3e+eFkmZzOl8JeaoKGT2
PZyFfsPaWhGpTXMiJDweQI6YMFzp45oUP1pqydNEkVgOO6/aolHU7uKxlzMaPv4k
Rvlu3Dc8mAyNfgvdO1yjdXo+vwRxehq3DsoLjs4Z88rtmN/yBS3h8WmAeMB4fDOz
WKXqHR0oYcVyAb5HLhmdlG8+83+PoixXvYTkuhXuDQhXsA5yoKkt2zsNBdWXn08R
wVcjryYBXIUA3+UY7RX05JgfXkV65HF2ZgeX0Hc39OnWXHeQD7eQL5IfGD2bJG2+
dDHZbI109AlaZr200OwuroCiea2vPui9EWOgTQWP2b7QP3IQQfpXGGzul2scCU+/
I9jkK1nHedi4biOFWAXg0F0L00bIFgs1Zeh7QqpzV5YZlSa0zUD/tDY02u+i3+SM
7MpMx+O4+PfuHuh5Qlr6feovbTIeuBfAT3z+JQPR7F4UMJ1xrT85nQyS6czgCYrf
hlwmks7OkRVxbBGbO997UUOcyDFrX6S+xLNfsunvW1XiY5Y9y3VPFz7y0LQgIiv+
+lpxoy6AlfSeZufU8jvUdQWhf6tgg70FoQRGKkfEJNKAUbwqYuv6YmhUT2Sr2khF
eRAGJaMeMo1ytYHtFmg9stBr7d7k33Y7CS4CcqCTK0HE989AJZY+Po7zhxizQz2B
tOVH96AxXGyvylCNjZvB1ZTi9Ai+XxAOu3fTFaDrZCg8pFxXx6eZIZyFaP+oEhWS
xM43OTLxaCqidh5Lcw1mamW/ER3WO811hoqFJIEjmgI4qp69tmc1TJinop/FjJGZ
b9IaBn+Q6H+LaY1QznkWZvrLraPq9auVp6dx5qNyTkZECygFsgUstt2W4Nemuk2p
pRD9+YIMEBiSGlpyIS5uY6p511eSZD4BhtD9OECDOs9idi4JjGbZRC5lzgWNMDLh
IbAMewbpCjVKw1JBxWTbzKyVxWo6NfAUvSUFk8FOGehu8DmlhEwY52pnecQE5wR5
sowdz1sglUsJ5VNC3oRkiebtj+2NI4E1bjmQ8iaih5X+LPsVlXZiq7gL3UweZkh4
6sU6QkTfLu3IrDVrnD11LzhuSkFo0jDyGmdfWvW4ljhgOOyp6YdNlFjEBW3PutLZ
Y6+/ddiOFxhSFJQhuTOWJPCL364A1Nw2PDLmGT3iuY01uOYhIcpu4Sr0arpQv273
1+HOxBaHObF7lSpqtuv6hubv9wcjM7yG3pkoSgE0EwKeL62VZqrcsOqmBP9xyGtU
wBf/tKtDKkMIz3+qA3pVF4SytFvgSWAl3bnAszXD+4rvB6ew7drU7KHm+wti2s8S
ilMzDXbPOZinTMDSjazWwYnCe9IJwamKgEH2dH1f33o4zJG3NOV/+P7Jx2ifzVVL
7x5nTwAAS3i3tv6EknnYq+lgUm0L6culFMqQmVWn0NQgvqU6NAk5G5LJdl6WnyPj
/f4nC94QUr6I9RCjSmssmocPjjP4HOz7oW3UPjnfzrI/rsNB5Q59TQZuXIqHBaGn
k3bEqRfn870pMPYnVGfIUBv/p727zOHihE0+V2Z38x0qs22v+EJaQoecXnHJ6CQG
g98GQGJajGYOQNuaz2S269Wh7CyWINCEyorzRQxSPQ891/+zFOrhL2DRPXIEBOc6
cPBqp45N7ACiHhwTaKwUWn+Bh+UmcZ9UOTSRoiqJJA7XVmaVttzuxNDROTO8fDbX
t3FI9VwhdSehs6wx3xwUW2wCgVTKQEJA1LL9x2015Zu/XhX4tmtJy7LYsOeTg1zg
8DRXNESnROYudIfqBWvXO/45pvryg8bczYCofns9s9wRB37iXx0EH1jrHgGEdCKP
iYozeHOXCZG+pJO+bIytm/RnSZ46dNN6Z8EQ54eV/ZB45p/cy+VVuj1L6SaG3TGP
cveiGksnpEDfsU9D9TcKhKIochpwg9s8WB2yygcBoPysHOIyInj1XHJuP9Er3RrC
GXGLy2xkBlUQIApAYBt3k78ZNUP92qgzjUcPrd8jdc3agMcg0Xcy/mK9m8L+SWqx
RJ5tRT6H8Y6CORUTyeA5kWi/c6Wf68hd8P/frvlvdQidvuz6ozoyhPWnYdghlww8
3X5cecBfcc//BUqgQmP5ZqaRGDAaSwiUrsZ3n/u4WkIMtrqfbsDbPYZ468NMqlLk
FJcL8QoVLYjDWkaMd2PiPfrNf89Z6nbWYy4WRmE/x4auOtLPt090y/SAIbLlNw9P
u0GCxThc02hr3nIHAUjWqcMp3G7cxBXxTCDXMq5SyhwxlFWgYSH5LNVpgW6AM94W
sMTowFNYGTRvFrx7AVOEmjbTg1wPnLskLLhIPOR6jlEPuLUARf1bccPoRrY3dEq4
ci0bTo7QGI0vlUtpvIWDbUiMr7anuuUM3g+gV2JNqzbl4HpSG5GPWT69JFb5PeCO
jueU2TwQurQl4MahyJSmEnJOOdivOYQZrmzonY9YCpx27LImwnRJQcIWKn63hZVw
SuDRvMq8V6izpwiTd35lpjAoMUwHKeh2Lr12Ya3KHpyedE7c6I6DkE7zPB7j+x2L
JOWSAgL7hfJJ3vjAooGRE+HKAvGGWb9b9ZehrcjRPONU0MY80Vl8wGwV94x8YQYM
LFqt0nYuhAnhjif8u1Sb+jNLVDN6BXC4HFb0wK+MDuDF5SvrsgAgl6BafiyBM4F+
3dwVItfiSyg2eMCJKKPnm1UqaFm49OPnDaqlw/OpwCyqNnZzw1ykKOpQhZERZpXl
R0WS2frHkfCzybiwUd3TAmHaUtaIGRRhjk7sjqhPEDBEM3p2MKI16j/R6n/bMznE
W/zO4DgXuF+Lhp5i5Sz0Z+UDIS6Eq2t/26IjzOrdcGqDAoeLbBmtM/+wyHPHAvzX
kvX7H2zK/aXm3eBm5j0ujl2xpgTbPR5MVUGE0vhB2yuaGJuLGK8hfKuthPOnNASD
iEdmWtDed4b+8gKIrcQbH+Qk1toLhetiFSqZ1idQtHLweQoS//xZWkKy12lynPp7
SAej9LbXu6q27Pe5VDKCwT6MjoyqXvLEs1Apj8r8Sm9IgDPIw4+WGtrDOyjBFFTA
TBFfDihEvnUuEjNxMCIIQASmfSg5ZEgtWQwUaRHHiOOjtZu7SB86Y271zGue1ERx
5uO2t+LyXZZA4sOF8FndMURaJI3RdbAlkmHkKjIyvkTn/ZHAolmp8/ao/qAObDzB
gnjyKZKppKzdXxJCOlXDHBL7BZCgmFS7qQWShPfqlRXNfSEh3w+Ena2AW4TfSWbn
e35Rpyapa4QuIrYfZ4jzyNg4sD4wUXuWc66Dn/cxoAz71746BR3aoNUbbZY+978s
W6wuiODzk1+sWVnIarnnMU67Np+xe/7sDgpqi6KxpYRDKTsE4LZD+O7W2iquuv9z
hsBxqixKWrQ/xoXqTG74d45/xCZX8IFUhEu1jrKGVhHP9CvaO8roBqwjroduNbce
JkaC0ApxH5UiW/YpSEFq403Mj+3LJG/G/O69W4zIGwencBwJGWkoK8LYMHljWBYV
jVFpSJHik45Ug6yhtlkKcl/f9/2oXS/yGcJfNip5udaEjxk9lOkCuBrpmMJ0kLAN
XUSDyLJknr9g/46YWt+MmI2F6x8f1VmJGaxROYL3Pd9gW+ejEhp98IoVkmoq7O/Q
x4bZ2LXjJzKXw1B7yLuCHqT2SFmgyquUPxA+wQ7Q9pdLzlh36Ly2oBucY+HzMmM0
4Izlua08U46qfUFpb4/Y0u815Tt4P4u6A/fy8EdUcr8C775E+T4ien1akBeYtC7O
38vj6hQhABv8rq70v32+s0QCw21Lc2pCtA/+IWhrYMY+VAYll9cLxFavOqn86ccs
jZtp0Qqt1np32V3JRKGXsO9DJqb9MuR5cuYw9rhhFY2Yn0OMoW4PABEeZt999Bhg
4zbozw+j3XxKQyDWIlYRhAWdQ3OWNl2o/i5o+QYwYbBPornkI5w3fFKebVssFO6e
hNj3dwve9XB5lXcsupfxCnr/i1WqR+uFshH5vP5b2tvwbBAZ6hHPK5ODBkkvEEmC
DeMsr+ohQJ+KF8OZpD5tpqDuq5CyOXr35EiuMnochzTG6rgEOiuxXs/KXCSDbT9l
2lahJPcKTREW8f1VRhPDOXHnvxnJApeJNCiFr/zN3xczV+YDai57ICxjzc0XMylX
N8QVes/iOUsGrRkAH71Oci9VQ2DCfiS//4S66dlk9oUf84/8sdkC3ufFWgz5bPYN
sVVSqIbSMEFQQtvRYxVGKGFRKu+omEsbabDYpWw4M57zTCXpqnxhvY2h/yYqTvJi
A+u7cVeGJmDgN5pcEY691XyZhjB09F+3JzE9tnr0W/E2bGLlPd2IvVmAPNVyR/rv
5tVpfC9Xb3iFBIkvcaiVrkOcXTZy5/AAMNv6UfJlZ6PGdOngA3e9QEemBcuqrBJg
GqWNBG2G33LNqoEF9jwlWj50PxU2F6rGdK0LlAOR/TGgC7nzd07t8C2CG76YXOGx
puZ0tgAX7AaSgiN3fNPlkQwl6r5WGy1RZiCafh3063E7x0V/HjU8MVSdyUKjaX5Q
94t9/BMqYfMIeyrKb+EPJnx9DrPRIppiez91JiUXQfvb3b63a12MJxeu3brxFD9z
g8FZifEXLEWuGYMBlOffQ8H2t2VaGH6bOB+QzaMAh1VTBufw3J/1Y6IXh91yj0X/
ODfiOjhc0MJI0h928NFJoKtH8Tzr8g3kIaiqEoEPFDNmCgBiZeUeteBPkQDVRXij
P1OU3CWjISN1QXFrktkc+ATPPCYxTrgDwWeukOrzVy7NRSf/s/0s6pd1BCxWX0EK
gQNDpEPnUV23jEpNKiZSWOnVmgu+fEQ37r7o3nqB6/u0DgEm40tc6VpbhXl47ctq
d6okXbYEvQy54NcgIRNwGMMGpVezau0FiyTU3vV264LIOLjmh8Ynhpxn4fXPM24Q
iYF2TyjFsbWX6ZLyfn5cLi2WpUScYNBi9DIRayswzqsY+MyQafvbvB/GsaOD+mFP
v1qi6dgusjTVhqJ6+rUCgQVymkB7DAT3sRPS4L2bcsSLaiktNqhnzlLtcfU0yV6Q
Cli9Bzn7kk7yrnZcVF9jKEFCCMIh9GrOI6A+ih4C1l5glnmjNpL5Nc7PkUj43tCc
ewqz2+gNO8OzNIGIBR3eb9mPiZoKhuxVgUQqsDo+mTR9S61rkgIV7Ss2XdIyYDMD
LKOzHhMsQ9pw3V5kgGTLVcFcPUkSISNpCZcmJ59BhkYW5J1RMd9yKr26yO/w22ss
z0gG5BN2/twZ5D0k/x/FECokAJR7RjdCtqgquMwbWIut732/ZFN7fP0TvhLVPvvU
XHnv4T3WGrCR539HpQUiU2XSijiSui7RKzNvDHtpJag1w+fQ8+xgc8gsxXjFFz0f
g6GRuxDrQ8RLPlsQ2JBZx9r1oUUH9FnqC4M/h1M3uZDzqpAlCgYadPYXcKm55A0z
4ws3EusRIZIOc0FsNTMoNkMiFwe3C3piNkqNEl5elblKqLuGKHdUyTYipYFGRN8b
NPCbPLsej5vOyQW2D5VDJ31QhDB/834IARQhjD5QwYdevrFgSiKRtMRFYjVF2wVs
MOmjTPOpAu4cGIOkuDHWcN2cndBtrpMmYWML8Zr87eBxMnsbytCjDbNElfixmZO2
5TGibATYICygnWdvD17xUC3Bfbn2qW1BZTBGaVoTEOEcSHlvnI7MYAdCOG8XFPQy
mzcLlcoRhs0knboMAriIN+pl5g2ku8cq7gxMzMxNxGSiRscY05fFwMiOas+DknQy
mC8tz6ZMsScbn87Y7MZEpJs+8lmQjtckdx+U2q/M9O9I2o4rq5qFDrDLZZlEOtsR
3S+VPpzJtn8/Y/ICOUpIqswh3M+nGWzT5GVZ0cA2Vi6asEKpbqt/mZQ39uVuMb5V
bQQhbqoVk8MthMlej6K5IMve6oC+iNy4fWPLajyEVJCx6wM29zmF2YydJ1sLiPeN
zHQz50D694Tze/L+pMUr+R4z9pboLmcTLlteBmEN3MpEhdJ4McDV7Z5Zpuj9wXRP
i/pjqu82bgcctlEwPBKHJF8njcEQ4cLJOq0WVmceW/sKUhsMlhkftUoLzW86KiFE
AgbjxptAb6rSLsegi7utJtXCudy4k/m+u4dxsUdabMPbMi7s5B0byIyyHkp2r9/i
Lc69coB4/EKO283mccZaJp42uSVPPxw9HG+nVI+SxvFJJXExCu6vBy/ByvC5h7Ae
HIRVUsxEkj1rZ0E+FcyIAfY2cEPmQqFVYnac6P5OPoPyKwHCaz0PVs2Ux90cqcWi
0SbLJPSdg1LzO7+/QB5BlrWchvMeT/aqdfrR23gqz0Pwet4smt2pMHYk6KoT06PZ
NzMbvgFPP0ar7ncVek0adGQEpGrQvSuG3yIS+33HMWP8LYN5/mSXpOEGwMhCdmTo
nnpnwqKp269o6m1gh/NH7IZol1M3jZiPyIlqmUeLmVTz8Q6zbcWGYJ5yi9ynZp89
eE4AzXcf8N1NaK9ykZMSQ1FYnIM2kgkDMuFMbAxGK8SGpBpoloPOsFv57USwYKFw
lU4jBETfm8Mo/9aplAE0+rbvPKcGHRu9mIxoOUgGJAhKZ0Kgw2TFk0I/frKiT21V
jjkIO8I/efqErpnJdap3p/yS0NR0l0RVZ6rTLXMSCcmZzua4qQ2H1DJHdd8+fRhm
gCyrXfRteUoc/hIcXPfH04RvZxcUwlbZo2rf+JoZubMm520R4tQQJOE6jEvRFETp
Ph36cRs6encbwoZ0o98mKSvFPso7hvdcbS3kNsUta1MyGdpKBVHk2Z68pwYZvyLr
/80KHL4R4/6slIM7mrAkQOFnBrF3+SKbiyzSuYtCs2jqgmlB+rCqNecha8e7jGIT
+QHypU7WE0PzDFyhba/6EDueAy3/LL4C7U7v5d4ufAyAKiOFR5rKhEGWVE+On+Kz
JMw4rcas4QX8lOwFE8AyDuqBGlI8LmYwndFmzMV/aCZSg40vDe+4anAoHq2M3wGI
IKUAPhAiYaC5MLP6xH+syZA/OXugCtYsyiDOccd/ADb6uMiZDoNTaidC79O99UAs
y52U8LqYQp9pwkauuPwohhk93JdWYN+OjIogEKkF+TWSGqdIbGNhJXE8Y2iNeVbi
qxG18icBfnD3u9tDUsQm8zZMDPnqP6/caEGK7DVgI8Yz/UA0uF+ruMv6n03lvv5R
Gr0QJNUOiTuGc1JWGm5twW2Bs8baok/vktndscOV7wA5obhtkkrLgyB/xwenG85F
4Vweu70WQRj75vFI0k+LJEo2kmYPNdUKBY+rwq7J3Hc/MFmQJH2rbiVhGrwT832o
paEBxYnFiBhyGs0hy2XoQOAdkTVvxRFQ0XKijBDwbKOh0ph7VIEfcqBepR2r4t40
7T8UwchzM5CNaDxpR4R96H/FBteXS/A3hPtHMvAtYHXRrTUlkDGdbLaKbgAUkj/V
n8HgfGonvXB19svsK9EQV1p5Wbn1ruqn6ZpqqyXQFKj9sTw7Ymt3YwFgxaZHJR2T
ldwD/1+797Bj/Bq1TbBgbKoX5/ZVmwwaByH6SO4vKk9rz+hRfB5OmV4buSn/2lHl
0u3Lednq1gC1z60wLs3wSjWV+6QBZiypueRS7IDHzX7zfnkalB7hXEmpEeXfNGu6
cxJl8m1wMrBE6Xan+O42zjf7qG8+FkQQXCa7sYcibeRUH2xovRaG2FEAOv7tyBcz
Jwa8NRYaWhXrHYMbGjyk+1o37aSn7V2fUh3kYxGcJlB5jvu6RbMGenK5KRkR9P07
pCft/amzPkwU0Tp0HGo6IDZSbgkI/gkx5riaODNn7Yn4sCCyU05NEHXjijGmO7lq
yV4YLWIllfEwOKo0ki20axXzrC6hNKZ4IPU7T6V1dNQznyDQdbkkj3Vbegnd8cCe
zlI18lYCuCzDDOXTAqq2ODCYtzVbPGs/ulGHZmF9zYIzCxLIAOuqzPEgphAKlsQP
WpPeAEzUPNTZDh4bMPFgBa67Fenurp/QOX4GmoQA9eYyrCvU71/LvMRab6U5zdKd
ISVIoeBR2ePVu0NyjEnM/Qxjp+I839pHmfF7NJ+cCq1EMDaIAYiLj3nR8uRFObId
56HbbUlj5CU+NUpT7oSIpmWO7W9eDL6iPZ9TrgGrTwWYWVVrZKZW4w1riB+FZQ27
ZtC82Rwt/F+dwU5PaML4LrlcTUA0X3VASO4+mEcnRphNIqhqS6YPch1EVl90Pfpo
e61zoGf7bhxhP/3Zli019zLqIx2WQc2fcn4mnXHzDuoSwY5adJPSrZkSDnnLmiyR
yScgRDDrt9NiDscvPUHqb7u1r9RQfAGiAYEa1HUPOTNdyMbICTyMmYprCuzCujUv
RwwuzDQCwnwv4/DdHzMbj5Drqltn6JE6PhO/VWq12GuCK/sHHRZ66Qndf1LSYEKG
8gCemdmd2HSZS6kAtKs+GB8lJPcIJAPZIhPnQCVIui4RzrUACq//ToFkfjZZx4Xe
s/diJZd3bI7F3D6xBWVTaL8VVV4z2iyprAKakPmL3cnmBcSo4+f7f5WARwzSlW/n
XIKVyjkAALaOJKcn5mGAkEc5rZIhUtTTPPZ/Gf29A79wZRiXPnJM+8cpWHZYjayF
ZVwdD721prxsxRrPilZo555ThublR2KMS19n7mQcRVs1O76JitfZu94V0VTtsmqZ
4ook4IgLv5vp1P3pJX2/e21PLOHaRZew35HQ5Cfkk7xMo8J4lXIHqwi8Gv8xfyYi
9vi1Oq2Jo1wA4T5OOqyexHUf6pr9NILG4fuW6ANCl9L5MmEoW/6PHOZ/b+GPmmEm
6IRvJLAWqHySMslxx4csCmHbBrVzEKbMK9NHDbocNOxTW6Rur5z42ZStmE8+fUgk
p2h/OVDj/wLb79++IzPIfcrNzDa0BuiHg3NEJCRh29eY35BUWuO6XajMCaHY5a1C
MsBjyC/9VFAQrnO9uVSaQnslS0EYaF654F9RPiYVTz2fiVNTuJ5lddwGzcjEuloA
yBxJowuENq5KivK/SkS93MqLONVCzj2uA7KJ/Xtiau0RrA1ZOPMF3t9diOc+8miF
ttoV3LADBS2HWOqNkohyIBsbGBux00rtLW6lDoG1NS+Qc3piI5X8INpfSaKyVmxy
Q4O6mIY6lgz1BekBIJDK/2xfnSZvUvzLMtcHDNUuB+HBOVtE+sQatF2PMqDG5pYm
GEg0KGuV1RBJ3M7iTdAm7NFcPC28aNzrmgy4MkMKlYIGmomc2TYYceulePPio5a4
pd+eGCULNcE8f9OAertyFceWmhpuqaEi5IX2mA/Y+PFDSni3N20GGEQAS9amSb5z
AVd01ernLjq2Bo3slaA7NFkNM8Wv/LwS4nOWR+LtXRe4mJtH3v4y3ah1thAWZjbY
Y8hLSZNgAbJJ8ngPdSnKF6TjpLGaLb9BCWiJ4M4DN9SMdcejpYG9xmgZVeSJVezS
PYJ59i4U69hgYRfsa33+rDZQH9FgGUgEYYbox2qpuM7kAg5o4kTfobOJjkKBkMlN
jS5/4wkKsnKwurF9qIP9O1Vj1nwJwJ7PccPddDCgQTeVcmGdEQyeDRLmJAnWLgvp
saKMGv+QAX5gst8Z3Rvy35/AL28zg5FlZdRNI8tPCJN4CSqyeelUys9XWMsCohJG
4FcM0edZEZ3OtmzCuMeerApfI62dxGtK1s+YhKoLnqckYhf02OHBN/Ilzw8P5d23
daDQ+DQKTzG+xmGXUdvbNTQdAfnjYaXZA2lfzvebGcXua0T5ZC9tQ9P2XW1lELhE
hpfLyIGMwtnK72LLMfslD657ro3QmTbL3hk4Aav5a/vI0PZU6Q3xssDu7HLLu2eG
JPl0RKCCjs3xAZwI5Ug55Tqs8m3+iZ99maMz30FsyT3CFQ1otP4gD0G/rH9EzJt0
/cOwK8cVwaQUKO7A//9FQcZOw0ykIs3M/hMffNHKV+vFVyf8sTqPrr1BOIhwsgFY
N6bo6YNK+UZa6t91LueRyoAYcELd9jGKOezXkd0JQnXfoeJNyEuYNjElFvkApGuJ
2DRJMdd6U0bT2F8hsTtn6CUkrHwpKsgDcpHv32MBkNYh557I12dk6Ee4uqUYT2J/
WizVUO9ffW7Jg7onTush5Iue4Tz80z8VMK1Df9A2ZIJluYK8vrWaeRfaUN9ZX91/
PqBq/SElOe4ZgT5Lj3BMw4N/sFaCFrVmSrkDndcJSdqzfOWgu4AjQ23oRcCfGkha
gas/jydWHFcUxnpW2pxdLYru/Su8uwRGyYZMkYAWLXbwI0YJkHuPgsl9WzqcMtjA
APYcyVxSK6avsP8Joh+p3pIQlpaLsKzCFw7S3S7L7jRXAudlwvRLFKZUbr7VeI2v
dGqOZ0jFNRwJ8jQEYPE7U5vX7Ab0BFpFkbT3EdwdjGEmmW2ak0utilL5IPgPTBjA
VxXxUew+BfmbnI6BkskOwaLpYwyUYTh90JChRn0fftjBS8mI0D7F98Ggf8WenRA8
rsgt7uKvh9M82RenDmhudHNeZZFehwmTWegnX2z/3CMy+lhQM+WLug7VJifn2U2V
W2h57wEOq2INs0vzOzC35kS0QhCtKUdx0xFMKMsXNB8eF0SrlN5eqJtaSlMTmPiG
xJC9Ts55Z6wicnz9ABPobHbZ9aLs45+j/Rl4dH0Ip42A9FAXmp9+bH/OoRLK4vRv
6cwpVffkrlglLv+W51hQnoV5dXF4SdBz3CtA9E5LvWUGqCJJv6AcOBUvu8YM57qZ
RFw789B3j6yIz7p7mitwA3plGVq4uWdeAdPq1oTJ8xjatAWIW3L0LfVLA4msQ5aL
WXnwL9m8tkhlxSo89WAM1VS8OtjxpKmLMwly0IpuMPvIYQojVmUWrAnll2/Av5FP
ZS2aCrFHuW+FyIkuwcEMsJnzATeH9SPc/XFpPiNZJlKUK3Aw+L127/mc5DKohm+G
FbbGpFJ2bmj4kr03Nzmgr3KD6tIKlLQCefFdCkw2R+aRWohBPgVzobwZjviNc2V4
E9+sg+v1c2+iuB7BBVqG9m/w8jkWdZTkx9cqZ93oyt6Fo0OWV/Qvy2N+vibc9cTF
r8kPiOXHff1gFM8DT6L6+wBYALd4UGJh2EK8ZZWL5Gw33dHSf9ClZyuE8B9OOFFn
DspwKaTh1jCem9wZxlIkTcvgzgSotvZwlIQHe9TfSPcGvBgbQL+763zzNdVlUOCC
/WfluecYFhQ1sGdOhnsn3Dvtx+L5J6wEUOqDVTmyvjcEZ93EkczfA7UEZ6nOGnMM
4iZTATiG8rBamT9p/9Fx/fZBqxLrV/J0clHXk7IdgmJLitqH5tsbX1PgJMk7n0L2
DlQDGu1bH3ExLmjNEyLpF6f6Kikb7vcO6kudPv3SVzKerRrr3WT5um2BogZuAu0f
pBs81Uung/o8lLnOXGvIR1EMeiRdi+QAyWVXRgM26mRXrTGMQ8cLoUogB0elLdZ9
p1ZLGk+We5rh0xABejRM/yqEDWcviBmL3Fdsz6h+kc1U2oDv4y7q5sJ8eBnkuRcV
uqpKT8bFf0AYLSdOKdOkScRd3puD1oY9aa717bCVj7vMTa750XBUav9BMN3Sdjh5
h43YLLKdtxObP01zSAvn9BieiWa6Sd+AYULST9/fwtFox05WZlkwVvoQEGabXcIa
4bo7SnYeh3qNEmzUhbhtmvtgrVkMkpC/ZZQRUFiSjXSwWeaOuEo4oNrd8XnMXe8B
VJWMHJTovDG1n5QN9wrfGFxY3n89Pa9f9+5ig7ek8loL4mcDGEB6q4iRHY185sIX
TmnOAOVpeSDug8Kbkdn33sW0J0yK8VRIw6CL5yy/nEAnIGSff98SqOw5XG2q//IP
rHMKseB2vCxFl9zNQsdDkwm2YvgTv6+r9u89CF1mDZPBVj6t92hZVTBfuKM4U1YH
QI8ZNssCdBjALfspnTVuSkIipj044SgJHXdnXyNSEPO2F4PT779cZabpwdLf3ERt
p3sNCsvAcW6oq6e+Q6yLGpDBAP61f44zcynKXgKvVxKM18rLbUc4C94LyRrFNAR0
JCR8cNpq1ZIISAbcVDUFqIlK/HIlwG0ZWlKeHrbhbTMS6RDC2RvclB4DDmFlKs2d
gLnqYfhrFpSddE9znE6iHEpbgbiTOwiGsCK3kzCBe0g8FvDH4si2l7BNYHkUJzo+
cGWvG3QUMJuYF5qBx7Kqzz+aAFGN26ft2kxBxRrPRiWsraeF+KNwB12NuFbGUyPt
yJp0tCBLpXbNSyaEhNLw5VhZ7b7yC+3mB7sPralnsM23E2brkftSJqRtOQik0t8J
HOOeqzpf043nw6EDXB7bpN29oyU+kH05XUTJcZlAa2B2NP5bOy4RCY2TOMudLy9c
LiJr07c9ygiY94UWBBUbtFZzvzseHJIjMNeHeFMEddrsjP2DAvcriXnKd5HGewWA
SdV0TB/QoWhwk5xyEiJf8yB2c4k1WqMEx7dJeaZXYbfq6wO96hHRYBCK+CxWhFKX
/iUVcPdEEYyADbN0li1X31vUUMKWEk4GWCugdghl5w/MtaBhmHhMLIHRG0wgKS9v
WvvqMl5zznQzdz+sIl0uDOivJjWD02a+6gLeOZIlLK8dWv1Msju9rthGZmJS39Um
Px2EIIv3Ou4XnofFjKyILn7QPI2RP5ixEmCRX37ZoGAdC4K5aEjVxu0eKONnZLPz
7TUQA8L1s2cu+kNgvcrtuHy9IbmyERhT7+zS0f9c21VC+pbd1T+3oolrw+8WeLx4
awgO+9+v2wCQbziqo1Rpd0Lj9b7DEnPpQIR+Oqof/PE5FyaFvRnjb1u5+MeGYZFA
0jhI5wt4/3Q30wIf8w+sYsXeuSZmEZepi9VqlEAk+t933FVZagW5EQ8l2RH/t7p4
3/7xB0NdnMsBNJW12Z/gVzPLxBSs7o6NQJ+G3U1F1e0Od4eLSl3S7wGgENwoWE8H
vRJAhEXFn3XMe1pf1Brw+zhDF7q6MJefuAQkYIHjE00z/CwFaufxojkzliSng/GK
e7oDM9DOw1iW4EBBEPv0fU2dm8kaBnzcP+qVN3wnwOrLTJCL4pv5OCtOTUMCNvii
o67rfW28xloAypytexTSklkxeIkRO6udaRJMR9gSc1htGL9r7vwRoy8yFDjtzJ96
BHiWj62poA2+06V2GNrDvnHmAZhnXt2I2174YYqfsUgUL5cyvbIqNMN6eVaXxprQ
peq7svcwh0MytxtX5Hat3iiZNOksTotSQXnazIVuXDjHIbJ5xoGCrh0kaFtFBYRX
zKWjcSOxBH0lwohqAAxi9AkJJY72YQsrc+AqyAn0O3/u7TUh5/+yomofAhy9TOV6
qi9cfQK0xwfr7bmYmwTL1R2WGMfzIca5TZoyaAtPBM3LH+girZcyKNdzmBwQ/4Qz
hWqewHfPThpA8PZbHMFEib0S9QsDeLrmCrmWqrlEAsbpU7Gh/rjNVmMWsm1cWKXc
vuGR3i0stW4EzPUKtp03BaH9TAyBNiQSgFMb8HoNG3fiIrMTUg3RWnidqadRKJhu
AsFDiJkMjNPaUOEZWRyV/sA38zXnRUflyHtHcsTxzUglYl1v04IFOXN8LPguCZZF
aygR8xYnI/i+fn4Y0OempcjQrPBw29mPJS1c3oJxVYcPOHIdZBF99MJJhPyBJyXg
7ZXZ64ZgEfdWka8N/M78hbyiSLTukki4IS630lEiXak5QSjsTZNZrZiMDvYiCCub
oq7TFErkEmsLv18ofyVvEkdNDyqpD0NSt2/6p68A78A/aUZAS/oY4JtYGQEvHYjB
MHZqznorU+dYDZlNpV1213VuffSlLkXesz2BmNODIHoEkX7BL2giHdiMMvMgq9w/
eteGaLDaVxYtfv6KQBy3MLWJhH/jcP7OV0sSdq+4lTKuU42r1Ppmu4K5sunzI0XL
evIKbcGz6vQOThHSOK8c1RRPxtcc1jdnpYp7zZU4+cIsWyTswhnEj+P9TpqjMUNv
rl8jc7R6YRCWYis0vA5iQ42/tMfSUPgfMJ1EyDMJmFkO1bouTXVRL7aNyHod87lO
UWiqJs4QPQa5Oj7v3sAg1mX+yY46XxgDyyOmXHwHz9oZv4rpv4uWsUoUWxwdt/JL
dmJ0tOXRMvKjlrwCJy2zmYFOxooq3t+yjxdyNP8tquNJfol4zESx+z0eiVcuwUEX
LJIA/B7KuEzB5g+NIMAUf4W91RdeY0Awef/Qr4Yxzy5ubIDjCjBu9cR7RcgKfE9y
ZCBI8ck+WA4a62ss2DDTNLcIOYYwV4ss6q3dFQBCfLiWzaZh4d6/eWkYnz5awHLi
uGKVlI5IfieOfluKc9BDY1w3aQgVwR5Jj8iHZYMCPVHByU7oe98lWAyC8qKbHQDz
erEQdfLFxyn9B/RcoaenCYWdLbrCV0zKcy6kLOcZAN8S7CBkwnnyS0EAHVH58DjK
/firmKkX1z6Y94wiACKUSHjMMQIYvjJgRqQH+KXkz3KMge2aRupWR0KIeeH+Ceuu
9L6lYEyTvkj1LHRWmIW+dKAwwPziIYHhjQQYta6hbOmj1u+ZHJrhc2IJX9xp1qwL
EtMHUbtRhZxxfook8m9WKStRjYgTdAyUWVrBBCx5ptJgxs2jrGKvcvhy+CmDIjT4
RX7RGmKskl/qn10TKgIf1Ywc01L8Bq2URdIrjuCOekQVHOX2fvvsx1hu3cU+rS6/
lSSeJB5/6OLhLpYJOQCwbfCzFCkwdwg9EcfufpqtnGddTPCuN3ovS8cEg7ukn+xO
k1p8ou98c8XKfaoj/Iy1uLQzYVHrFkrBKsjutGRzn7xEy+Gmq7fZdu8S1OYdJ5H2
x3PSebMeJjXCSYjE/dBeuk/t+g5lUCnw5g5PtojoPzUupdEpflhHHMWTaO9nDr9g
3Jqy1u8CpubmLJXeyiApusIegLkwGfnTQb8A9t6j4LhSqgKCcKvZ+52d465zv8CA
/5NEq719fg0hbkTXjuhSSycYHlb/ryY3PDWVm/bJpBWQ3m+q/5gHeN+nA8DSwsn2
uLcxW3JNHhF6J73uUHGxCGz6UpZfWSj65ZISIx4wHc8AhJmCOPZOg5f9YtgebybW
HCsz4OAIjwHVsUq2Dt2muDZb7/wlAGiiyX/k0keeD3Z20ZAOiNTXRgiMWR+qNrvi
GuslIKF0Lvmwunp0ssvFUuK/XoNW4XsdtIQ8oDEu8e/Hs4dgEYuo3yvZcR7WyPWf
2go8J2Yx46d1oqS/0URCk+1wbwik338KBmBhtB7tfbX1eyWDYSkFFfvnlNhk4kXH
7SblI45czttZcgqCs41wbRTWoQxmNCGpDhX+/c2amguHmbRx3sit3hx3SaZiE7xn
j0k/ICUfMrKM+vrw+0fW0ACrZsu0brGFwclGV+1ZT12eWIHcnCjeRVHJ1qynT4aE
06lZmVgxZdomG6hKqeXT6FAh2IlWSU3aus2Rl6gMtZxzt8zemajNfOh3YvaW6SXg
afnZy6I3/2wwyZwCx6zbwqvHxI7lH8xVuFKUkrwKZafLXDVXxdeegOuBXvv0znLq
or/14Q22WEJrgH3NVZNJN+u55wR8RqXuRk4MzMV8hyD9CWBMsc5UfVHv8p7+B8ME
WgoER9tJdSDXVw7wdxuA49PVvJwTJTI9cvbWGJm58qewxhdL0HRVxrMXwr0hiuUL
PaVBkOjbvY+Hplo4HFU8Xmi/v8dJ2TmPAsKMu6an8MdOImxcxQHOiCVdRUNLOR6s
cCNomk4rQVmdl8kBSrIbTAVre80qFr6III9uI9WwIDQ2s07UN8J7Uw5Vx2ohrXBy
6W7vbN/mNlEGwgsupEM8BjTXiRMVPYeRFQtKw6QDmOLHX2t2G7dzLHF2LfVjNwRG
pI/fQMAeuPTfhUrQRr2lUdzYrjHQhQ4Ba592cPJ1cUbKoGdvIlwSVIlKzHwUVIGg
wJUtQFbXcqZ6zzGPUQbSBzYtCp+f0u869KY7xNLEllVrU+7DtAlRnBdZjm9MyM7M
DIScE8bE66huWy+PqSulLwxEq4LXtLGrlv19ODC5a/UCeGFYCwdpe5d1p0j35jDp
BVUu2AgQyJZxiObIXUYnKt0kJG5nEsqhqrhz/8w7bKX52FjYACskQYoR872NWCD1
nh9Q9kKESof5UN+ctqYBgtdQ5dgYQEe8ZK3u0jBGvd7oWZvYyXmUkoVUTT/wkmlj
HyTjiWVsFcXgOkixhYQAv2ghqxf0lwsAjFPmv1/Mn8oPFBPIOpQPWiqiooaap5RL
1kqzwrm2Md1WgQpyDYpK9oDYTp3/n+vIYsxTr3/xf/lFS3PZzzRTV11sGkhl8son
aAbCy4d7X5bRnS9XHVCQ7OVqRhSXcPVakTgvUGEYATyJ9zdP+Wyw9FEYkpQH2o0y
3PsKj3Qr886zw/zLrF+lRn3U4O0jTezlcZ52m9Gdt4r/9D7YvTXd5aCpdlwpF5A4
2HncfBVPRC2u5Fg44w4Y3fiZRRn5xWjkGGZeL82qm2VuCLz1TpcFUG0FbCh/HuSE
ybzCBKdxRMzkBGG3wvh8XbA7tyi64on/5UBtvDESawMs+loHkpfIWDvAV28IzAHh
DDGojt2GFdx3dqBnCRaXGkxkbgb9VkD8VBG1iSyHXeK0+tmnTVg5ra6zKLMKb2Hj
lsbEju0wTa2IW6eXClN697EufGvYapNT74Eq8Q7FGa74Q/0VboKG76uJr6SZMeUK
zeTI0PwACb3CNbiu5WojRQZT9ErYoQbjDID+2TRtPqBjcRiSwmhFxLbvmN1Hqqtw
94Ogtt00bTS7wN3Qe5Q9EKWZ5t7i3+iY/ewdoApOo4Qpu0OsLbUc5n7BqHULTdqp
qqVXm8lcB6vxFfweDKk5qASnaBy6oFI96cHgtcG7VEWgEM3lj9rzzRJ7anD3KbFt
B0SFT45+kX1JlzUjjuseBD3bYyDp8/VND0BSfwh7MpxsYStgMH7dNMu5ikWBkkm/
z3QopOc92mXAhHTsf1tPqQrNnetVVcDgKIqzSaR4iGm+EMUZpQPSQm+XsGEjuOUX
4JsxYXYo+GpOCRBSSU/9E8qbh3da4czC1PIAKpKr50U8isH7R7fRaokHA/9h1MGv
I3N5EO5ZwlEeP10cz2NzGkEFIXCf1GuWm3NDak/hV74zzmd1c1Qtb4SgjIJ0TVyU
7ljPAj/sAxtycbntElm4ZqxjDVfYxn98JEwgoDJ+VLSkDO/VL8zFo1vWkRt+Vs5s
w17wLH43uOq+aT90iKf0BOxRU/OVLNsUVl4KtSPrtPrsz1RdJPUjJFOHD/93A1zw
UDgzklfm4fA/XMTqhFKMe5+O+yaJKQLYWjFkM+Rdv5mbeIVafQbcOThLHlSegKV9
82PI3VQcHuvlQFbWQiHjzAM3vusYDjdIwtmopTFK0vy0szzNNPEp16rNaWaOxkPt
Pylo9BNCFL/oJuvD65CghUQ37gGABdtK1X2GgWappTLc/eiC72Omohb09ReReqF9
5OHGbz5Wb2bt5BlxECejfCFqb+zu5Dj3Af0uLY4YkKQ1ALu5RVAyy4CrA4ZPuQZ+
KsvF+jkPbioDnml2WRiZSgU0ptczET3AtZqTYTc8jilO5o1f4asg4KO2YcYZRJg+
yA8x2SKciIyEK5K5MOFt+cUJ/VSMu5haxaIZ2HooRXF68SeNYu4D7bwgxbjYmhQO
On4V7BVv5GOoFRXuJvSp04ndC0dE/fIRexTEzgWZQr3uqWY2vSIhrflmlcslktzu
Cc9LUwN7s093CHH0E8/dj3wXQQEegrp9ZasOZw7ekzpTy9v/1/mGidkxik/gC3Pw
64YhF1LI+8iSxId8xRNb0XDpMCvW6neWu//CvAoRC2+c6gkDzyP8tRK8KA1fn+tf
BYUuy7OVPkk9rr6vYSfSUWlOh/ZlSxmFESsD5+o1EGYlvMK0WAvycIOZEpa8LuCu
16YVR0kAoCAlB5eIW88vDhDOily/HFDcOKX6WA1mBIUYR/1T1BbWCJ8L8z6ImlKO
z46SviascSveEqg9I9F9OdC8a8i4ifsPBJ3Z1/Qu1DXx8PPxOchGgqFuVcX3y7Kx
hR4FJ7mbN5c+zs82JvPji8C/MG9EKjvlWd8v80YkH9ezUHCLfgokL/zxIWsC+QZY
PeZHmeUOtZiSmfQvjb5242h/pIg457ZtHno7NxRuGmDTACKWwru7lZJllH7e5Pt/
YEsn5ypKuWR2L3Vx+KPNyKOc3zXCwFF8lEezYFJZKiodcYSOsVeFL0NSc5EKYuVt
WJXAxEWRArS1k90tOCqj1U5g6NAD2OodXbo6oOtVyDzRoQcJj4wF+Ozsvtxiw0FD
rXWhPmZn9ngjOjhN+WCFCHPVrhQlvKNnd/Orozb2HpW8AmUiPhmotcGyfK9JBNCZ
+7L5nr8CywnmEL9jgaYDjNE7MtwAIU8cJ1z6iryEREYRsqTY80PO9XeqyQD2gaOx
FJ8VWfKhXZKAyuaQrb1EIZamC6Gi/hJH06UaG/trI4X3Pi4CjvjSYCUVpnmjlTEF
35E4zwQyaCxbQbr76pY+N10CIQXmKREEsV6+I0OauuAOSgg/CIgG40Y6uOt0kfzs
CLgHgiVpxvED2BdHwCSzS9iyGNV/1MLjH5t30S98fxKJ3up4emXm7AwS9u+u4HT8
ILjItwZq744KR0Hdcur7NOz7W7Os3MmvIVesatTUx1d0kgSO0cv0EgOnFx4Mi69/
zps2TjuvACY+mNtDW2wayYJo+Eba6ide6nNocLFOYOKdkdeuA5ndgiQA3E3leD3i
H5PBL2724OJ/tuUsm02TyGowBJL/zxGhLl7CPBms5YQOwCcPTNLTVPd0gxKZDP1+
xuqC52MeFXh7FgJbnAMP4/6rqArAzshFqrVJww3lQXKrYtMpIx4Viw35ECbRz5hr
Wngjal+/pD6Ag5ww/Z9rw4OLyGtxv6IG8ubMBirt2KRtGIhzUItTLRL+YHPryHSj
ZoTHnk80oKRKdwXpzQdxMGnvDQuO9MzcVMsTtGZW8IL2w7rc6T1vj0AgvKC0POv/
wPbO64OnHbLyIjFmDAVzsUEocecrcL+bzPcGLlNyuwS73Ki4VBRqDLgYMAGvFxp8
R3X3oyqBGDnbJaGEqh7xTy/GglmWGwljsdi6T8ejgL/aDrvC+Z1/ss+8IywJlqpF
QRsw1bvGTLaQHXRTF0qDh1BSO1eFLY9Vrbf0X//zp8k4CIIg+MU0pIieArnDUaLM
F1ekI25piYrsWIxJ34v1JgZlhzL7nahUNfUSabk0ypmNAGqleqtkxHSEOAc/kdUZ
AV5wS5bDTRlXkbThgoS/Nmx1Hc8b311cdppg3S2Y8cgRUkqw/zlefLsWMTJKtjqj
m/WoZx8PSkmIsHjSzHn4x3QWIwXVYQzWwSMoVvLKcjPjupNkzG9ihAXULRA/OqP0
rFwOf6yAypvRfgtJCwCzRaXhHXAAvijyu4uQJJF6ZevoXTraeO1s8IMwYnOYTBYw
kDbwuD3GHjncNDxyPRp6JRE2z1x+FNUh0e3le7H1tUlYb4ASQw/Fd9PpAGIfM+8k
qW6kMWgEiWscbOiotPenPq75ypwiBSliPz6z5uXOYmtDfVvMo7Cw5K8lLdjwSHdL
k+8HKJMgHSESLYvxSiZGyQRAcIuXRyN651wwmxumoq+nol3uG5s/JYjKQIgUt5a+
lENX65Z1X9XmI2cnmKza1L+aN+cSb9RtneAuymMb3qFs9z6hNf3hyKcptQL4oEsX
Tes5eLUrOPTdFk6cVLbNu7thiCVbfqVVxh7EdxVbZC/D6cxHfj6eU/BWUiA6b/nL
KmzXcumaP5vvAAHRX6olN+mf7O/ourPgbDEY13jLJnwBhPw9IEFUPvZ0hpZzMkl5
U5BH7m6EsqyingEhuP/hJ08hIr7y0T/ACWfBPE/VLYmTleRErQ8x9qH9HHGtcEKI
m/7TJgwykM0lNum6gSxg9qBsMnlZDlyX9falxPhPmQemcb0KFsWOZTRdq6lpaAsU
JN4yz+Y33GAG3zlx5Xx2D/nW6N2AFKqYcJxwy3NVMWtyCPNmflvH8GktRzvcvNgE
TqjqypVcjNT0rvduP3IBjuRy7iCWC7Hrp8JYve9LOdtOgKlin21wgK61edLDJReM
hhEUhmPKhcVtZgsaFhyZD83SL3LCD6xvetThTl8A/w5U01vjDE9mh340ytlQsQQJ
0h+poxyBXc88kJi0ws0rSOci4LK7TqI3YnPedx/GD4dPjqIwv9GP+P5j5KICanVz
PPl6jKcrsYQyA7NGjovSv5G61b5jtM7O2bjzRxB71ALmPSPR6TU6Ns1QW1CfCipb
uxwRMEg9IehD7NiJ1fjJL7VMFp3tj+XfbiDAjeD6EyNd2FZkBYk9rqdEvCrriAan
bB9eigqKGXdV9us2bZ+WHNuJUUZMzW1+ByXPJPhXQXpq7yLeXW9wn4Rr4GMR2EBm
KH/Wegfx8Axq3apEsgBAU2z4uVq0XmcChJLC01FsGBEieGUgLWJtmhoCF9wTOIpo
WcqoKz5suoueAgkVqyYitsBFM9CMSzAu629FW/37i+XlzjOtRx/wcuLfoW7bP8t8
3qIJHS68kdR9cz7yxUtuONuZva5N3+r6p4tODhJOOQ6Tsuon6oCa9D8iPsEQxAIc
W3S9DOg/fS07kBGj+hwLXt2JGfLlAllUc8k+B3VsI6geApmU8DDLySK11ASYJKOy
Hu4mq/pkJCt0LVCR7ndktVD1RDMEdunz/YIrCLVNOaFRdgt8hoPA+w2QUW270tlX
+yDK0TDEjO8si55m7G2Z1vCPJaLFoAj9D3GUtsJsqnjp0yDi6vBmpU4fLzCxXvFd
/6H3iraG87rQa/P6M6vGvDlZR3Y+IKbXhKKCXCxqa4FCymp5ueOAqYE1M05kxF1h
+hPp8zch8clXAxsyiDOIECmz3alr49xVtLYDj3urgo4YyjW2KZSIKML5mohK020J
+28c+WU7J2Pm7NTZP12VD71ykFGw5cOpTue/j/cWUomx8U+55lUy1WlqUw+7Y+xf
TsFW9cEnPRcFxTvoG0Nzi4eyAUlLvboN8EuiQFDEGc+JmO2Ojq6rgyXSiod9DJEm
yHWLfNLjk9WR0npChDR/5X9HBCxcj58+/gbALT8mWRb5Qz9ejUWrBtsSmBMRQyUV
crWeLuMwzGlJuJFARVPnrLZB1Yra0fgNlFO9vFfIu9mEWUD1VaX7eW1EGj5j+Zlx
URohq5s+bPX2uZu2YO9sIH2WpIo5wSV310VhxqUgx1he47xroEKL6pwOmTj29nhc
aRWaqyp1J4z8M97aVW53xY+qx+OQyB6a6WR/y39mve64liUSDmyhGnoJ7RnwbsKy
vNT6X4ReKzGw9Fw28fRvgeE9scnfQa8cRdY1LBWikn/YyT0/B0ghPD124Im8Ih4Z
j70dHaxV5aTlIm3j3OsF862KFGxvE6gUwocysJozjPm9mothPP64HoGWvGNf5xbd
SV4qhKZ7cEehguTl9ZU7/O+86exWdeaxnh/Nxn0G/g+3sUwo1rkMPEGNy+GoWmAj
yoVmRoClHeLa30u431c/8Eo31URGSPF0zriNoFIQFFZvARvV9I8R5Ja96pcOJPse
R8bQnuDGEtH5zcoUDk44IHJuFczawWWLdryeYJS2Ngkpq+yDxsbAZDsK8faTZ4Y2
eAo5kbJ6QY+O4hRLYpa6RZMLkvTLwiOtCl0gK7sDlHcl/k9M/K2I6RIh/+oIu8iD
SrsqGazIi4FnCYACaBBsVf73nhuQ9z5KLtoigw/1LZrKh9IMWiogChWemG9rSRv4
ZLwf1fIJoGgUgl6m65A7OX8gScbKXGqBwCi3evZbgugA7Zy93vkhNEG6ijIKUuK3
KwmShC69bnylFinSA/6+/sT6Z6yE8ssvcYQ1Bodza5ohXbXlFIBlYS8WUqrp6jMf
UD3NnAEDDpA9u6ZTRh1/b/HA3On7/XYK6Ci1LFnX6ws06zzlqHryNcHmav2Rp82G
ZOEU0NR6rSHh6ZPSzAKeWA+ktxOcpWYjdDW/9haZW8wX5j8RUawOxtb8AHgqF+Uf
UKpVekw151Ld0GC+vKNchtMOby+FIPAzudmuy+FzMYndM0Yi1YXKdT/K2+VIh+Am
xI9Pfh/Thc5LEaXVBuP4m2fDFnlNo2FwPLaQdghcJWpsCMGxEg5j6Nrpity2KcgP
V7A2iZrp/hng8bAWM2xmnYJxKNoQaHl3nRAGg6q2cc3g0TUNaZs7sjtITqvMRdj0
DWKS6qJPAK3fdCeBHEGZU7L0L/rkEMognFuaHXhT0VntuGhFoZ9zcMYxOLsHGyZm
XCxBUaQYMsh1Zv4yErXYJaiTi56JHJ9npQAw48C7rdoqz28hu95Ckz+qWkhgO6cP
wKxIyRPiIaEpPxVQVFVdpvjC1P2TJIfr+Ve4NHNhRXYuffOMqqGab9GgFpPVTepZ
wjMpFmZv16FCs4QEX6wvoqilKeVS2rrOzXIxe/x/L+ciPY4W06dKAs6+SldpizOW
2vJ3Fbx9lg04z11SbQQo6G+jzzbSI9HBCXWYPvAg/7afYpl4ZLaUDnkKOO4maptg
v/nafgRwZc35XZ1chlQxHaKZnX7YuQ9py+10jvbJefZ72nqu6gMucFsGDxD0+JNs
mFbVHE2SkRcyu/A/2tlRjttwndqZp0tMMgINql5hldfOM3axKDXtmbVUGJXtufrd
DkW9sA1ObQOvkJiK5SBbePq3BftCqLtCq1/knfWbAty41bew10pLc/MMQp1AXeVk
6oji7jUvsnFsp1P4wG8E6POfVp8EvaaRupiiIg6eVAoZFQn2kM1ZEk4hJFLBxc6/
Zf9E8e8litu+XCROUv0wyZ8EpMd6HxLavUwGsirYcjp5wwML5P/EzO4Iq4rgX5H4
4Xami2UtvQd1c4zc9JuKvUaAroaZgV4NCy0oNkxO9K1x0gJVA/Gj6J1w+XP+5hUC
Pje6ZI8b+TaLU8S5QQY0Cw==
--pragma protect end_data_block
--pragma protect digest_block
FwbGE/dcY2raeR0uf+rD+HjfL6U=
--pragma protect end_digest_block
--pragma protect end_protected
