-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
BhcB7m64rIK5c/+5B+wodIDj1EQA3gFTGwoSpM5LxAaSc4Vl9fdmqfeDp4uCRxWd
3K+JV8PCkAgd+pzGCNJrtL63Cq9m0/yeXr3BXRyAOoijBHnMSjm43bxixN9AtMeN
JK4aT6hazUAWWhMfIW5gGl48oL5kpAP5N2Ye8zsdzW8=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 20576)

`protect DATA_BLOCK
UInlhOLnt6S4Tj2rZkZ8qzSYDvumT58DQ01I+iQ/b62hWCaEpQStY+d6k7b+wcpf
2gA60f04TbrINIGIbIKBUcoVh1WKmy1lmIsNcadyZUl78Kl61bgPT7Vve4pJY4cY
qf7c/+h2Re4rrhV8zVgZKQATEuDx77jBJ+hci4sOoV/T4qNzjj7ieF7OC1vijrF+
/H+dR6YxvvhQvlb79feJMDs05WNpq1BbM1hhelJsk/J6ttEZWw1to5Isb/1MMDgU
kcjWW0VgrEZ8gJdY2TrWe2j6Y79m63DWiedFOqPSrZIKUFu3j2uTk920+dmxtpbl
85Vfe0uoikT8pypCUJYRLNN5BWRpTGqcg9/NqBPvqACuxeyCdySKffO166AF6Ugt
rGMwhO3yxzg9d8tDJ8Sjj+HA7a1Z1XeiDIlD50FQ0YT8CIajlnk3KviyVXoYv/mp
YGh2BRCJVe986/riDbVZnyE3XJlGexvycSY1MiSvTRtYib43nHPstUWrR6LMbfwi
YR7lp8IhbGiItMQMe0O+fjoXDGVfJT3tGqHKsLauO+TtGb7T0nnVkPWDxBTyr8Ne
BRQ5K7aDVy/PPgFMMzRxxBW0wQ3nhorwagZD4Q0uoNap2MpJwKzEIT5uITdMbABD
pBBpbIQqbV1SPoSzjFKS7pnyw7P/dL8ihb29ljqQ2IjCxn1A1h9UoI/CY4GF6Udy
IBcDqC3H3usYz/q0wbWwBlR7a4E3SP9prGh/7UiEqK700Bko+7jV8ueou9MQfjmD
fZOKELzY77xbwi9iGR+T3fuijwsP9dUCiMKm4PCRaQN0GEVNzVpOjTrBkLkgBYQQ
VF5OsJMNYoVn/3ijjJ9KmDHYZ9UW7aiOBKJohawly5FAxb/3h3krruKvfMZ7ZjVG
M7uk8yXrPsNQS4H3+/TdJXmaSbHdnqMQV4t+PV+t9AtKsAMvVIxmhEZW7OjFlrHD
cpi89udygSvIP810BIAtISHrUI/LOXzxHnTVWJjLWZECNEQ8qaNNXeUN7NW3KFPL
IRSppi+KFtgjBrua5TB2lZ8MsuoXo0sT/aPnx8hcdSijlpd18iTwu6I9Z5sJzWs3
myveVOto9amjpt4CICAkCwDyrxeaEIPVbi9lAeOp8xiX8wXDfULCoquovmMk/QFT
TRq59uIw1OBG1ZRpKxG2PLKRV1zyXVtV/CVITUOYj/5ErJPC/n+zoDXqob5gzSGH
Ea7b2Esl9QwceTGR2nojeKi8zdOTmFFxxzvrcVgng7NMizxN3xwOdcYJEfhyvoPU
2/NqG5NUXRNyBlskNDkx1DlmjnAz4/bY/q7DD3a0a16NU2a6deItVPMb0wB2G/8t
B/fEzXB0bYCIKX2rQJHDfZ4p/M23UoSnL0fv0IoSOQibf9YxPrUbvuXf1HC5cFnf
OFEL5JepdTxe1dn5OuT2b4S8xZXDQsNDf0Svry6XO80a69MRmOK/AbT9FYQVQhXi
pN847u4Qs2W5z2kQBNKejM7xrFe1nQ9fYAX9+zvCPSwIwQWmTyzko6m/UuxoE3uj
BhoQMJ0Gz0sB4mB3OgDTXW8AkspaDbY186fJTFqBDZhfhMZivg/f7KVna5vRcVHv
aH9AFIXbb3/8boUgjdRSG6jbbaum7NRDesTiQstHWdBlTpH0XXdakKQOO+q+Cdfb
jXQRC8o4+3Bjz8UzuIS+u778QueS2LUzUET6TmrsTAGVNExsKsGMMfSUuyFhSROo
exvsaC8GWcc8LOJxWbwT7dwwchDsrz9Us5QVqQQEkFVijPIZe8pdyLaNEyPu2rTy
dDg5oCmJddyBu5EQ20u6E9azZjulvfJVT+pm9j7uFUwk780LiaJJXvVePcNSGO4B
XViJYSTiHKC7ngp3kPDzWxIM1Md31Q/EuH2fC6tHMJBGz3QXIPv73X67Z+vSa5wf
etIMJKhc4E+LqPUTZXb+Q47FXRnughiiM86Rpv+gj0tUorr8x5bOzfuUQp7eP9MR
VHUrZqy5COYsEAM+YkwN/ofRU8MUu1A9B75aGekSDseiu2gYRLE7cTrrhHBh3Fk0
gGCKkngeB29LZpIq4Oq6y2rTkPKFIspA5N0niGMyTI6C5q19MwvagP0Nl6ZwboY9
2JrVl8wryaQI63+UiGkBFD3dGHuZ4KcLtyA33xpwz1ghJOBFQkhBBrMr8mMOuozy
kPzX4dntCzDIeHX37WAEfUO8o25/64oJSAaArfoIJdlggcWUD/yNLzfi5RfHrqeS
ME7ncg9yIi9Zk+4qmOAqb6fFzhuYKVNj02IJaWV0QshKtAN81r9/jEhjJ5dtJ9GP
RRV66adK0i29i8jOltAxRMfdlAyPlqvYaI7Vh/tIb57ZCZpwj0NuM2y6wiilhoQY
CfBEDX6XIZKeD+PR3c2OEokkIM2/C/iL0nH+H+xFjEMv3K/WQHeHbKL8gO9Jc/pr
oML4CcG/RDSzD/5hY1ciJFrmCWU9wbe0lTiNKsEYuRSqjB9IrloEgyXIHkLQD0bw
a3hiRKMoseAY0vj9m5L0TtkjjJ87s0Rz2gmrmdEqOdWiFkgCjykzXtf6DvB3pJ7E
0ZTjC14RVIi7TsB4iFyDlzKCQHwYv74rnuDZ4YI9O9IBi+PHBQL+bQYDRUfhxrlJ
o3BEzJtWmN2BEr4g3IQN9+9hg3upHnurAn2Dg4wKr+N1v3rcVzAeMZCWZ8OqY6ng
orpO9fr1pawCvJDTemQyIR9/3ER5/Z9iv83vFnNiueUZOcCYQKNGRVAEwfvTmu+7
1OelOZ/HbbSczk9HwaP1+orkeYaLhXvn+igUrpVvydSQAAFQ8AWsk4znJxJFXbDR
XSAY8mfZTzzm7dPLJOuUik2sLsOrpQPZ83SOkg/y0hWeqktTtPSOyuxTWXsrndKI
dy48/eqOtiZ91/rEfYGRJPv199Mq5X5ja6AQRSEnAp3TbGmMyYgcHblP/qNKlsIA
uWzUyrDN7gStrbbTx9Kp0Qq4W03l1VDpxOT0CQ9eh+9KmY5IyGXc8o4D9Vkdc1S8
8kDyiByYuUuSHIwkmjD4F8TmL8QfHEZXrJfAP9AphjBLMwQ56Uj+D6hBdS1eFlOJ
0eMbmFO+EUL/XYsh/t/4Be72xw0lLkAPnX+NCjUMs1aL57ULpfsi5D4xyu1J7Nnh
wf71o7/qh6Ac/ylHNuASyqkZpDGAF7AW1zE4kIZWX8aOmDncSskCuXGjrGNmnRlh
k01fIJxlV/v5Nk1kpgDPyeulrBUc3HO+Ix9KME2yPbs09YKCEqMk474Oo9EbM0jh
ySgCFFfp9MxW6p72mM13oSkRguZFPu8DzQVdrmQGVEejtB8dTMSro2pyUzhExOeU
/2TbswkUS84gl0CxetTihJHaaCM1rKyTrxS74wyx2dEH/wHqN0iKOeyvUBIzwooc
EMqxaRygevXJIlbn89md+VeBIVDbmKQxE7XnnQhVCgIobq4xoDWFu3Y+PgDu9//M
Uckc8kZoX6ZSKmXiyDSZwCsaL+I7I1rZRiqq7Qx9mXuiUQ8z32gLsCd0Bd94IYPA
qazbucwhjiW9eILTRs5u7v8ZT8cuJsptW0LSXXdQoTfu/2GHm2OZjOtqLjK7c1vt
tJupiZAG6IBcOwErAitSSAmR6f90aloESZmpV/yrha/7DGfE06yAcGWi+FhSs2VL
iKOQheFRr3U2vOM3KcMcXnYEPxjhV2TbnWKw48dO4v43zKFiS7PxY9gY5xVz+S49
g7Ac944sdZGbTBa3ZWqdtiDX0TtRdxsvXl26LpESowDdU+m0P3lKfiBNFooldwcc
842ywXHnGY4XnBuogX24gsjABjkweCngsL1830Mmhs7ufarBKJYMRRNkAqzBRcKV
Lff+NYOTL8R/zi8fm4iZD0n5bOpABKirric/qgKsepCXGwPSQNaGclcS/bO30GTj
wjFLj6IRMyCKpGpGeJkRKzIElg66v/Z2ykNGs9rSHFv82j+BwQYY4q2CIDfFx6R9
7GdioCIRYWJxVNDDWdqiu8PNjQH40cLkLapOh0YIfj4D/u9CBqsZ26yzg6CoUXaN
QjzpX8mec0VpDDDwl0+uaax2sxGsCA8Wio/ZIZOaIv72vz2X5u65VDHgW+ZMhV3r
PeETHpMWw3YeqPRSpL6I/dyx5GGPuGeHkFIh+tD14SWkm4QxFWwcGQZk3vJt0uz3
ZNfbYNQmhoypudBDlRPcW+DWcDlkIFrYN5yMewjKLALlROgL9UkLwxWNSq7FYEJN
kxL6EPzrmYIub69qM3IEaXdYsP0lSwKt3R3SdJ2KFxHPelR7jNAPT3VMPjFuFxxj
RvuJddMPTdvh+vp5/fxD06V+GttgKprucCHO/5+yCFAHxR1LNmxjqTUHi5C67oOB
FKQMqjrwL0ULaeTuUCnYq9yruOiPojCJwo3h069PKyFVvtVdNeeDmP2XVjrL/u+v
DW+Fl9RynVrUtzeQM7yCiCxLcWRuCwNdWuoifvkKjW5hyb+Iq51ObUjscp+qO5iI
APlVrPUOMy5MCY63gP/VPl4xcGnOzkRXuDozrCKJqTiMiQwJ+qJe6ETwvWqfGC5Q
VmKSviKfZajkvEiqU0TmGWp2DDZlYIOmIhyRMq0pNKp8aH93sJXXbq6UQt6EOPeO
ZDaL+LVjR1vAYiWSoDk5cCdgWKBN4p1YtofSU7QF2oiRENkvkUiHJKk0EhqgIsSQ
47FRCNfX4Fuu6Qos+F0vzqjFvCojeyjmym6Cx9krnZh9PkihJWDUvgwVv0211nE4
YJd1nysvymTHAvS6OH+gdWtIR/Wm2gGa2rihokZy6YFm4ImOzQLrKPTRT0eq5LNF
h+swysw85efYFNkh9OxGh73JEuFVFDuZZiQ5SlY4GZ32VL3qkXg/+eU1aR59m3ys
ux/Reel6MSSzFpdRHcAht1K/9EVsg2+LivuaGWFcu/aMb1AJJtCynAAwQA/9ZCjm
M+OnDaLbgoHQWonXSb8aozlRFzLLOcZF2FLl7PKJZ019KT/y9ZuYMMOnwFzNWnx1
6M3B/7B83Wc1K6/IsKuVRx/Ft02cfSNOkbWeQPE/ENV49WuvjB8y3fTVHYBrWepI
NGG2LfYW9naogtBA2ZCdZzTelffmAlt8j5BzKkR513q3yoqrqvy2KEqoWTnIf1hV
APwGkRGMSr5UZLKhnJbbbjmenqPBogV2AtR8TPcblCWnSYwvvqMDO0R+NWeXgRf0
QOsbi/GCgg5/SPg/3YMA1g8v4CjkjrGH6+r+ApRPqfBKTxwrJLkvQSfZRg8DA0TC
NoE8ebFmZ05voB1Em9iWh/bnyxkChU+mtjZCz0TjyIJyR2Pmf5DmdrfFL0SxIsXS
TlffKLiOlOgPHhsZjbBFsv/0EYu8W57CJWVtM3CLAczV4VEDT4/3dIq52edIpIoF
BIRIx0hUM9e8LCYe70LoG0zr1Kl+/qaXTb/fpg1BeK4uzGKm1PrebFJm/Hp3VT+Q
AxrvdLh67yz+fqGkDetMuic2s10KlBQc0h2vpHjW9gz39Egq+c0bwGbpNFU6bj19
eavvgznJ1e4bkkJ7WStO8n5yunG3ggyImcbWLEnei7gB3byzeOtfkcdTkHEoZFrL
H8Q/VxMhIDsh1idhdpn2HbXCgUr1wrk0s8NCV3JXqEJ4OvrvEUtGNWWIsPZTWlwv
9uaAa/HZTyNALABsQ/HIp9oIwNTym4SjZS484T9vXxH34nsyexnjOWsH1D96Zal3
hQkiaC59yiFEGcq6fvdiKNPAYC2PDC8Gv4m57fBv+VCA5sbEeBlTS5sM24ppfs0P
8CeKY20batMnR9ChY8rIpZO7EBOky+NjTYJyi3IJRhxDez6K2u+oVjVVqHqXlM+P
hqGBSp1DSG4bD1SNdv1J+kWQitoo4xaWU83kz/DpxPckyOAwfy7iMFAgneviqbd7
hnCleZrcJd4wCXMzbaD17ccIr4CfFmbN3xvr0MUj6PqGYrhq/4s+H9zbutENvCvd
Qj/liSRdRShYb2rj/6z1yPVS2Y+LKk0ELx9civo71A4GDwfRrhUHJERY6e4KM5j3
uZZCzdPPHVXH1Q2JTD5o9IOqZk5D4OAtyeft8lTaL4qdfpe6h2gr1HsyllWueZcr
96XYOSGnsJlZF8caP1YUcl2yGqpCcpa6VrvwPVKjwuPcH6bywcoW5LFLTkfF3cd+
Vlk2CkovWH2vS5PYvWnAAGIextgJVDIgd/eY0NzCRmho0kO+HEOZVv4dynD4wKkt
pX56W8TCw4vv2fdWotMYLvxfUNxB1AgioSFVz8495SJXOuw+PO8m6AZHtKbk5mWM
OpQdw+36DJZYdS8pZnZHT7AfUxwtVmYWa+QlfhTLCUptfYeB2cgVOys6dGSjb0qT
U2TiSgdqW71ehzb3VT3J8i6pFR3coGMo5QNrs/TCjn9gAdh6EXNaHj3Z4b91XJ26
Q4HaD9301towqx8MU18xwCpNPaIkFpNrkBoyzehdL7qmgvP5OgfQe3N2n2um1YbU
s7PVAab3uXB4Z6Z8plAq6h9R169Kw3MFFxzCp3IxEYpn+5pbciI+Yx/z2j+BXUpx
o0yYYlEzf2x2BhYE2kkHSIyeTq9HWNCdsPNxgOrmigvE25YxjvM3R75p+ci11dm/
cImyCRUIbDMBt/LxQZLL28ke3HK4sBpKhRN9S1XX5EWbkvhN+z0eFTyHH+hx8anx
mCBuyCwQR+xcuCeDwmzncrDNWNP0PVAijxj92B9dOO2jq21a8HxQaobjjo3JgJNX
PTj0GDumLumyxo+uJoSriI87wZeQaqSZ1Mqehwdda8Cc7RAophd0PWLMCnsEfqus
koQ2Qd1UDr5ls/prVRKCBF72fy04EB8DBOFUvsYGVAPh/NOuiTr2PTugQ8x72e1T
pPCBj2WHUZrjls6x9I/01JDvhCSa1P2zmviKorWiXPwJu3n8XCacwY4mahLNxMSH
mlrlMB01Z0YxYVBWlFFUtwab2FBy6ee1xjBiZLlTy4BprbnyGzUZ9X5Lg2W3cjkH
SlzN+Nhw++9pYWgrIFjByqZoTbGs6O/ImlsZJfgM9lBL2Y/r4l4h92UgiZfemaSC
E+p3dA/3miuVsP52w3l25Wuj1omMzmXudYhWTgiEpEyP/O3DdHtxw/iinahr2cvG
frBp46zAfnHThl7RUBs526FoMYAE1AqPgm12ekiiV67osnmRfTPybY2I6vvysWzx
XGvA/LZQaglTOTjns4nPAoOmLDqZuqgHScNo87pLy1OWTPjyMgAzN1MgYLuC8dMs
lshIhALGBiZZVRv4ZayOXzgD4KLIQAKEX92kHeuy9h4ea+3ibSl3r4D3p9XdUtN+
MDrNwc4Z0RcPAQjKpKg/HZ/Z2QtLoomxxWeq1LmeClbDt/VJpdJ695oLDrUo/xCU
DViMfKHyDopaH99lVSfTHM3a5k8FVa+JDEE2Dw4flaK1mWe5JtjmP4vLLEqIg/89
8UQFjokYe5IP9BAou2+RqqH8i+3vDF0SXUkWHOZbTCBL1FnhJSp6+fh+g7/tv/kG
FEdZQvtcqNpbJM6MYictHcsI5ivKWBVze9JL5PHKc92iOsmKCijsGlHbCCzeBQx8
pHPIrLA7dqJcx3B/Bvx+wYFlL2X2PD7LyrrOTrzLgEjrAnVRz/li8kRr773wRFzv
Y0VZEsSOkP1GdN3eH9IiPyiXC12YOY93ys8L6fMmy3OWQBWr04s6bzYaI2QU8aQW
LbQZFJ1ltpIlNqBJxyxXhv7PdhgshCSqTL31IdUqQHmA++4krCpAoGgNrdLU1aAa
Bpz9jw1uJAHWAnEiMg4XF8PstFAUVysdzfgOeS79EMbyW7ETCsqRmL9L+BMHz/FM
y8CLNxb5Y7RnxjEZ/TlaCUZb4Jw1nNa7g2Xc8p55IErw/6gwrIxP4s5ughL/x+Fl
uGHoCRImRo4/1EO+ei156eLXhz/w7pQpMq65/PRbjFt6bewk4MZ9WYG/sI5EDUJ/
y2SEtf+ncSn72AX52lE1ckmU2qCnpOH5Row0gzFhcSipwqNCawtalQVwx8YwWHAm
QfrUOULDn0WMF4EP/v8dgqh6Vmm6AuB12peBzSD8vFsGeGW1mHRzLyqN/517v4bb
8kKjKMnGfKU49U7qloqoLO9M0T9zk4fPqvCM8BCASGldgVj+RTLDiw7QA2xgFEtL
XcUqrniALGZTVYoA60ZNgHeVkkdhQsQ4Yha1JtcEdMcIBsnDIhqePwo447F3G5NO
HkorVzJBRuzDdCRfIesww8r8zC4TJumV6OY1SmMssjeY/lqUuBzXle4wn8posyab
IS0iyjoi+SQuZjPjU0ORA7dbKLZwVzmX9BJrIoJZg0D63rxteKNzxaBukyL6TkTf
+NZgCoGsoll73RiLmCKpXCgQhNRwIiQoD72pgBRFqmzxMEHWI18FyipBDcSUehTJ
QceYj6G4CETCyLFjdFIizzAbmYpfdpimRAKlyDaoQ06//k2Rps8sdD1b7qrG6S67
dGwsyM498jJ5C+S6FarTgs86X92zDg+5YR4QIE5WB9JFadt3eCDujzEHxrvipKAR
sRI/fh9qeK/jsAS615Hdc+YXbBBDbFtBr/lPLbTW9EX/sEQC77TRT318tPRpFcOW
7xJ5pkEP8adTbBJCi/SSLacQBg8i/hmtGt5HeMmmfRgeJbWdBP24yy5se8US8kKy
K0fmAipR3VS7npNURvZLV4bf459PH3R11LgZ4yhWGYP9nmgakjb3ZsisxcHXj6u7
63s36moHiHb4hWz+8xMrYtS9LwRzUIMDfZp8jBQW8qeQM/6ZdIbuPyxKH2C+Mbxc
RQn76pvJ5jYMiPPD46aOD8KKTKCR9C10a2TvSiRHsAde/Sl0qguLsJ1fPr3+WevK
+pJi6YiRQjSUWM1D+407REw5VCIqR9Rfnktpedmehai5tq7ALPEclWvBDNT1/UAY
Bo0EaUeC1XaHf6jPeKtO8z5JZU1EYSRZDSYOa5pTrHN+VDkJEggTlj1zq2GtIhhZ
bw+RDUx7IpxbOQytR+3IIUhrLqf30KV6pjSJcCTdlU4M3jeV5TuS0b/nU5l5XTYj
zH4/5OSdCnkPNJUUWY1nM727z/uvR9rbEX0Ds7cuH5CAwasN6fFKbN1rcyqv8KVM
bIiLIi4C5DEvGQaS7BZz/OYsV/ejgeN2vNL97WKygs4Tdb+qFLd5bKAhrI8SsO/8
gyjMVRoaIaP0xjUh6eRDLEZoXvsYiAypHFKXSoRfAZliNkZYgSfgPMMFVOzMHcRc
35z+s9NOpims64KQzRw8CaFK+w73HjHmt5RGJFadsWmPa3PjdmXL6zLzUrgKNlUf
3ri6h/Lcmd/3PSj6VwzK9fdjuUk0EckuH60sRuNgaPU8lU3suk1Ipvr5wYwsGb/H
lDrCYUptg8E6gkV01Au+zgCCtlrogac1VXS8B/qjkJgaaPfmk8Y5w9+zAnIDNFmn
AnWDjp5m/W5VN2VcFHMxmO+IklB1yawYq5EGoew3TVJ7k+jQNWCpIVGaAltOuH0s
vKiM4YOY/9BU/L7eUgYj7YU7bq1PqyPu/2tSnNWX50uk5SN/m8XmUExc36S1sMPw
xcIxXl8JnotGErDWsW+ibpMixmg2f+J9TSgg07nFXyf/MUqMuy+tinhleq8kun3v
gnECutsMrRA6WmB08UzLE2S67+42kh0c/Df46afc2jewotEzCOUwDZ87s9m1Id7l
vKTI2KG8j0nwkWrt5rlOKxgT0nm1KEkx0FVNDwNsTitVm/RA/ZGUylODycczLhaR
sTyFd9bmo5HUE/Vvk4DpnmpT3R+QS0YWciwoKf1a+hjPbDfjMSgmydEKHfBTlHyf
0olBFgscsM18T1N6AyGdliwy6qMvTi6CrZ44JG7os5rm+A73siIoZ9CKEoJkockY
5lwkk3cHL/hrl+I8EXZUhI4vePJ93oXFCpOQta7NlgpgLsM6Bi/770CwGgFnqmEx
KEzbSsHDxxov8epxfSSRiDz4iYqe92gyTVmQgCZr1vviQsz3Jkso/qXdNqOsaDQ4
BCMz+3on7UfCCekG2q6pVDT8PP3CwG3DOLDdYT0eJvgc4jPJtatUuMF+mcopdhG+
XUdqzZFv0on3toRrZbitn3v+HwgcLQOCTM01N+heguHeXh3qsFBwAG5ilOtRv/b9
Hqbdelb47btbsidQHoK3u+0lD/gi9OiLsGt8A9VPXZ0dA9FNSlSM7Tfy1CXxzj+g
uZt5cu3NuCbEbczFBJkXCD0hcOTay+kAJA8JivWoWOEslWrczdSJXk8tBKJ8XX+9
3wDYh7rMyEejuN0zMoyZqRUV8u15RWTMr9wVzJFUdF6uplc23eCEz2CseZIn+OHp
K5Ys3zK5Zjjvwwp2c/OjHa4tl04C6dVIfTJwX3aSaCSLViFfT8zdvB3HcMlnpwmY
+n00QSeor+Hd+5iL9HWbVzPi2IZ41CNjpAnFrs3pCjLwntFO/jAN3cT0ZmPcPvH+
oPn5p7V9SxdnqhsGUqaZOoZ5c+9ht25sphn0dnLmYOvJO+QwHWhC4o20i2L7gKpP
8AbVqnW6JeWnw1f0Q0jpkBDRJbWdC6UtBBjrmaZOgYQVUjqG859N3PmQ/bZcEYFO
nGh3CCXqbT+uE8KG7me2lVmyojr+WtsW2ZZWSlqHKww7snr3VJ//T5/aZHCdiohX
Z2gt77TsRfY1TNZ/cfGVqesFChp3kBCfUbYw3/iAoHokgT3owRci5ZwHyEq/rozz
/AGSjt2DsyWr1wNuJmFVtR99ZPSZA1Lu9uqS8BViDnH3W6XES1bXpzT9eJMW++pn
7tTaB6e9N9sMpr/bYKTGRpA2ZSloomlNV8Vd/wQpGzn90/VuhTCHraqQ9RT4zhsC
YhrA4cs6Zy53WyuZsumUcTj5g3a/6UlEETEsVLTDURe43b0/TvbDmbhIlZHn+bem
w4C+o2saJ/9WzxNG6ifKgTjpJEYA3D8KWeawRkiOkpWtYoG/3qIuzCt/+dSQ8c7E
frgy/+PIK6Frc12Ip8zsZ8XyP9WQTN+aRqc9IDahOX9JA6rvqYknsWhEq9ijAnyS
53nv6V8ijAsjOER+5krVyktUpPuldYULGJ/XhqvmoQ7DJjHqmST/rCwGjIWJRDtn
ljh8TrzkaMdOZZ/uJIUsFQSwedshDwHuviON8BPQGZ2XjRYPL0i4aHYhjHULhILE
333IoIAAsUUhCuZS5KgG63n9jMrB1mqh9kmYuPZXMdo9o5/ORlmrLZzu1aSjiju+
qj193qhc0qZGEKsLeVv7Cmds2COkT7vFClXV//dXVPnK76zGsYEMcfppe32ZZY5n
AhsD+GLVB4Pq81YqO+qxMjcRz9DJPNl62Y1cMBxrGeIbiD+P6ovitXJrwuk2GvIA
MSpqezDyDqJM2yFFr57f5LAIOxCV0KVgU1p0Nu9NbliHGk4yoy1tWHLiyncxm3j2
JXsVsydO0qJ9g+UVuBMm31O0z0HSXSmizIZYVNtlWgQ5Rf7sTWzTkxSRbECJZRQF
vStZyOOyhYbFsC+L6rMa+Ty0UBK+JDEpT66xcwXemIYftpH2vq+rfPKBjcwYdSEk
L1eViA01QREfxXL/Kkmvkf+PqM8oQ6ZC+CdsXANyxfl1AF/RRWKY/zlLuACy67zK
q6jLdkBGi3tN0sCbH+MoMXy4iANsMMDY2828qGAz+A3yxlDS9+oV2dhU+fzZY9Nw
asAEyGvu7pXFz0xaKTVy+MJmqEjmXDK12HiqVFdwpkmhSLnPEAxk3AE2P/gIGluk
mhEv2VxZMCMQ/S4+cY5tIwKZu6nsZgqmEu/88prQYZ9Vb4u7d72c4ig52OEpt696
sb4D/3F+Nwp6p/oapqvWD8TLGWXeNF1mZR6I9LiQplHYgot9D4lirjXhxe/ndUqz
+N4/WxqLNJZh9B8aOsWoovjGK7as4XKRg2+aTtc7PkD6wwN2WeuiWkSV9XvmDwOC
2YvxCuR/RrOrFDfgj31Afass4AGnm55W+/wZzVRsG0f7EH4aSHoqrNYLemhoxjC8
CXwbsrxIx/24nQ/eXatv0MEQgElN9fN7wPxrIfdFoZudW732UYm3MvJXT0YN944f
HQrOuth9fqs6F1mC3Ljlszkg3h6KzPqVlCG1JbLoYRzQYckUmmNFvAM08CGI4L4I
jdShMxEixuhYu4AoQcTebypwBPyTEKSSsz88L5MdSLJGeq82a0kQRdrf5vd3RdQ/
b61WIBSYw/DPiTVIRVQpUcUufTNZ6ZjJntChlKN7GdXbwhqtok+Mp9HdK4jDtwzU
iy1eeSLjIspIv+kcf9jqPpJL+YjnvdH7gbovuDeebAzbbJCITY8QmD9dRLBQRvdD
98omPRjeXGK0y/AbuhrbqlpOHcyNLWZIyAO4OCcr41HPT/Mfmke7rCQ3M1XlKs+I
lDWMhH4lCcVetL7GeEMBNDNrDbiYoIFqaOjScDOYh7aCztRfvIhywaWnDzYpUp2j
aPGC/3eFALTBSAjtjwx7gl5LKSKD7DeKX6RUXXHk/YUeOw/We4U4D8cxdIfuzJZ4
kqnXOnXzdDg8qp7osffECy/SMLUL8Pcx8xL1AYaEIfQ4PusZp/fiwoXj8PVHsB2f
QY7Q9P9FF/KRcJWTwQOJE//x7mjv6K91vwqrPDlcMeQJee4LdGQHLr/aXL4B/dRy
dXLaO6BFLTUhe4w68boc3uxtkXehMfExHu4lk8rJVq+W9yb8PqdumjaXqIBXSd3Y
gG29QS8H/PfEv+nDfmpkz+/DU4PFUVlWgPggY6wXLtaLvg39OTwtNzPb/DF/AWH7
ybJCgmD4GMXxXrtr0g97Owh15zQeK85IjOoniihZLDsGmTu7UtTFxeWt5dJEiAY9
bfbchhUET8Vs6nGcvJqhQoTx51n+qaWe9bk44m+2lRxs1LvEnT+NU6aJ2yxkrnJ0
WkQfGFwYKwwhoZ8yPc/Wx2Pt3ZamBEDBCXSgCeyq66ymDxsMbNAvCvfVGZmFsmZQ
xGLO6DdV2DJsY2Qg7LtCpVkYtfYciw0UotmTqrZv/ZyEnfa8aSxQZ9qjhDpA0tJH
eERW3QQ/Yvpwo/BBNR2pzWC3oZtbQDmu9LA1BEEGfdabBSKFIafNpG18jh1Ofo3M
m4uJwqzJxZI0BPeNYw0AP5Q/7PXxpAU3d4lEQEqTviYiOV2FO5LyoZP9Mhq/uqVH
KWQQJ+4Lhg8EUMxMnoT0mR9RA1EKY6tSaosbpRvKoYRYIrQyxddTSzhKxaETmOy8
uYW6eQNp/JjFlLNUm9G+YKC9/Bxyvh/yITTiwTeNFaXxWN3+ra+a5HcadXQOpngS
yAkCc8ZyyQPmcxLaBb5ww669wlG1TGwK8TPwbwrDuHBKuwT9iVk2Lp7GLChEw+y4
1/VWNjm1qiS0ahBC75a17j5IPt6zIU/mnrDC6xbmgVobestoExjNWZW0tY0GNR3B
/JYQJEt7Un/kjbWJMIwJPlWCiI5nh/h4ohDQczth9bpQobjxWweqGqqykKbpF14H
QT3/cRMtZk0cY7jbZVmhDRjmlJ4nnZC4wLGKDS/xE90ZWL3M8QpzeigCtWyOJ+K7
aiRN+0J2paTBZWG5Fz9G2Gy9yQfmOgfhBtshxmm+tUDTaB2pnqNUDufNpmRi4Q6B
+yFS/CeUNpBGxznQBINVQL1kXGLteilbE1MHhANhycTnFJ40Bbx3Zy/4ORn8d+Ne
C3xZlH2Emm1w2Hzdj17VDl9kzzT4Zu0B3GFWLwp+QX2Wuh1odNzw+T7WLEg0/jiH
3QJVtJgyi74zvv+zA4ofFnOdPyRvMEZgXjKt2c0T+6/mILelOj5qzeQD9owGLP2Z
fe7NXoqVpEbEcMolQQ0FjWyngYVxk+XNEmI/x5TfWd89Rxwyxp+yqL48cdcvXwr+
cen++VZXYoulZ/p/wlCVZvwK0FWPTm0vsYiv4tw64SV0c2Tua826suiUl77S3AfA
Dqi6ITSczp+wSNu/N9K1VmTgUWA37jtloZvWbFc4qr1d727H7dzPkSZHGbpBv6jW
O3joaVdgbXbXie/UZzDzq5eSJc20ucXWph0RfPWClxP5sYeXsA5K0OaSIGVeym9H
5ZrLVeJqKo9Vz8uf+dy+NNrt9YOF3A3jiO5ojWnyie6uLEdWY9Xqy2ML6QpJ9E4I
7/2XdXcHR8Eod389kJESjZhKeJb/1PAY5l+Kp7XJOJwRh6O9uUPnGlinb27KHGzB
/+YGEiOSLkFK4f4ug0lY0A/Qw95XX0+3UqWOCQEjdfIxFWQdwZwNYiibY/qpGmZa
oeh+w7xJhGGuUq8/6lBgbb74lMZw6VtkOq1wvlNnJfWl+SSSEplLYRwFMF0+trMb
AoivXEDJ6219632higusrYsfNhBuu4Ch6bqfrm7INsnJl5O8BLy6NL0FkKpnabgt
bzbH6jPX+zWUQlpwE/rtbW/JPYUDHV1eE3pvN0hSImioVY7sGSWEsIs6sQcM5UYr
uMnChr9jxuQdCqGWEQx3jKC8NhkB8B+lHuYxXjJd+PXQ6wXEM0wgP83JpsQzs3tV
kES/DsFzbUoYc2o/rRmtYpj0k0q3TKpCF4paXPstUxN2eTTKUs3TTwGJhAI0p5jP
CEoR8D/8CKBffxMQB3WcFMzLyA+zXSChQeYiqDcwvBKAREoZ0leNlOUhXGckAFrx
ldHcQBSziStKNU6slUPSV59rBBfxNiuaV5xyb/thy8L3o0C4ay9Rw+4Rng6UM2rA
5nJObLl+tpFunIXOGOarfyfKxhtIfG9lAxx3lV9IiLGEBXiOUWu+OMa1bGE8LDRE
zxFR2VJS+bOIpD9r6h5XhZ4V3+4QLW89ES27FIyJmxs9XZPIkOzWmZHLtsJM1H4f
ooDvQRX4kMmsjfeTrAkrV/sE36bhnXyj01/QXMaC5X4Gx2YE70dRCom7TKWmZI2t
Mjq5pssdIqvBdtWes1LLAUVhLjJxnKwkH/JjqvqqhLAb7OIColZhZTM5xCiK5C5v
PotjPmvyUi+Pvu3ZtteCE03Cf5N7a80UkmdJ0//uMzkCup17Xr2tjKAOtmxSxGhJ
7bvnV4GVqisCVnNN1J1lT17m0gsEBIfgjSb7AWjsEig2N7MPz4E+7Yk3Tvm778HH
89Eq93RCp+draUfXJtZMV/pT1QyVK0EiTu0E4qvJCZlPsfUaQcVpglTDFz732eBP
VY9SM9Rcot1JkDTDQ/fGTdxCW7nqT3t5F4dP4HTaD6OBeZNHXcxdaj1Eo4mldv0q
CLCVVKZ6pC1TUIvMpyKQmZM+g0UpCBtB1ZB2bqyIq7d4G6KRKINk7zqjtCnU2ETb
+y22zNbGNcfKC2cx+4//3IPgSLAMqsQr+mRUsrZSuyGAkrwzVt/3JnAjql0d1aAl
iVU/bUIthICLmnDaFN4H154O5ZkE+RZ8fXA/5NSOQ7dCPgR7D+9QEZifKmBV0aUc
U+LqJ+vvQxvORRGhMo6f9l4K3gPY/3W6Vrj0fX0KIS+NplVkRl3ZyiRM1Xz8pfJz
YCGW3aQn5SJ1gRJlqg7Nq261GJ8vz9btwPd8gHRAMLRw2PRl5Z53Kfwzoh+qVNq1
JiA+qqJMBVV5T/5xTpTc6LukhXaPcQITgW8rCX2/ZS6wzYIoGrEk6h2hpFxHUL+H
jZCrZpMc+iBpFXWIY8EI6TM6tYrtpWgwm9s+DRrO3UQRIgMvSLl6RqXq6vgMjGTN
Wm5pyTCdkGUML8+HVOO8KGG2EXRsely3ecbR8qIF0LnyQzl6A1xgnJY1Oi9GmwtN
5Xsr6W/HpazqEc9OsN5RKjrfC5shpQDpquHG/MBmctpx3InIo2mOi2g8U8dwmN+g
017Gg9ekDgAus0KlUWmEsuohuOAgIt+zeBvTQLTpNLIZwG1FKp0y6Snsp7jblMY4
ZTUuswtp6gvNS+ST7YqolMmppbH8MOdHFmtExfbbkJvowDY7FvvlnOmVtEM6jPem
4CXMT4GIxXnLQP8fm9UOLb4CpUe20n27F4lnCsj7FRjHjDoW3TnbXmOt5UTlYvjG
Tkj0cO+7T8ZuqxJfHOAT29tg/8GgxzCPxwB14XmtXyorNa61/FfFZ+9lGWB6cqeg
Fy8f1cCsvtxblAUhOIYqDwHl5EJjQtwAfGG4ifOzEXQVhUo0tPAMxgZApO6gGGsX
KI6ju9XlFgKMpIArX3yq376HBMfHYZ9NDtDrKA3U5fF0CViECOxLWOF2sbEbcgvx
jtWjYf9hKPJi8FBWPn26/OTHhrN7VzYBLjLx217QS2ZUiDNEgYcYdm3wsTQVOsAP
uoa1CpoCjUIIEs0fu3y7vFRHyQynoyrJkVBC7Ipc5tBw4fP1aQQw9ZOgSdXLP59R
e2ZMMr7mVVMrFFsW04eoKxcRbqajs8q3fw1UVReG/SfMu/kZ3/Ez50f0z8F1YU/b
t5T1rxuYeZtEIQ3ogMsm7x5cSs6qaNDSoIf8h9dX3LzsON4R7xielHpyiJdPKYSq
mq+POqRfqtFf+LSLcHazCBhu8CLs0V+OSHqTf8uMMkxwTBqI8T2ujC2hdSftVdiV
cjLu7R+u2ToSbTVFG5V0R2CC+oY/B5c5EcvOnga2qQRfOcIgLdp7b+O3sl1J4aYG
rYAkpKYo4Cit5ahafH0GcmypB4hmtrr49ub9ZupU+ji7T5MGfSyMUs0L01QWuPIy
qqcnUoWcGIcoe7EypjRpUyCFbc+HHCZ7V6SZwNSVBjDYKJFm2hv84BptMj3zsoI1
lNSF4bYaeNdl0rE5FUvt+J0hMg39XQZrz6kukJX5lrMNayrwSK0sD9tQrBi+IxEW
zIxoFKK4SjWvh/0cmCUDPjNhONqLxeHRUYXTSOPquofWGDsYOKIVzvrZy6SGUAQy
iuWiVG+P2xgb1TMlUL2v4WsQCrKyun6+ohalMn1FDFUJiNDRB6N4OeiRYRGe3wEL
1/RC9fTfUP6UJFxQaQ322ca6N6Aqv3RwCkQ96W8AjynTtcFCAj9UB8WrIiq5l2PK
LNwoeoiO251eq3lOfW4CGw2ngN5GImTL0HYe+I5iLxpjKgsz5mx84xRmvfD8S432
pxA2ZvtI58y+Tu7rjmfEvUlOvNh4tiBLE6QzRWLGASwG0qbJOBrNUkMvsewFqbl1
8DbjDHZF63cKrbMJfzKvssJpmp9t5fWRY9OSElyQ+9ktu9RuspC3qufnhu5ZRMog
zXZeuesxOQOKFNfc1T4jzwYJFeZjGIxsS/Bhm7KBb+Uho1lsAVO5v+Gy5vIRjQjD
PM1pDKqq6ts7XNeS8zB+gIdwZMtpK0jMleTeWgF/1ObzeU/WRcQCEvYmjlTYB3Gr
kfNAC6AHS0FNc7dqI/+oQjq3GUvwszeg4uY9L8iP/Mt1HuLoltHPU9S3YseDmIou
Bfcl88bbGP6i7KGU/eUEpZmIlOJYA7rJcvbK0MwYicYRkUZ3GGVEX4UJv4SzbgAq
+X4clRy0tLKbeGffuqAo22ldaP8mp1G6dxUEArug7pS4Xzs8VG8nPNrEoJqTZz+e
B5Z5lF75820psDCzwI3PDYbu8HLEh7xJs55qebfS1ItA7a9XSp8ym2n3QRsUIsre
HI10PVhvevEDhuwNo1zpP/dLsHYzfxRD6N7YHta3EgYhXdOKCojHd3ex5nZ/2vJG
QKkzKF9+fFeNL4OK8EoEf5exBjSCrMQIKlsCYJphtOCCsx33EczKQq+kqm24JIYI
yQLQ/uAPU+DQGwEqhuJjVC+PCaP8SY5jps6qcGNMhPZ4/y9UvfBIluuFTn7vEsXy
xMGFsceolvu2QMzHA7FysnpEqb7X88B8vUGOqgUti7qHXoPHygc1x0ML/ommhKmt
QtqVyYjEGzCbYp77GirBvSO147ohSLKfl6uelsxGjUVMrSo19TEc2LR6EARcMfaz
sW7sInx4tgM+6o3p30W1IzlTSgismL1E8SqkW5RplXB75ISxxLOcPdE1hXqwHB8A
AiaT7PNsTUIuZxYpl0ibOy1oxWRRF9SyT3eAiy/21vmBtOlnurfexzuMB0lhL7vv
Dfgd+D+22s2sAzHOX9MSMcrPwJC2hqVCWeW4TaPpsGkeXhdAhFkQk5sv67aS1bLk
lJjz3ElfVsOGOkR6Chpit4xcdxLRXMEww1l2n5XoP33W5tN4SQqSI0K60T6SUZdY
mBy1CaPq4GEvBPgCU5aJnB+2M9IUiT+5viyiyTkdMKyGybRCuh9UF097qDfuL9kM
ooOyTN597gmZAhl6flD+aLTHgpzLaanIEs3HYsNiHud6B/kofYj8CpPkVs98Oylu
p3fhDhEAEd2GfQJxLAB+h6mr1Cvd8RVI7fIxb5UQh95DDKZ+1UMelV+TiM+kgvQH
gcv3vO6ayduqP7LABGOADbAdfa8iNYQC+u9gzCQ7tUSHyvOXjMeadQ+s9FNbqqzU
DuxMTntQd5lIxFpX8m2E6rzkQo1qr1T+UdnXfMousKL39Yw+iCkDThzjc+ad/hVP
c4KaXEzkOTTdoQefb3Agjr8zsIFyn4gPT2ZWB60qv1vNK3Ojbt9jAgTiY2thtibA
K4GlsFixW4xsXq29C1w93qh/wT24/7rwVv0zjOqzNRkRVLKyYgsGtn9oXQitSsXd
GYy5jpbBKXSqPuhZtg+aGacPyNXtL7qnyzLDTDEfWluL6MwSdfLC21bsvik4RTd3
TZGNTS/oRkh14G73zqMe9xEgolziqooSau6Bz/aAZFoqCH97WhXdwbv2z3s6MrnE
L28SilcGBc1CsDUHlhSA7NId5mqSP/1fD7HVd1WTxeUQpmKCw8DsUtD5KuLiXcxU
TAqG9f32GwSSnor+jtcp279NQLVyWXBCB3hUoPxfQUW0QWMvXz1NKazox1GL/kpO
k7c0Y2DsajkL3LMYyiDg54ob+tYXW/t+4p+zcd9A9+3xTQCF6qpOJfCBCyXpAUsR
21f3y0lrjcZ/Ivd1pJtiBp2RRDtffk79BAgK1DZMCWKkFHRhP2i7ewzVFunLrEmo
R/zhleJV+NGYtsA0gKpjoHLlDMtsV7gnmyOseXx6cQ8UjYCfm2xKIaejpd56oB4T
WU1p+lGBRodun7HMJBpgTX6EcFqftLdbdNYJ0THEyoKL32nSerpVxbSgl/UI+wfp
d3w5UUoDMpL6BUMvKTTfRIJny9pSx3E/ULpgeWVNjd18PDIFdJlOhIijmBISveiO
v9hn548lgnJ1fBIGdJ2PO7HE9KJSWUCSU+Z1i/TC6eQGpqzkgxcCZwOLLeb+xQX8
Uq1H2aQqzrfjuREuCg4WcZhKOfgSwXu1ATo2DUfpyMZmaNUxJ+n83rRBxI29fMR2
AeqMwToP3HmvMifUnGl/cLyrOWrZzuiz6sA4sY2ySV2zp7E4fIjTNGMXWw/hHMRZ
dR+mDmWia1OOYBhonGUbIezOlYZTxeH5wf2wezk44rxJC6H1li/xq9dbApFR9Yoj
9D85OJqvELM0vRXiHmc3/zloGceCbgjVQPSZLrFd0j5GL1vXXB2KhddhhhX/Y/V6
s9NiIcfPzfTlpO4yUyMxIiSzqyqOt9OaVqkDSC7CBiJaV5f2mSQYt1P0/PKUwIKD
3l9Bkt7ijJxhyUfwLWchiulqEJuXRK594FH+3P2F4CJIWAgtjw1y2DqQkob6v/5h
wKQJHH8hS604boNA7v7YhKuwse3nZrD/hh+BnQ31lettkh4bnNJr1eYJ+ghhjbEN
ziwhbuDWJhaTLhtMwkeIpqbx5glRvGWTarwMiTh8WpAMpqQt1OfX+VCVXp/Ovi5m
RIwqFvAHsgGrQY9RyibClRdB7bKDTxoxssPQ/+rSeY50sDzX7U2838m0cLwocBzg
V3gSF+h/YPl4uwAwxy5HdUWb813/Zq5JREhWxLvEBOSHWcUcLn/6wfzsH+1+INgh
HNvDzj5hKqDrLVO6nniqCqpKKwvifxXlTKoruVBCGUhNwApuZqzUeurG/7q1o8Zq
OaCcFLa/GtC9FGuNj0avh1Kisi87xvxYphUGgPPyXhs9pWeRybrCflw+BPE68Jsj
jkVWksNHghvlR/yXZ5lyJTMFhg4X7sPkTkjMUn837M85KS4bFDj7N0mb6M16vDo/
Rut4FMhfIMT5FeTF/xnUt9lXuo1pM0jQPMzKB7ySR/GzpgNuhpzK+CpaT/5OCN1H
cb3HXWSAt6Ew9Y5ZARtYMoW0VGV9pgCh15KqDjxktWymz2FgYNT6gcOI8Y57RS08
9nE/rrOHLnaK72xv8LfhDAaMX5mFZ2jpeTzu6V4XHL2hF1yQn93u3o/+B91oSYT4
M9ZA++snZAUZdGK3mTNnqRoiPoW13Z0CBB76R8lsBMkzbSVnbe/JuRuQCNaPL3Nq
tCGj7cb1dDOusvDmQttR04e8wkKM94jYBt79e/yDnJFYGLjk9r9am5Pi72GeFZiv
JG3bW9lC1CdyfuosSc7R/vMh1CvPBF+l5hNj8VPK/ibVNDQ5EADvg51C+b+/jzmH
0NoeQYhrMnZ9ZI3ImAax7GTqOT6pj25ZrCBlE4hmS8w7BLUXtBCfYLl1V+m7MMVh
/C/3rD8bY7BOAoOo0sgEdR7iDh5LgVrbfHFNZ440XaayGSuZyxWpvhuoWRsY4y6C
/XjbiG8JpmrBsu2v2dyi5FZO+YagIBymqc5x40yRKbNtPymk2BE8oT/iFsWAHb/A
hjzHsXKgDnMtUgRydcnKve2mCkyOnNZQsuFKvAZ+DjX1XOVDOCObyC3TM4/xFFA9
4aMsXp/HpV6M09nbufyWXfFefxVIq8fUSOYmpA/asYUPE42TOopzV4q/d78YaOoI
iSUWXRHn8Y4YeGlzM99VLawaIsaiq4r9+fJUZyDK4DmD/wwntfvzicCYUjxrbbUO
WRamCRtSkdbt+51tFGxkba55/52W5SRipTrdn75+oBUITOgJ67KagBYCiE//UTez
QyzP3DaDjJjuLqJzcWlxLY04elVJjMNh3QDRjZ9wH8wMIn+cXS6aMoJiVK+Csdw/
jv53QRY/BqZDEtSnWdmBeiVcUPIuPFVH89otE2+4FgyZT+mOcgaI1BZQ8XwIwX9p
PFDULaJmR5PEDRhWoO8NJGS+3JsV+RQU3TtEeycHQU1yQH2xy4Ckbr2ZL0jmsByf
0A8KcqsmXn3bkR9Lb2CsxQx3FXaG5gJvjp2Z85Lym9i+6le2QQvXTd6Z3UyPXIH+
gIO7v5Rjtj9RTeCdceMcV9nnYMLZes4c21w/kPKh/nzgQsgFedV/995kd/B7fdHP
/iHgUY3cJOkk7oHFT5At6bva52AxoyRRGb70YOnjOqNHOIRoS58RGHxG0uuf7A7O
jeEYbRBP8ptT//JYSx6EHKvYQoI3SCFqlNhlRX1MRt5iSAi4DYXOhjN+UsKgerTe
RBfHUFkVfn7lC0WPOyqxHyIuWW8o5QBwQ1EFSor2pjIb+EfOrWdknMx+5SL6A+Df
sSHcpd3mQ71B5ZHp1+l30l79BhQhFIGlmfZhSbJP6PAkeXEldG+Fi1Z7iwrkNirR
yx8UUoSzFWgpqMGe7y6+K51vs8gTx6QE2nBAbJufSZWjKXO59p9oE9yCBHBA4y5Z
UgYjqebSCUo0UJDmgzwqGjcru2XjopewJiade4j9f//XRCm7opHjMgG2BcjE0be3
JxTqisottiimjMwE9lZcHH55gtTh9y3a2OA4GDbTFKjwM3uE3F99jXzhOuXoYjv/
56/3UNYK0nF10gwaWaDIbmsN3ELLmAJYRpeGJ0HbrOcmg0BUHpFJ1+ePSALHI4f3
8zA6emcUREUgtsfeGxzfDsv8Pp9/plR3NnGxRKnYCyHBmKIoBSAWd83Ii44X+zIa
vuT/2CqF+0nJYMio7jIMIsSX+rJ4TjKjO17+apCKZPTU26eyKcpdajZ0oHcinkWw
hg4GoaAk5bjRKZYHH9nfwAZ7Q4WDr9S8hSw0fYiTl29Kcpd7I+MVc8fiuGjpp+tq
tbWEojmWmkdCYZLmsXlm84ri7gc0H5Lr6AiPFTkS/NxcUFMp7AwiuhaP8P2uWE14
kB+hQNDFh2flqkl5Q1+DPQcCubiq0DqfUpT2tCfEA3ANu0jHa7k1r0kGX80ZAU1H
gzQfS5b617mNZ91CQF3ZDxHk1R9kbRCH0pLRoPaqQZ7wyMPSqyur4+QZiF/aJ3nh
HZYNMMY8FxXETLtux16M+EzJixYrIkS5pwSqKWWL/B6WXR1oJCtvtgTwIYgktPAX
pFNNLgUxmWrxhExTlboS5q+JCNVjX2ELkr7rM0i2nOUGYV2kCcWr2IsYLELVVWLt
VdSF1u1ZOhX7CbvByFabs8oUJwvUuN3OE8FKFKX9crkC5Ad2S5ClVEMhwMNUWb/m
LMQiqtgRrCR20/E+6y0lQuFHJ4SkhRp66NG9Nx70VSnkrefyfGvu3MW9TjVe0ORI
J0E5hrCfUUJAd+Kkf5ehp0jumaGKBuukhN6LHmp4PvzlGoOsFFokWHdymXNLQrDi
Zx7SEEPMfc0ejlAWn9bUfUKXyjG/PfkXLv9FunL4mXvCGC4sGYYfCpWzcAYlKYxH
54Tj9oSTOrCOnuc+nXYpzAmidKI4jEufcNVwvAKcBk1K9jZ5/IjksvfdtVKHpuoi
tg7XyZ8J3fQ/u8t2rm8hk/h/YjqQM21LHvp6zU9qqGTrIWMmyFfLetccUU7nkEFy
I315q2DEQ68o7dc4BbiaekZaQYNA79WDEZHTIENvE3yMXzjSV4PS9aRTLvX5eE2j
ds3Txp/S09FQ+JbEwJFPfLiMl+Agg1/ANeXSLi+Cm7elHXAaor1+gAmwqNuCVeE0
WMPOs/6DUis4Hx3NISbvM9PkeHPNbuROSic3W3FzXDUxFYbASGqtSeshxZ/ad63l
8p+upuUnQoahWGBcP67cn58wwtOAMzpU1DspyO0pbjJSFuTpp7/quInwACgOpqCo
ogKRScQl0Ju8VuiZO5sn9qxLbCaLmQO7drv1xtG8P3Dy71R9dCVDMbBK3x75hV9k
01lVlZ8/dwrA9GGtPzp19nJtMGcX/uqc3PpXzmOOQaL8dM5+HN3O61gaY4b/pg9U
GwtWt+dabZ7iRw/RgpsgbDl+k2Xe41o9WHdQm8V3+4HnjyHkq5RbFj4zndmeFIT2
DiEU+9f0LBCUD20nJp+ErarZFNv15yIklGfrIR1NHcSj2bKoQnMFxshBOBdyKn/U
/2+WmxuDaJofompGDgbqQE3N8NXSRANeMb3trXCYKcUq33+hStz5e2tS8OKk3CwL
sUOG2vJE7BCxsvq+4xCEmi296CgEkBsdil+TuQA1caQThwuZRxLBmFulzJpY8ogQ
EdwuvuDKL8jPtzcxj0vbUIpmy5ZXocjkAdxm93KwrIqlp0kXyErUa15953zfmqvy
QLGwO6FQvCZVDtqEGq6xN23WGwhzyffBCU6x/C6wYlUUPL2ftcynvF15j425RPFs
xbh9E42yQCaRyb6DRwTifD2wEfBZVssXYg5ASX5FiwLfWDG4L2GHmcmG2t6pi4Sz
UZlran0MttFUhSFMDoaGHQJnuHvWHi+EWAj3P7l3fMYij9SBJ7W5Q1k2wLRrmgFX
KxGsnIHSRBg/UtFWITOqwOMuMf6MyHJ9G93q/WXzAeuhcDxpEUi8tFNaRdwPrzoh
luxoe0d6gYHHkw887lzs/XPa+U/Lh2SAe2VCkKMU9dNMpnBAedKtWyO4JBDCGero
ydfV9qZb6XNCS9KUlPMeX89U8laU2NCQH/rIlaDwsdVrEbhjFUYC4hYOpXhMwB+G
3ZqgE1u+UgmJbG93zkiNO0ArcObEflm1sHZEDW+kzKBqNk5dGkLauQ8WHqCWb6i0
C/kFcMHQI7cU/3kB4mH+OQI14y5k9A2q6dIxaEZwCakocQtbYe1XN8J0CAOMYw8t
0Z8+CbwzaIP1GvZYGnD+F6d1sxwYmcgfMIdf4wL8FOJdnZRF2fSUI5cHCkDUhWS6
eBWSCQEV/TiVjD21m0phx0/yx5DYi6RAgRww+m2YXyXwh2kwUolXJb/d2YBJ7v/S
RRpFCauAaSmgNUDwHxi3OGL4nSWzN7R+lelGC+lOtCed06AZ/uVRz9PPsgld0UmC
oX2ZiRKHP2HgeiMHq54OFhSfj8vG0MISSaq/qUf4eYpLrXbHfOJCll+Xw+X9jZ8S
zEoveKI0mRRcxTEL69mM/jlCG7+7R7aOeUyPyKwzeEbNuDG/4x0N/WCijieUEe9u
pnioyEXHCQaxTQXimkK6iOOzOpv4jeNfpmImoFo5J69R4RwfOa41mmGwxFdpkF/4
x3tf1p8aJxIYBj1KTg7cHPLWLN8eu2aZL68pp5eTlij5RnRFc2bL6w/oVepe/ZXj
7xhndPbc7DfE3DqttJ6X6fmWudgBzQ2/quErocnHr3OED5Aa+6+7WdXTwmn/g7hW
8eVTAEfjZHtLYi7hPJkMlc4R1SJEX8aCHye5DYQBs89Emj6v8jf/UCjoxZ/cM+8C
tV8TAljf5Xpu1lrx9CxeYiOAJ9OLEJEE4dFbx/cv3L0kvFEtCwny7eVbhU0qCIeS
m2rOlwtoIvQJ4jC2Smi72QEXWwdJec95xGXJA6+O8yxleBUJSedF1M6CQDlvNCqk
OD2NlLyMSTf8Yx71AZk+WCDWM7oEF0sNjd7dnJ8l9ytdcVrXIb02X1cn62HviyWv
6YJRuEWjhm5FJ8uywHwdY3qxx7Px4WqxdOuYr2sQEPp6QcMXHHrvwf2Zxk9fRAWx
M+bcv5qtp3gk3V9mYXl6h+NFKPtGEpGg06L0QQfhI7+vs7VnZ7unzSPsf2sZ6bUm
E2Pc7W8D9MzcjQad7XAvditzbwQ0LtMIg/EkIyGFU/prcm3Ux/XL9h4CeUcGrxd/
iQTsw6nIK02+xZRLGeK5LmYR8vVdUpoMjCO/APFJ2Dl+qVcN6jiebEt608JLSf8f
2+zPhK/NtNGyDwGkyuMnkvBBFZbwph3oYcjBHrrIGZ7pxDszCil7ILAxojwCGPx1
6nIDk0KcYlaVk+RY+S7CjQ5I5ctjJL5e2e6CK3zoWEHstjunXRdiRNieLvCySBEr
B3Muwsdi1AWb4twG+oidirkmpSQ69gWyVDAuhnifF5Z88eiY+3vgzARdh5IWmaZC
9+4ZZEvJl9DFaBDVI7OvfNNbHy7m58+pHMuKB1T7AxhfaUW/0hrTN52W5MF0EfBZ
7z9ZttLF9hxD49uBY7QKwzs/ZBGyh9iNOmxarnRxg9Iq7k78ZJ/RctHoS4Np315x
b4hCBGe5sWszUllc+ozzyj6oZ3gS1nS1ymESuMLqpKoSObUwOVDQ+Iw+UEtTX/MB
Emd23GNsuEQXqCrcHNw6zP3ypX+CjPB5LEJxiQuN59E9u9uQ0xOqkd74yJRTSsks
j350USg26SJ0Sey9ItuJdlgaGKqGgZvAEqE3HwdNa65wp5GznEjqSzU46NHuw31R
UEYwmGCbvhrJXPjKXpFB0wso4OpMN4fJQmCrHwIvrhx5VOx/Secupfpo9rRuCB3X
W1e82VQxHvkDFqkgzA1kzHFl8rTlRGk+BywBvq7DJSz4HKybneAwO0LPgT1rO9sT
qqEoh4ThQCUR/adwylZoYO5AcjxXGr0/33Pg2caIRxvxFr8B0/86xojc0nHwn/dz
StUBzU87WpRbLKWxUwo3XD1+TZbFnOzd1d24YYoA6Qsml0ehh67qYguYn/IyhJhi
kO7u58ClbX5LAUkodRAZEiY0k5UZJQBz0i+oHtT1OSoHqQCDv/H9Jd2XdrJIm1Jd
2D79b/DbCYYYe2m/5vwlKItxbT0MMmwJrsoWbn52C2SKHnSGVv7t/pnHujYxZC//
eCAzXzGysRlOpVUzlRgws0MX0nSqhxahW6jmirPftw49Ze/zpckUMJnTwmxickDt
lKAbMiWkk3ViPYhpMQz5KgI5XMTOKnn50YJSSekCfRMMIcQSumhAJNdrK5rebtvM
TcWN79jQB+PJmka9r3Iy7CtgO+UqpRLeKamRIsltkp5LTuU8F5zdbEQPuiMiYraG
556dtB1iTmQhctmWjk7h3xriWRDtu8SSKFtBdlgpI7wrgXbzVBKZev3BJliTZCny
gLtsheNfKfZCBvPlCc0OYUSA/Xu7iXKc1t8Ua4MpG/LELxHDEjbDqhL9itRaztb6
cT4Cs1dxOGxZpS37yI2Q+ac2+mhO9lcQI/JANXRWQnyMqsTujzniWmrg/InMwp/S
bnCogha9UfYKFkpfw3o9AH72feJatWsCcFS+KOE6k9Yl3NEUVMzazxW+VZQGEkpP
9cYWAZgEo+KeT6ywg6LYf3mWUHq+Otfh3fLzZupI0rDY8mU9pFqWvYO7rQKvz4PE
o7431GF1DuZDRONARP8g48/4OvD1nLlZORtybgpcAQB2TndyVBm8rttH59OaaXUs
MNR9bP3+P32587Q1C230mKPAL34vmWKFxzpsrnRcDdXMWwSggdZHyee7FcuwzGQ1
RqjUSn9B9mb45gvCtnYyMBdOAMniA1u5VmBMuBgbe0+unTE433lbj+2mphhH4Gl/
UdhJyH9vIT0vZg94GneU0NBxKKSZdfcww3XzkBDet9KLjt1fsoYHkrjh6pummxZd
FZXTjgO3WX+VyMxZvNQaDEjecXoteM+sz3lz8A8AbYz9x6LYB5Uq6taLhfAXurJY
RTJi7pWVEFVFlIKIvOD87ZlQqnJWJkdxKp0nk1WLJwCnoEt4jyncZ2kYOIWnDsRb
1/8PuEaxCOz/h72uogMTUdWVs7OHlY4OQ0i2i0QJcPckkiHpXlT5iCsaTHxlXR/B
yXfr0ff9VxfUOJXo9DO9Mdt5Qde8ynkiY8FoQqOlXGG3tUdr90ES1nrqkm3AzDDj
jVRMWmr7xGW+N8Y4I8/NXknY/5qvLP+iGJA3S9xRwpDd+mXtAdR6DRfQOZnrkLHl
nCkNIGr1wL8Hahee7vvMnrndgD7deJi484sACgAToN/RyHu9W/yws7IMGaC1iC67
gaVuMs05nOGod2aYBg5llTl7pg4dv5LwRNlRpJA8BIwW8mdYZkOffSiSRyzKNfg7
5iRDILwF1Fo98YWALO3sQ+KlM7nymVjTEFfn4VT5AKriOETAA/ZfDVOlPzqEaxq/
FNQr7b9eHGbMo2c0RRERexom3ZxR8eLIol7ftUYYy4/bQCPk9/u373hvj3Om8Hp0
3CYj3xa78lzSHg7AaM+U0UGcHoso/RBYZ+V2ob26Mx6KgL2bDes97EYAm4KlVgSu
GOoLQGqu5VXJvyVCUQnkfY81hYpAEPgsQjLyFjLbjciWe/YXNg+0lABlmgLCP8Su
8C0L5au/rUA+yn1ufP1HHyqDP69BUCvziITuTEo/1/pRPsad6jI3rV+bNsJ8qyqZ
d47V+rAqg3pdtSPgzN6Ju7MxcnKHqGlAK+MDGQh6H2XYBEfQ7dyAeB2pvhLCU3n7
gm0XiiayT8TmdnsKsJbnRIgfNRy4R8WLIcvxGxEiYgLUJ3c166bCIiKSBjUHiC1u
9s5OnNcygaoI1hsRkBhHIkdl16kOa6B2apE6r6XAG5y6cgxKxF+aVLrkq/Fp3hD6
vND7/J/2K3Gzw2uuqMHbpqdIQzYsoZu+LxC/QcryHmwmPiE6XeLLywXnT5umHnDw
8HcxKQ5YU22YoPav8SjI7g==
`protect END_PROTECTED