-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
enKCXfxitZHQEx4eDreat7J+CYJIkRx/aDHjYEzH/WxvCAVs5BpiNGGgms+V34Dn
9ExQzgzaju1vMNFWnhXxuJmvZi8V8hTVwR9xREP4KFAzmuzVLgjUltCcA+oqb8Yq
WlygNf7itgBGolWeAoElsKBpl3oce6qBO04l1LUgZEw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7585)

`protect DATA_BLOCK
Sbw0q/kPPq67a/RJj+3AlJld5Bo+8xc/TYTbLzb5uJ5DXprKIv2/mFnPaLEs5xJb
xJjQF7TA90K4ffrDsmk5E/lO4tE2opkzhEskmsnXxlEDvU8jKwiIXEluG68ZT43U
eJxzmcGhKbRlqf5MlGeNbZ62PrF79k8x/yRhoU5jI6tzdZi+UNFExuSztHViK0wJ
QfLvuEuw0gS+CjILusqLKxBSzC7wBCjcsjA/C/NJSSXcI8UB2VC+JtoEesw4vJ7O
CZWvsV7hwpASyQO/+XEIzE21r0qVNrtzd/qFzHBL5hlWp5ukhdYItVNLXIX7EfgD
FqwsA9Q0QcABXHNQAFGE0da6HNmbQhmOIM+QqgLhWM4FktHal4TMUMk3dnoC+CYb
3SmQ+4CDDQHWH1IQmSyvuANsW0KIUlNPePJ34rredBeusSbd3jPN+605j6IeLcWS
62X2BLYllPI++VA6bo6kDXLVUeNJuDqmLjyZ1rYzls8VTa04rCSk5ZTGzswaA6dm
KLysu0yP0UAO6Jt6frFd1unMb32JnTI97NR1x0b8GbvHXVYQW+/LcIYESLJQTmCx
xWaqSx8XWMhthAJTWvaT+84Cce32h+r+RBxCU1rEnl4rBYnAjnM/5HGBSjGAfx/d
tmtrUsBEm5grgWrb84rwRfgYeHuxdwwduQr0OPC8u6xkvorzaVjLEvQ4omrwnQw8
fFVKz81RkFxlNwaESgyFqjZGuOyvJx+UnE/xn8pgzefpZUvsR1u43Zlo87hOipsD
refNH5rVoEpUQmc3JZrBKGb39yGrnKu5jJ/rUmH1OKKF6ZPAgFnyw0v5gSccGvPB
xnDaB2r95EZ7AI5GTmObq/zfn0JEil7jd0R5QTVJ6Bv5NMEa0mOilKFn7/UcP+UJ
N6Lr6Oi2aV3K2L8y2dAZhHm1ctsktgT8damCwumk5sPPrZ6GTnRuYQgk6c8IL5B8
DHhj48D8rAy2ZAlktvdkQHQauSCFuwhJi2Go/NNyl+QEWmH6GlHlLgcIyF1oTCtV
3XNDi+PM/wEUKIJvuTPdGY4nyvmLeLmUlWIGpzoJRN5+pPSDBLduyPiPozpjKWm/
DL1Vje38vfJQJV1BLOnXr9FkzZolRdBv4QOctZffPZrrfS5dyzeC4W/f7ZJsRLs2
rvqFdPPQ8aJXLYbPbrIxmFLOjWEdZ8pMTKmESY/RLK/rtrx8UgbTmzOjEM2HIL4r
bKQKTDFB4Y7aK1r3I5B5TqAtOcHq3jpdprIRNnqtvqLnN8fKbM3bJtPezCG/4koK
6h1B2t/yIuuz0Z3GWHrxQCced2FPIQhT4b0xIjvz51qXEFpUM69XcR6G4Mgv3ifN
ysTMN8QRonlcI2QzmtyD6OnE3/KZ4Un4HGkvtClmlIw2PoWhSyOaVFRJz9DxTx8R
uqHWwTfed5jBaanjQrCwSN2uM2IoZ6LRaOdEdblrOqLxxi3qx7rlp7F35LsZ2zUA
6bvkZVciuUdhOglYgFB50xCeamGt16fmejwk+S10/qyPeOpHmh+4yz2ENiJJ8XcI
qrJu9lIjfPnFy78yvCeXkdLCmWWvjSP5axJvR0B/2KmdGkKJPDm3seZbA8jouQ4H
qSNvoFHqkIcs7T2TVD95C6AnQAMi9lzYTa52JfWWDNjY6aMZcDHD+NmCD7caItrD
uM186eLBDXF5Fia5YyQM3d95j/MpvKRaCHmzAcup26s3ExVaHA/+7MtjMbMPj4nD
PcsMwtMObgceyWnl2bL+CgzRSW4CuXuoEgq322nKIAiXWnlTGYqslgUDF1X8g4My
m2pfkVad7Gj+WhAlyZERtneZazZPLnIN4WKfN/15CYtVwO+h310vTIn7F69L915v
kGe0Fj/ssrDX+lhAfUAeTuO50xQrQ5iRRIGpp9q5YRVV0f/Id9rMe0uNU4NM59V1
R6s1EB8T3RpgsJtVgWXOgbBRHNNZskM4UiVbsTyTh83tbyXS5HGT813/ij3l0eHp
DiA/Bhh06KDEEmns/DYYP1kJt95RXCPgmKMVciT18HrO3a6N8TPtFP/8qwxRf1P6
Bp3vSuK+zSkbVu/+F3aPKfl7MkQlBlEVaYtd/Zj8fyfj7q+JvpJUfGGc7yHO+ARy
oo8XKOKmF1y0JB5iWYQJtaD+fupyIxuVGu40NicUoUFxGHL8GWtto0fh3Yx0qIsE
YoahG/2kbBKoCmk18lOLuH5qt2A+pKvETgb0BQFzYPya9Oqia9oJXJNzgnZZ808j
PoJa7r7Zgp4kyrbxvxwfM20MDSNvcvWVFEbMra08OvSSyXM8WwcvdJpIkgOzVvBq
FTQ/Z2jFcpeJfdZA9aCjpf3CX5rvmKh58GuMcq9YcAgCtXRJMoA61ggk4DHe6qzy
WyfRaTKbrMQVHBDeZaZcdEFfPIggUyy9+64Eb/ju+9dZ0IoT8WQ1PG3pf/zsxGOV
avGDxdWezFeZsIj2Dx6X8s1mLeTptAwGARxTxbMWaiHX1KAyeMtks/VYcGvQAjhg
89wH5nCg2FTkUT5r3WVMFeYZ+0fMDR+bSP01OpZCyGSkN2SFhMZAPFfBOLzP2t+y
sNHmFndt5FdpVyBmWp5S7luwM215UoAY4h7N+zGmikysh9OeQhB8AwO4hVkvSkJR
Z4NzZVYHuSsTnAi7m7nJChrcU9inWoorbTRxY08YH5YI6iOk4KuP/4s0Fctlv2YS
7DjJ0w6A3+R8qTi09YcJvT2Mc1lViVONeTdN3ZE4HIHOH2yDNgGmH+gJMLYdeahc
XgGjF/kgDr8jUOYw7bwJyLLTrfAZEjUk6XXrFmiyYIWSXB1XV+C5aGs0MyxbRV5C
zXEnzUviNl/cX3Elwsa5/dl2pb0kOBax6eEGeRpm7bHGwPy6XOWhoGifvT+JkOZs
bDtj8EQ+6F8eXs/qmoPWuexFwXTR7qqZSEUOE0LbgZB9Rrzr/gxstfgEHf1QUOGA
Tf4cPy688uJvE0cPAj57qwhKigujprTR0pU3Zuf4KcfeuBgmQfHsg4B9GYxyIxYr
TdY2K/2LswjeGCU/823kY6qQto/9wYgj3F2sFH07H9FVOS5HWhXMqU9NLISmlx3r
pouRgRWnnNvQE8LuKhxs543xvw3JKQJl7eVo5PTj2li/yDY4hmcmNwnomestDQY4
B18C5De4pdq/aw6ZTMM3XQpodJ92Knzplv1vWZOWaD23SzIOQXxstRPIVqpJLmah
XZU3h4BQSxrapdN+APENxHQXc+xZJRdNY5HEB6ugGdIeyi68RfeMcJC1EcCPwZ7C
cstrG+5vpScnd5CoHR9i/VWzTViSiKBKDjS/xK/ACk2mOtE7DVVVG6YDvfh1uahT
BqQt+ULa1AtjEVKneGD2x0CeuvpphgMc2oOiBaEJwBWFb8bEVku8vLNXV4hQib+I
rIUwagVfnEVEtoHLlnrIukOABdQxElQGt5GpqFqiGYLsy82AIutJzFzH4dANwp41
JOPbbJggDUmfFORddwcD5y+1ZemQfhR0MrxL60/YUjknKbgSR4bC1gTe63nzwoJH
QA7gxgoQLhVE23HBPguHv/30/beDDCjGdk9bBlgtPXXEY2eOPa9odzs/T00iPDW7
mMyI5qgqZvT570jbzF5RCV2awBflK4KW5jXy2A6VbAPewXKmzhP4lwe9Ord/bGnN
DqTQfUIawY4voFkPEzk74iwVDA/V/c8U8dsFyoF0RZ7T/VIMnYltcR47uI6D94St
ORKX+EdaXulwJwOypQ1MzaoqIYYGzKb68wpfVvl7i8huAJlPEA6yEyE6k3khbjj3
JCVznbL51JVTQYKJ51l5ua1Pi3bECeMqgCqVdt/pgDB3G0IuAyoDOc5Ka1AQ/rio
2PIoQkia5IKZpZOd5OnwL8JNf7W39AWjZoR74gRKassaNfeogXlYVj6nev7EbOjG
8FrUdE0s1OWfKOr/fvqoDlI0czOsnSJQemAcBYKHs9JLr8Ra6AQwN8aPq4yCOI0s
x5MOr35qkj0VGpP3k8iUv+iJt1/RBUNHEDQd1nQtMuxb9mZxGU3MP/CDMem/yxm1
t148MsCZTO56mromXLOXqoUB82FXyngTZJpzUVE4x+/CFhPcKjE8dfHGvMKzknU8
Wad4MQeHQlblP5Jl+sUKmQIFOdUA7RaydnpAJXRu4/85ULpUhcKX3Bc/IJPf/YrP
b39QWI7vylyG/US9bHL1N56+xzVABqnT2Ch4Zcc3m5P34iKsBeQKvq4NfbVZGLjP
rnbSiQ6Y0aaQNOQRYHWSWrMV2JKqg48F5S0yxlckEzLisolKUWC25iMGaO9hLzYx
CFyYIOSHEQIOoCpAKzYjJPT8EJxKaAOqxDEh5G2HTtcd3JCzqMxb9YE32xnYFrMI
bt3nthxE4EA9A6NAppDS/Wef6TYxR9U1rH1oGuU/DGlLl/F9dBd6tbFOMwD4bLpj
NEbEW5bIxWgVypHDPA3Se/9E9HVK06D/YuZpQpswKjUql8GOaf1CRIjGel0lCma0
pY5A6UiLap7WMK4NlrfKdybNUxdeENXNUdOIRWG1kdVEs6JjQivIwwx5gQTgSarU
5qSekk65FY66eDNNMr2n6//650cUSM1oqDBkldV7Awm5va0PvPDLbSWbCaByB0Bs
tkxwFUIRsnjeuG+krJ/cIg6Eag/yFAVGqY/Zg6aogRB/mKUxgq2QiBkzfU2ffseQ
2A/u65G+KhHVOlv6JfhTg3c6lYZ+EgZGyvY/OS382/1KfES9hUoI/VprXQX1w9ww
+Z9H4P7mNYYrelzqu9t5RJ/C9PTOhY6Yw2we20xaIzajzt8KmgG9WyTEuhqMgB20
5UVZVIGQfrTsvZLbb3qu0J4fion1Jfw1CYUS/USWgca3pqZoqyoR/0ht0+0eH51u
ndaeTUMOVmNNqUOvEuDC0yo/10OnxSykoHTxyJ4yhyKa8PQGAy7BN+8re2/CwzMq
GFgh0GqhcZ/ftsvEBTesdI+rorCDPIppTRhHo6S5ZfQZfTW7hwEE0YmbVmn25aDr
Z7AtN71e8wkDvA1JpBoBNKnC+HDACg9L6KCBn4xOBD2zAqe0OpBruFwS+HXci8Hr
4zJDEALqIMSUNpmDxv/Gqk0iNc7jQkok4y6ThYcvXozMu1bswzkZ8Rw8N4GA5Cmd
cnHFiaBaxVNPHTkM/GreBUJN2SqkRt57BmN9dBBy4NZr6O7a6Oj1PD4Aqcv1D+GJ
2AmlxmYztwKOvBHPpbcOaFK1cHWtEgJat16T6HhjiHubzsCpVXYwtsEzHEV2J8LD
zAk7z6uyXx9QZIp+4fmg4bqPl5u+8slyPJQUJvDaHHJlrIWOKHxA6awrsdr3emWZ
QiiHqTVAbm8GU/YKl8YfFvLSGcCbLxfzuNCWiu7WBA0PWkABc1cZ0gr9ntvxRVVv
7vVPlkxblRaK7SY5R60Iq+mqsbvNYGtRCHah41gi3FB6ceQEwPLnHLYiBp3palP2
q8ADjji49Mi/LTIqWix1R4xRA4goii4zv2NTdzeghNlaP1xbRgLSnZM07ljIJZj1
8pqF1tOKVFdTGIfO2nGyH0nVKd6njGSsj9eqeqtXmlnI/pCXyX/ZDTOjBmG8FSh0
OLG4vbD5eAtGkocjVqz2ry69e91QYQ2ztrGxkM29tbZcir06eVGcTf4Z5W6HcPt4
LTiey3W9gq5nerAFnij6i67qKQxshxBepFPF3reOI12rLt1lIMm83ZZLNCsAH0jB
hhxPfm6/FJxUdFao0YmDvKcjHRNhNwb0MN8xJgiDlrGxvLU3/d+tEoeiLpGgX4zI
ImdifWPT6HxdRQ9AOInj8quNj5kyOWCZZkPpbH22pt/e3h6S3Qrtnxq5OU1iJez2
JsHE5qXKMC+79utSbUklzu/EN8pc6hvLntnbQXX/gb8XkIHNsDUvjb9uUa2FFwVL
Zyo2v6Z2YgNHi/SxKLq1nIjdc3NTz/qgI93/XMq58WxqQ74vLHrCfJf+8xcSFNeq
pNvXOQGLnp38z5v2s7toRKYiUVJL+mxjMiV1m0mm7Hp2YP7DgEejN9dA1JZ7iie0
oxhk5x93qXr+HQj7OvTFdH4lO+UCAnpbIZpBGcLLLTX8tVw9Xyy2/NAsVuxMtTO9
SD/vQBvrU6rtCwx50TKHKg1p1PKQSUC0J+yNczc/qTi+/Nw6nrYhDzPs/wM3OVJr
pmbJ8ZGiY8V5wUtceV0s5AVd69XrGvZjVJU8cKRgF03VBLAoxZFQ7MPkiToJFf1a
Uw3b/A8TkD7++Oujp0NtL1y6rfU4HyeT7P+FeRsD1LtuYHeHrC52la8BU9cwRqKy
oWifRfkAb75YcdlMdWh8tK7KCcqsE0M9X1KPnL8pU7Nb1GjKa60oYjtetYhemFyK
cBqvuSNXvtjhqvQVFezF1OHdPFjFWVVg4KQEMOGFe8X27LvjGsVQc18f3s0UXqbe
6kfW0GmnmC21pTyDkJEtKJCRI9nHeT4IFGsuVBubKh9rQtrOJWsLjoyd6TCus6ov
hOY6Jtz4a0KaRabR/ElbLFZqU5i8HSxjJrViyYuwqK17nSgXVdrAkqjuvF1Mv8mb
d4OBo/F6von8UmzNa0uuZCLSiSxc6LMaoxnGO6Ox9Er/Qd55iPoU6fNtIL9Z6YZs
mIoo64tmOmNxtmliIp6bLFfzI+1TDxlHA/w14SgqaUMRvY9dCc8ZYrGmbrQlqF58
gGle9Xco3sihq81FK1U6OsWLTy+kKmSMPk1WLUPqPNVNn7UMsOTCY4K3Hju6N4Xu
XndG9ANz9njQZ2hsxft7etpmZmEWKfDUcCUMhMh2OdBOVbbAh8im5gD2lCdKE5Rj
W9AKkjO1yK3cXb0M5ezpqRR0Dz4pHTaTcq5OJyQXQeeR3/IJdBg9u06OrTWqEszb
39YZsJbM84Owl/vUGvQGr2KOJlirr2UYul8sMnXAQ8RezT1ArGaifmmD4hjHUd0v
CWuZS8gDdtWdI1q3GYUCpL0ObY8upk4n4npuNdc5y/buOcjehwSu2OtWnkWzC5tC
hlHHNndr1R9kYyCNQR/f0TaYLTcNQxICVKtwqKpdWIL0qAaiLBxJw9n6lRrlm8fc
gJYww+Jr8GWDDUacDX/lB2+eAPcnExJ01eLHF2g8aUKDA7TcTcgAckYLwnfCeP1c
pYSvDhnFTzyhcw2gzwLgeLDpXBCm/QTZVJICyvhts/SqbFsQmE5OSofQFrckS+JR
ta2PxR95nxSu90IHHKzDHAqXS/YpLjzuN3GS3ZJU9BYgA3054ZtaATX2pyEZh3ru
ogwPw3goPQJG6juzoz3SOaNS6kiOVKwfEH5+h+8wYnlG+lEzBOlCHzfgG8riS8sJ
9drSd2UYiVxmB5HjwtNFgUJBUkwXLmiyYZhJyZDiY3bcbcU+l+3geYWAkmo50wz9
xFWHDLXy+FFjz3REb84vwXnpJ2/Li7qHZhBT7ulSLZb3ndHv7rp4ibloKpbp3Zla
/LklvscMHP999KkMh58JOMDcyYzIco7b3WabLag4qSrQ9QDB4S8+dk5tGLjhQfvF
qFlZZXZ0zY7gJZZOgPD45r6IrfskZYh+siDnoDZ3T4Z0dgkZxSEJeCTOtLJJenE2
BuJrLYWccRvFkRUGP6H+4V/v0B7ErDCi9fnd/7+i4PEJGi9ty5u/HVUyFiA3kBoz
X4luVUEMZcQEa8c5N68ERug3qBPkOAlQ4yn7GRDZwI+72wL6tV6QROKrEcR9lqsc
0R/PaDDwgVJVmampSBKzvZc91iicXQEzVaTJS/nZFGtcmjMMQmXlwfsudt4KBw67
voLLG/E8059paq/KVbg32C5x8V+J5Sd384CNSZ81nF2ZJIBIqBo54H4bnIqkPX0v
m/MMhZx+q76ikzfUVgVAjB2neR5xqFPv11P/BUExcp3NF0yfKZIVC4p3jxn92Z0F
2yBxM6T3rcobrd3gdrWgD9qK5Kwvw7+90VXTvEvQo+21D1BQeUqoF34bW5QSiBqp
qwIm1QyiSfbD0UW949r2ObDTEcMHzBSiB1UsxKQMEoBg/5njnQwRv2wnb1OAB0rH
uGvbykfRZ4ixRxJX9NUg/7xCq9Cofa/zyVReNRKtjRf3WsAedTczoyReAdjFPPQN
OcK9KiQh/fv6EU7UVLjWksshkx2osbJGSJlHnfFKlfG+DkEix4aFafvzwEgctdWj
ehw+WFgqhCzhwZoxANVMaX80nbDOiw8H4gPA5ggykjArqTPuinhzmw5gE6siaDwH
wviXJlxvXJGlh/d0aLrMs65PkaDy5RU5ANJdA0jnbfg5ekN8+/GH+K5X2VeAsuEC
EwpurRuaDtpQEYD8gLJgPyDBypy1RfuIXB8Tp9rWxYA34yLgY1iLBACV4NnyQfAG
0i0DfOByNlWdsUXzsood1UsoyGJgoS1kPnaSQDnozuitQtU6qhd0xK4pu0Q+/5l9
S8p/wdCz/VmvEClHVRjpTAMgWMvLLyFEf7574keH7pDY6p4qu/G08SrDQXfkvlk1
Ai9oB0sur0cM479CXeNS29g+hUAwPhRXL6KIOCtZpsH0BsUvehWfyouzBoClOypO
5NQJEZ/uzE9G3CWD7cXaSu7ib72DrPn8pFO8ZGC9ukDigHfqwYJs5TWWU8mZAPtl
3OV3yO9j70T0nrvPAr6RavuHX7H2lZDC64Fweu+Sv1F8JFpufgZeyYerCUCKDcLb
I1ZCi+cKek0tIPw5aoBTl0YySlUMbMx6aAHfpt2sPoe8hoqyWsaYoWWNmVYImvnS
c4yIniM38x+QYkCJYzU5aYf0hwZIRNufdnXkOgr2/u0BR/vaBPTAR8lfQOxV9Ylb
T+/diVu7Il6gOpZE1HYerNkBQp6CUvBiZ7Uz0GQfdWelToTh2ytG/k5DtPGFDcc9
k6e7vHuZTtXLnFoAXwyFA93SKZ4c55OiJvhpB7ur6Hkw2zMqXkGc7CUa5I/tF1WR
u+goQ1vxj9QUIRQLR7pMlEs4Uz0VFnP+q7w2Vp+2k27dhYHYltab2Ewdi2hJVCke
Uz2z2RDeByiYc8O2twH+zshfIqtgPvHPyDCFMgEAF+qHuwNPxGWrSHODJOXth96+
nbSE7o1HqB8VQhvvDWjn+C89tNj5W1b7WQnVLbvEbzPIqeKnTUtb1DKva/pJj+LH
iJ6shp98W3uuP/mMqx4ZjjRkn3i+H68kudAk/xTGkPl8EVoiPS6bGxwYwEPFtFrW
ZBf3xvD/6tzUSXW5RO6pPLEhe2v0nApGZ1TCBghn2xhNSu4UjgoKYYCibXj5aQWQ
mAtKQjqpwnk4PhoRnAxCpGf8N7d2KKBSuwBajqLIkrTlzIjPb+YcoyMHOMbfkCda
U8Z1j8PAgos9hCmFra4zYN9KOoXMmCJTm+Jkb8kMTv7qnWexJH2piCA9GyKqMU1i
57dzab8mElJ4tk0QIzKsWa8luUeUrPkbXMLe3ZsNlBuvy9q+kP3l28HhgTT+vN07
YnPaaARC9Gv8+dqZYe3U4H5QHoCZ8fujHMLS2YvhSYUv559uuSB2P/OlCWqxX6Mv
i0cY7CAb2bdoreS2POTolTdj+5udvXo5HMzaop7QuGKxQQVPA/zhBSDFyfR/AZS7
CXfNq6sQHyYtcFG7hj3Q8k4khWNc5pgLyKKsf5JdCMaubf3EDN3Pz9jxRFEQmv2w
8/wf05ERjMQz0hgZFzUtbdZf/ZJyEJ8dWR42I9of2zuE5rVhkaz0TX2psMgVb766
gIBgLBXDrdussARkkgiyzHu5qXJxeEJlr1SMx9jmNHpnoBtVPTaW3PIfcU7Gu311
ngRt0dHxo3xbvFMhf0C5GRIZFnLHHR1dIPBqw0xGU8Bao+D/OViU7/bARSvkfe2p
xiwzY6cTQNOd1d9T5uHfOvkk4bt9P69N8t6KKT7ZZtOolQI1xPXMO4RQI7eW91FM
WdzRgbt7PaxZRrTEE/vHT1uSIGo8r2NZD5vqB61y0C9etYijQd9DfZtaYr4SFfrw
STUKYXnrDLZvfyiPUqJ7voqn6MtSHMzdv0KL/pDf+KWl/mcmqnh8V6vIgm1suuv0
v1l0Fxli40LW5N3iQj4YzvqFBeS0caGwTwUEzTT1cQ5CgAI7kzIVsiOJgZMYG7yJ
ZXbWVNOJHl+h5a+mvSchNowbhhxaE/YlxMOhazdgA32MNTLv5IEBBPucIv4Dx3CR
ZMvdZdIrdMNzA5bYUuDtxJsy8IrM3IfqvZasl8KIE3g=
`protect END_PROTECTED