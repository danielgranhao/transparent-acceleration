-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
V8PWXAKjG4lQ7KJvPMdZ0ZbiwbQoJRfqWj1mqicvDWAUlSAFDSaJOxiWO+9LNKnO7dB1nqpu8SV7
MPb4fw8VaAJAn5MsN30iQatEi58O1IREMct1t9+21+Isrr+EkL+37iMKimQcXZoyKd5Edj1nCRYd
opuM/ok5AERc/yfpLjQVPz9kzHm28nppqkN1OK7orQ50W5xiPucWmrej5uqedYc4xNid7r6b6Bm7
IUN8fxildxm96ik0BNLnYHfI46rckOCDpzSLiSt/SxKYjlcJPw6RIpmEr0jb+xkXweix+1Jkwb3O
y5tr8iaQbW7ai65iyhtdbwHEXT7wZeDiHDD6Pg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23328)
`protect data_block
UAGExTACRt5ncf3f4zrHqz67U9EHzIjPBPcQecrFAo/oj1zbR95px89lQ/+7DHnDODqfjgRvdiBv
W6Wl1wyztorLPwnWtwRY4ztOQBsXjic0xkdDl8JzZqbfNG8lx8J6H+F64jrQ1HR8RIhy1kihfS4F
a9W//EFGIiCvrD3CwOjNuSb4yjJkp1UutombrHsTjRlmPc2bg1RLFLhqc4kkQV7HVu2hqYtbhhDc
cqyfY60mN4gRy/kmOCfBEPS19fQ9/PW2YqdJml5cPjud7NnHp/4YWENEv2xIkorMdK6zwUB5J7Fs
rNxniHeFcWTu7fLgG3hcytcixmCU//ar+e1mnUxQZWnF43ZUGZSISVY+nR6urcCVXoecQHG8e0wL
B6KyqzJiMpsBU2eeFaxu/+uplUHTvTqpz6S4bcRovw7w2BBqL2FNJMn82KFhTfjXXBNwsZDmsM56
PlkXbuGpppG3g6DD5Ydkeavkkdr3+UIvZww+c6zbJM5p66Hv7TFEOlE/tdL8am6fdxpJV4Re4/GD
EDqRJ2iKDaRG8lkzUo7qoXn/kfSyP8LjJIHqayg3hHLJ1qux0yUvU9uRMJiW0g0vHfGvzyF5Skma
SMhBOJBpOX7bP1VFpmeptEE6hnibbErzwBDyymW2k1q3IoUDcJNuPf8HS5LfrQ+7FyB6DGldY+ND
zL8IlQ7c80AJRNuslXvRwbxjzEWwwfKu6D/s1vEj6UUvxFsk6tR5c4FEtW7xU4Y2/+Bt/019dR4K
iaORXsCotb8e7jgqmvuW2+F1N+1c6udC7SYHs1w9hGrfbe32oLMJTwSRnC2mh/nsb7FePbdaeNI0
S+nZM1WEKa4tgBFQNvR9QzXCrojBaCs5S/VJ5BKyDgyrcfOq+Z04DfPHbfx6/CAAinp3A8FztIAd
8iqDla9tJEDIoEwCOB9ZzBbsBTNb8YSBOMw/VUrBO9nmGOFRkAEz/aKKNhjTy25E+tZXDo761vIo
HOelSXmb/tW+kaX2dXLLJmz4XHwshId/pPb5tIOHi8nK8Ws0SBLnMS2d835hB0wqEMgNguOYHkpi
1kuneBZ4ZTxGmDxi1qYpPskGWR7LcA8Jm8e7SIxNpDZ+wwH/anwdS2TiENq5HOgFLKAzQbzJG82L
TwcGyAIeUHedQ3st0yxLrrnCh+YRIhkdRzUX9aBnzeKR2c6r2/F5OqOQ8ByMkmSwqqcY0jgfqhWB
30cWBo/m8fIGp2smJt3ZDAeusYxBr3vnanaNtsbjKLTpm6vu7SurZXw1HO89y9gDcXZNMvXpWAQK
D5WfSOCBKMhBLCKnG7xyYgBOBrZ7syb1s81HuecEDD02JQJIr1YEGkrO4Qc9fk2twru3howVjvMw
MBTx8SLl0lJ5Ftw/07aVtwZRjHsJfON22NDZL+1bsVo3SIhJS9cqyUsRPuAuf9aeWSgpYxdCf8jA
D79CV/emwm+wQYEwoudiv6LaKsY3v/c2eEPy7zXioZGuI9ng6qGZZVKp5N1ZldcfrAtYtcUli49R
xGTnRFjf1kB35SQFgTH6Oea/XH2xDYmn435R+Bi0WOekQcpvWqWMP063oPrEdeGPtBqoGdb663un
v2sn9NHiw/ZCclgaUaLoSg3CJX+lUX1qhF8OSw3xvrQsS4zKnijO4RW16p02fCVI75WdO/DTjUq6
91svUBmr7RM7GxRNNDYPkavs2oJSNZdkRWGe4tnukUA9B8+8Nr7gGvG4FX7ULlQcXIVZ3SR+zc5T
Dz/nEmk2d5e3MpUv8kjqCdCtC0Laq9OqKwtE5qPFpWtcmUDdkRTQVDk2x9UNVt1Bom8WLP70oonQ
Z7+MEk4cfjxRjekG7haE3d6oJy28ME5HXGhXvQn/Ndp9O4OUQYimHvh6Bu37nuZuQD1rBqmC+1T4
KWd0qvXicn3kIyoAYz7gyBGeSyHtSWqlIIrbFwZeMcdbzfbANKBo9pl1lviZ81QgcQoiD/l9oazC
f1vTOHjpyk2+OI7IZ2EPXsublP4gL210TNHQPABh2qkI/ximlOC5GNxSoLoWBUBavQXTnXCoeEtX
39WL+Mp+zUItCjFCILYJcH/vwbAz7dOs2CZl7DLvWjCOpDo1R0LbtqeJmxvAdqMcCtUpJ+e53PZr
vPpUkjMOXWKO8RQxOYbQNlpQGy+5wvtAszF8vzs9vQRFlDyy1nnEYm9zf6sEmSWDaTsgMnP+yLI9
xfEpykDENJdajIwQT3QM9nLjc9DQF4U7SYQeA0WFPBjc2BpnqlbgxQmNpbkuy7IHfmriN7M6BPmT
5gT+NHsXAzvznStRv542CBLp03y40OFHfgc/s4voTtM6jmCVsuZF3h73EMehA6nFfmJTLtMMVliG
Ok2FIoBUUM+pCud1bSCtNDAbGiI4IQV2b3j1LzetzBKCT/pSbrPY8BdD/1zXymMAVd5SAnojv59v
n9O8Ggo20t1fsLNkHshRu7oeqK2pAVJKUM1dG7X8togBsp8Ci4QuniGXbjiVybVqLRlp7TWBrHM+
0pwMGXxecSiJPdwyDfe6NqsBByPYlKaDRzzkoiSZ10uxQWy+8v3vnz2Mf0Y6mvBDcjOS3woXNFC4
5DZP4l8+GLFEuypCx5DSJy7DwkRo9jnSJh52df0lJ7F5hfDPUjWPMf42NtzAe0C8dvaayMbBqF32
Ao+1hS18BE/PITBjuvTKM7Xl6WiZVNBvLH1KbgA7fLRjdMqcvtDf+5q0UPWRR8GC1wb08Bv5Nx7W
8SbNNg0xaQeR3MaxzuttYEmo3eKJjIWsWzYCKkJ6h2s+Xku+Fdscc+VipNYegfU8aAn/o2wj/l7o
RXqEh/CDU4HdISceAu/URMJ/zJ6uUNK35LrbA7JwurKgMJevuuhDDvNWDPenPnQn4XsK3l0G/qrk
IM7lijXqdh4e3Z59ZnzQA4M/gqK9sGXyHz6vj9ENuyjRB7AByRlD4S2fhxuQU/1XPzHaYukQcSeb
DZLY6waEi+8WOGyqo/8Lm/NnzblX2Bs9ZBTO9JfX0ORPWwAIpfipfKejT1Z32bfyXVBADTAVtLIy
KFxKLOmVSCAx5FwriPDwL5WQEslXcVwtlvHyzbIPxWmETG8soZfA+24s8AJsUPHbRH9GLHopPZr7
cZtnHxLC4rh/UfkW7amo4F0KvXHfZPWfhBEvDBqch3mVW8Nx578z6QmYDcXuujig0R0inFX/brdH
Hm3bSGR3j2TetISCwZfk7OyDQLA0RRUSMIcfThVhAd4lhKKAufi5BUf4uupskGJWuJ0EqxRQSreL
EV3YP/oLJ3g0INcODBVxhmSbzNaAxvCM5l9wpzIttyyhOUkJlgZfhoGRYByOY89Z/w1qQsvzCQNj
XkDqdjIPFTt9jELOjqDW8nEOJN3a56QWY2SHm3KaXxiPDoG9Jb352kZUfjKnNyCrnbUummK4h2Sp
tKd83rgX4X2Wz5Iy1Byp6lRQ/K2HTJokFbaCWcXuAMydNSx2ErTtQQjxUKSMPH8JBt8opsgF2U+T
HG9mGw2zC0K4NBtJKxWY7fOLSL1E3IwfUI8vecGPhF4gKOiBOVPCfnf47BJSsqY3mL3ut2wlUIEL
DLArd1JH4luuyGzXbAD8wpL0Yzbr5VoinuGC8wJiRKgC+faZhoQrgoMhL9Y05GsilyO8bUfwJtib
nPikeOuP42sRJNYWGsPMzMaaVidllRW6oWCpn7d0x6Bemc0j/oZoN3Z/C4AXXgkYIzdwStqqOOOn
Uc7YaOrec+IfkE2suaWGJ3Jh14CdNGX2xaUfLx6DRlbJiTBluVpY79cNs+EHwXjXIAMZF8SnQe/+
1qLaP26zYfndloIVEoDXN6PnPh+UD11YUedvXB1NfXSQHfbma3NqFPa+UIuXHhVUGnJRilHpumxM
nD9wsCEmp3VbSrqQnRRnN4mJe/H+5LII0bOTkc6hCBa2qCBDTW/18M38xruYxXsE+hhGGeApsEPo
yI/psjGRo3ul6oLZXLl4xfgknmrOK7aQFRgLFgzOPxahM3O629Dp36Ig7vkZa4jGWSUM5zthc5n+
ODJ7p+RDAQsWq1t+9LdOoj75JVLzPslj6vttEDwiTM4vPuZXsyKzJx0ap2HXf6WXonQMWRKdNEFg
+BwRDTJtu+GS/OSYncpdZPWWSqLun9WhlaPHgn4WegNlGTHvyeQLmDDR4IOnJe7hyz5j7U3p3ccl
iMQ0doQZS9wrrWMT7rTemKhXxX6yyIPFo6dLsxfLhG2ESCy5jNAYpakmpJNEwxy75R6yLA5RDcEy
+R1DNR4vbT5D4OrF2xKeBprImQ25mj+e5TvvNTSxvd/oZHJ/2gZyS0X9ClkglHCAa83AGVWbiMIv
PzFvg6HbWzkpYc/gmWFQQsTIYqW6mIyU67mfGQVhA7uDi6bx9t6rfZQrHZTbpBu7OuAGscMyiDtH
nQnGoVAD74ypqQTT4fyzI+i1OXzaO1cNMeWVVjo7tG2h2+4ywVpBzWSllW62dj/SyVlC2gWEs2Wn
05xx8zfWDxhlbwN6IQU1oCNaorfRHG3S4PvE48/eIfJhoLM3+mlnFk4Gs+wbCJln+qGOSR/opO00
U57sw+GLHNoxLuekPi5JWZ3ebwnMkj1LrM8T+pk5qMXOtthyTfpNTCqtRRXNCRMbmkQYNhJnb1Xl
Wu3QzVvjf1+fRe6dcxPYleSbAUjFl3pCBQ52kU98Jyzzf/hh+SLUbEahKPHnLu6QgOiOAPVd5vcd
kUIas9zY6/52jrKOjTwTlajf6w+7KsnD/UtTMtaTt2dHJzIVbOQNe5K6l2o3/+1xC9s9XagiZRwT
80j7MjhIz1OFB9xwPmK3Bai146/aiBgTDOo84bgzuUGL+IrOvLZwJ92Ktb2cvo5pdFRi7ILhDnEa
iFl8tOtnS05Ai4juuamEFl85iTfww/EbrVDZJytcVZ7cz/CiJXaR3paFymOYkltTmMQsWMBT+G6r
0hZgzgzOJKMNcU+wB3he9f7q6gKaIG9ZzlT454TCrHeQZcb5WVYRLqR00dgobQDRySBMmktNaZAB
fJ+2PgU48by4pav7nhwy2IZ/0Aa+Zo87uZ5rsWINDxMmnOOruVoniqUlOuKpLVENmxzLPL1J+PM5
wRA/tYENCeBZIh/hsUOW7ClZ3YlUlnw7dEygLrEFRc5BzWbB48AFLKEeVuFOK26VqE/blg8XKoDh
J3ZIHFio4uMpU6TjZdCfWe1GX9ZX3Gg0Znl87WxSZ2neipHkYUo9f56pAHK/GYc/EfgcYUmU/ZVw
pzGz2cy1GSBC2YXT0ERBi2rIxrELp9LWd3Jm5S/YAPmTNnqfeLehzSAKprGH9lXmU+hXFZJtLZOr
Rt2sNGyFnvfuY8cRl1rosGsIEpmSOQzHyh0ue44fxipb6w6xE7HCleVEgIiXp3+c/IYWrTGO4+dH
V6hv0B9YBoC2N+uZDBvEZ4aDPFOZ/1XL9iG1TgDeGhyq9dVpz1XDvG51iy0cU+4uz0eFjlxYme7p
CWGkjBqfp/gYAEE9YiOUEuODAR0ZKoKN9s0m5Hyb1WwgwkevCz0YDt847dMZMb4B77MArM6QS0FJ
iuckRfVKExll0/7WsW6CzysXnqzTcGjU/13CChOaViOAJpl8yAOeYHFu4pX8Kgqq7GjrYRXQzffd
9DMULGzdcXH69WLEZcrSSV9chgLqSyf79tRe/it9yQwoMIClqRiybWwurOk6o/ofDEhmr6hotAga
J9Ing5XwZxoxS/QaLJiasS3QpnC5UKS28kIUdmWnzdUY1Dr860mJh3579roFVN6usGp/9KTMJFeM
C4eT3j5AJAfgQ3xgcendzUWjCIVGW3RDhExBgwJxGm8wm6dIq3yqk5xuLUUQ6G0KCT8bW5QIX8wf
KYcwK7V9U19bhYD88urUZSbkHNVopm8/nfTprUItUJjnWgvYOGVqT7jW0xB1W1vVY2Ixu8Gb74CH
UX48tSq27rYvCBunBgjaYnKrSrXzgV8/q2WbcTuuNBsirYiRFIu5tDtAIO1Z8w/3xfZvryjpYBrA
q+NOs0joOa4XgoKzaTcV1rtOg1xJ60o46zxqSohrCraXIscnncn/FH0stI3uOnk3L80RVoEG6Rjm
YHlcfYRk120I79mt+Cs9u4/Pn+g7BEB+7pt/eeRxj3KlgqSTuZJ5wFNEmm3mbUrDjEmhSF1PjCWX
7DU4/DKv5gPN4ivzN8SleamJVpvDMhvuKEVHrgnil3ehqQ5ojAZ9qmS1pabQbv4N8we+wwk/ydpd
SbcYADPyyONRv/SBJ9AQAAVwMTY074FMjF843l/EJPwVjQ8plb6HFkea93XMpCNgSZETdc/rZR7T
ogZfDt7aJbT0FedncC+2g1GOvTFm99WPu47f48aUhQlVNLHHqlJMV0ctQlAS/STN4BEvYylj9yLp
lnaDt37E42pbBlPgt5slxi24IzsUv7irbOlMg2ZKY0KzniniL+CPyQ9QV8jVLpLeiFaulEJ/cVab
On9TY7W6AITsIwzdc9hemWTEa0HwEObc/h61Qee2RSw5dLX+yM5eNTzpBddvHBaRiqtTCFN3Qh7Q
94fnUuKILYn+KOiB2QfN0K9WtE4Ei5IQ1hd9EWXTn3HPjuYR8xlznIIofF/BZtYA2g1Pr2NHTzln
eWu6dTpfiH1ecxwSuk+GlxFYbKRBQ1v4+bzfsMV10OVK95I6RXpyEKn4avAzBIUuwEm39VF0GfaO
RMnHBffa2b4kXBrDgOkpUcNBu759Hxx3NZv6jmNEwirt1m+ESna1A34cESXrd0Q/RJ+h30h9kCU0
N7CJsMneHGrh09n1D+gqo5dfERXC3AJ6J/Mpk6WK1DrJt0o2Vgsm9Z0vlmleFMHNvTfWcSSdzfQ1
ZUxUW5/gDrVf2XQyJKRjKJlEqRCsZ1pokGQQ+RHy7/+MbsHHM2fSnNE9ZjlI/70HFuhdfK7PglqY
QNBkmrX4cr1jy/aLWJQBYPR5aMXq0TzIYVD0RXMTTwMN7spmcjiljJ1mACNMmwczllUHJPpjh78o
Y2Fz7TvW6Zp1LYiqs94/mxXHjuLqHDsOzH7zogZn7OpmBhfVxT4ur1qWrqrwplJFiLK2FjYX052Q
mXIJsKnyAB12GiXvPul2veOrIEmmEx73V23GgyKCZ/Qxc9V4WQeVpTslvNew1a0fDH8lgnAib9KN
DeaX5XX40mS6kjwv8OEPahk5Vt8BtLY/Llz63IASTHZE9ZuHAMZmLbL0za3lsIAgOvVjnl2cQ06v
/ZwMPskkiVJi7X0w+hBJFF1y82OWpzgHA7BaEB9tl2EcoirqkTr6j+MvisqhkHWP/U9W9IYjuPbn
gckmrNMz8OL6RY8J6opxWt1en3rJrfJ6CnBpc0lvq0++bG4ESo+jCwF9xd0geiiLPLqlfb6lEX0J
lhRnlsN8LldZZxiJlilYi4B5e0aKJUnit1yrls66krZ30wY1lee3THnP9motmSLD+e3x/4RKFZaP
UQIU+X5MSD0G/Z08sLkL+SeLQT+Mgw0RZcaYq7+D41NZjgo1tPb+d/o3EWaxSJpIz2ghOzop6jJy
9i7JyhfZwUIKySIxDDgxeT00640+4R3Gnyjf7vRf/kKf2EEW+8atI2g6gL2trCY8PDuhwWcSi0It
1ieqERNq69t09y6JETVSUgOszEoRuDDsqqfdVy2OON1R+4gWIaJRmiDNlycypwSVqMPa+moQKeiw
b5ZpL1j6ITqBsfxBPdGv3LD9OrOFeEI9MG5Kph9LgwKE61WHkwTlp6factoTcHdUI7xUeZCFmIhA
t82qqnqiWdPRrw02oM8v6464Ie74AA90lfcHSbhHsYzhEV7g0HuKhEDzoMUsV0IKlFARVBO5SHcc
dG5w8C5A4fx1j0vrtgS3d0jcgadDjnC3MCUYIRja02kuH54YfOWrqhU7Pk+pXUWb28R+d3mfSJ5O
nG02lzTabDbt4WAlCmZj6jezu5JBSJ79HLmUdM8m7rpQLQ3ToHomJepCROnBq2HLir9VB2iMDXHl
XhKVNr+zkuE3y2Qm/y73vOAZXqPhUg+SbLsyeqoSIwuj7XcQocbXCrL1ONMsZ9+4dJnDtblON4pR
Ni1Y2oCdq8cKk6gwPs+Ts1XQjrIKYgcFp3cZtuLEF7QNECF302T04v7LRiHtDnNGvsQulfeEOlik
fRGPRm9sFigRmhNq33CqzEk2Ybl5loA3GMb4dRCn5oNs9kMeVBAfrjT9dd0fmNCZ/1dkJ77GINl+
QaNbDwGp1GKoz3d9bjPQVTrQth1Ijh1nDAXLi5BmnevM8p7gMHi/saR/TGlYApd95k3yFNNSx20a
hrKVVxPEMM6eOokxYGfkWFjeUwTYwSe7nJBzzu4VUGGA6S8fDArlkn74t1AW2CbvAce2bRGUe3Hg
F5r6qkG4+Pzq4MHfW2ug+ri95U5jlacjuA76EGqVsh9u8Tq0mBKxqx2N0R98LNzZf8y/tKzia6AJ
AVWMu0Tbm/82yywKBBDnlVC+xhMKoOLWe0OtTlJvDQnnlx2VrOitCYnakVuD4P2m2owtnY//bUUL
Z9e8q3tcN5n8jpFBVgchULWgoSBSwORt/GSnJZUVI/d7X9Aw01Uy0r4IQBaEg087c1lroc/+RhEK
wdiqsZLKNv1Qpx00eA0cUVab5VRpjq+HCa5Qi9Z72DO3RTfX124BuT6j+KiSZPyC3eMplErjDVpu
KUXJ0Kpl49niWa2Yu/oaJuA6y3JgPqpx/NKU9xNNDdbb9NCz/iUUt+xjBSHG4lW+AOg9dik97Rna
gH4kymhWr7B/Xw+piruNdLD2PZz3+ZfkezlK/nBj2eSUzmI01reUe36TC3+pb5PXqR2Sq+ze87vP
iwc8Qx+VAna+wWV4yyIHIyVj2yA0FyHQnd7f9X066RjvpWDmU+vi/Se/jrrdyPEVubGVaKPBItCe
iNwTGJlFS7KVRmC9E/aA/4qHLhuMuyGRXGqg6Tz7f61cIiGNsnDkhr87WYk3HV0VQBdPTj3//B9g
buLbI9sUeN4ppAxBztKl3p10tNIGALrD0R6Cbh8dYQhk0hOZcG64mcNwUJC5cm6TahzAH8Zjg+oP
8Ytkbh9I3jGa6zHZpGflV/pXVmJPTgVl9fER22DVNjGXbAOLiGD6lqoMObf71e0kZXB4zV5D2rGn
kguKn14cHtingEbVwMu3Mf/sfuEDAHHZzK3tt1FXiy7Gt1+ZXJed0+BXoTaCI0keKz/l3hOgmPqj
v2DHhzavbb4mjMdyPzkIAmt0N+CRBcyQmw+axsf9XTVIeCYkBa5FuvomdRjYZ6MUD70imBnfxl/Y
U8VS/8vrIPltNYAcYiHvbfsxZWO1HCc5wA+cZKFZtIKZDum2PsvW+3YvQ4UHrTv6iSjoDA515uyo
J00SjhKBhOopUBNIT2lU3JAmxzcmU/xgHe2V+BOoJMIbDgQlYm893Apkfr6D2RkHvl3mllZtgvk6
60kFdqKPeu1ZOmq/mFwdOfg+GC6nZuJwkkSJ/HfzPWwn2otR8Rf65BV/8qWHS0wqMimUjPFyGQeM
1FXrsGP+iI+71Z0PAP+yvT4lvTNFnKMg5k+rx3xgtrAcPnGEXEv78JeZZ4sOCk9ymgmY9qrST01S
tDItSG8VEothgcD5LcyySe6YKsj1ZIcJq0ah0jxCXFoosuSVAVHgZg2TMqDA30ck7slvM8+fdwim
pwON+3wi8dWOtiQIAWvdOXAzfl/260/preTYKyXOGbwmNNQeviNGTUhLgQnN4bQx//S1tDaTzVrC
z42t/4I8UvpmvX4gUnNyY0bHMtVTT8Bdq4fB8Ae9qe3vMFpmq+Y1uZMwOyk8fsvsn7Mz7mZemN3j
TFcvy5x9QfpIYOhkM+w60ezHPnza8RIKXGnZdwTiUtL0Wj9LPC8X1fYlMfcie85Ur7QgNN2IZgn2
KZf7n2Yj645qzRawZ/exKyBveR1AJ9EG1qqpL+R/3Armx45WKZhUcxpFrKJV4vOTV7pGSyg6c9cL
+a6zA8Ij8Ptk9gowpXwBEnO/p2qoYrXZVEN0MoJDjf7QghEM+/lk7T8WMA+p62nQqDWPEhHXIISB
QNqmi/zf6dt5zDlpfx6jo8p6g6oRQBECJiBkLDQgEbZcnxsWNTeRIjE8m6SPzudfijjMmZGGUjpa
EOg+v6OT415EdMrrmyDtWKGQUAMLxKNYq3Wo9NFWSuRDLW64G6+hIIl0YRErVOwrJX0Otfxi2+GU
mcAXatEEGWS1JRzwydDVfGFhrtkGGkk0zaVb6HwSoM9LvfYRvldD/fsw6AzOfLN800Pf/qOXBZn2
RwmPEH58iMBSucdYlEwU+LY70hB6rHEKr/0183Wa3go5x2L1S9D8JsjchHa2xM4FSSgtMQMEXGRG
sLkMKyQwObSSHoa56NE8tFlOuJN3gkMu+4pCW57U1+4aCExaSsMTC97h7riJQ4Cb9P5i3tQQnxZX
yI+PcXrNCPSD7+2CJql8A3IgWyBL9Rpm5j4Q8G+8AeQMA14UvrpznPXOwmQCsqqNKBR3nD8cKYHd
JHTVVmAMT+d9/XMxDssCH1G8d28Zvj3DStzK7ViyXvbrrb3lwmsCy1RBjhcZQ6F5xGhVkDeYpDDE
jAcNM14tEAw4kW39MUvzRC4UhGGQoWdMd9boea1pDndxWfIwYV0Ov+YUGxbzpGkPZVOD2GzKhA6M
Ooyj5C9p8plqJ1NizopPwAeD+YThFH+XGtnkKiFz/A5wHDtXinwOeCK8Zo3BwrhmMYv2fdkf2D06
oT/+4WdC6enbqULqqXzTQrujBb6UYIMom5xbUoQiR5oFvRPTM2KF1imy6tLyAQKuTRw7tVlZtBNa
fEn9BhTWMAl4gCjMdnNrH3zlSdQOYqmA+alzkbhQB3CYEB9zlvC6gv33J0teSoW8IpxxoXWfaLly
wZOowO0U99NW5lMpF8es+2ak1xalF2NdiW+EREELMlyYVcqBBloTsqyRH/cZEPYV+9ODDP2pgMjI
iSh4Ggagv4U47VhyToI7ox2HYMj5DlMwjhmnYfjoAVH3GXIz42K3SXMR4ANM0Wo4GH/GsvyBsUpE
IxGXTNZYyTdl3pZwW5bOqZ9K/Kzmtzyy4w2uiJJrSeyIam77Pyz659uZrcffVfyjLRqOfe2HzyUn
xDGEukSbeuJwdijo6cIlofcOfbDuNUeji+gc2O1QnXqraaUJYP9XVpDmO8CnKN1rl3puQSGBGdNQ
ExFO4kD+EFBvuG8moLYSPGhvf2XhjLN3vxk12eaqp3v9F+atNLa4eOGB3b1v+/Bd8swfN8UDuMEm
E4jpbzvOzHe/zu5/VebtoD/lgU1AXwAt3mxTPmfAR9oewIz8M0YqTjI1goK/xyr8bgIthqW7M5NI
n+A+sL5JF8DKu7tqXbs2R7X3t30fDkkZ/PdRIlL38FQCyV2zOBUlg5DgcWqd76nP1F/BuCXd3pIe
DjIVOELJ6Mm6fkt0m+W8KeOc3XaPuC7O9+3LJcdZRFr1wCptMk2LWvs//O5hUwFTFb3fELkE98Pm
o/iJIXd0h5rtg+st6s/C31iRhhas960YC+euzbIpzYp9Ddx/rjAK1AjGMcMUSJgMK8mJICKwtgx4
3OL7yYhw4KQP0JmrptXv1EMojWhKZ5kTPZb6/j0XsRkqzWbfJj7MY5fZ+zcQEF4SWPzcmwEvtGzi
CiGaJXu3onT+G/GcADXRk5V7+cdloknr2rkNWoZgOUdW4e7oQ80hM5nzFrMeL8Jz9UeRdphQ7e6M
MZYC3TsHiqQxtYXiU2vYTQml9xkzerm9h8zJaeiNklb3fKSRAI3Lqe1gv8QzplC88dM/40+KXswK
fcymMn/5CGsULP7kE50d3h5Ey74+yI2pfP8JJsd+lnlrbO+266k+TIGZJrOrQD70Vc/6kmq5zc86
abfl01BEGnYj6FkjuOo+Yf0w9vvVDwDi6nZU97hG7Lofqs2BqyC8pIiAUmCaB3ATIaYj182usfjr
0O9n/hu4vquzjpXcXsteb7ljpQsD9biN++5g4ur+erC7da8FqjQV5DdTlarYxt0/EIteXnFTUHvF
8eVZDscCsS+ah2nCIclGbWe6GDK8X2+fKbiZO4tKR0lu824xmkEyek7qoAkq3NQNd3yWeAM34ZHR
C6ZvMO2iDIDeROOmO0Vz/xwMGjRW1VscZZTAWthrt1CYEw3dNETj9g1ri+qeldnDsTFVN4ZJDoEp
iB2ZYXHT9zG59J6h2+OPw+dq84xcvaXKkLAbmwMsIxYFjcnZiy73xTsR/czuCurowh2ecndzOUx0
aGmnVfsy8MIWnhkISVb5UxsKwDwSAvL/HJsp7faFBgEmgy/QSKd1Yb7XtjSuECeQ6uLqUMYO4Cp9
Hwbpgquwm2nuPnnkoUCHbt1jhOsmOe+ubBOI/ROUgNO3dNWX7qfMFDO2vfwwNes6VGsCUscmNAeD
JgPH7UZHowcwjmYKW0u6omKkNb5PFtSHWL4vfCRr03DdT7zKqrsob5MYs4vdjFtsgOPu1WmHSpLK
6E51qzBAWXrl2n+rwebWMhv52B3l2RRrVme1K2cTov73dFDNYn6Rh+Y6fq0G2o6IBH006AScVzM8
L3HwnnEN738B8Iov7VUPs31TK3S/XgARFlTpZwKKqV+e+giuVMYhebO46KbHKEY2/F28cds7nf2f
AaukFyPkBUT0oWVxieWXp6a7wHGcKkqyiyvLBppxTSSMKFXV4tAzN916Ho0ZPd+DDjFZFCW7+iAI
HItxTYhuhhQg6TN9LoFcKD8SJ51fPfK7q411RQv3E0ebL/TNkSD5ObcOMxs7VynusxtH16yiQuqY
O0JjRsRIn/Y/0emgiHsY9MwEgNY4KKEt0z+CpIdjCqwJPutrbNA63IZQ1y1TArvZpwBCWLHi+ci8
0g7rQfug1E1D/dly9i6HroTpGaEfpi4EHkY1GxrIJrbX9yjBvnpqxbSo5UhyyvTHpX+4cUfQ7ajL
vqxyO+O9x+BZyksr9VedS1TgnX7jGBum7+awIMoyIRnGeLTHJ8joCXv2e35HAusH8jOKQISUDWZU
AfEDQmJSxkXmIMKMSz14SP+pBTChoupA+RFfzuoyMrDR72Cb3arJ6SM15kXlviaMeZZ0+upVg1g7
jQilh7vqNAbc2WNlHY4VLwURZkHU87nDG0LXy4kJe7Tz4Ld3U5D/IjjE8XGl59qtE3PY9ODwKk6d
hb3/Liss+0w2DCbo3WMdLdN/QROqjlBumznJP9GpSVp4tEIS/PrTdGBA05igYuGo28JB3OflL/Q0
d53MOXKKQ4x7iKGsCEZRIZJW1wBYZhD9tDipQTkZapisbGuxAUcI5Ndj/DN3GnWm3PQsfpsCwi7q
vCRxi0VelkiiiGp6uamcUWy35MHQNrFetbmLFymMP1mtgg6MF47tFxppObqw4IOGuRih1PhvVkOs
7j39ELcnsc+NOXsDpXs8OdHPFRDWeHpPsowyXzXUU733y6UavpL3bZAW7qihuVrFTOi2C/n9GEmK
wscQ0VR75VQjVb5wJMm5fh9+j0a9DtheKQx6Ic2kd55g0agg3eRozGgan4EsxvmNTa+T340by/PU
PMrhG0fD4mw65442W86FSy9EkKxa6VRSh34CuSMIhIStjor5fPImloiuCYv46D2x80g7DbTJCvR3
4kwgiG6QYveQf0qaVxLq5ziWfDXLrlZ+GwS6CcRCtdzBWYfJqGseH9IbqMOwdUMBaGQnB5bnt5S6
x3sBxbvgyoy7HwBLKdabPTtQ4ar2t1WLLCcXPz8ouAzmiS4fulqIJEsrlOBrvHSVTXt14ip5mqHa
twyvJWBQOrjGebMlhK9w35sybqL0JYQr88PweDz3g76gmnCh0FMTIvM2lEiOM9EGDkRGH16D5tt0
hymrmF2bdpTPLiw9VQEh8t+bejpHTP2AxX2ANJ9IOcU+nq+DMxpeI+d+BXaXOssbwVQoLhLIahWa
TdwoLuRXmJJs9rvwrXI3d1hyaB/FSwnIESvV8TwFHVakfjLop863F3hhweo4ylE4iQTiMlG/ptYk
N8QLAdGyvYbP69mO92Zms0OOAvZQTNbRcfEge73p4cH9LFR4GRdYH3m+l3deRjUFGaQurMqUU3yy
Q2ah5WNZpCVfLHQ8ls9STea1EqM/t40wkZUqWHyecPnVzH6L9w4ZFLZd9q//Jxecxog+jjL+PHis
zumQPmAjRAQd+JX0elrekZ8M4D3HVHQOLc78vzSsTecLvhUKPwJjDwI4x/TWo8eMJEb9A2n0/3Ip
rw4KQ58Evpz8kmxClf0g3QFoxyXoEP1x+aheYt2PWQqkQE3F78UCbkNelBqUN33VT75mWiwVmmI3
tEUmEynzGY9UaoHi5uT30KF5wVfB5G8ZSiTUVZbPrQmwNKynaHXhcLpIxnyk+nlsFrxZIPggCJ0s
MR9B6dd4RfLLfNcO2laJSq2eJ1hnRfkeR5xjurmp+uZCJRZWj8Pak+TJbUwn0zzAOXZ12xyRtZ6i
jWrByEl+mZHsUAiIbtjYzsRmpvjSwPTfeiV4hFG1MW/GTeB0Sod/jDT7MfgA7JPwleooBpQNC/sf
TH7Y0CBN5428SOORCu98D3WUCYGkz1wkhsoscKv5dUn7GbGqXgo4FLceRdyjkctaroBjiMDG4GxM
eNe3BwhwxjvRSv6yVFEuyiltVQiV1CtrrlRf/TOD+Ijj8xMHLvXBHcewdzKjLXRw1fchKPbXyOlO
c/Wm5VL1r8GcdzZkQrBOOzrWRxSnNfdybYR7b4TOYVdtWNsVLkp4vLqybzdDwssYTR9FBTICQiWU
RJKrCyyP9zShsD4X6T47HVCB9uD2UEiemn7kVRK4xsvZrtwoO+3mQi6fn+wZ/3d6RV+C6bPm9bUx
aY8IoF3Kr0GKTgRI32GnkIXEZ3Q6Bh6TeDwZfGvpV1iSXd0/QeV/hLyn1GCaqvTZvFgGmRBQiTLS
u3saLkck83T8hsNRG0OBjT04sTeHHidSFWwUoe83wy2i3YjixkQm09fy1qw1CsPzlErim6XLI1qu
+3/ka0lJHItyNGKSCIc9XMwt+x3KBt1dsfRIFKcJd7G3/dYnLQH87+lPPUPKirRU1SkX2YiAaOpG
r1Fx2GSr/9kFCK8C9+xquBK8nFuXau8lAVb02pyo9zIVo2i7feGJSLdlpTpKU1YHXilesL8nyLQJ
4GLLrStCOYA4Jm2tKq0GaR7NFVsobYsrTxTSWLwKtkf1dOsgg99+fas7XaTscd+H8d8aFkY8tdXx
BnN16+c2wDDCTedgdErJQvtbDFooWmsrZIhWPl03wW/Qqwo19U+oGWoAOc2rAYEVQcI1sytSOw0K
C7BJ4Co1ZcgJKAMm7qeEXZAaOCKFHKOG13rprhBIFBrWJC9MuDVtJ8QZdhFtHx0wmaOk59w4LUZP
kzz/r+wMY0Tllmtr92PsZr9V7Gv2yBINCpPtFO7EnzkjIflFNlvw9tmKszdEQMFY5pnYRRVQwnE2
TpLDZaoO2b/ug+fZ68USziG8IyzcGfDSqrPVj6igqJrNiNY522ci+zjXNswOzgxOc4A7yVxTGv2U
Vg1Clw3txwMqTP9VmYkNLKZ6yHp7Nh3UY3gD+nzw4YTcWXu+UBzP7E7CNtXS7w3QR8GiTsXXwMy9
dH7bH8c1yB4kaQ/zDNX4D1c4cvat1v06m2NpcAphA4kgcRNxmDPinyLXJcyiIOpggTReEd/D8eHa
QrmmveMMU60uzT0GUabPGgcGjkQ6hCDc+ewZKpxQoeCgvry1I5tAo7eDKh8uC9WI9tECvKW0xOFs
nK1KfuXoa8Hde3zRV15Zhe+25D9B5KY1kuJl2ZDIVbOdDm+gdsfdrlZPG+DIxSB+7RP5h6dksqvl
hFm7c/as5eYzby4oU020SuuZy5bxbc+IM5AzNVqOHP5LfCSxk8stvbJplYlJihhHALIPw9hSgVys
GRkNDYhcYd+hSzzpCQ2LJqCBEq1NG+omJLIZoiAS4YnlxX0YGRiemIFxkztu2VhdGUiJyqploWYR
YC9EYA9MLqK2/mNfVJ6QPuocOyUYO3jIDYQWhGDl0n+SiTDGoCGBBN7fR6fiQUR5aC/sHGuzEKsT
JflAF5x8prirphMqfWyxSMqX34b90HQ3mSGe2W4PBlsvyM4hZslScWy5M1zxtwpz/dRoe5d1kOn+
6P8pjpSU9Jw/29Kn1s+2N+mhUAbEqV9RulmiXAWNRKBlugfZbU4jmRQawNEovpIfNCMjsIxWdJU/
Ku/D+sdNInuNWgJekaVt3iFascP0dPMNzMxOLGwa4VialPopZPf4jVmc/A8u4kbPWVIqEQifajNV
/wNckkLFJGV5xdyD7BncDe3sdvATXxMt4gGAgoEZ/8Vq0Tdt1biOejHO+Flg+inRol9L67WdzVBk
TLk+aYZKGIkK1ewralGeqLEOjw4CH8QMFgCqQmZIiEDjbpcqEOE+p4FnfUetpcxvteigz9P57VSk
qN9BAK3/HzPA3o7wdGEPka9ejmWbn4MgX+ebUYgqIFHuqCKFS8eDSpGeBQgE3z02a3+tQzUaVwOt
Aiy3M8/JJTd6RZ6wZxHKy7Y+5xtTZMMvKY8KnV50utSyVenvmbMLO2NU4E01qk6jcXT9bbIycfBF
hMA03GtCMAbR3aZF6D/1ciaT9oS1M48FMTdh2uXmKp+kJhCzRDhbUYzy9iSTLNV4aLoblMC9a9uJ
NxwYYR0yINyYSMxyEh21qk6hcz6FdTq13gIuA7+JerKOhf94smu54y8eH80sNZC6gbulRMYVbuRD
xpO4hdzhcT4w3ytvOLvApGF18Me0QmDbNcJBPbo1ZDcnq9J6+sKhz50PUZJ9524LbvYm/WDAnQQx
d2VvyydgD50FP0oWvaoer8vQiTK8y5vjpui10mtk56gv0x3ZuEToJQU5LG45O+RkPGsNyHA0/XTe
c5oG10MrlgFC4B2lPWdgg8Wm4W2fCCs2MAjb41ebV4lWvxzudDRnbnF7uyZP9xjYhVSQLECVDDdm
UyD/DbLVLRVUdv6yB8YGv4CuuWgIPVSYUpuwyG5igb1g43vqzN5cFqiwIq4yX7VqkMQoJxVaiYJf
nxIFgI623pJLhQ4h1lPVSlxKBVkUjZIDJE42cvSbE7X+4Hl4OjaDTONk1UYF8NahMkNEp+QlpKf0
Kduk1JhYilkQvNm8PH2JfQQaMS6GDydxgj9Sr7/iC7LOtNv5V0lPmK0W19tATJ2ZDGRpbmpx56M2
4YemGLHXk7LPy/NR1EaSTXoy3wa46+1CiQfzqPPte5fA6p8IMdCPFk1JqPGvRc7eIRQYnQlIfEzC
cbCqQnnpnm47zD4nOCR81c0u3ZchBCGm+2FMNGFuCuBGc/CXGEwy/vuPjzP/MDNhXaf8WL9mB9Nt
BgfuYFINL7YwuAIfOxvT/66cGP8u33lk4MSqhyuVjZjWsTMGU1ifaaIUNEjTMITiDMDBugPoKigQ
vSPQmU6TvHEbQPJ6ej4UPKkCMBXyqEzigPM9iZvY7FT4k0JC4Pbf/cC1nvAakSEahaTAhHAW2zgc
gyqzGyjpXHj8VN9Yk7CMjfFg9mqvhhNDZxFGfduMrHPGTfX8cDQFy3hiLFxiSFOFbVlPhMSQUFu/
bvwwGqXWCpoYV3E6JGbG4Wqtqvu0tFxDrptepWAz0+1dAtdg2LtOoKZfLSeqAgjCykYUMcg8e+zx
zpTPcoAhWKYjyONHtT1yPzVysx0bPDD08ROTLM0CaYR5a4GpoQXDcIpVNuux9+4a5xAj2IigjGin
t75P0zIOGFaBE4vjR1KxYUl3XP9peeaqH4AHINkU04d+7OI4nUj3n2h6Pt2MH5WaQy1w8vAoh/qX
4afpxEKs5wiI9wQjlOk39SHKNVr5bUq4PN5jjwkD93BQDwHVoutHufzlUvQRPI/RT+/K0/pOay6Q
cGPy/yUcxvsu8yo7+nMc4mQGv8s/sy2PfIe1RGDzrdKp2Q0kQVaCQCNaC2QOUuguafceMq5rgb73
SB1i/DkkYcDLM9aQyA91w81WDZ1Eixuga8VHRur00x1tDrcbZX/iRRCmmAE7bKf8S1lkoyg4aK7r
2DjKL+mfgK9lfROMsLzGblIOr3bmhcK0wbH/uNI2tLgevveEqdaKdpfHlMft1bF/WgOEMoN8AqU0
libM693Vc887T9c8vIUE2vldFtdHEzirtnFznbZ/0cbvO5dNw6tx/Pb1wC9ZVaOpH5ROvhD27Ie1
/r1LAvJQN0a2Ld326734mHyeU6mZm7A1EFjywkAmGIlZcH//KUDyMaA9d2SahZzSpOmKEJ6b7Aor
BVsxj6VPfeyrbSZV3y2LFjEGhNDeDuOEik4bNIv4rhTFbogLnFJydm69gPhV7JdwU9OsIXBQzgw2
fDhR277dR9VkjtidAgbT0+GerjMZPuxn9XChTS5qEiu5f9LaKxtc0RuZO8O8CpSt+mp2Qg3YFedP
Mr05GiA/1mpoosXhdbL9o0bNch2E6Nxn76iRVbIWdQJfD+FrK/7d/UwNeNAL7B99omBrhE5FdkG7
fxGqVpTlOUXaR2N49xGa9bO7USfPA6ACD6aezfi+LuU7aP2ODrBkKbbdAhvAJq1bRaj3Rzs6Q8ic
WQ82v9T9F2Uivn8qlMMTpshdhXo0WVZw9X2ydkrJ4pT/RSeCd1GmuWBeeVcAMPCX7xpqD/4tAcq+
s4uOqdgqh87U97TCdyXtHm3NSCVyGJ00H7NkvWxPS2aLgFiA8cmLJLyPaJ/QGkIvnt0qwwzpMWdb
qCwlIN/iZRlLpmrEt+JZpIsKYEDleAbKxv9h5q6JkF7GnOYxO6Tj32NGzAxV/VwW8Kt2JGNA1jbO
5IMVxMzvcD3Av6QBrLh2B/aEeQQUPXkL/bMNUewa2kiFQ86WRV6+tizHcAF00BPgtsYe+hXZiR0L
/mPkAh/b7MhnKPmtP2FIuSMtm4oYmjuZZ4jdcCQ2Fw/8mDfGiu3mapJlZqQluozcTEWakZ8HqNob
FipCcdh//LBO58Jsa3x3fZqsLezH22TOOJdNPwvwNbQMPQL+epdARIunZz96308U7gqCyxRYYU1L
JQHL+qtSnPVV3+TSOkCGZgVXhkGEZ5XLA/ovrZfgdqTaC+7FReh68I48xOgpXneJRBoAfVT+ejlp
JhEzanyP4N2M+xqMnUtR1wFcxwptNkebhPpoenDRqAKIep87kfX3DozfvO9RFRJUK0pZubZD9z/t
UTzHQaSITHyFxzrcPDorrvBY2se3Dpj/3z5YN7omR+a2l0T+gfxYhcPLMkD1Pfq6VLiDwdrm/apI
8miXe1Vu78K8Y5P0dOHtomfenKrYtpGOgTZuaf8NrgsiNrz8HP32CNirNs3uhzu+Qb/eNKngRuIh
QqrkDHLJHRtedP6nfZwH6w1ld/0lzLpQy5UTn0QnD1Wxk7zqKzy95P1ju+XjoLJ6F7C7J2DcvkJZ
qXKrIBVi3GyM0IgOOD30XF4k6Q1cuI+/w52h9JRfEO+xYywJ1uUPgG0M2eP3N2imXTb8bbziBV3t
oKG2OSTbzVEZ6A0ZybPVtdKIwFBDQiqgUF2tBoHtl3RuM7Y20ESn1MtUTIDCNHWzfYw/Pq81ks2x
R/kkBpZcfgA2crHCFxvl7LJ0Cn7kk8jjFaylEHw6ozl2seHLS5ZdL9vYHXkmogNICXTf2TTY99Ya
FuwnAtzf53k5DUwlX3VhHIg+a4w4k9No0ADzAIiMTG7nwVKFly6ucm9vnyWVGhtSpGX6MO53HQxP
sQOwDH5tDwbWLLWbL8SchGnDb+WVGH8UPN1Jdh3nT1LV54kJIEo2SjanDul7mbTtH5+hU5eMTDSb
dMhKfpi+PnDV+aijucsXkQqS9rxiN6xuZUIpEAFHaPGrhGiGCBAPYZY6O5GkPoLm4IqF8rZz5+gi
SHXFdLuh6kapBPyFJD64Z2QQFT+qpOOHK/ts+6OoJ0l8iXgAqAL3ibwNlxeKcGpNd3swBjyCmR2s
emIfY5zZ0vHMtF41baljej94kmg+PrV3by8DJErxi+kVAf5O94HidUTQ8xur4iUcSycm4se31Dhx
dcdDxf9wNermvcSdl91cxUZEOqZMWYieWonJ1LW/9wl33MgrFGk1ijO1SHoNU6vfC8jaqqLmTVRX
hxtTQoNyE/rH1Zibp6hdHMd/aqeEnXk7JgSDs0wVAfxfeb7Gi5wxvkTaaS78ODKxqR1w6eKu1MLN
NH9UJG/uD6asYV5zUCk5Mz+S3Ohrj53XGlwQELHuJ6pstKhtrBvY0M2B6WqtUrrekEMYYr51BDCc
7lt6yyL9zFEk0NIwpj8AHtB5xtAxJKLo0R7Pe8YBcBzIBMfDSJW59xKkqy7NvYn9UgyJgPQsudHH
RkOqNYBxv2D8R3JZKzdNAGPFFHXQ8MZ5DP1Y4lNxtXlCYF07YlVPeyHHbNUlvl7Ce/miS18x+cLg
aSrHeTxHkhhJsjMImjWqWj+bpBU0lfAC3Km1U7yC8/7xkjNoKrZN9lvv3CkoeuLRF+kSH1E6/Lsz
yT1GTNDErNwJLtZZs7SPSkYCPH9HDcPkFS0qyN/jWVAe6odHs5vekoGY5FB5MytR/ci49OK31wu+
GVvtM6JJFS0WLyujjLEK3YZgEhGwYfhIovwTarInu+zKHOrY0QL1sGxVZDuYLHFyPSQfSZcRu+1o
gPruXuuAZK6ZrFFvkQK95xOqblSVAoYEowkwh7+0XpClzrahSJFW5f9pEhx3dtzTT+jActn99j88
TDTQbMKfYv2ROepP2JSt/rLTpO3oRyGC9imirMyjRtGw2zI+O6dgZt/e8tjDH2TTbDjuuRnbrzqv
M0s0hUbStalMZvbh50D13ttk3z/tyfU4cri1cBDRyhs5UoleKt34nWg6LjRxHDvto9h/DA6ru9Uv
hxG7vtSDGD6sBVyV+FkHZAYQCuKaHJ3FZCuHSWnUvaZOU/tqumq4AxWb92jqV8IB9E4EEpkStuBp
FLEUDDiSo9IBv7pID1Ufm2d0YKZdFvulQwB49vV6cAQHARRfXBC3DVPiC5U0/VFHBWGEtpyng7IX
mrR4+pkYU8DemfVFHEZlyycH4IFo5bKkFnWUtYJ32LVfW54yw4QmCXy8ORR997ltD8ynE1s5OmFM
z0oQfDsvZnGIwyAgOTm5EhRKm8IioSQnf03T942hSSRtSBsTZQuxudw/kJYRiC+fCOHFypFfjR/y
oL+8JatVG6TvGbaNDQbR/HKIgIf9A+E7iB6US1FkHVp80jD+Y61iisCEGy0PXaR2pr+D98JB/wbG
VP9OqQFiA+I/2SwPGrB6Kqsh8WUyATVVWN6t2rbpWzq8pm2AFTWhFUEIuZMG5o5s/jj/jnWioIRk
izMbP44yVck7Ew+9LiFaHomoNI30njoz8GFZSq/6QwILVO2GCAf2WZbz1UXazmtY1JySvpJlrLbB
Hn1X3LLIadWU695veIA4TF/nAANfVAd3W1xL2eY57veU59Ryv0wOqZGUQGjlpjp4Ej8PjH4eblZ9
iWaKz24qgOVZS3AcUfsMUUW3mB+5rZP/IljcC+D3vEIXgdxJtES574mb+Z/xDfP+3u5fYttXzC8u
XnS2MskzojohrLUNetpURUe1aLXsyHOdnTdgei65LS0zUfZw2VZUUQaEX7TQKwXrH0OSq6vwLZwo
YaIG2P/LeKzoJwjHMmZhXSGXqcYe9w7hvpsGj3mYshFCO9B7GEYIZoiJSUzANprIu0quSxRP87+5
5MSX/PWBeczxrNMe8D43cscWoUJh3BznTA6riEHo/Aw7OD4u4RtGnxs9wo7KJmM8QM4BtuQZeY5D
JHgYvcX39rr8N1Fr5HiWcPTyeCNXgzfdpJpH6LyctSt9czgW1F+lvx0fFMffdUH1HjkUlK/lU8Zp
YYccNPNms3YLoF7yqO9SKNmqdiJnt4n13ApcBdNsG56TOronZ/cebJOXDtbYNNCo1jSR87KfQHWF
vQ8tJ/1oaQ52Ztvi8BKtHr2Eev+ClTyQNDL9H5Nywgtw1L1Y4HfSOMdg0SMbGWWXwp2/qPCHqzEI
MeHX08oAd9raj0AvRW4WN5RC4jmOW9KpNplVB9rrYy6WAu+FSChdjXHC5fEjTjCq8gexpfGdhEu3
9gu1pACWKpXzHp4RP73CI8GzpIvOcGkHAouWkiw2X1zZCJN2/PTbUEMis2jmhgpIobJL0NVvPDQ8
eXkxG+NB5zFXPUdakg0x4jdwD92WyX92mdFNRKfX+/ZGim+mAU+yxsoq33AuvR1MTYggR4JpO7zk
1Ze6pJgd712zsE+YpI/9ijLrEXyfDG0U7t5tJeWcyKqmex/+kMYmI7eUku0SDVellqejXT1T+Cg6
vfjhlyQq2YpRFx/qkWiCerv1Ocer9C7c3HMl/6TRMPnt20D6coQejPUTE8CMqWvkrxUmO53YmLfC
CXz6opKx1L+5amFYBfPElRC1qD5vSf3UnyRH08nTyQbao3cC+4y6LblfUOq/uLje5RqG/elK/RsC
6fNgwQ9n9b3d2dd5ajBC8592ccLypS3af0J/mMqx5ZmA9ZxeqlHWXQqQE6ngglfXK05XSnTEmjZF
jmuE7SL0AJOG526kUAHwRKA6IyXLWCIfKg2nh1RagEBY9fQbBn6Sb5P1N8LtcY6AH5EeXF8oupd5
3Kx6xcnCAVIknbPlQ89UheIGNx1zXXUNTIFbzTIlCBYLwJ1rYKK38i/O+8ICgJQDIJtTchgRtQ4z
jT6i6JHKg750mYP9hmgmKY2siwk0J5VkO8whAmKdRlA3fKtnYUq3qCem0VXesyKXeRC89XKZHS0x
twfkFD+8kyNXbAVQogVXD0FV3S0nODhhGp5eb6AOqw9DBCySu8Ga1XeePjJcwMI2bKviAWnFB6uz
YKZ9KpyxbXj/1Fh9gO1djOnTZosd2MNAbG6zDZDpX1x9SY7A+xNmJ18wSxRPZS74QAM3kL21nSGv
EnfdQitsCSdqsdcJe6sDZk6BPn4p1rotJFnd9HAs1NvvON64EqVlImUwb4aHQpSFCjNRIec07RqG
Et5ynAQO7zQB4A02MEor8a7xfr2b77xuerBDHw5gT95Eapc4DC6Kw1XxSIQD7CmKp7Cxb34fshIt
4XZEHNnK+o1JEo8l9HsneKP7YCJiF6OyCdFw2H3lRB2ZsXuUCX8rGaJxZcvmB4Wi9zxiRJkioRmG
1f4vKYfGGJUIo1Cm8WTXxWWziG4/5BoDyUFssWw4T0CounKqOPNNid0LGqQwyCC88OWS7yhAzlvv
tJ9K6yUSLasGBCg9LZ52BasLlQ3/7U50UV69meEQwBHDoUfNOVW5AlPf84gHyn59Q3NNZVfz+BcT
rtkeU4lCB4j2dOoLODXBmPyi/de09iynlQq6oryKuM+3RL+OliOTzgqcxc5IbmMcGocg31boIIZZ
v4SaCsYOjDM4bjXaQaH89J+saA46ZwjLj5w31YSsUB6ffm18onPKaNGAyZ5bOeTjVy3gyzA4F1Ou
0PoYwiEprFM0VHMxmSNnaMyrcJF5MHUMnPfCn4g9aN76mKua1MtJNLeFPg+5ClXx9Nbnt+dbtc9e
58DHmHeLR6LZsyUhTFEU3jROx7+DOFdN8K/TUmWBeY9Jc9PG8wAMr1+scAmjMFtNt+SlQ8Fay/JC
przI7ttmEkgu3xIgTZWxBO1PCPd2T0G9eQEKfZ6+4s0ush8fFwY2SM2N5BieTTZPnlR/5cFJpaKY
hz9h9r74FNSRRAGy2RreS0HJWYoaD9O6x+jQ9o7c3TkGn9f/iO+urYhJooX/BlPlysfMl4SL9ZVk
zn2EoO2CbejRdlVL2GGoX6ZWs0jJOpAda3jEIlwY/kQayM8yi72ePvjmM7g+xXC5y6r4Mp4aBWzj
NN7fKJGkh6waaYWf2TlJzs172oJeQyfV1QhbqxszBsb5pXIYE3RONIzqXriapnP+EAkNh2GIVYLe
xkzYOPrsLnDQqmdHh4jCswvgf7pOlf0RTXVfTxqqL5V/7Ks8TVx+pR82zg1J3smWexA5OKWUX+bb
0Ne9tArWvoX1usBGUdIdtcHl/EU1ZcU4F427k04mESMLhD20U5+ri2mtlUb+f7P1nfJgmqf9QVmq
kxS6hyHEqJxGDOL1osVwF34sR1w3LvgHBwOjEs/GwwvtD/k0Si+ZKYSFmcVPs8VxeluASHlfJrpL
DrOVWvRJMa5W+Lv+fzFqXbZpQ1Pu+eQ45KL/gN+EyLawN48cgfpFqtmzA0GgF7dJDXuIXEz6DwQo
F9eJcLSctXDr/Lg3djxBkDiA9k0DOGOgGOPiBnQP3aq72gBwGOCZOJSymCCnr767DuG82vi0etFi
lQlFy9oesk9C3sJ1EcEQ1wySqaeGT3rzJt6TQ3wCWZX0+LKFf8xYA5Ad2dDxEEHMGdhxclittzdl
M+fxjWW7CdCAaQagwsifoHAh7TTfRMcKgTjaMm9zy++nks57pMIi3fOPKl69g1qPN4+KXKIZ4Z2u
MrefFQv8cmC7uC4XJ80e+TgksO6JGD/N33gVvcSvVr63oZ2vCqMkwRqbcHNlCkEXjHBFBi4NA6S1
INW8m1VBfEZ6FhAr44gA+wUMcahDwt/89kZgdBJJRWKx23K2MXaIcS0kdWSCjJu2d+lm2imldnNS
MrsutO/GfHpjx+n89hnNphxc2jdACFivc0PXFa7JjYsAkwGMMGB2gCsv3DqH2UCUdVreyiGb0Hbs
GeFYHUIQ97uX1gR5Gh34u83VJOQKAKh1Nw6+OfBHxcopTFF/5o4/iJH/xR3hw7w7bcKqDCaUfVrI
83+ySdsjfBPvFeMCz449x8xjafc6rALDZY6PpScd6Q90TfSP8Ff0T9r0ZydWgCscamSy/KUWoCNE
heaAWSoOH/NM1qXo2E0vktOqmhWt44YJK6cWHJyFfTB1mU9d6tm5rsiiUolcrE1q4qRMF74GwK4h
umicVFZruE73zIT4dnX3aitJrwvS7hp4xtKf84Qi8AN0yvFLbRmVGnGWvAPaiE3mat/1+iEVf9nH
w4Y47iCwOjhO7qYTWkuV6okNhKvCfUEzo3ySYiaRdhK54O03m3VA4w5khFL17E4GO/OeWtgwrpjp
MOWuTgMN5rJSYqyE+oUpEM/hUFzHFbB/K18H1vWZSEfvLfMNjIPLTSz0h3qTU5KEulbZfKHFCLp8
5HuhN2qX+2nCgYnWMGf2XCGNOUXNtYe6TKwpcQxQwsYyKVAJWbpmA+j6CjWyABtefN3OYJJzInGx
9TLbWFiPccRLltpScVZFsxfXz6yP37y476vCFIoQ0w92FjizoGZM2dMgUUuTcWTPrlPHlDvBAE93
7E1nSzOiqBh7Vh7/VF+DCqfE7Nm7dnwnLlQPx3X8UI3U9yZCkV8lQa6JYiBmdRnL+c80zN7mleBz
pI/l2Qffu57q5Ad4e5CR6d96+7PMc31jwPapT+SwiX63UErFjt3OU43jdtyUAxLocT/iQtPcJY95
WSmIlS0kHlYu+5ljYuM5wsl/m9XKD727x8i/Z0p7R4l1KdZjcHShENVjXGRMXf/HzbcCBUaI87nC
j6SM4FKc9G9KPNQtES662uZlfqWXgs67/K1diuUVdyuY00mVKiO2QQ+Qc0ZkuZBVb8UmqFJoFusJ
5g/u0vNEXW9GAz1EmAsMbh63jJR29nUmALxZFXDh7F1JjxRHnq/2ZnhE+H3MB7hADN561yejNGNX
bhmWVSbhEy3pmWxoOba7+QDzrEvIB68hISssJb9IPLV3nWASN+ziwa05/gdRfaNU2gy2bpZ1lNAH
0dmI3I+hKp2b5U2xwCCI2D4aHqRpwhaOl6uwXh+MwuOpOmL43VxPixjQxlehZtxlz4fNDzhx0tW1
CKRk5GgZ/0UJEYdqjAfzjH8xOYgNzdc2zaBoK8lM5r07ZMq5Vc1Xty8FAYRq+SkKqA6J3PO/rqmn
RFkrGg2Gulg+utwoBKBO41Lut4fUKsf314OVP835Miua7SCBFxgwl85++3kgYYZhqBL3H9oQzXA7
wEyFoMlb0BkfWGg/FEUPxlwASRPXEWWaXz+KbL6/9wWzYTjkjRCzPMBXsQ5IK+Uw1ud3rR4NUfoP
LZ19EGR6CscFIlTRZAogpTOnMSxusAP1K+Sqy5/5li7aviMmdDdgZsPSyd7H0zU6sL/S4LB0XesH
k6vi+HHC5WknEiFughh6J0wYr3eNV6XhuSJgAZjqPwLi24xh8KdAIVwyJtccJFCiByBKxW4T/IJv
0YgwCBmscr6TwTba/h1av7EtZWQV3W3n1iOKTs45ldQ+pHFMcizgW6Xrrzh1Qe/r8Gx10k/MZXn4
1mp1+Gmax833WnZUkDikFIDFxZyrQ5daa2sr6ZwoNkieyX7aLvKvWnoEc39j0f7aAGYV1DW0JEjn
yNNxRNrYDLFcPnvFsa4h5VDsrtV8AJjU0Kf588ptJeUYlUUv36W0WeuoS1uTeXwEmzmlXbt616fN
CR2JZNwuxf9gGSN+jUVBYwfGvv7Jrv74PsQKk1XSI63a+/j8HbErdeNGoIiW68tyOGfaBwMZjcHK
KIYk0bLqI46UQS1ynnfrhC0JmBx7g/CpOHlYP/Xnu/aDs80AbsFt718/IH3fM5PBTH7bxO05LhT+
T6uuJ+PQG4pC2cDC3DP0NbckP07Kh9zyQQW/2qyaa9PQ5eLHwOpdpgNNddsy5+7uvaM/jQNKTe5Z
tn7VLijK+WGenQ4BC+8a0r5ec8+E01oIaFiDM4T4h77KaXK8Wfrp1IAyKoPsaeQWhovM5h1i85Pt
FKBVcG/mUQCusjNT6N3cDU42IUonRCWnxyAC/B0aq6LD/bs+gL53TjTHHsautuiU+RjV83oZl/Jl
tjAKAz/+XvdoySW93M1WklwWreiCZQsfDbCZWfINqm/gILinQhs7/cVaz3unMt0k+0KL075lSf5Z
u0dn6BtIhvGCwiUAYZqio+DR2ZwhCLK1jARszAP2WW8BLjzKzXQWEWgf3Al+r5JFB0SnNJrFiGgE
7r8Jr0N5AFGwH7l+lr2pxxljgEkwGM9F8J7nXX867O0oSPiAS8IoFxODw0Amf7RmSxUcKa0s11tQ
oOZ0s5kDA1egfTNFAmmE1fL6N5vnXJb9jtplIrx2c39U1pAkG/qWxlK31kT2KB9uIV8YxUs4EPNQ
4djt1F6so7CYnfgb3357Q/5R1+KjQp0GXt1R+S6rpBZJyu35idt6Yw+zrY1zJjnJwhaIWYVLaUF2
RQOVqXlBYpWi6TMYKsEg5Qzt6Luw0lVvMkeBuuaJT4fuLo57dVfkVyhnBm7QrM6doySCp10xVrzs
W5D2+El5dxjIA6IKBrcGTTi2kWNwGTOcRu4fJF29q0JkQd3esqRgF89vL+E9mzpp+Njv5ToX0inr
7nahag+lzfRLiy+mI14TuRd4vEaQM3qiDMEnlk0yLnejOrFuEnnAM1k2i6r1MWV5EEDMJLEv7PDC
lqsjlBhjcg/5sS81BU1yVTOiR35d70Xox94d/AXMcd5jC9zL0G68InLN9X6+1cMHACdvp9QVZBUO
SzCF0ybepBXRwtSxpSdC7Y7yu+w0v1TNNT3ugPojlak9Qk2ecXJEGjL6qh7tuQqdtqdmTWJQcjHJ
a1Qi+Po+gEPw3klT9BBtos5yjSgRcxp/VuVagSrO53phAC6Ht6knjw2gW7MgzZ94taTKEZN2ZDYM
fyMCPyLg/zaBG2P/Tn/R/DexUrUqfehUmzAuAUTWMSlEaj5+klO8fU0CZAAo4iEiE/9LCdChftEu
HXsIpXFBuK0FDZuhRDB3GsD5gXk4FkJYH3qMri3Gi1nzvEc8+Kaio3QWV0lAQ2yRSLSivsBb79L+
Faplhf1Al7kdLQoKyMV0XB7ne+5QtG4mTM1t2HO4Bxp3hkf81N+Mw/cAxSof8yNw3l2ofWr9q354
cpSvLzpXqGIPHKr9+YV4s3lGPihd8kCmWLgf20jpKY2We8wvs9gtFXEjkGy0acIM8TiY33IrhkaW
nkbgmuBEIdvTd9x4IOz1W4s3dLz2IHFc6nADV1mZ4xlzXZZw4QAg4FZiKszkJvsJh2gX7utNm1t3
MBuaMrw94h9zLzZ6rHom1+J6Cp0PGDEshPqT4o2RojZxl++Hc7DERWHWquiE0SCk9wpYEqm/MiQ2
I0NJFUdrIdY0jwbnc2gPJff+SaRPw1xowP3+nyjuiVxEP/4htbXzTjK68Esc3AjqtNDFU9nDtJ2e
dKs3uJLCRF1Wps5t45qQgMdBxvWKRFZh3fb4TiCrJZsS/ipRs/N5YJwK+88W4TiJtIaAEFnE+T7a
0Ku1HVnAHGsmjsRhcZvC4Ls47tfVt2+3ncmqkbeGbMNlo17EZyJS7SdF//fubaWAZVvtMIEwSdIp
mXJs5dEB+NhIEGKdoY96z7lNpZ2XBPMhnG8u8BV6kRX8JRglx2yPxVqcoMtY0OFFPE19twKOY5/y
WkwpBA2qsoDRjHajemLqjyWn6PfqhI+e0Uh2veqXG1zdewvW0jc+75C9D+xXDMRZY+I5PfNEqx06
UYhoPuKyEMnKiMFTKJQE1txUhL0CmCILfKANJkYW5BAi7QdxCaP6dmI9DGa8/HFDEzmO+b4lokvT
LtR7fp5HFj12mFOv2sauVA6NXfyq5UQtZRc/HQe9MbvD5DcGgymhUc9SEGJVzn6aW7GT6HKhTQr7
JbdnZtVIJJIkeLChPUD/0X2rTNENwOc/C1mhHOOMVVMNK/WrGDJZIJqyzcnD1Z9fIctI5uT3h5si
B1syHOw1rzNTz67/zbUro1/THmD2k6Mll9o5bNk7FjjWqgGINqgKa+R7cfY05weeHl6ohajeEB8P
ks5+UBFGgbUNIkZBkz6zkWR1pkqMH+trMxg4AhKlccO8MyYUCusiakjMddZe4qBke+K7VM0ZQIi7
fZQ5nJBfJA18C8soUaqHjZJicFhlwuwVWt4Y7AZinSIpM2/Ot0ipnQ6kxc2CNMJykS881JjXlkLM
EC/gAXtuCDYa3UWOY7WwCizKJBo3FtjgOvx11EkWBU2UIX8J7lxFmrX06qn/YwNw1l2CMi7C/ePS
deU7RMoWXlyPQNWqzDmsxdm1hhQf50mZmy4kxvGEL13EnDvloNZ/PZdq2ZJS8bLAPz9YqQ2JroCE
LPdNejfhHIpmBRbkWWthTkMYoD2zLxUuRCdoSAkR34mN79yAAdBPYdez+OA3deQiMY9wNPt6CRnN
vSqw9OH3W7nud1QJ3xOoBLbO5jJ6AtXjGKijQ3f0ezyRBw97qLCVEChbyx9BMNAfBEM8ARISmxEB
mc6KwArTeTurVQqgvIKd8vjvJv+arNqFYDLjS/ilq/zNdsQ5DrH7Ubqy9ng3FQS4/cZ7bJd7Km9f
dJYesjsoKn+usX5kk4rQvi1V1+ZQT7Xj47Ux99h+wkrKzOWv2usBFvOQ67ga7QGxERApv5150yiw
wkwzWzY99/e9cOyEC/I0hTmcNhDmsQsrDDhf9+eQqjBY81cAEfAebYvnTWQkxStM07S2MeCagwCe
kNTibDZtCODJWgYLNFIJULCmyagc6PySCgjoD2t/GwzKK5lzHN1FaybrXteOiLsFcMTbAu7cTSx/
bpYby24PGCQNLWBtSnbONlpRP9woDmkpLv/mn6bSbz/JZ7NLAA3zV9Qtk4pIDiYoLp+S9b5zissv
djOz8hYe6UqQX4TIc63u2f8i8R66SYc3hAEparo+gQ5nmI8knJBsAT+dWE35eqaochvGlDS9lUcY
Zt014wvwwjAVxBRqjlBZNFETshRNIdaMvbuWIy6OHo0VpxeR4jvyBkG2+jgZcvg1ZziYJkbE52qY
N2Eu5VrJxikbsPM/5iTdkEm+SzdtE226Kwhw9HeP9fn8xGdjD8+cQH0xzsLbNm1u+EPP6VOJ6YlA
lfcs6p59b3Hlt9SbvPouLACZQvYlN4GRdzQC6TQlXlAARgBHhd0ruweXZokgpya+rDIz4LcJGYmh
Sce+qSoVrer8IZQ4Tfnkmlv5pK2tUtkoq260hF75NS2404buFCtiJFV/OXQq8R8J6yDPUqEtEzPV
qW1/yoTkU0ScuUL4VIoQIAh1/iPlYGIC2TMqhh68k574yi5vdgg4pGdbsLqdh/UGbit90+1U9/5Z
qUWhdObuHV6+xtSD1/AeEbBgXAvNOzSIjyEr1xDL2XggfpgmPHT5M6R57zzzARQReLxVv1JWVluK
GTor22+bFOPO/rI46AAYRX/eKNz+AFEy858Rxz7hJpVa5gg6h8MySOY3IDXLg7aA+YwDoEaZ4iHZ
ucQ0ZQgpX24MlM+lx+Kw+kS8IwIctrBwbt0UkBpunG7O/jDRlShy6j4oVQ9AkDVJuvCa+Soub4YP
rpTsieZGKZoVad6X7MIGOlBQqE2TOBG6k8ZDlstRA5ZRX3C2IUUxkXNBclSpB45fGZU8uqytLyyS
b8wmDsIjr7R1onnCoxZdyDiDFW9MP7zALArLA14IZWHxrpjvuOtLJ/wIk3X5rU4Yl3tUVeCWBErk
iOgpwM9WXevAmp4tenQ7s2xlTDoA1U8GMjD0ELDqevqEW8sy02L4G/HXzmysFNmlM/TreKATrlWz
eJYwdqcMTMADFy2zvBSafHSMwPzwyDTA8oiEpluSWu3PBoxpVw8GNq1/ULBcazFApOf9taF4JUjo
xb4snAcqPaK2LrIfqn3DjUmFXuH0ue698WA35Pvb3czhrsPTssHh8dPYorRF4xEKMF0hH/rkN3HQ
T5RTEgKoLfYT4oK56QGk4UX5l4gG+OS6awa4fjGjmpFvMtqq+BCtMChNOaTDVa9+ir0kJb8lJw6+
ep7O2OISogdslugHnMsuYkyQSPaa9T2AMCcHlKS0pKkxQ6FrFhc7L8WmdEUrbB31gvec3wf+xBcY
xgvdnmV0/ZwBlGgY7EDdy1bZbL2RhdK/fgwJsqxpnPvv5mRopNlyLsAtCfrZnLs6G9pL3h6PNKHj
ClnajEZ9jaIW29f+HsmKx6tTQIvIDbQrVrwhNknahfPMf2gKf7mjSfBLU6B+pR9p+bVrT1wmEDri
V5y3ETIE1HkraTriDL+xxTGxMY0A+VYyCnY2581Qcc7IzrP5D1mDphf25F7nUgw+0hfEhoEKc0fG
btFKV5Kf6dOMA4pIrdxqvbIeCkz6c16RnfWFCd5onHK/V8/oONa6GIuyEyx9uHLdLRyVFPN45/2d
dHefvmGcENzJrETrimQ0
`protect end_protected
