-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Tp5zgvAu9jxnpMg/n12bbWIlhxDhskHmUsEiP526FHU41+s0MRof7jq+GcFmUNpz
Fpw7kbYK+ctpnWiAcviYnSkdoGleVNu9WPvyVBqEDdZb+AU8k8It1sleCLwTEm6R
RCWo6ZT4bAMdK85P0cwde2gKBx2Owk3nnjqzPbh21gA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6016)
`protect data_block
A8nchRrOFL+7AwGBHrs7BXchMqviGX8kJ6014W5RUbca5RW3pOg/yD+Ci4Jc667/
O84sfqYRpS8PGM20J4ye/Dz42jnpWVwO3TZ4G/1OCtgBOjFUZHxgxWk0W7iK/Eym
gy8u29PSLYhPBqg+w0VNbb1fYAYMBt27ERWpcLNQWh6NhR7WFsFjfwd7NvAVwoLR
7j+jFmLMjmcB5vyWOnRuj9U0aye+G211DPNM2bV0TyiR9dPfsilhBDUwBiketv5D
ldJMvhMyQbaZgY0kGl6FPDV3VUndVLiqHSiJTCsOOGjL659v4LFoyCtZV8Yh/9a+
fvLw+ibyQDjjrumasGdq6hzlH6ZjVJ0Wu0vX9r3sL8WWMqpue3WQCzET9ML723pm
zZ9eF0iotnV5l1C7uQzZYPXDO9QYLwfrzEs/A5y6TsMPaMucpadiFcyMdvSmuZfF
F55yKUmGjxm/V89FePWr1sbLU2h/uzyVkOUPKs20kbEEYdKFEqm7mBAFKvHco0Bt
7LtyBj679pk27kp5ObUIV+Dgg3sk9xqcOVAgwOh9m1Z+mUEVA5ay6mf04+63vVGF
f/dfONEyvm9hGjnJ/V8ItLPaNWNdDN1LAUe2X+TRq4xJT33jx2gV1CyR9e82a2+b
cJAjFk1MALW9vaEqKwO0ETWEFx028DtRDegbam6OcHqLDjNNyTZYcVZGYNlDtrOD
YMtp5s5EH6nY9/NlY7Ypykgfwr/BV5gyEvP+cgjI6O74MuOrRzcLSJ9bPV7Hlxzf
F14fmfs4QuJ2PCUw1iLuQbBgRrDLULb4htBhb1XkpPxbvFoY1FtqzxkkJdHeI2wI
UbxdjDNfwqZ80OR7B4nkkSW7Ug0xfgUY0qYWpXy2OgvoaFVDP5BApSyfxhJ6oDf9
bKDV/Q8TipgQHw5jGAY9O22Uu8FyRuPaSSNKkHoORx46ejnc91rFr/392hhftomG
9K3LyYJMnQKbTivnYSabt95fkjnJp08UMNyzynY7OXREqkh0hT9L4RC4vpsz+R0j
Yb5fYAw8NJUkBat4K/SylVsdoiGycBYTZP/wxSNlYOcyI6pSqaoGwBmA2hxhtPJG
4E2XWTzQbPKua8e46pG1+s+5VjmMSFApo1ydoM+cw5IPXA9ICGVaUnYsetOJ49kX
6P1V9vQTNQui0Ao9qt61BiwxLHaM1mngQI6r65qm3Nb0aKehQ2gIek9/uhr7XpmT
5Ub9xPe8DwJXlJxXy7TKYg4LpNn2xzZlavTJX4KAl9OiJkzOxx21+eRN19494p73
m5lR2ubsizwGigC6kcjg2sf7EwhR5xawPuer4B9vA5PPDAxTdLokng8HRHcr5umd
vM5PU2AQESul7S0GP26Mz3UQRIA0jkSHQQuUscTFk9esSmrWjNCUdanhl+Zz3c6z
HnzQTSQ1/WKdUz7pR6HU5Uiq6vDae2Ath7j+u0hfMwcxTTNxE4+uuhcUBWjec1Nw
9c0uklmhrdsOVbtiY0r+T49q5E10d1/Xlgjebx7DciuGuznXKzlajnT46TO5aeZM
7gSqcvEFTX1pJpY4LXz92TuKo6qXZEaQo1Izg49edRwXAyNFtcXVngkaTN/xNJ2Z
cWZEJ+AvNUIugNXB8L3QvOFTVxRRCvrqNfih+l7rIdhFtqTUfLDCv3ErV/K3JoO7
7047jNgKKC7Vxo46gqc/LDIofHncpJaNNvP5G+Ezb6qlFjkFa3LdFqEULftUamZo
fiCTOSWj9p73/cxlEgpv3PelzLOcmcuPAjGzU3CEgHROu3DDvfDnFa0tQe7h2Wsa
YyIbTIrFhe43Z+IDyiHwnewvnYuUcwr1O0HxHJ7J06AeNEb9I3aGuABXPPEgYJWK
gPkaPjkdkKnVqRbm8f2Q9KRLB+UFJORElngrCCGwGb5wGxAutH6tzbKifvOLon9R
H9hWOGkfolFQz9prCySgU1e/HPF8biBfKqrTDjpCQLNXTBH1d5kXLictc5PGJrHW
yoBtMMEepVcPbcsk/+Fds0BPCOvn4wei/QorV2Jx5ah9+U2QCkm+m1kKgBs7vyHA
+ZripLWl1rzlfEbX60aLR+pBvYa97+JRziecDQesTOabY8rdDvHY/zKSUvElR5co
CvhCptWK4aYlzcVkswYocYgWCoeznMY8lcie3Wqli6nnzU357DcyOOrxEu7ilutu
Wau7LbdrD5SLQBp9+06+WkE1RS0f0BjF3zvVkbc6eRFhHdHzsgcBFoumdYGojgq1
hKHl+41jXFmMjnXYwnUuee8nNBYVZ9/ivhuZBnIoaJjVe+vP4pMlYpZjuPTXiqK+
dhNgosAZkxY0gg6f/Ev0U7BVFItm+Dw6NA484SHqS5YhSM6i2qe7vNsiJRYIhYh/
tzF5QmZUECWPWVzKtot9XZflbAgHf3SFcSM938CCUbAhb7x5c8MdZsRz8sYqOgYT
aLAjH4d4EsDBusJ7ezl9Cjx0aA1meL1XW2nvYf44x0JHptSDezTr/5sIDJU7R+V5
nr7MtrBpzOhT80Ho66CKCnXwiWRptI9ijmkdi/1OLACJ9lvW+N34rxWqWQxMUr/c
i1r+6PSg4KRGy+7Tf24LYlutCDqJCIT/fAP2gGH3Gch5OydvQX9tdfMMhVxTooBT
DBez77SUMCAIoH0kQLzp7SLTV/WT8Kvj+GY2a89og48QCur8s74jmZwl2wZ7UMA3
BysRNVknBDotyfZGOhNqaRfh+tujXvmzZjt7l9z2fEr7L5/5KrSP3Qn1kREuLv5X
Il+Bs150zjsQrSK07leQG87MMCbAkBXNEJhIlhp9WV4vOr6Eo+fV4gsHd3fx69dW
H3MT7ZzfLAdqXxdntUnri3ooXvt9i7E3wLPMY1MILXpzg3ObfGdhfBdX0evMUOwQ
i7SOnu/lbDjWlnB7T7fxD/Q1SA1REiUaO+xyn4nvpAShUasHLjK3gAyfi3CBXAqo
36xdmRYK0LiS9BOTFL3o9Jvo+9tFwUgD3ZbUHVHQzFXzwA9guZ7RCP0B8ioT2v2i
TATR67776fVwWwuXV5rfeErZ0xdXE2micNpLOQVWLKvvCh8BWchIKL3W9sw8zWxL
hTJ+CAajP3QYYi1hYlzZ+2tw0dWeapR8lX4cNVaqje7YQRd3Snurjy006OcBNPzE
apN3ePI0TG1I3ohyjOinjCS/+VCsJFpJ0unoffnSg78WCm7Ipf0K/tuuAgOSxk7h
72Ha8vm88Ef39Swz0S9RCJtQaFG32Wxkdg6w7sslPYfr7qTBMATiMfDHvndTfa7h
ey/A+hm5aJjuJFfHld75IGgwpxAiD0Yo8YG6K0WPsW/6l1+/vrufHib8OVEwU5Gn
ORVp3reNvOkoc48fiJdsYFWYtVheiKGVHQ3OTQ+S7xvr9XMvnXWXU67B2SFDDrvZ
beB1q0B4WVbGjhXIHGg1x3N2JRJ8W/3ba9OCjOEi91CWbscJH1eyaFjEAbTl83P9
uN39g4GhplJ0hg4aht5ziI5TM1fo90WrrhpCtfWMJDDh6PDeKdHQe4JZUwQ2FPJF
w3/WQsTZl2TMLDCGIQeqSyqZiczNDFQ+TuoGCeceqldTsO9bA1r8H4yrxD91217t
ifZCRhedogz1jJKCEThFYCd2hQehmBvxYTReOeOAEcaZgpsHXy3BKGxB2Hg5zPgG
wcNsYIOibdLvbJ8Neddg5GidvufgrYSXZyiQS2E9KAxnv2VUFhuILwK5EMS8A158
efvKuTSjkSguhj5gIhoUXF/gLIvaAt28Rk13UGjCRacYEpAlcHTZLUGpx1iOk0WP
cU6swaFO4CX6JXKa7mKXIdetYKVB3VGjeTQ1NuSMkwLf7WOklXI85iVdWhd6uE74
ukzWhyqiq1+v3wyUst5O6O3UA7FuUjPSB8QkXStCs0TiCT38H1ki74Xf9Ib3oln7
c3N6KwHPKKU7JdKY2bgyyPdElxqBJaoI2QISOZ02dit9Y5a/YEDopygmvmawRmJN
MtJMBPfdD9zIPVYQXaGVcU9TFgiOQntlkRAAzdIMrUrn7WqZXAzwD9+w4IZ6H4Pu
RP/Nvc82cDmXmC0WPmF7BIw5609gvDvmrigrVIsPwoVK84vQeYeQPa+/PrijG+Ie
O8GmfFvBZJgUtRBKVyDarPSMqxGdYJluWGVScdH7RVd5xR72/+NwndWLMuLLj0ll
kWEMPRgwXOFJ3RmZntBE701pJbsH0f5qmr3pWvYKUFnnxjeeC+Sp9FMVW5ACL1GV
TnDR4lru2baJ8dLQz/Yx2WGdFE9m3V+WT871kDnb95nKxwbJJoGrhgr8xHEB0QuF
x6ZjjCIuuy2Tyd8hSdeeD+a9e/vYligz2DpfpRMXF0Tdy6F7P0+rjAOMwUPKn1Ey
ApMbo4Wwlzto3nxLZjAGIrazoDhD1aADkuSIowXOeba96Aei+MhGQ61SgCKmebnt
F154ZZmiU36gRVs6D1Eds9mLJ3jCzpB+OY0m5urC94EaIEsykTchbgMZxOEXh+91
4j4xuCCiTBuMQ+fQyH9ZdhqO8n751t78Sf6i0jYHk8/s6SPTwEUXZJsy6InyunrI
+5ffKoN1qBGJDqflYwk0D6HeSZX9m4iSKmQasXPbCcOKklUuvNNKjLVe8FLd6yrT
u36HzHsDJc+Tqu8Dsc+VYJHUCxVbJ6LqKSLaXZ7N3NlgDJNaC0ZQ43NNs9huSokv
gw1A56ikJGEnM+rMPIHA7lEH/tMPgMDgD/d1E2OEkm2zayUmbVpcs+NkI3DaZBZK
jjFdNFFZyvoEKIVBoCD3NDRx0l00MBjyCaSHqEm/iPMAkO8y/ApESDPLGeKZnvVp
t29V01/r0SHAk6FDf5MsK2iVuFT9LCblQzeAL5boRUWRTEP/AWI5LTJwOjDLKFY2
iz7OxuYFH47Mqa134pJdurpcuZGthKkI8+f0puItXu3I/phOYjaAABe9mMAwMTe2
v+Oyj0bQSEPyHLj2UnGRUK1jkHM0y6xsp00R1Jw70GEKD7kEMA2RCZll9Rp5FZS+
4IqehBCrYQEP3og9v0BKi0dn4UZPPsrOyO1N+tWwWC6BJJl7txDr9kDeG0BB9Px+
FVZke+jCS5Ah8OtpHSONPB9qUq+rav3GTGJNRNr3fLdfzHXBT4q/xoemzNV4F93S
6b1vwMMsU0ao/L/EdQcxtyHSKcF+7Z3PaaEQspVIk0ShDpYFeB0qPGmHTesdRt0j
byoRDnTN8WAM6VurNE1U0g1NuxD0e0H6G3pgitfxAdcFmm26lKdY1Btm9CnhPEjv
sROTz+XUo+ZxFvobJM8CWz9uM5VrPYHyF2xW8THeuSml2ph3iPq1T4jPZKGufJz/
KyEso4M7TB8ndqJ/5rDQRP448fIc3znxsXPhm0uw1fI+d6KtXBjqDXSke8F6px7F
1zMXWAEw5DmiBRQoNyizsYKHsM8iDfFdX7jPq8EshakFXLEtQI19AI8UPbA9hH76
4faA4/+U24JlbbxnldwfV0/3QFzjTcqLFAI2CKm66L2Y4LKPUWj4nSAq5Fqag3X3
5/zP+H8xnctHoofSb/PCR1a3rV66CnT6pkfErzlWhk9F2hEsSFiLtcyfjJG9ZHc2
sft6z/uyUSfLbDNaJomHJDtMe+y6qbzYf0QEkXcA4RawEZOSDyh8NwIMf6rWYgyy
ZXkY7f8y7FwCEKjYuSlZZpcgSgNpWK3hNou/Q7sYEqH/FA08RLmXmqaG4ttXq6Nw
Ik2Feo+Yo4zmJ6uXmammUByaw9ItwggUbdv1CJueAv+/j3mqu1FEcFRTBuV2HHjG
I6URvn1RFcy3hW+0W5qD9RVDuFAlfxufInu+r44MQtzDZIXH7A8fup4OlMtx7zQ1
vR8nLB7lLlD3qsUG9Yf5/Nabg/gFeLJ+sScTnWtgmnW23Ai3GSZxBFRM0x+KaM40
3Y4GRXxSzkBUwsaPQ4UoE48lUUs5VVLEIBW+MnmKoBZcImHh6pNCe2WzcBU8yeJ6
Cjf/EbMWMf/9A8k1BJdeGVu/UXV8bW52ciH6owEJoygWIOyTQxIzniK60uV56Dae
r6QdYNroa1pNwEcK7A6DqfkMf4E++y8M0V2bzHMyKPCAfdh1pDLdb5mJc7ovMr7K
aS7zT+FLpNZrBopUv+J5W2fqYf6N7xQMCIqbKXI6Pe4lF9i/EB/t5T33jXwTTyyP
zV56a59tjssppiFem4Tj5iWE1fDG2fOEM0qDYQN49wjReBCNwRuOyQBPNe/4r91c
v0uY9XCOQUrHPemAGlmkD5ZIqAzygoJLXmN5xXrwSQv0m6AHPBTMN4inpkqynrPK
AMvYolknqMp4KRZl1dFLqrPfCE12xWexBLERyONBdbxtEfX6EjXZnThpfGpJNG9g
VdgsJVcWC5ygIYbhjnbo1kNkk1WA70b/TgZcpUlCgbD6dDpDqqXNaExiEhprBNvJ
3SlqHwZhIKr/+8IhQ7ltNatqrQj9RyYPywkAVuhxXEKcbj4ymipzQUGYTYuFHI1E
4NOIOjj2tIFc2FxvFu2aAy/iUJ1ZAdYQ/lwv2tdCO6wuRCwYCT3r01fQT+pucD5y
cpkn3GIRWx0iLyBlxiga1w3GeuYdDDAEehI6lHb8W0S1IdkVxclGmq/eLNFm+zUU
pzExr7yyZahz0FERhJGKv1itIF+nRJkELcVg69JX2F5WviKTc2afWjpeOIGyvZcX
SJ+61vpQX5Lr3FfQpysiM8e7vQaNAT/6yY/s/RvMq5fvBBj+HM0b+gYNWZ8Ri5wY
/vcRxzqRKkz35tjuVJ54pLdzHx/jXGKeUM0AOKeDKOEmW+Guo5fTXe9sBeXVCJ6g
fRkajCC+2j/lUGJ/FiZCjreQ7a+pDaYURK1qGdYBUEj1lpiFa1ReXdxj0UaY9fPW
MxAiEfkeDDSCG6ZJdCAW4Q37cJSiTa+Mq2IAMblxPVthyaV1oFxX+pMka1SxMXGt
wn/OWzz2YF1QyHQVmmiZD9mIp34IAtMKiYmgNtqlm3617nj7vU0t9f0cg3sbca5w
vEUribJ0JuRAtZj9NoHMPmNrdEh8gv2XzVpHD/2nn28t9juEolUeUfA8kmzbHJkK
f3rwsn3zOR+PE5dSymyzftLU8McULiQ8bZSbD1uUrOGCNfEz6OFK2K6RLIIjEimC
INLBWhBaMSLgX++TaRT9yoqvqahyhVK5v3oio/OYDktT7ooxykrVnvGTtWj0zOpX
lzSTJdLBmeN6tSI9DjLwW2AmkP2ckcp/tMdv3T/b5qGCPhRic92Jy6sxHrXfU+Dc
+xxeHaekUKMwO77vKwEPfYfh4305SrBp+aNbXZc2gB8ZKZ0eqC+eNXsnzBv/+tmR
iPDl9498fmtuJaIPb1IQ3CGAd0o9M2DE3/OYZm3NjgidLw4+vLzag9OierPNcjzj
wE8LGUW2cdzKLo9+wlXgW2nUihMWhQVJALyw8aDFF5mfcAEIRWVrLpHPbeUwXuzW
FDdMxQhjUKTe7W/d1q7f5G7jzY5p2T7ilhu2iAqecjYQEbSsxTMGUbx5s1IxzeKv
SRArPvMwjahbcbsM7vFFPQimShEUphONE1qcsKAo8i4HVgcB5DdWn9VPQDc1yLG9
hHy32cewgMGTtdCZlSRJ7mdhpswY5rTa4HVjEXuPm2dDJWTHFlX5UmkwpI33jzGa
T/xbZir8JRuj+JUsu5zYsJvJCZxXs87fiuAyka1L1WrsD2WH1lQwNBaFpMEM+IfD
xVZ62V+3+akcKmJmV5z03UV0g5Gd1urJE/Ou+h221dP7zq+j+N1YWkf20g5Uasou
BXfs1QWZoKL5iqMuTPGEDZm54ODIjUNvgfKQu1t/lnhxKRJnphsMz3L4kd7uy5zA
ipJ/joFaiQq4R/SuCUCYvk9+wbPOCUgGWuwTbs/4lnQAef5RJfPHCFzxGU/Ncinf
qBv3qvjAQbm5IwfjP7LsOb1++D2HaSMtosX+iWPDwVg2zXs4Fo9WfAR2mFVfGOgJ
g8KKkQXTQduwGzx5oN+ESAM2XEFZkzTmOgLae3NBpC9dCdfcRbrqcus2WJxOmG14
t46bgpy0X+ChqIciG4ahCQ==
`protect end_protected
