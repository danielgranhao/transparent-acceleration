-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
EQhb6YHL6pW1T8TTnxNBg5sZzfhN1RTuR/l5ggTqFYsPiqEr16cIBIgUE0GpLkme
quLoghFghzm8hUD0mUB0lvkQOH8+q40vv1Uqh0Fx9JTDVgCLaNNncyWfBVLuKRs8
wEUcgKXw66C1TrAR9D5vIYZhTzQvoioUn42d7BioBYc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 49769)

`protect DATA_BLOCK
Y+Sj8RyITYkwWxZ4kRi2bJY3VmHKEZigH81fhE2kBRG7P4D2HX7WsmEMB7peDqAK
IyysNy1p3aH6djTMa0W6HGtnm+r1cDdsDOh3ajX17yva1qajcSx8TJ6vPlRuKsSa
e5Zdi7LPlMO5eu2DJXHk8nD10ZGec7adAYnud/Ph6sIkrma5RfjcmkqSdLHHamya
2BxQhxJukQlmeD6CFME+T8u/16Gz2KZiK7J1vP7x6g1raEe8xZ9Me3oQ9cDPWWaG
B+lPEYKVzH1cHp2H9YGq6ULOPvW88VOTzMonNcB4kbdRQpfCC5/sa3XqAlgoycPg
PaNYvPSXUpAnoEIf36NttvLIYXMV2DRx9ESpYPTNN95HKbtyGMQcAsBrmMfbgn5E
YQqeQGqAruPuPT1kxwHtbVP1yWhBgwFVZVXGgtyvDQtI5m44SKrv7OHx77CnMMPe
E5OU5X249I6McP09Yb4QiJ+HJwRUs2fHqAChd8u2YZlU2EgVlNL+6Q8IOqmG8Zdv
A1FKfZoO9WLUJCRGecy5GcV9x9uP4RvPYwL0aOb34lfCZGMo0mbFYNu+3CYCkfHf
2uoe1lZ+w+bwDq4eunphtJFyrV7pwS+xjjbLtFo1ONTv8XPzFh4Q1rFu5PG0ocYN
PW7RRZFhchAT1OD3oks+YiUai+fQi7ZpZjas6ps83MbMuIR774BaCGZZ5p6IqmDW
wFqHMb8VK5UBNjyGactvvfx0rxpavgTo3U8zmedQbrcMBMVmNOpn7mRUaYr/duYy
x1CBXfpwvPRY7ZwuL97/O4H1NnRJt8YUMXHK0LPavO8698LYHjJA1VodskQAiher
0QR3EOwuOGSGOrONBNxAnzA10BRuc9WgfYr4yAcNQE0ZoonZa9jwXgIr1J8Nvvd2
O/s8KiqU9+JaQZMto1jzrs1YueJSt6MlSdCSDYv4NsiDiNr4O70glktFUPZoEIdj
nPQp/x8chH6hJUXSRNslBX9XHQzOkoU9cAOrDeFmSRYzVIwJYUj51EDcHij8tbks
9jVM0BSNtk63aXK/Via187urcK/5VU61gZnppi+CXFZLwsM2bGoLt9xlTwbJZa3I
AWj8Lqyfp+uO/n4Cp1S64/UEFyaedCyL3LGSQZLnLVHMZCO4Gu55MNco4YSlx7as
kW8xCm6fIt2HlTQHyEU1+6AdS1TAjIoy1MmSDMF348LZqpIay1E23ZcuGHjwx/bp
42UOvRm5SOi7UGHxSZT5kGNeOeKJf1QrCM3CsReMVUR1L8SPJEGKhhtHOYOjoS8m
4WMHjvNSS2L8ZbMj+zwbOcEZJQVmRfPH72JzlQlFeg1dtEqQ+Cjge6tGGLQqJLhB
RGijqCsDC0pKGGQfRfRxN9YwGwMe6NLnCZPBQ9J9FyBBe5HoJl68mF46N8KqibZA
GqlzDf5EvwE1646oubgGx4IqjoT2wBNWHu0Fhg2GUklkjEDKSn/iujD+zbDgV5s7
iqnWP6+YgABqDeftqY/texpajhMiLaPMVuR67cTJ1eb6uM2csPjAoFVH21ieZwqC
ho2WF5Pom/jYrdB/fjYr+ftwOBpfi7ygO1KwvCTnlKFElQLPsNgGLUETll8esnq8
T5FjBQItBjNshMDep6GQFgvLmhjkNQILHL8RBn5zQACdKmj1imrumtKt5P9xDda4
f61foLPkyNrwXVNaQmL9/9LqtYttUyUzT+QlwfaFGxZlzHYQS8eCSGz5GKHaLYQV
UrG+L+OvoPyMNOH9GX9zMlwhHpQBv5RnxaR/UyI8Uv2+gslcie7ozXhB30JwSGb7
DM3Q/2LsGEMCrqak6AwESuiF0dwtVRfMoVRRxS08Gw4yvAxP7brI+ueiuyVWMYxd
yajeHdeENQ69A5f+b1qktxR2At7sJagRxcW5YE59tYB49uji6hybZL3NrwR1GcAr
bO7F3KhFOpNne6HG0rV8YVkjKa07OuFzi5m3m9CZEGgMJKBZ4o6aZS0vRed/hccY
cc/6NMiMuGze3dyAYdsDUw9BIbvLfACBAWNL6+PLx5nwtwq7rQRdfJHihhqjispQ
LN546Fxv7m4fAn38Use5cESQU1/bZsjex2N/OgwGfLslLbo77BkeYs76hapWs36j
9lnVYtxzV8OaP3MQYOFvcmCqsBvhnTldQ04PPCyVhHa0gXI+tO5QPb7c4VbqZEMN
Y55fMWdoXC1meGs61Z3YntVe538UgwoGw6CWAbviMxyMrJDCakeoySsEOS+t1S4O
iNLSDRghDi4KtlknAYMEujv0ewtsV1+u8l8IdZuu2hfJso0zW6kwyk1VWucesdqH
By1RX14hO7Dism6n3f7/sI6ZGVcVHw7/qv/WpFIMOH4+boYovgAxg+KbJVlgzMB+
g2iq7YZ5veDduRVLjTxNDBpulhmxa5WIvEWG/1Qdanr8FO6eXKU+nBvlvMtGBYfs
8k3SDgoWUoBTP60tELwEilSaP9xgbOjqy2SeC1/IE9QlZMiROV0W67KNit7tvl24
cy/Tk73bnPY/0CGco3YnZx7muobhcmSUipgteXygzWQ4mGpR/2cE6IQDo0jKwmHR
hkRxYql1e1SsJE6Cp/3hNrWAsMhhO2ZFG0/5uNI+1J3YYJl8Ybb8Y1fba/FsQX9F
RaYMid8rqzndtC7hzlF6rLMJ/w5EHXNYPogtR/FkATxarO4EB6QaZ+i7+GcGNxIU
WL+OLpIWF2UjK260OrQEH6d74B1IATTi4zS2PjnrckFas3k7GGoW1xQBDF4epuik
XtT6WhN4sqrp1bT+mK3vyy4DK67gKWmSNhQfWjhCyNP1diXldbMY/Um84DzNuA2B
tkjLkNv2NAmLktOmRKP2CCtIHMjcn67AwSMOQ5xDx7RDZ2RLl7bM7m8D1+ukxZhZ
H7p+VAzS4xJIhB/T1E8ESxaxqA+1N1SnF2g/sA93cGoCRYVbct6+XVTqyKwp7fFl
X/oJAxiOeDwkQPC4rI0B3cT+EiLPfRcUkf8n4xGICaF8MY9nA1ueHglCm8QKCWmG
wRkckshyIETd4jCWFbvKWxs2DoZOreVjpO1KLTr5AOTMBfsqcrIDISQ2HH3J9RlC
BzoFHtO1DRfmpAc4ZTT87GF+srjQjkVm4WczJCUPS+gegoOqfJMBftdF9QlrFM9F
0UpRP+LxNW4IkA1A538J2yv9pEw9ssgG7OriNXABRuqI3nYSCGaTHIcVIdWclLUx
H1iiVpJ+ex2FRINngnx+NBwY89umOI6kfxyrPAD6v8sHjcjnYHcIuL9C33FZR5MM
hooMPChZwqgve/ZhG4N1Vp0gQW9X/1NnkuOazFJ5UA6/6+ZNAzb5ON+dyLuCuIF1
K2L1G5ZATUsm1YehUfCJj2NZpcC+xG95jzjY1iyWse9RBl6qeAELbzzd62DFlcfU
eIvUHsFeLSMmA7c8azjqVC4D1zvYgugSYbahYDJFDC9QguV6ci86ivzPkChEGDNx
I8d9l5JWyhbOFQc54xrRgofcJsmTtM1/A0yYAhaoFC+lYSBFas4jvdmXS7Lg9bP1
E6T5K6sjyAq6jXtxOk/MdeEAZjYzncEZiDoA284/QE1FjLiu8wE4hLBKOYNPZEAb
p4hdpNhK3IOt27QuHkMOAyNKTs+JMX1Whbrb0ng4KkyYzMdvn9u44dk/KHwVKwav
9J+3M/+sVgthcvhjN13njGWbXL63KfCOkncGlFraPzIYx4pqp5dl2NdWu34wbrU5
v62zw2YShBbkJOjw3/wc5hCQNhduq0gYFTzz4IMf/9DanJggqcGPnFEvFbhLzQ+8
pafD/TEfLMEODW4frhuKqWdV+FnxoAlmWgIflw1vzDRlaJz7RTl9jX9S5y1rj866
H//LJBGg0vqDqcmNMu9QD74AJ7ZbTkpW1Iw7jauVwGtX2+39Z+xL5vxm5Q6+6EVr
fBXEgWW2baf69SGwOqZf7Ti2Ronv7GstAtbhQKyYWlmUulDOGPZKn13xlZQTIhpA
wnQLKPX44CakWAUq7S3oCBOihAW5VGfzjZ9IQDfuEiW/K/vhrTEA5/yWvHPO/8uP
mku5bvFrdztX1UNY+40QwS5Qe7lJveyC2d/O9w+/mOhZzphRb17V5SMAzpDneJ7B
3E+sfXLuQJreHkkmbeYeYhEGb+s0qo01AwvAXC6gUerUqCjF26CNtF0srYcZ6srT
pPiS8LtsFJdDJdKUA4F4Omao+tTPdXVMY1QKoeeS/pBjn5BtvIKrhvg6g68lqBVJ
MJjPCFE/yCgPacUoN888cvU8qUS0Xx36+cbZPz0G7K1rMd4gChxOhEe8cJLUeylT
KCfnlxUXHdmKFH2D+IjYZiLNQNb4IIJRIpRyG7xqfFs8IfClj4OLopJIoFpVIeeQ
0O5PqqZ2PgDXKtQPQ2+ZSXCwYDWg8G7CAfAp1+Y/Y7mg0kEnrvFs7BDNA47DZHkk
hrPyEp9z7jJiBsxeVdjN+Nn1TIT6oQShmO1d5kRRwhH7tQmgKXWa1ABYgygpIgN3
clI6aw3UOTappfDu9jbIHTNcBpEilDFhESPl6+lEik+MFG512d6mV11+623JmHhX
8lV8FfyadJdT5WprtFsEAO1BfVFNBdW3t7Isiu5XJhko7X+IDuC4tuu6VZv5dVB4
fsCiXts1O+mjX+MCEFBLcHZva4U+x6Nz/U/nBjVLN76XXsPyRuPZjfr5ZkNw1LcT
37FxzRpvp/LIOk7RmwF8QPRjVyFgwCVa5X7Lfai2GdMwIWJXu6kKMNOL9y5FokxZ
lpFmZnDo2x7x5q6XwMS4FUe/FUriC55wOpwzrIffWlYc+hLZFnGMskCAhq6sRAXT
5OuD1Oj32AEj0UMVpT1NVpuawLaE7OvLuRc97pthLYbc3/zSveyikvFoIegOjFbN
xbq/Y0mOV/gM+BpPyniTON6d0eg0Utqbz4SBv0hnxw6yh8Ag3yDLEXBLPplQDYg3
1b2BML2CrM2yqfHQcD8xczExhRzAp0nVgOLhnFp6EZgJVz1X/1OiBxahXhrv2g9z
hmKcCpxmE7x7tAGKdsnO8D5cLd1mKHvxSV3ICN1ZTgtUN6NNhf+4Z+CL4BzySck2
c6lUckxwMzZ3gSnLj2VVPb6laFB8R9m99oepx2fmomhSf4xqGI5VGZfCaSOJxi6x
dZjTNjupfqU6/8ZiXboVoToyD6uB+Gy2saMsierFjbOa1J5Yu84vf66s8VBDddUT
Lppby9FQsGsHkTWQK4VASekLqqv/LjYGYQJ3G4x4Tn74nzm1/woNj6z9VCchxu+4
tmzPQu4p5eTDxmS18ixQfxC7rFKdl0+w0wT+Qj4fKTAYZw3waAMBu+JNqW5kxcCy
hkRFbkoFquGoBz4qxadVvfEXIcv4F1ourhuxzADRu3eslcKGeHXLukyyYjBVALBQ
6TeNNWu5Ahef0ddHG4BcacEYbVJKcJy5jHTVTLOYSLlKwWXMUy/BRL1vBp/136hM
xxh9PhA5aQtiAMCIUMPpRzSbA3hlmSY8yEU1yzuRuE2i72Dse25KT0BIwDzk8phL
szQYuMDsHW0bCoj1HUXY2SBc5FgkVVLEDA1rv/tDPg/P9DRstAMW2xWAErOAstga
C5iMBj9vmwHqf1rvvzK2QM06Dl1L36HN4OcpiXj9VAqTCeRanbJ+XuWHTvveirIA
ymcGzqlkijH9T9iJxYQsUlF7rUhYadYznv/vHPfRvZtuod9hQZfqPlPpOJVBhQIi
ro1UsPoL/fFWy1uVx1kMQwAO9qJyq4ZU4tfhEA5oSvysWiuQyV4Vc3cvgxKWOCQ0
X3UMwHHr1Lac4oiIZ1nFgWVuKdRbKjkO0V5oH08mx0QkQ/vrK4l601BSE7nfIejN
oIxs5BjfHIiojxJpy+4vMTeGGV00GZGqG7XVTR5te+xj4gcdjol4kY5NV9QHb2rH
SIUEyA26xkcFAZhU9oi+Jz9gOgN8BxO8I6FCYvJHSNPPSmfsn23hiL43MIHGd3VF
N6xhlx12xGqmGaoO0qo1pigKTR7YwaEU1hlYXdkItDwS9IchIr1Y+fSsa3SZLL5O
NXq572FyNY/iZfYd8ufu2AaHXgVTBL8sw+5tPB7GeQw8Ty6a3hAZvXlS/Wv9YtoH
+Atay/wqBUmGS765g2271e2SHYjrI7hmnRkOa60OetGGwLjprSAoMUq+++AMW+7V
UvIMrON96rGNuUS6HOA0Yj6+2pMrdlX2JN4469TMSDVwA/BgP9GMj+M3Zm4xUrwK
ZyZKd6SohDCyJfrg1TX1+OQgVu2s5Yxm17TAgCfLVVKnAFl2NVBbhCtKRm0jfzoq
wV01+sOwHMkqgagCZyPfQs5EPKj5XeU2XHYTVYscNGkBUrop41ccNDnpFAL9xa9G
b3V70Q7CKKRVIO+oPYXOlJZ39ewo5PvRbTnEOlCPpvFBcfyldQKH+OPyRKg9gx0x
dxveLtjruJXSsCTZm/e+U/fyLCIJeSMJz6dpP0zzFgWbez6D3YbqhD+dsAaGEV9H
zGpU1iWqacIrsnW6szWcFos6WLxdLFnN0Yyib5ZkaAf8nfP4ne17jExDsqIsng4k
NQDhpWjJ4C3e48HSYWINiScT9coEZXa+oxlQG0NR2QXfR3npwsNa+/Qj+OKqt3BM
ED0e9HKIimWSGJBAlittTuJX+d8lWkmNlodyR2EEQvGbIcV5eGwpLzIKOX2rrQ0o
Tmb380zVoYgjvF1r4elz4Jr02EwFT7TY71DOJ3Eymhux6mZ5eCBVe129dP9faGff
KUUJAz8dNVfW7HhZiIzksARBF6ejczpGY5qBLgAT4k0poYc2chJNsUyK0cI/mS8H
063lkTD7464UEl4S/JEQXYO4TrXj88JP073ykFBNo35ubzecP6Q0OV/1yUl1biFG
Gf3xwNXGbJhLIpndzXJdQ6GP7QZdOhvy2H/Da+6ebbZOVBqa0v6V/KEt/CluflNr
Aloxj4a5h/GZPEXvI/Yp378r2OrBXEz+1zKQxSyG8aM93aSCvW2sEb8WnSABlA2a
x4QaD08Kqj0G2J/XTl3yDHWijNkk52p2krQOYNpceujl5VGvPKR3NF8dwsYrqFcO
jPXIHf5Vj+qC+U423k2bxxA1ojSslKtzryF3fDPa7Ip3BbSF63NRpyDSs/g3CJdD
8fwaeMvxruyn26lCLOsDqO/5FF8O1HMv3o11A1+G4dWQDnKcWO8vBGEj7T+lDoYc
xYDATpacmjy8AwKpHjZfmGSt4T6PB+2YrC7cYnaddpI/GPmJsr9sPboEDRVHt0VX
r5+bV5zaKloyW45zRfU3d9p+hiZ4+uEPYBNXWzvq+k8u4zAXZhly3rk9NuJXO8yO
CuTAtrq4sazuQHVSnqRhExIIh+P08C8H79FK5AYqUsTTE/3BfcsttCUd3vG699c7
BY+P1ImXdaisNMEMrrQb6zmzPgsoVke6vhVNYVBY9bywg6Wwe6N8wcvPQ2wJifyU
8TrzxzNGTPezDGZA0o7TeAW26/QhAmMnARF++QhDKyNlduTLiu9Y+RIn95Ktjj/J
HD7ka3Qg6Qr1nDw2iyqIM+5rBZJ5Y5l+U/lipothIV23NTPxp3S5TyaAZDBUoQX7
dDxHxRMl5krq4Y4n+NEyBsYUds89Zk6b5mbNhnfL2MAy1El/qd6pQl/QB4vcrO3f
++68pNtR+kyjucJG/L7jM7dj3eb7bqjRY7Y2ffXAiOOGzChmAt4bASG6oi340S6d
DbCG3LeyJuHwS+QluPv9Z7NhkqGvp95slcm44n00CkpLnoPtChObzNK5Q1l7s0C9
u6n3epyELA0VycEy7P0ifJADr0+VhM9Ic0j+FAnGg8G3qm3VKq7Nw48ja2rAt3yV
mTuIkBlL/HWGmhC+XSVOcc/suv9S+eUl9dJD7wqKeN2LYf7VTej8wvfqG4XT6vq9
s423VSM2SiytmMYAs5j6shqGk6/YVTk0ZJBhPCAI4ISUV2N8YSKo4WB+sumUIIxw
d3TtpexFoTA4rnWHoGAw3NYujCC6iWMJ67HGsDYMdCZOkck4+/wkhBq56FWvWgOF
vzMj7ju5TI/K3Enb1w+e4kL4oLqFtKLIwEZTO6Zxp+VTvTGWVatpAVeIk6K0kINC
sUy/MNbRPgg72t5yfIN0N+ra5dNx1kjCmQFVtXR4+FYOk8ZexiFWJoc91rC+vPx5
plY0a0iFh7iHZ8XygxHsx3X+DLnmjyoqR0WKOACykQgnZZkUktFtVtQ4h+t3JvNR
XybZuZDL1zG7IUgOdQIbpWih9gZmFD8d/39vCqWg7IF3fCFyWi5ztwtCaZpKgfQH
MsPWmrifbsnZsBCPnBHL8MSOICVlMl6PyP89Eyb8Oj8HyplNJ0/6o2WHnA6Z2upc
ijH58uB463zez67jskpbCo2zMiCONGjfPAS18bvIfbvh5xDNictO35khjOqImyQA
uGfjhFKDvtJHmgPfHDf0cqr4Derp0VU4+v8+AKbMnFuqVIO/u1OFlCLMDV4z2hY9
xFmz2zOpv9N+eoyqJNlJqKQQOuLBp3HBHDsYMDxzIg8M5JcJVZsuJsi7VAkfyT/H
N3IEoMspkrAceI3MgvVE3D6d27i/wD9UreZgFIKKQLZPVO2G5d3zi9ikuQIvi33h
67b8LX1GZ2XP2JVl1JHDwl/sPTwgL846VsGDLSG6PcHGGkBp2Rc2Clv0HEr3l0Kd
IpTSViQCJ56WOB1KU1KAnaMamc3pjIhRcB5MhCHuWYkb8Nmp52wKLuozYjMCQpQl
EadLpKrkNkMiI/COUbr3CLpBywdfdYqGvu/TtWHEWjwOZOTrofX1VmORJsCX2Jwc
47WBn1b/p8sagVasvtO266g4S03kzhCriHUFUdWb/QDjn4UgZS39D6tzRN3ZOGsY
04x7/Ikt1IfhJFV+dY5UGwoAUrsPyKo3mrExAToy+XKceGWo1hODFHBwlLBS0u6/
U9Si5JHPbtBz1tLg0diCZrJ0Wv3OsP1k5cJSpA0slfykWxEsWiPV+nXqqDy3Tr4K
eU6bboQgHVXZYYKGwRKnEwTFs2jykBd8iIeuUazaaIovVUgAveCkyh2L4zRlFKKO
VAvPeD2Fl78BnGeLRpWaXqcIuONjZYYPHWG6gV8KCbCoi0hTmGazcPKDkRE477jH
8R8Su1AgUYfFf6yyDFvDWjZJU4Ijt9NWAsH4Xwlu+wzfb9xJgnjsXub1FLVeR2TK
0XXh2GY4AQnJFPT448z9U5TgQH1wKs9Q9ip762sJTOGXvBTnThu5kbUu5nkvd5sB
UVXE9SVPeotnSkdgJ8ObKv3qMnox/B8PXKcAvZvOH6qicRPxoZoCQodUvpTUqGkk
SEIQOMVHuDEFF8uDyku6QVYmfxwJDTQsFLVxOgXyvwrm/dniUj1vKZQooWVilDHI
FwyyhV/2ix9HBov5+fA986rSIgDWOamEOPB1HfcNqdQPRMfoMuM1qVzJ0UyTMGzu
wj5sWScC1DECOFaxFkhffyNMyE4AJxUTJ+419sED2LBVbFADTYFo0gwcdCB77Ns8
09Juh14aI4kvpYj83/jPCsO3cTUll+yeaZo9M1sVfGrfzUyq04RFGHMy3WtmlM2k
zUMI2Uq6NvM0ZbKLztEv3R+l1bpqWBW1yNvn6hOIbQNhLoPvKEnPxStQ4X92XkFg
lcMy3WxZzmF08vPJtT3dUMIAjYW4f+txr56+HgjFcFIDTUXsSEaY0tt6ckBa3Ytj
fg3W59K14/IlYdr1L7DPgixqXuaZpyBeAAzdZjElDmayBteOkRQdWZlqHvZw0DUp
bYRG+WXaqKJRR14pYFYydb76wutQHtcjLsVlgoya+EqAlDRWLWJmPS+ADx7SHCxe
ajM82y13Pk8hyzwHM83944EsAL93VjyuoLU/oaO2y2P3mOKMQGX3EYD0jSjPN1qn
ZEqv6VfEuCVu/THzMOsNi2vWhTomSuNcEAHo6kre3KvZCSdRnemvlPRa5jYR5Wmf
CbB61yEejEFVvZJoVezK/6gu3J9GztsBwwPO3oUvhKlmemm31aqPLomJBdTuAfrq
o6dNwYOtjF6idy7LfH60uY1XOyhfNFoTACHQjE7cSuRDEIy6Sx9ywLBnmCv+PLYG
vcLvYwFeOo23rPfj8UlVMMIr+I0JjYiQmCRVehysQAl6WlfqJKG3hmJNy1qizzq7
X0OdJMZ0EN4LD0SBmYGvbSUI/NElIOh+D23yRxh6TLfN91y2Hbd0iZx+i+pQ5Vrr
AaOp07hXOMsZ9djUTKd497x8rolm935bskGQxtpe5q2fAo8WniC8i1GJqpuLFmXR
j+q7O1TAeME5Zrm1LQgox2ONiBFl2ZtZ3KTtbDpJ9D9JanFuj5FuuXGieY2sEc/y
z3i35Y1XNc9q1hZIevtN5EqOiqW12dkKrpnohCLcveAK+nw7GdlDYRIxj1bb5bu9
gpcLTOXO9NoMvBf4V2gFMU/k+wV9A4J4gpps+XxV/luJaYBCQ+rRAnoY0YO3rRGr
wE4TuX6lkYoisKtDDCE7krfei2K5wFPKWNsFWTjbH0Mf+cDYYcRwUz+rnbee/Y00
4zz8adHZyPu4Mkh4J5SbI6A5RLxOmrDWw9FZ4d+fH/SaG6MWc30GG0gTqlKl9O9D
suMJFW7gdTKHn5wQKmPDIYHS3OaRzYPhJBUWKxN7/QKsd2IxPmC4ZuiIAgR75yo4
z3c/YoBvZRTH3Ma6hXKv5LCxx65PRFVM//vjuuhWxalKkPltFhvFjm84HLPjWMvc
IQnN8GHXIKAvIfWskf9IYOG7BMghRhZk4I5sAYlnrcb1bLhfe7w7BkUJxFr1e0yl
cxVOkvN2UD1O40uygGkyDCS7/krzldvltKBHvZnM4TsA8VsAbmkT+eeXQvl4BcnO
Pesz7WdfhogpMAWyLmFMDhuBmjNfOCjURSl/Z765CRtunmWLdPy+ULW/7Wts5qjm
G3eKMlVrSCWzXZmGvAQMeh5dTLBM7VX3y30iiQS9mQbO9cw2lOxZdwNFPyXvoAnt
OjlpBoqR8XwSrjt69HP2aJrZrMLjxOrzjHJLAF/fq3fkJquDWnHWtf6QSS8l3Y/i
KeUsefuEytW4+FxJaVVfcvbS0RN/cz5ls8p4yw46+4geArGeSGe9sKZNpeBJPDxN
kuInrRR1By+rjKgTcqd3BWcTBYZGxFzEcmZAwvSL2M9I2DfFAXtiwE60ERnt1O68
8aN+JYobEB9PaD77ZcB0CB78ZFM6ah827QJGtwZCP/8GvSFCwUMbkiHNmFXK0ji4
8yNO4RO+qcciNaGaLXkhp39I9j65g7Akn/OiGaLYJyuAA4pwTfgHFdEIGT6pfVxD
B1wgOuGqCSFm8Z5S0Lz3BRBqDsaNVTM4n/5wIKBoqQNIqVl07rPr2Bk4aef1PZK6
ad6jZPEawFnYqHld1pdcyyTqC6s0IPWvSFVAo/0HS3zMBrtRTuxAbANELohRcAHO
55tHdMEWIg8cZMAoCpmn8KK56RCycMfamnpng+fBL1zU9qCYz01XIe4FD6QxhHQ1
eJpVOrh+1h5fGSaEQB+ay6VUTaXUXPbb6D4os+nHo4PHo9ZYXx+UEgNEiGzJzl8a
LnynCvx8aLenKXwGYj6gevPiCTapdXvOB7UX/uNmrAkZntQPRWyTAMTdeKH9FNv+
ik8SlKlUpR25oVuTY7ZUZDc75EWS+8ADNxIL/80iYNfhN8FO8XGDJ7iwTGKyUx8e
UCkCKH2V/YbQwKOh/j5h+inrM0fLLnqncl4QGtthEPnyCkATXg4W0HLza98CdjZH
M3jmReGgcnZJHnTZlOVX3RqlUjBmAOye/oY3jXpyYxTMo0i6ZehdHvq8V+nTiqGt
lqYdud/4claMcFgZGO1DcvA7y3iHHJl2wXhO2ieyuBx5TjPGFjYcsE9ybGR5yAhf
aufHBc/VYTDVzw5RbERR+QLTi4t6DCBlH5uEnwNIn91YpyaU2M3OKrAHjMQfqNtS
2jq7MUyXDdE+7e3v5wRHIhmHERsS/CoG2Y80TmLPTpG38u+0LCnDtmKMEuCaOP2c
N7e02Ni8RUPBcPS0J7puuSO6wf0z0wTcSet+bdnzX8OZKcC2ok8RUIsWlhOQ+t+j
j77J/GBadYSjNP2tpa87FW/Ws7LbQN2+r2Mzp+6FHyJoRTlAcV01toL+pB7lWiFL
i29pvDkwZrMf/3skYo68soq+h1gQq4Mj10ppa9TLaZ7fuusgJHRaqRmjCl6GoRIx
yf2aGniyPVy7KxSiREf471Bf6WVlrmugcJjDmQ3SKn0IvTSGVrCL2R+kOWkUr2H6
bVuy3tFNDwAgpEFK+AJJKRafLATxZ9BzDc09f5wKvwH4WNPjY7wvmLT+RIWSlJ4i
gHj0AvhpO9mcz9gHTRUUAESpBCghEqkbFqysqmcEnojIGXZypLPpkO0wEvg2wS/X
CWRqsb+TNP9ppeR/wPOXfke3cX8LkvbsiIUyqjS9rHNRYtpDzXODtxUIYZhH5Vpx
b5JarK9fokp/P9zdKIfHeZKJf3YlUiLm3VEBLvlm4li0dlDJ4WHPcdixJ+9z59Ao
bVrPJ8BwnYlodW2VSXnr9WceyqxzmTO2xLpXZjzA5a4aAlVKGH/B6GCh2EedIgCQ
dViNPaPfypYk4uz9B5Bzga8W09vP1JM/JAiBc+j/w26QgOt8exmftjGnJfYtk0rk
Q5ADXww/d9KtaxvDRMIpAvvX33CnfuA62eMaZkzCceuMTNfvLiSmv4sLZSShyLnJ
tQPFysrXSo/O52WzjabdN3RlgTMunGbx/+KUqqohQTW3ZQZrlNcXsYilDNf/l2Uy
pV8NORhvnkLuSpAcsiuKGvYebFsF/AXVEyRKVcqwyzG5urvg7RXCUwWHuAxUdXHN
IkQE6OgjYq/1TphKbB8DfBuxcADb6VOyDDbYNAusGZTsu4Bz6dkP2R65bUZ/M7Lv
9unOez9VwfMIbXSzVcLbIUBOfDQXH2SEmGsbLyvyAiJnWx4lLr4XgQcPz9RJzU6C
DrDk3fa2moBc8gJWbiDd9CjBaU1KCKYFriJVPiztuyrnx+RfK16j2LnmCq7+KzdA
nxwrPFd5PtfmbV9gEJkP4MBq2KbaCbbomQlfvyRwZFKfwp5zCEY4YpqX3RwfWGrz
ed9HKzMXCoUC1sHlk+jSCsbJC5hBuG4rekh7WAUUPyoVuF0mUWQGUJdRBxsLN9YW
QMePs1TT8A2HBdoSTns8Hq6un7KVOkhWs2QfojAq9RbYkaHR8kvfyJcnYR6uDbRX
XkwBWJizTh5fzf808qPbi2vQN535w6LgInmNTVX4SuSnMyReBcZR1OU8C/pOQafQ
kTw1gZjNllMuk/ZHq7fxBP6QsRWF5i7djBRlrWC+amFMmMqTwh8reCxtC29U/nSF
upku6JDLKP9WlHMcSIh/W5bi4UAtEvY72ydnYLXJjM1KczcYC2gAG+3BzNP5jnRp
AF/8omvhcQE7KmZysVRikd0kT+DGQFyDx6aR/+4qkfbwLp14GmhPAVfuWvCmTf3D
8JC6E9IcqTff4TX8e2iaBVcK6GvJQkND1rgLWUs4XI31Qb3tHVb0/E2mRCLQB7eQ
u1LcohI/aGS18A04g5cSCDDlHG/bGhtbbcDosH3Nziq+VP6zRnUzhFO5jUKxz/ON
AlDrB33eptLb0EqKayuOSyb6AgPmZ2QH0Yo/YZFREGux/F8zFdoCwRGoyfUceUU2
iFBr1Z+7R0ZkHMAM2ROFF0YLpQCGK2I+J/ok3MtoZvu3atY9PQ8fiMHG8R7VkRs0
xX/0XDQhstwgrahZI3zy2pupnVevH84DeuMz/RckwzsUD5C9haFahWxdTGVr1ctG
AAy3gd3QZX0HsgjI+AcEmEm9HxLb3nBYz2UKf8UDfoZF/HF7ythUuCK2HhlF44KL
ubxA2LuKF6ukIsmYifQaKa2e/UVQ/lcXsxiuYc2Cl6hTVUJowthjMtPsqZmFjQMi
6eQQH/kpgYTJNjhpfVB+9CQ0P5KT0gqB9E9+okabJ5htkUKmNR8w3JIBDXjHAPrZ
HkgZo2bgqq6fEszHjTKn11ieRnZC8a15ChkGyiUwPkyTCzFs0vBhmOlWLdSDP6g+
gCGwd0tC9nuamJoN7D/yCsl0d787fDerzUiLjmIY0+7gou+SEFkOX4ZSWHA0e88C
/zxufJLlG3ZLqzAJMSseSM3fp7fzHFCOgiKFxLLuoOP68evL8Cj2vvQN0WejeMq2
My/s1QspRInHpJWHlfieUY4YpL3hpwQm8YK1uZ2mi7ZeAt92V4APxz2paFwhKYsB
ptq/W/tSjzHd8EZo1bIc2pkhOTHhHkRYJG9UIqSV69wAp0aBHbXa13C0eHZIoKdl
foS/NtCj3rPRTupYHV2HOTwA+y4HxXTqHu+zEV8heefVImELX6Cae41DUbV9gC6v
OhIW+TajSZhCDoLOMVBK3uW2djv+IUibJm2azo6q0pfAoYySkjg7ZE+0OEncViOM
cZC1Cdt+NfqUmAQUvoTgQUeg4HNX275wimJ4F1lwhQ9tJ+ugk6eiXQdJmEnZ6YtT
TrDlyb1YETgJlvZtTVU993ldMHkyN9gG7xoRYvknC3hYT/1gyc2T37SPWro9t3D+
nzBl9bzZsIcwsgufduGVpSZntKW75ldl/NUY+pG5cXXfLbp22tHOQVBs7qJb3EyB
7dzit/2XY+7RN91uYxgbRK2yP8Fx1wZYRUNMsVOqhYd6LKJb/oD7C5w13KHiVrgI
oY4sk7h5arXND2VLUC/bNPY4oNG8UYtfphl/LIhVzUYWvFHlHm7vz6+P7Z7VoLqn
0oDb2s/yROkXAT25SCy471WdMl0ik4ZBhMMKQufK50eoZ/8QtxQtNeBzQwkP/NY6
XoZDsA1s/to0EwPC0i5ma8sgJCziEpW1/Y2c9i2Pg6ehF26HE7S2490lw+hOPUxN
oElSyMYELD/H/G1GnXmOJqYg3Hu4XuYuqwy8qeFlNigvETyu36Ovz/QqQCAQOT87
vk05WhyI1EXKnmKOxqOZP6ta4MRzlaBn2xKPPWOik+ATZRxNcqp3R+DpRwIfAdtC
wy4Fceo61vnRsdMYPI4G4B4jfmFmTS84/04lbllYjYIccf5D+l/eu5zxReLNwLSP
pCAXCclf3Vl5j9DHj9TSw9mzHJOEAWS3nFU2PQ3xF0jnyClD/Mx9at5MvhrpIHeI
cF72/aCcAEX1+E1KKZVLpWs44twNuOfMJhGUbHXgfd4bZRDN6AAmKWZxjjqnYLvt
Ycblpbybjl6HJBVaMiEx2B2+YQLephpeAtUNgSVGgojuHKk3U1XYMCSP7oHUiGae
getBzrxd6gHHwdZVuZygBQnyLu4V3LJkvfW1LD9yQ74kwUAE8G65AWTwecfaHBtd
aOdxp9T+v9U0UE6f49t3EpvDe52RGio9GBpgrHYYRCsT7auhTUzoza9hNvu5xs0a
nzhJaZRK+f40HD+1u+miDyk4hrytvTWEHe55EZqXQ2UBICxC4oX05mm88PkglySy
s9ILWT8Eb3Vg88f8p1rFzrw5Shs6knjQOB5jYxiLElPVkfDUbwVKn3IOVCUZAAD0
9JAQf6XytLrt0T9HxNigPa9heR+8coAeqIHR7hyvzDIEfgtmfxyMadgc7hVyTDST
GwiNTdZdS5GqmPdAbPFuGJ9Ts3c19/x52fmpQ6FZ5qSGz4jpkKIx90gcAjECTbYU
0Vz/1k/uvCRoKYo2pKKPfAZSEJgWlgcxqqjjJRbXjWm9LLn53xfAWohD52Mn2IWt
WZ9JfMOoOxEklXQXaZo+r3Wwy1UmPLK22OpOz+opJvkkdiBGdAemFeFVSXllfU7+
3v64twp2GhVPWyJWcsxUVqyasEHBCIxC0kyr6q7iBclA5rjSizqUaaDTYdl861fg
SYANYbcwVZmcVhazvxBJ7WcW9VhYjxI7qQPaHf/+m6TrWnd3BHmH+UmM9NwqZEsf
zC+cBmeplvZWkSKrc87oE8VoDz2KQuQGrVbXS9Qh5oCy1ozC9TFWfKCD8Sd6dsur
h0tinYdu8QL9Wt38rUzy4SgiCeqt1zqAxgSjfBuQE6GILXnqgAR9x2cp/GhYFol0
Xpltnyvs/wtRph6oEPzIp4kGaJD18xL83ydPNrXrqDRDsIvXV4334C3mP5nW2zDf
cgGwKyam4hKUehobTP6VB4ud9kSSo4gsxA4XwTZo/588EOVh5tMJ5MV/omAmWqtN
pxBHnCNPYJpwWtJJbw+l1yCW6axAaEfll+CPB6rgjcOVpIXThPZArhUrEHWd3zXo
RqVBvHqGP/4iRMrZp9m0Q5f5wYJfnliIwrOdTP+PZ9hn3G/Cw3OstbDYeWm/hXl5
geVQgrJ1oAQJHkm1XnzlwU41GXHHPysQ4A2rK+ne+ZSSbw7fFCh2ngp8Wf/u2j0L
daNhJ0SpboO+SGMuL984djpskskI/EwGEmzJ/kFvFh8CtrmFzEgqn7R/9Srm0sE8
DpjfYs05sl2TuiSaBNpm2HfLbT27mxyd7TKN9QUXtKFMq9SM5SBIOs//47v5LDzs
oohBaVpYVk3Ko3yolx5vGMzSzNTBgXDdkMf+BLxboYHw1axhsPVXZ4wrYYOUd70g
dJ/mszWF2glMnlNoZeg6U1ATgXKQPfFbTY8B+aJpUYjdox+fE9QBRdRiWINjoEwJ
lWyT5LSQo1B2mLvFEXFq8Tm6+5CCHzv6+SZGv2WN6MuGp9aOYVbmAtm/aQiRKt/i
+nWknP9PKiGrnK356yldVv0knTB1OP4RB+7w0/vNzQ+z1Q6qbVY7llHTxjNq3dID
BvbvXtQS/091afhfdufOWTmzv3c8+7Avjx6hbPOCNdi1HVtYxknNA95YQQBbugbR
Jf+K6OqsoipFOFQYvms2q3DDFyEUb3Yf5XK7i3S9N1ymct484G+WdBB0/NRUBp/V
Ci1dnuZ/XXzmZi6dsb1lVhjIKZykArB57eZhzPnDRwYXZOcoTn6LjLwyJGJcB5ki
LHqxgaiwLXHQW3+jWERQf1pDVyCmncCcG3ZTtZw3+IQ0qtkS6giBpugPLczWGnDH
dcJkeL+VQsViz+WrIWJsf0AHuHMsXDY7NRKa35TSnlDpgLN/5oevrJVYyYScYapZ
mcybbDhKR6xdBz33Ne1dcdUS8H+xZSHBgpxdqMu2JgKuaLN2/MRaC16zMEH6eaMj
6CFHEditdhBXeb+oGPmxeXiVnLs6HBnt3ocPUJP1Wg1DpD4QNRBRRCxyF8Pk+RxK
kqU80la1OcHocQjtnXiSbbK0GhRWTiPUuHsSG1HNntkwzrqrfo+8KCa+BmDsHzwi
Lui7pAj5oRDIsv6Q2+ksLDgGrsxidLZyCuRhF+1rlbnqS9ee0Ak0DxXLWVx7PaCd
1OhUzjR1gaQikLgyWGWilzZQYrgVt4Yk4/N5BZ8iBDaqxIEoL4atdZvc9VDBNMaQ
1z2rIoIPNUllGu6baek/sM7MjeYEB7LLXjm0o3RVwyADHGuuPoBt5Kit1uY829QS
r9e72g5KS9OlInB9VIz+12vR4/TH/Jn7KUs9CpMF1sHXzYrp9y4ry9RxexrVCw0z
6H5e79+xyBBYqK9E8dv1Ls22w8IojIOtSLsZHoGpT2sTN9isz5rAhtzJmjLW2ad0
wAZaYY/LtPmPINz3H6NM58hp8TsVOvteAm1LIzCIaHrBfDS6BL2GedQF/wV05SHT
kzmOD3Rkw4LLd8EqDFW1GJSZwZU5ycSE7yUklVZsHYLdSkYBytsCebrCO3A4JzQr
D4+puLy7UJMg13/8s2ECEmQtbUU4Dn/6/rcbj6jHsFgWy9h/b+4c5ZBqRokK1ErO
XXbbAbUtKXedIU/8wtAu1CMGFkUmre2r/u4xFGci0CpJJNDgbWolN7Mc/2+fE7AR
mh3sHs4jW69AXaFlf7UBDjP4HvkncL2oUkFpUd74reNmmrUiIlZ1Eik7wmvzNCaJ
L/q8DwSI6esxDYKZ7ZOxC9p7/DngbT0hexRG1f13Y4Zr/f0lpq+87Z9G4hB7hYC/
sKnIOvjcsLiUsSUh+sttuMOqulDcZ8DV0FLoTnwvFyM8muXufpnKZf6XOA2QFcHg
DTDdSO9zWULpf1iIjtl5EzFjd42qiDATWVcM3rcaEFARibkaqMOGWit0s39fm3w2
Hydo5SEPRTvynPP21AvOC7kc9M6lSTB4OVB34dEYdDr+45CUFJZ+fP9uYoKrkXoQ
8gtATWh835poQqUTpLGrNWeDRAqOpbY58i66C7ievJ+gwP7R+gPz8wMDxacCBCIz
jc0kpiW7UxQ4tjeIDIafmKwFg339YlbO+sLW8MpK5dWIFbhTY9H5MbDl8t6IaKIT
fnfhaOhRVucxtNZTjyBe730L8gPFB+pDzq6NOByPke+1bClEZttkHerb8Rp5YoFZ
PncuaBZqft4M3XROsuSGNIR/CPlXfoeROjhA2t1/bh7G1dtWRjXl4cqGqUctkA4f
XN9/CV+S/5zI/prO7FHyAzcB+QQwQQX6CSqVVkXxHHASVupH+L9LmZ2JTOF5Be9z
+JTerk8s+03yhjsOgq4aKcjMw86zykizgzZWinEghUz99n+C0WD8f12xGA4xsD3s
UMOzIrupF7723wHkZZwVtXdwXnYVWqbBsRGcG1gPfihzw2UbooKc3r3l2j5o/+em
SSPLFN2dM4s6CkSsh3e9mhw3moFlPbdtvogM9MtHsiTry6yf0wPv+CQ8jCVe5KH5
2IIPDqWfWKWMP2s2RcmFzdY+jEFxUfTNXyD4S+f3jbUQsspzo8uUjVJ8X7CWcQp4
fBHJIWNa+TuAzZS/C7dAgmpsdZQ0jJQHqrFRAxZ/rS6B8PydZxLwEkc+wACekET1
cEth1pBP3AI9hnl2M9z2llWTydMS9lfGAh/w95DMzCKYNCktmJT1R+1Wah0qiY8V
iHgqRwxuiDHljVpJHP3dczBk8MH9kGZjyRVOEOGRQVztS8k/cMvPGT36vS7xQe4r
mPAXJnIrMEvPcT7cNpslYuS9PWmJUy+DU0eQAnT7uKmpB3YiqRVI6UrMldWnjrzM
/aD92cQzUJOmcTsjt5O7Suq1MAnCvWaZNN4D1ok2G2M0kIFSy07OO5Qq3MBN5ZmM
+z281qaGSeguAflN/ZVDW67svr7Fdtt/+Y32a7IydZUPtolk84g+gmk/XvsSK97l
q0f++eG4TDG+nPZsUqgEsjpc4xS4T3DuslIzkZ9+uFpFF6TUE0ZNnsZt9gg7/8IG
8QiaiDfu3UPsiOYWUhm3NRwWLEMJ05OjmHjydb+wvt093PCP27bbAIwnBI9gL01b
PU3H2pixuCD7UZkw4uRJ8MpoZbfV8U3tb9rObVHB2fxquDETU1SDbxcpy9GK/Kwq
4EZpCE6CE8GksQx8IUd2WMjpI7mrslIZu+54cUOtJAo+KVodg3IVxBQGhcnbK38q
zNYCfYTddIIM0ALr1egZlDizJEECdiHHbcd9DbdgMk8dGKPtZk32/UwfKDFyY7E9
pgQei8kEJe5t4UXPZKP7BJdQj+dXL3oo667LpVDM7pziq4izWq9A52PGicBnu0l9
w+xfMY0ctS8ct2keeREC6zV/cjMIZtvqexxEelDPMXxztDGuCH2exrW9fvWoPTrP
LcHb2rrbdOZG0ETeR3G3QOM/8jliN8VM2LfS4Fsg11U2sHv/AGBZVWFB2gk5eImM
WDblnYWzL/pLsVqLPx2CRHEHl8/neIwPPf2yY12VBACTjrVXvh24K3Q9WS6Jyc13
UbpBYuirsltjDF3jqFArFbt8LEei8uI7KQzS325UFwQGi3seTCXob/85Yw3GKhFB
SQf7d+T9Ter/nOuMa/VL9hbtzirURndp8qPCS16JTwMhmzTieb/V5Y6IsBcQz4mr
3rusSeAnKcZ3W8OyDsX0JjZwUHaFHTpsFxMpPFqBGs9tj99qgtUXH6/6wM8hAbgO
gD7W0eXJEDUcMJgJoQKFISG3ws3WtFUVGCBKm2J8f1nR3VtydvFOTbp2jccf+9AV
kRomYWfip/IvgSLRx72gxOvIY6OLJStRxUDEnjt0cYtJLh1LNHPjGArAjf3JRaXK
wN9imkOOeXnPIMjdNVS83ZtNi9ArH9M3w/Nkl8FA4JwK+48m56SZxSrhlcs7zNIC
1k5cU5NSuy+di3Sxf7YhGjGPb2X3/rYGwzHKuHGFEWPJVs8/zhOGPX3LUEu9nVq9
45uHHCFrtmtbAVQ1zXGtVYH5mLVBMaw+Rzx58j8M6hXcZZFbiRbcidEr5buW5vIF
zx4B5AHKp9Q4zMuBdbd7J6YH3negiYYI1TG9hBuM8hDkOQPXuYG3rjgJWYqqlGaA
BRIa7qMCmGvOsbYhGySIAdh3faL4rEargLpLPsWZifJbjo0/4x7jiILlOtwxrt06
Qb3OQVY0k+zWrTWfYcwOnsvxzXW+levc0leWeDPktOmEfZbu+flK4wPo8dfNA6LO
2mXMCwBd9DzisOCSUtEW0Sxtxmbv7hYubcG9V2skm+rpIkbNIUYSDqXpcEQRAZCC
6xU9RWyzlzz2fXXnzqH8gkmEbrPzpCguKhnEDYhQ+Gncx5Yu7RWDKrk60+vcpFBv
cN2w60PM2V9MrHAgsyFnXc14a1wRQnUbV75AcUq6Mit/z4TGUxuA41edS6jRSthY
F9p2qHXouU4XxvgFfRATl77XezVUa08IBK9kbrnidnTC6IdlA7ax4vqNVpQ8HR0j
vHpE+OzzRE9CmxcFsZsyiPEV1HR1Jjh2Kk6F42A4AYmopOmvMipScTcyztOAMzS2
cWA4sNgoBgKKrJCDXbE7EBye8gEftraOd+IbBiGGJyvwLpA63UAJic0brDZ6+zL9
we7NDeEUVRqclNI2BX81hX/Oun6vkbg26tgyegeNFE/+YpB9u7iaaYAbrBbHeQUQ
v9ChP28Kwt/jI2QUEy8nhPwKrRNpzEjaAVNFoptOElK9m6xeuOW/24sZww5/BsLc
eUiUB6uPrzySI2ejurFuseIWtCGiCYa/X68H6LWgkgy6xLtPU145B+cPRzO7a+jX
SXbuci5DRdZlUhY+fPG75IvnUq+y2RLESivIfl7xyZumI9jyZvUfUq4rR2ncd8jq
6UyZr3n+pDd0PDJCYVjM2bVbgDGlVxPGzdyirwJ4b6pTlwGqoDRc42pHVzAZ+dWe
+ufRFMz0pIXjBfIQ9ZfhUxXh59uLd+lK+BpdTD4kFSNVqDexYjefZRFv16ulecNA
t27PZ9xTSDP5/h0OgPlAo0qL7WG51cFmxQTTA3eaGQ0ooGKZUIm8ubLBAJlbjsWD
P7wBTy8SQZQLvRqzbuTYBWehmbA3ni11LvCwpIDTFx9MMYNLqeqnFaSbwSodTzwX
G7c85wTv3DnVdbXC0aqXeDVaJ+R7yrqdmcuAuph02IwSM4xwaNBfSvCExKpH/ReK
UoEPu4LXZZb1YqHa8aSNvt/aTVkh05YV59bCmnw4Jdp0Ryb9QRjaZZ9RlBoJ2Vky
MatTPpNVjYET2EWJPitgp3hLSGqFiTDZ6xACaDBEeOgi5vN0EOSomR78kTkyxSmD
6U76DCwXL3Hrx9hk6OGKOQA8Z9t8i+Vi5+bFR9Hx9Q4lLwPMsvi7pcjJGMG9BMTK
B4nowLpa1b2hZoy1hYSX/EKLkThH3cGHLvG9wnY3+3NLP1HH8b56AxRL48XNICfn
EMEXFNvTTlmZqHUMM9YaNQCps+S5PdBpPVV4EMegt4qfJeK2Akk+ua5ITfGyKjIx
CV0VtEPJv2leguhsfhuyF0p4MW+zWVH+obSygPdFTHfS1GjwoHxwu7PGjbDYRj4A
6JjF2t2ufQXmmG/S1Phm7BiRMoQbGVwDZRkpSKOIBvJWjc8uhfiMPKOA0gyPR8wG
l7L63dq1NaEufov4DsQ8zL4sccRAZckGoJOZGOSYXnXEwTjvCbUED9CHKHTsYMPx
5pk5iiUm9v0y+396CDnePByl/J1SPfgByGOThqRUQwt7k1YR9023P+0VGCFLrSv6
4UFaUkgqU8XDdCPuwonn3bd1YhZFDFi7FjZy6iPBRkaBIyttqK1w+Uzpt5F5eKiC
EOQ4ISgNP4Vf3hVh/7uazAyddMuZZKuF5U8N0As4HjccfYowdDQTyhlN3hqH0ckn
hVGxPq/GK8zKi7eWsg/kA8aF2CQsv3f5GMAIP4RfDo+s4OtOVL8MURSrGyLhgCYr
4n8/fogAdexCDBsZiizF0OZWW1+54CHzSdWyW7q093xo+KAmpvZGeH4Idh6XIqfv
NGQhtOhnZeaX/cFmzYeXNNoNtongQXpVXl1uPhcN36JKoTvkydFAYNztzSgk4mcZ
+OnpoowS647wINVDt1k3yg1fcRiIOql846G6Cn/e/neImxVjy3iW+Kyi7rduvEjh
ZlJP0AjVcXCF4yJ5UZkZGwL4RRrIfCuG98n5KxRXKPUItza0A+9cO1W1Yeq0P/oo
teBvXZnHHRNwWD9rqefQTvOcjP9Wt9xmNgdDQ4s/fYv4bVjzNcaFYvJZctO/9KUL
FeRfnGbRkKr7efZXJ+L1eczabkFoQ6I17FVidNF0YXMeAHlP5p5IgObROaoTm7t6
qoR1MGEcImVtZ6+y76RtsvkmmgjOxBl9mzbv3O1UNvo+yVBGtBZqaP976wvXw1iN
PCMWd3V2+3iIx78okP1YRy9LVxZ6rbZqiSKgnhqR4UwoPKttsaEy7mU1VldZwq3W
bF4kCrJ06nby/xJV0elyI/UZB3xP8kIyZLObSx1BTjZQVBV8pvpgK38eQ4l/UqRm
qWstK3n/2kM+0n5VSlEI13wmzWGdnHE9GTVl4GH+i31beskOfJrmMcfxAjBO1Xvk
RjQIc2JfxscTusviRsToQfLjLaEp9u28g78FHdNllliWwE4UCWcfqzYgjqa8bka3
HJisf4vfmegk+UsWyAmUtnW5yjVfcJCyB4K39xbZrywd7edBPjdEh7U3raw5kWrA
+TU3vwRa0WgrJRNxqf2bVACncbymULYAmnesJQM1V9LpJ7/5tAn7tABgbOOF4ZX2
9HflcAXU8y/Yf92mtJh+/cr1ISYyaa8Kyt472tL7uQwR0ryhAU1/ZLGANUUvp8i9
OBlBAJEeJS8hhjkvf7l9SlD9+J7jzNY2AopVvgZGeaXGZgC6eyFuGbY9GJntGfaB
XEyMLUlOFM3vkMxAOnDNEGpEUGaMk3hH60k4GEtxu4xJGs1DqNLVGyyV3/0b3rvH
JCsclGH5COwQgJpLemh5ZPh4n28UHAMFOQXfDbHkgeVwJpzEX+d7UhDfH+hSsFOc
Fy1lq0OCrdbuXg33WX3iJAtrke4CszpegIpjjIbhXUE7hSImwVfyCtHitPQ4nBKG
PTdYg/8L5zFS7FXjRPoHunsnD5xRTNMQz+Ym5uSpFzyDOBenrQUBIx9QyUxrOtaN
1x3RWMs1q5K3VtvK77Pxw44SoGl4/EjeZnKgQO1AKaVtUkpGpKozhmRidHLQj/nj
znXrBwfP9KRPHHg17uVJmx8tmDH9L8NF9Ou7bjPfHcdZVTcAxB7wODidOVC+bPZ3
PVJ2ZmCH6U7n1aR0APp5rL6IFQB5HGtGpYZC18ol9BXW13Emxl7gNBwhHGtjMXUH
NiFRCAMQEnDjsoEExNTLfYoAuwA41zoSf3LJxyPCQlpRpqnZB6VaxmPMKaJld5YG
FP6K/CEmq69d/5dDkXhbKO9vCGanRSrC485OaVDjCVePiGhuh0L09ocx+gC8K1G0
k/G1iqxCQLN0D43zAz6J0HLbnd6jBELsKeDdUvfEPAUFhmQgFvvjVl91C9UJeaOZ
vpRg76tA2/x8VO2XJHkzIdZad8/JFHMbjKAtz8htFy2eVRDUS9BW10M9nvEV72d8
g+0KNoBbyZbTQnI6wCHquhSafxE5mLCoHLqWW5LwoaqgueubF5fM5klxRnJx8Y2C
HO2dtSOG+88Zu1u11r0M99TYGARpX93SJBZSusLJB/Imn59RcQGzNB4vLaIpXiVx
CGfuuBUkL39BBWF7uw7hg1G+EGFFwIWdKL5eaFKI1We/4kdPMS76kr9YU0y/xql8
JkUAYrWRIeXp8Y4aB9/4XQK6ZDpeJ03eK+ucJeyubvcuCPsIB1q9dcCG9AjPJB3A
OnBGItOBee5kgtbls98mRSfEZB/n35oG+vI9l+yydCohqBfsaiYC3vWN9ILNBS25
RD8QbQTsL7m11YZ+DR8TEeE9PaJeLPZkfX4iY6GntqVWa0I1QWt/hN+lNLItCUs3
Y5HfuDtL7fKkedARpY9ldTNKvWSdYEyLluaEiY3JDH4pODfnqHIMp4O8hvtREo9Z
UP08V/l28+Eca50PBlhgXv7/l68fRrbi5vfLomdLAqPl5Kq/NfStLr4/a8rAV2Zz
TEueNjzGjbnD9hwUgtwzyzOEgg0We7Sc8J24KGOcVBslQdaamNzPounIVYjXCWYw
1oVUQo8J5oG36+m5GofBqnmTPnQaJPhkSZfbhrX0lByacESY4KeKM1AQtkpB9aat
p6bR79tiq7gpofTOzZ5cuUY5gAgFoUG2S1bUJXtEsbGw+ttrX9mFuj6e9XWv1evl
C0B5uswvpGo0W8i1WkM5QwvzgyPeDec0A7q6whVDP/0UHoNNP2rCp00XIZiJLMpT
wdvI49fDy2y7EVbxmuimH7OfzJRgK9laeDiRris3mtv/qDF95zV+jn1FajW4mNr6
OVMtsF/lbWs/pCIY9nUkspesmCZL7PRcrBfOSOU4K4eB1HoNcF9nCzwy46SepiYP
zX/7rKons9HxJZZVh9hKTk7p94U+uaxPxcc2B+RY/4eclg742JGmFBVfbeDh5Olr
knqK5+7TK2U56tXUAOos+Z6vEz+kx1aDpbGLKrHkzEYsLzCBU6eA9MiEPI5wmk/O
s1ZSNMRZABwxIx9pADLzqqUXILpuXg85iML+4+8XKDilh1MGR7ZyCGzuRSdnN9vu
yebj6mDL6QcoDsuF7K/HJ5wKa4IFikFX7vg5ZuuDw+ib8SZhQVO9V4Ta2TFgkFHa
VqolHMJO2uSlGR8mf/n7GGRqchlT6gEO/hrdi1KzlhTeCthAN5+cEp4jsllZ/OUv
yQI75QFQVMWVCAbDDCkffZnmDZeeKbBcGivbMACZPp/oTkrwb6YTuM0SvFLwlc10
jhgv25kGHL/LySD6yiJoMki/VQv1cZh7oNl+sMeSmbE2dJ5hYTLoOSOXgE/CMaXr
hNaBWzb0J8R32WzQgy1AFOReRn5g+EjyxIaE/qEBB7wWN8yuONdiZD4RuhIjsJOe
Mpxzoz/fubWP9zBRmviDzBcUBV59zboSTT2Fzh1FjBcudo5gpMQNGSsrp5KpyfN8
sEh8I0SIwP8cx9nw+uaPfjQ0UAWPr6kpAEZYGqwW7EVLCS4EdO9JQNPFUKo06WSV
WOqBihgNSmN3jwTK5crDTXoy2luuZbamdZcQEYZEmpaK2U0ZT8vqNCKF0iJIzaPb
ty0IlCTmZp3LV+XjS4gpK3F1nYuDWCAEe2+5pIBCnC1XikAo8IfYSSSa1/8vfnQt
p6TTjlvdZnP8O3jyqtKV9fOQdcTR9ps1e6nvtvAA2rRWs76XeP63WpxHSwycPkmC
wvRQU9LxGgK29jJmfjnSBPAmq0eT+1JLhg5k8mUfD3i+8DdGSNyBUB1fBc2TI8eW
MInWKzoxcKbadNx+XpM8yvWvKn/ao+FunGkXbB3n2sZLl7MUZZbzjuGKFLYytIR4
khe3pwUgzcqjxY7pwrgCVvfVuvndWPKYyLQb9Ty1TwDTeK0i3JQ3NXnNC1Hbe7m4
8U4KTEaoLGsx6islMqX2uDXu8Z8ZI9tYHm5srOF9pAsVmbQ1MnTZI5eyTA4lp+7a
tKVjpDb6GJlb15JZeVsnSax6c4Y5poZnDAxiPHcmlmy5OVMR3Sv+n01uGP4hevh4
jJybd1u/hqB9DamDIxqXlbA0+xYek2Ol4B0MpqZuDxljSoTDu44N8WoWJSUFSrDi
V26VrRuBCw3Ty2iRTFcre/h+JuKKiK4atCGIzn0f7e4/LP5BbI1GU1BvyHhk56EF
VwvWnLjxj8d/imtaJVqYcrryxj+TzHq64pQEeUpsJUQQpS/Ybt1bIZ1C+LRpM8oy
6XkDidHLP+27Ty3WubND/D91kq5cWWXbYz/pazHBkKgWHjr7zxgi1wQHuRf6MnPu
7KLTtuRODCY1ZHLNpF7CSKN/7Wn8IeWr/HBjoE1+A/Lo5Qw7TuzFuXn/xIpQH3lC
QOQpwh6DEpBYjcmke5Q43RjmrK25e8KH/z1wuJaYU0mgDYfLf/WQOCExhHg9CBto
08kVrjN58dMh07dreM0FqVW6yCeaSOiQWkCBauqqxi3FsXWQ/LkiU1nEOSy0WR3M
Ac1u8WMxOf9Rt/a0zAoGfbYgcY69pVEWgmhNRLi3aw9NHJqg76CrHnVA2fJ3dmZO
jEkN8uTflyr++l0aVcenvj1CsReaizT2y5ntF9e/Ozn1ttYjXgvwqNr9mXmo4AsW
BANcNXRNtM5ymSjDdfF9+vfFz7tUlDBtlDjLmBTU+jsNc91FYLF7Rmb88C24oi+4
MKsqbllt708RggaZhpgPXPBgkXfC5tqyLynLp+IhZmHgSlITdbuVBINZknN5NoBE
UMu9s1Nt7zls6iv5IqJu0nAjQt6ZvFQVfVYNUd+I4LvcKY7tOIcq0+6iF+km6URm
eJw48mYI4tmnFtVQXJLhGfoGbHJXuH6d1Eb46t6pQShknAEBYymWr064v1z35j5l
dqMmt4rXZH7K8uG4dvFijMEAlXiF0IZl5lOiw9a8AnkBDA8lwQAr/75XyPITrm8I
l9cfRE7GPz/UMBxVMrC9Z2nfNE6/RR1E2WguTRNPGvpUhWkujoDUUdBxh9PAYO9w
QHeT3xgxTJbs0FCBiVv7gAm7xxHgFHTjetxVAWmnQhWcUCCyr2hx5lLtCRdCNGFd
JwkMLVtoyVCBQQzrjZqy0ggxiOBwRRD49Ig/D38Z0Gis5UTLR5XU+WlOBv+u/m29
lUdGQuysUsuSOSVvWVtY7F4QB6NhhNfGR81sVaEc7C/6S52v0kHXljsKCOFD1UzQ
zy/GH3KPa8IpswgWxX7JnYn/UcmPV3XlDNK10A+jVL2tVX6uFm78iMcjzYFlNHqV
zQ+2efvKBgls3nvAh1njrJlhvTOi14/9bQCDQgZ/Asf/dH5Y7gtArr73KlOeWztw
NdsUtyuZkt4jmlAITk89X6JgTUh/zecLrWq+SDYfTUrHbbJ9Hr6hy5lcMF4W0eum
F5NLvSxoNmILVzKbMwVWZnuoGM8Yw0bFlE943YgI9apJeMum6zxJGGelSEkbuY4D
wnlJ7F1zTIVeermKF7l9ZkVbtOcVEYm1qKeIzvmYkBbszEIsbxUwZWKELMAy+vS5
eJTyEgfxf9o4vwoR8di5231vPzwFxHIVId4c80iaedFoRcTaVGbGmV33rtxsvnSU
X5D/tWp0Hk1WfoacqKB87ygNnowGZg58HmrNrsjFukcVaTS4T4f3S8gIAzHzOXVU
I7yKvnyFuI/Ar2rYk+Gzp5vax55XVXqKspUkqYG2ecQZdimorDxp2wXNYSjfU3o/
wu/MhVlm3ujwgEIzqBUGHntoUO3H7Oi649maMIhT/LDfWJNbbrn4prBV6iJrkEFg
ktBEeKPh8GNjpHhUbzyI+4ALL15mtO4ukJkU/8TBLHhVfIPUsR5IlTpcwtsq4NN2
BTzLoc7UzFFCjo7xpTMtQtiC68YLxML+jYx7K7ZJK2nYHrbtqOcxk7dtSVyw2byL
3tVvE4TFe/nVGx/EWZ59xn8xpcfFQ5k0+jnPbV7doxJlwaAnLbnITfKES1AvQKlR
1qTTw5HlmPiQx5g/jZboWIYOvZpWMxSLJF0ufN8n0HEYaCsTlBDiBnpcQYQLalBr
muNt+vqw0fvwb/RgIwd3UgV7jhE8SIxepPnfrBwtvDfkrGRdokfcLnLjjXAixwh+
5EyWX3hBGnDPVAqawbJ+zraA/k3i1CxsXzy9/ycV7fqLVU+VBlN4BzexBAOyUaXe
nAVK6zhzEv5Y/IH1xxPZsb8F5NjsuMvE8tDBX8MUR47qygbsJsxM+T4aXjWde4iP
2LizbG/+wnwFNLryv5B6GeW9jYafQejC09OHrquAcYrivJrciXFv9Bq6JpmHgcyM
yWTynoh6VoJaO90Acl/KtIlVuKu6cJPdgx8314duoqc7Dr6NPQxd1/z90j3dIQ4Y
8kwN4T9pzbgas1oWoQ+a4/KbumqudI85gDhm9AL33Xf27Vw7orE2jK2aqmaQ6zZz
e2u0y9cxn3NiSXl1YHAdQe2J41Sa7S/ObjlBIJf/j+QX7PTMJYFx6BMODJ5lFfY8
+O0gCEoThlj7kaashHXqMPothJiyht8fuuSFTj10XDXj5OL6JQE6ho6DQYLKt6CX
H7hGA6pXrWMlBC2CnSuwpDiT0E6RFgvL4J1tM12l3yIdPPMN+mKb7mOuzrX3EibP
A6jgqAmGMsR8rnNCUnR5O+fFKKRKal96ICWf1mse3plBvKeQ+XsQKSVDuTO1sJFJ
Wtra2mT3kuCUD9BBcW4XHDX+cKeZ1PCy6MnMr/2M7cdvRZG4qH29BQlYsMl0EOF9
+jA6CmEUagZM21UuWy21wn7iAM/OLS7RanJbrvxhjh4UHDV2Kxndrq27xa9dpROE
VTsVirH+Kauo4MEvS9EbSzRINOjZlqakMVmLBHF7mIQz9+sFLYylwgWOSbXsRxSS
gDhodW9sjCSYp/9T6t2qAQ5MmLD6d/ZNhcuHnJKS9bJ2Q0nEZqEC033uis9qsZIS
iKZgfjm8deZplHjYj6nSH1/fgC0kKCzUZtdD2c8yr4tosPSrpB2Q4FTVNEkgmVPJ
JloZZOfpNYVskaSU3fUzS9LUelTS67ohBvXg4noqVLO4WjipGTDwh6QQquF4WSsT
qPU9aZ7k/pPtvSdUCWM7e5+puAQ/OIKVv3QQuYTqtIhSMU/2OKyv2KA0GHoNYaBW
ZnJBVjmhCq6o0wMbTxhlhIHE0Z83B7WfM0q2+09ePu7oweGagBn3ySy7Tb4lc7bW
nOsJfUlJZS/m4E97tdD8nEPulzO3wwv4CEnd/NTNf303tzVcAApJ8OjHS/Y4jWTh
tHWIliA8HJBLI49/W13D+OgVQfiT8rHFSAaYXlBX+VfBgT07xBgcBaVtvOTJl5je
1RdqX7td1f7y3wt4KHAY/zkrof9XeBBFXRWtso1Gz0Wnjt9fl1oD3+D6tNqeL2c9
UqvpytdCfh3mZAyelUkKLqqM1WZiT72+Ca0/Dd2B/UYeqs0eeyHADNnvIbaa9jqj
arJBNT8eiQn4q6WGGiMr02VbJ4KiD001Eh9wXx9bIStNZ8954tbV6sVxa6ikEPh/
JtVe03du6azyeEJAo2SD4h1awmmxiK1K6P3Il2YFiWJCHcKzRdebvLUa05C1PCdK
Enxwhhw+E0bb86WRdd3MuicPR9k9bPkKy3T2jLgUoTMor1dFk8xkgNsWAx1nB4kB
jlL1CuCglbCLqXC8H7mrORdhSF6QvAkAs3q3S37hVej1zDuDXbSetFTR95vo8g4s
o3xD03Yr2rK+DJrBVVQfQ9BbdtAEKUNsgF/Gpi3PQymZ30NbwIByBJP/dmAx486L
dwWtk8AWjguEbEHzCah4i1Mq2S1ooI96dmCZauVlFms8H1feHGHfvTOTW6f2dLka
0F1FmIcdb8nN83NK2PyLB6ezbE+BzMe7zvmPCqMEnhs5Le/oL9+EphDy54wL/3Ij
b4gbXtsZJpOmRgUYlFJCOqxEZas8ub1f+BekLJ2oYyvAH83BnNOJzZZLxOjoBOoZ
tAsjHnEJqUJJsyZN9B175hpNHOS25E+ATd8ufXIbFOQ+lyhqKK8guNcPGl4B6TYf
IC7ofzOA7tYiG5jmOn+FjYcZEcZCeRSud4gJcbK5cT0uS2LF+mbZd085DWmOpjui
rTyajqohrqM6SdehUvXZv/qFfZRJeCgwG7WdESgJlzqKM6+gstGmOvb+2U5CidDT
8CLMdc+Bg2sj2tbzm2PoDkqkXcaUb3ZgaOAVZMiU8sRoAOT4+aXD+k5wEgcERXrt
GNbFy3GXWXMATmtH3wDRx91gBnRyYP3TPVHYARbWKX2fb3SvrhrhtWrJtugb1Gfx
vUIi4Qzm6mPEMnNfirZRnwOKOF3IYLPRz12qPO5CkFwV9jIwxu+0UPrWCAQCVy9W
rH3kQKcc7L2fBIj7tSxvNDsw+5/hP15ERdwqP3uKEIly4yMOVVoNeiLvsIkwUCLF
kT33MneGEzO8Up68Acuci+aDwjpZ4+tf6a0iqbk6kRpJI2c5wu9JDmiWEm6RUrCO
PzqoPsYEwPrlhRh+c7Qa3PsEhPJp5VjNha763TQiERzeVjr89zl4UXjEXM8XE4H3
OnL5c9Mbf+7tuSAyAGK4EL269FwRDKNPWLfNhy0IRT7Gm2LEPWms1OK0aWbaEFU/
Vtj/kgB6cQieViJvzlJleYl9QFw5Kvt7rfp6yIQs+haTFD6Fd2rK1vFM1zAy1Au3
G3Sx+uX2zpmrzGSbn+mBNRlH52iBNyJL0eYIU7NJ2vwSH6y6LTSdgdVw9X96Ey51
0xNTq5OBOuwNfofvl3Jw2nSjo6fhyLDjEkqaekpa5PmqJRLJQ3clb2PvshW3fGaU
PdZWKSnGYs8Klgnu/zANkH2Lf68eb6xj6+meJt6htHM2q1pfnx/btTnvxyEP+mm/
/uSlMcnqV6qAs8U3LLjn0jCl5jGi7vOvTFbzFDIgvUGZp231nz0AVSuU78PchPTl
NVUfzwGlnHE1gcalHRK7KsoL7FDpqgs9rPPO3FrVyb7m2jb7+Fzzqg3KGAPKzcaT
2xAgRZHLK6eeWiIPK332KYy/KbrrtPBI6c0SViqZrh8lC2oB80/iM+6KgHVAkuDZ
PzJvwRHQx3hCqmP2GF5udVqboshlojZP+Eat5RwhOE5xoho2IBqk9exE1dEjY23G
WwPbn9+Jd58NY5D6bsO88UkyJHiyez9dbFmXo7GVFZkuGbcSLmy+85dztGc4ph/h
e5FbcEwTDllMSYlWBicA2oxdSuws8qAeD2SID2n3DIUIlryxmDbnLNuMJ3rxPavq
33/701u0fNz1RY7uZnswPG8SBRlVFqUyNxiiomEJSNEEszyWEmFj8dQfqJO8eDGa
j8J+BgM68TCMIuCFjXtQrxAe3vVC/v3Czx1MZMHhVH8md0fWAfCtzqj1vHx4r5MZ
/I/8/wW1olQtXbk+ax9BYWMu3h+SKO+dbBKK6LF2S0aLTWYSGLafltduNOE2efgz
dcwX0dlPSv8c29cVtCHHd4uBnXuidFBD5t2nCg99rx3nOTnhAJAyszynDSoBtBQV
W307NOBizSHAiObVW+/kriXK6h/aVetNNK6R4h3vIsSuvhyXSzFzur3OMkSsZbNo
InZxRcTbrVhI0x/KYaNQn+YDE7OxNM13KJBlmI0nw7lVmHB7L9N6xAoV5E7bKWIQ
ssYKtRjqqha9w4drlFnc74jy2MuCJYUFge0Gjz/5xiK9fCsvzoKnPOFTT1fZUUC6
Ckj0obLQ/E0F9VGy8NsAkknXdvlxwkdJU3GY08BhNqdarVzUA25ZsfwM0kffoj0s
6B5oY4D6AgnAPOVECqg5DJm8TSIPff0hGx6RMI+O+mgDMB2M3ZmPZmWE3m3q7gaG
X9V+iyiaZ9Dl2zDZuvm2GFEGHs4yQ4ggpqocN0Q77zSMoDPZB1Nb/jHiTiqsPfpK
IomxM9nZFEwBeBD731UUJ9dZY8C+ZIRGTvh3ce6MNt+0hFwg9W/uK8vt8BhDZqcs
ofbeFrKxeWyIeZz9OIWQIxvi3+XT6KYsbI5bl32q9n3b4MNNfGtdblyLnLgQWuwf
mArZOi7nEo2IAXZ0dXX+zeNAoBJQfdYBhx/3+E4G/MdjNJyA4VqdSjxL773A76h+
+yfCZG5qJ+TF+lbja2K7qryff2XtMYR1+ZQZDyLrPBSYxK4cleeCjwvRhm/us5bk
2ziTH4ereZ+AnhvRFUh5rOqf0APpPzcg84wPIjV5OvkKQ2rHI6M95iAD0ecm3yng
0n658r+tZpbUfXwSzM2h0HjT+EmlgU+OWEGq7J0/xwPUG5KVzpwQ3L+yeZ5Jfh1b
rOtOk8pupRAe7QEmDo83dFSpwwtqCRb93Jz+toYS5c/h5RvEGZ1CkcJDWSodK+2K
UqNz2HrNsGDjBxVCYocSh1GXODdRTGcVYdZbfixdWcZxXIdQ07XyhSCLjd1US0iD
0qOar/S9SjMPovN6CLrQR+UrypFxoMocrUz0fnHoloZobzkr5hMmkfgUccGlgN0p
NZ41Diie76sIYJJqkpSku0GEOmdGcMHJKa76TvrqHjKNBh5ThrdBY3uJ7ticl9Tl
eA8v1upqWuQT6IoS3aGvbZ+Cwpc0bmc79Xg9/UL5k+1/x8Z+JsUXxqfN9w7uq2VQ
kpnzQmNxR72QFGDri3V0pG9TwRTI7XV5F7DLNK0AJQ8gFI8muhpVpnsHicyicO3h
bDjI3d2jtedUR9JywpYB0rJAhpyxMkPHDe0d5uo+1RZDGm80H4klAWfhy2Hs80/I
TZevZQ3/Wi0DlD99LcLFwwFkbBNA4Ftzj30qmBGV4eze80VA2tU7RNRd6mRdAWj4
tZeo/Ghhy0bT5HrBugiB8/2sc7FjC0he///YI2GHRM+1Fy+79AA8K/ZFqwBs3kpB
JaH8Tw65z7obUI9mZ+UEn0SbqocOJc2oUbZiK5TrcJBQmwNtCZbQHqkSSUH6u/XL
9sYKDVffx+cyENm5xP7KYufHdo2URIfqvVZuzc1LpjRDpa0+99zdInc8BQtNy2IE
zzkoQ923CvmXQ4q3sCeN6TBLT0lGXGsH5ZdZbOFr5YeTKWdU0O3puD3dfvdqEgul
FEneX8Nz+sphVuV26rfVh5aNqNw+BS7QKRZVeZzjlXh5oRslPOqEycQMPLpdVhh1
w4mynd/snv6O6aC5QxCRBeSbe+30IXmAmT5WTImMAujeq8O0KbPwNLWc1iU0rAmI
RDA1AOF0Axru6Vln6NG6NxsZo4BtUAB2jvquDdIfoy3hJw+/INhdHVCL7BKUt8vl
ZAYVOdAhTHpOAkjMEw8qnw+Vzp64QPujKNYlXccOC/9PibnZchI+gDOGqP/tJbLM
QvsVa+AgRg+haRLsFGIxDvqZ7Kz9GQ2cEFBP6HF42cbQ87D/LROk0/nLUfXd1ILD
AB5Hl/pLhR22jprb534K63iVwWPBu6PaL8C5bqygSA3Heyn/ZCO2pH1lY1ZDSecF
HjUz7LVSJIZxo9uWT4317SRuhtpoK2SEYzcpR1TA2dIcO6p3xszNd7Lqstr38LaJ
C+TB7OFUm3ZisUOMX0OKyD71avb+Y96D0dUBW75QEQL3HcnN9ipEym1ATt/HKZeU
NMyXU0CrfYgWTn9biaWhOy19Vx60otzYwDinBAUE0UKwa4HFVq0L066jSSDxcoWD
P1dRQE2IIMTKsdPAk/CL7VtzQPUXcnsjCsY214Wv0+gO2ntMv4Oo6XBqwwVNot2D
vifMUZhzwMbE8LzaR0dMcVUmmueRlpGK2SdJGb/FRPYgwShVhrwkStQ+kfHZDT27
Txm7uYeHSd8IK8737+GV1o6WKwyl7mSlz1awcnxMJ5XJh7SpozRfZYbizYrZhNR1
6RNqYghEDTU0O6Ib6mTtNnVH4GE4Y8G9r8guHLs6f0EsKPA9aRsQgN+Rqgl+EaPd
tWq9srIK7uqvQjj99jXeGhDhfYp0qCkEbi4Gu3CqGnVnUJYOgJ8jazCzOazIP8Eo
3Yu04tz1bwT6FC1U2wPrqrJHQmJe32ixfzHkzXmR77iySOVDApv5UTGILIzD4bb3
Rkgdqn3D+XVoodDtH2aAIyqhvdrY0avMlI7wRW2AA1n53S+2owLmU4ydTtqr68Ov
SbJvahmI/Sy1L1kwy7viucu8025MmhooQggZtK/8++Sn+LRbQOGIZ4ccrei8pX3z
kjimfvyK2JLryVFMlh1E4Z7kXX6YpGN0sHYcQ+sExlq0H+9NNp9khEZCAn4UUXCI
AbRenC0bm4qogHWacM3PD7tY2zATaC9aUwzTnJt2zaqsqkM8yTxeW5tuB0cQh/LC
YDczj39VFHj85Kxh6dOAVMbnBSk9OyHqwvcioylKQ3eRK+b4oepvfcd89vU1ZTMK
DMZJq7CL99fphvsCzMZt9DnwnwNWtq9cfY//1O1VlOaQJjzW3vJ00pkyfYsuDh9p
trTb3PKTfOEo67aU0L72pqgW2DBu91pu/3BRcIzHujtTNzvAAxOixqWpaEtxQ2ug
n0FhUTIh+lzo/+qfvA7X3dRtnkUJmvHHGcPPiyJGA+uSdiel7RiT0PDa3Rmvc9qv
O7YYNE+UxC+yP2ZVmnnXzcdJI73jaBsfXu58tgxxGYNHra6szN7ABvz3KHfh3QcJ
yDm8PmFl5bfLuO/JBkolSyrSDCkNqwsT+pqA/ATPu1tK/SOoqL2srTAlM1XGoyqs
v+PBETQQWcdFxFKI+zUU1DBBj10oUBytO5TjNRGXeURHDtlScwUbBFg2EoNg8+P5
I5SmNo8Ie46VmlMvOJQpGKniF+X3Kp2SpGQqhRX309qjdgJE4NwUnM6fDQrePZjM
1zhig3AVq7AYmBuc9HxtXU+3kiPmLA/xbwSsJ/YnZmiYQ47Qg6tkLiwvkmakUih+
gOGo4Mj34CAweeE5e+nzDZ7EO+Yo+HjWScwRAcNKeIJtWVWP3EImT/TgIVUyBL0S
4J7dhgjLCXjHulSRUA1zcjKzdBu2Q+qJbuKyu+q3ci7I4LWjYj67TEDCdGOIXDGa
iOsj8+nnkJ0Do8/cLxpHUF1Mno/O1saUhzrGgiRuBCgQhserIBPClEX6klREIYPJ
U8kRR7mFmltA4k0t0WQfK440o+8Pcnd0JA5vTermkPo2HAP1ZLEX+5+pokutflpi
OW7rbjz5qfjEN6kMU95sREvardS8NswmLbCFDzeWItGblMXLybRI5x64jdH+4yfa
v3F5QxDhUh4pZfy7tQ6bwPd6eXuS4zpFm7xbbpApFddxFGT6CilUqecld4o0jN9C
JCItsxegOfyRInCJ0WOete/vOYNZjOGVxANsu+fVgztzcNk93T4k3W1PgPxv9AZ+
qlyVnL8r35FtoUYcEi6wDrGxLC+k9twDVor1sCbkWVfcRlNKouiE+9Rj5+bpN9Ko
r0SCHP10uukcQ1HJXpUEqHDvkqObpSRP1TO8GUVHqWH+SQ1YFjwQJcdBDu4BOho+
y+9Vd8ylzhGOZ8eQqXWDhlFqP0s/MOuP8RDwn9vZ5r13OJZ8UrSeaCt+F7jxWgC9
G74pwBdjmffWAK0zcpjreT/q9FVd03xoX/AV9k7aberRlFB1SZHBLuVb3CkUxbPm
3DVA8UTRR8eo6OHIJ/fLWNqwUFbdhx2Yu28Zdln2dOPyZ1XHMgAJIuGk8X4na7Wk
JeR3T9ipZBrUCQhdLZ+juYRcuXGzXFuWIASu2E7e4Rqfw5dObw5HdpO4B2v6O4Pp
IdstJ/KpSsd4wLUmRt0d8YLdDsrii0VffsXvk3KwDCAlqk06enZEJGTo1UYBcg72
/7owZkWbvffyCL3DP3GghH65S/RY9Grz0L5R7LzMbtHaAPi/1gKpQqlVRNf692vq
sB7u6oglW+FhyXVtKSOmGZ8pcSTKHXLnlRPWKae91vzZrK2iAar2idrt1rmsKLGH
kdafdkiSyU6W+i8UA8a55cx5a6BNfIb8/mlTUdjKYl1p6cWraR3ihZrSOol/YjyD
Rs/RbSVbnZH4EeTn0BVILZ2SXvfHN513HT++byEcU9CcoR8eGWMYTajt6lJWFxJo
742soQbdgNSzNMlOgsJMzeKNIV883RKMwLhidRlpPLEfDiIB+GyHLzIfZ/5tFFVI
3QmGyp3XOowh1SVWsIbCC1W2+RkJ1dUxKpJXs5AoTqetKoy6Mdj/Bv9yE6OEk0Bm
mJir1TMB9jdvsfNdOnZc/IufG9Khq4wkSM8K+UuqlyKZABbo2QK6B8K5ojUF8ztE
otlulYZjGAm/4VBn7c0xdTC5mNYvYzYt+QJqjHIEnM1g2McEJkKOT/TBoLTt+hyQ
Vo7mmLi/prJEk8FjoAlEELy0Mf2ShaqvM8bqVZAf9aezJzDrNLTZvtonjiGvGHeX
pAG6nYzUcFnl4B2JxAAvKvnto4k6nYG6a7YKCU1C5ROJNjng3FwIPw9gTsGXf+Wq
xqYXwBRCufibEKdlSKR4GXEZwl6EdEgsm9oH24xkXBQTGwKiqkQd2OvVsJH9oyqK
TQNlufxwW5fgBx67hzPUmAPPv6mCs3kCMlq+Xou8ZjbReGpndGTc0y1f1yhicToJ
GVgEBF1wdy4+uUvgMck7NoNd5UIIeomz8I3B/mzf//wDVBCJDeTYYVw64xsyPzy/
i1fev2Wroi6msqGrh96GxFGpx7j3YF9YaDotQtiAGsuezIUqhIVJAzKljJSH18v/
Fu3OWzQqW1V2KEYQuSJkI4fkBGDchaYxyCCzIfkvyCZRD1h2azwCQ3TY0Ux/GVHH
Vt+MXKiNur1CzJBcqSGWX6OFzEVSMIvcPhQwWdd0MYPFhDd4YrSIpMBGI6OGmu3C
tenhhIbIHeBSqp/ackOka+7vSnZf8eeKgeXhW5UGZXjX1TFLhiACBbZ08Honxgv9
Hx+6GspaNYmqusC01km3NdHVJhVn4Gn0LvWLkag3X//BRNyU8sGhiBsp6fPhqV/q
0U4+Xv8BBU1O6RdhF7X4fu2iHEA0862XbX5CVMhRGBziXK4RUMLy97LU7Glhj0MZ
3KAmVZ6imRx0w4kNMwNoFgdtR55bBNnJe3YvI1/OlWpMaal87tiIGEIIVkgRYfkd
9TSWqdm6TQANpINWzFDzmR5B28Xqm8q/HEa6lZjCdSmxMO+otoaPlONyt7JopsHd
F47AmOsCWfmCcayZ4sD85YzwDxhQvDed2dfwUJeV01iwOfQ8uHkf5xx0dGviA+6l
MAY6+UIubk06Z/ZKKVvEUY9mn80MQg2RruddAUDkFPL9Lj3l7z3Hufr5OnoKX1iN
q1/0OJD1682jDOZk3Y9q+Dm7PRkOXPY/61M8ICXuvKtx21B4/CreGI+h9q6yEkBS
ozYAB26mVLKLhK+ZAT2K42ARNoc1iBBg3SfLLfyBH7ESE8wpbaivOGe63baK0iiW
sd73QZ/TqIsfLScvtsOvrhG9JDmVPA7y7wiOaxSrooo/Go0/1d3QXsw92NYAk4is
H2GUPslLwCZ1YBVLsMQKOL1+AExPD2XQq4zUYpXxvDX5TJtOJLtuUR/Sl31DvpoJ
DE1sOsYP3q+CDDHOU2Foe9EJ0gCj+dpektF8iLe49e8OcnrgPaC7C+6gr2wNiOa8
1gqoUpAQ4nAzSydFFMfitoysO6nReoMACjrO48R/blcRMUFKAOkCjWsxPWKi5XEP
B1lKo1+57CCtvIZBoqLHdi4QnazjTH/XudU1FM0gL8YNidhHlFSAsRAcPXQF+Pvj
oDuXP1XxncFYIK9us+AR1KRbij2pAqoi5/U0isoUCdej2A6v/MJbLkO0aRwSwPdS
6oAKgBpziqRLYhJEmdUuAn7EmCoLaFBslAASnwZu2bFOJG7UKbRj3ukNegxYACej
wWqhzapNeP/hGHVbNYkIny5eAC9eWXAORGBhcYaQOe+OuNJw3dpHlUCA/wzXeBur
OHqiB2W+/1K2XQ79TWrVh1GxXpQqgM1ZQDfULU/NBgNnLWDsvVyuS4oyeQeBJAEg
pfJgKGdAtdmBOGo5HtJg+NYjVDnXAxx2RMBVl+lSyiNX16kTwtXU5NwmDtngKDJz
sfMFbolb80u+EJXaSOszBUgveGNCInT45hoyAbWH8dhBKaCC3MIqgtOKq/vCZMKh
YPCChLm7WHkDDKB4Ek5/17TvCmlICGOyaZ9Ymb88Y0xGQNwjxX11sqwAoJjEq6O5
dgbUW6kft04xMh1GR8q3xR5y6HY913DU4iYh0K52Lq/MVPSQ1hYdJvo1lh9rgI8q
XLGwIaKc7aBcx9oIcYOMNIgPYEWB8+BrhEszkyrB6RV5qXBDgKm7Mb8O+rTofZsG
HZIOceqmosySLVzGJGYzjbOdR0r7xByzvX8pXJAvEZLA8YQe3Y8fo76yuimHyK0S
9YQNvAGcBjgLTMfw1XU6jymvmhd5buYzCXDyvC67XtKnyBgdJtdcfWzbrnFN7O6g
I/1VV/+5ThMbuP+LYXWbCOf2+Li7PIAdMGA78T+OlOngNmF3VAsZrEynRr/TrCAF
IAKTM4QBmR7YvGINeOCDiGhpFkJut6S1McGar7wkxqqvrwPwSXLa8AzVIlRYSBdf
y8qRfn8sDN0zQ4NE4HQjr7bMLLZkVzG1J5tZZklSc3CqhHTAbm+qiv2qY96hqqT2
3FlPUl4eCMAhDPoE1Uw+1aJgqBEhyrjillla2t+lV4gdV614Wdtl5Hs5ep3rvdpQ
NnDmFNOqHYxCl202Wh2vovs7U912w209BzUPT62qJ4u1eYIp4iAycyFqi100ttwH
FjIEz2P2HU7mz7raUAOu52fvr3asDnE7cr+tOqG4WpP9vx2DVBrGJ3r/qa0u8nDY
pA9SH6s0bQ8pUG7S/mswIHYBywAY9AgvL0ovfXxIpmPoLlltA5eCHFI+DiYu/oM/
UfNyHbeB35srvRJCnGuNAjtO+BJcf/pktk3fzhPaohhTWoT24HzXVjikJ/olUGKS
cS2tDrItnyyNb8tTrZX5SsbHEsEr+2TWS3FXFnrk3gVXy6esE3HOv6B5tWlSPh1E
YqEGUKGBc09KdIeMcD+0lPdYOllBAtA9jpMiPiPduaFfk955U5N2aG60LQLrE9QJ
x5p7BM+mXssEJfV70Crspw0szhFAVFXDNym82z7muUSLXsaj/3OTMz9KEgh6tqvp
3f90jd3VeXXamCgBBrfBUoKsykAbATKgvZ/gPjEtS9GFtCS5GGo5n9uhR3+ODXjk
hRv3n/m7adt5dm5XfGzLRnt4BaqMbJ9YV6pLILAbRY/08YsHHcq9BRkwq8DYDy0t
vO0XyiAdwf+PL3xlRQoalOLdiTklZS2QGDJuI6hgxI1qvM/mB+rGsdG/ri1Zr85D
AJlolBpAcME3sfgMNqQu3nb08P1/gyUFSp0Zi9VCQbqxYAWwLJ+/dQCenALAocwc
tyBReakVZSxZW/PgQyPst4x8X5sL5vFlSGqvbEsoWP8+Pazw9apf8SqH5LDbEvgF
19LPAZMXyRJQ24kzus76dWnNufl8RUd95rQsw43BwKbJpVUe7h+9NF1NraHIHgBb
g4tgtnFwo5CeM+yQASoPDkdJT4bicar7nrpsbFs0jo/kZReopm9n4rLcXLUQJyXF
6WEuRZBzArN526yQ1HYG0cedCP00gV6gw55PLkC+1KTMAsKmiV9jgvgBwNwU45Ao
rNyL6ZM0KRdJ/3IZuYeBWeINecA5DS78Z9Ax49FB7ZzwicGvNvmcmGltCU/O3NdB
DglyYh1I27a0NKEcm4WSLuNpTDTPl1OLhjv1+3DTTKZbnbdabg5MXHWpS4rwRsBo
os3OHkUg6C6rZxf93n35K+ILyptYMae6uyxNpx1TTIbrVq3L6V7Kimx+dtzSF4ii
IA9FxwMzkD0+STvYb//z/TKAdyNxLSV6R7aNmQET9ugfo0DCWyR3ojBvqNdDpL5m
bLmLWhi88Iu7COeNUJh1ZBHSH7CzEOYCkMyO021JulCo/VuAogY4kKeePyRVOG12
e1Hf4g/YIubdv7bMScyFKC7jzVTw8xPzcBAlBCX6gg569+WFl+acDAaaKjYAPtg+
9zm3Jm6aTUOdL5IwyKEB05PwmHuT5eUuQAeU8woGp6+VGkdhe+Zyx73J41CIXJUf
C1m+AzN1k0halkRAbdEpRQIsCZfg9ugopEv0JjfRLX4mRlVpYFD51Sj2+ktgPFwk
Tp/P79t/Cm2jV/vdJhMblAsCFr/h0HSj2+CVZ9cLz2/dp9LC0fR/llRyIUywtzuh
HLmMdAzMmS6AjhONyl1bEAseoXpkpnXqTsI9WL0QaHMMPJHWU2oDvD8vIVEbqTf7
UslIfBqyznEiztvdsisAYtvfcRMVzio75YgvFxJqAMEEH/YNZRzdqLxXI911eRXc
QCca9rPm7reSBCttjZ5o7H6gdCg+UL+4A0E3hmANWTiLbboviTLTyPsvhASwceln
eqQsZBLFBtMjKJGlsF0l9/DEGTW34A5P/9+HGotXw/NFnIgnE3vOh9PCMi7f01Mm
Swwuo9x+33VCwm38UNWfvxvFQWGm5gRgzYxMKPFlsNzlT+leMKbjJuTZqjSEXSnm
eU1gCOqYvsQG5tgPbY4o3NWluHBavaTShIoaZ/yadIMT59HAOB6Bwme29JQpn4lw
+vnr263JLB6BH4bIaNxhfLrLHKXUmtC4ExqywOKnNxwf9xtGVXET3KW2ClgaeFhV
M9NTUzJDkCpXbrbjy1txp8Hc/3cK2kN69EkAeAdFrBA6U99AQ7Z1WT63Gaeunq5K
BqhI3lDGXLAoQdVdpeT72r/LBYv7GrQ8IlyhqCSfYs6K8x/hsvX0Z/G5Jup3ss1g
oOBhs4BL16B+Z4njnCbEkwhbQDXRH6NWHt8HtFTN0Ftt/GbR4V2Yg6lcVw3sLozQ
JYQnTIDqNs/Uc2rRfoS64+pSgn7i+4XeCID3nvhyan6ANsAdLNmvk5U3hRrcLPdE
8EC1xiibbdW3HWWpEQRpaAbyQxgR0xelFggk5pE7fq8T3LA1+2L8veSy8qte2YwI
D2u3g5GAScofnXWvM1x3KNeCzFIIpj9636RCSNnjAeF3Zf/C+TSKT/BYi0wmFnXo
Rn8Mox1FAnwGtQuqcP1g+BhfSu2Rnhi9EojMeBX1HxiMqqCL5bHFf0/y6/CNiYi5
N9sp1+kLww8kDkC2dqLfGtswJN+Ql2p997CFDDvS+ygnoU9ToNpcxy7d08Rt/YuQ
drMwuBdpga4yLLxdAHHA5AgkJRDzAAJdN37ZDwSdltipmSzPdEGOLD3seZ3TKA+M
xl9PRyfKXScK4lNlpkzVT63TVDN83B81LnTLizKAUVvlEIvHmhUJK8Jz4ql6C0bQ
k4YyiGFD88GcDpIzn65Alb3vB9/iciTxcLg9L689zuBJT7kMiLBJi8eYYaFWE3pt
ZgiWPqclP0Hfe3O0b32pbJr6TJKL4N7fGOzZtnOHd95G4LmeOkMXrwLxvbnLTSIR
a32Nu/oocNieKypdjRa9oqClOkAcAOos7swF/ZfA2dceXTBmB88FuQjWW7kNrMNp
qL7rFU7GW0PF98fpb83Q9ls5LKWrs7j50B4hOy9DQDd7oT1b6nMF5O7l/vw6hib/
Q4InPvPZeJN24e9EMXJ7uhFDWKGHi0ZBffrA5vh/7HZSj5bb/3OG10nYrkRZxkYx
JHSl4PQVngDJyMQileXbrUmo+Q20zkX91DrO1QuvA0pL1+ZRDsosqceYmIRxTeje
iYj0EaElZNX2cA4KYaPu1lRnAdCehBlsgSRmEt80Yt5K6AAak0NJYIvGsmwQEQ9g
jzGcaH4zqYDQsTWYGR2DYP2COQ4fy0F5yyMD5/HthuPLjjLFCsk81nbnbfgo2+1s
Af7M0HP/v7XAVh/yZNpr1E3FxV3Din9dcz78gf2BaWkZYNuU8Kg0AsG0IFcbD4Oj
UcE9ZW7akJAXf52YF1BcIVN+e1ObLHc3AD3LSaWgisMNSRI+yLOAx+2hunv+v+m6
SY77Mpt6T+3yTQQ0zIr/7JzlwMgM0vbZJPxjB+IN0Rx+QELwxgtEZvMHEfcuArw/
MkwsVkVqBX653Ul+I+FkxBtjxTrkUPjtQgG7zRQBngZveMr5Gce3uACf/0g9oF4x
Ar8Po2kKEJwv2TxrduviHLy4jQRkaG8l7lAQXRHJhQs8dS8D0q0s/3Mz23mEMoKD
plqR8AZKrEJrvMan8GpUsWZFPNCpAsmdvQDYoTBCOpsQaL2UD6FqCm1wG6G/HGaC
84wB8Ch9fh7gEBf7dZrTc7iM1lGyIr49e0khAIMM1lMgKR5F9aQNJ3S+EYHZ9F6p
a6CmBrfEb9NklQEDkCpUlZr85+2foqXZswlNfKpGdFsQtEUT07+IECYrpeyI6BY1
H0y0dAcWcQZbVh6uZ3UI8993+i2lq9p+gmR6jvUdkUBPHxtGGsZNMTW/G9jgNy7n
wXmvon9Mtrq9KQwZh87soyCHb3EDRbCTzOI+fLV+zXm5/sYBh2FVrsMwiJgIebNu
znrammmA5Gi3XojCk4EFH6kRPxyvbjqkf17jiabx2D96Svg5R4lFdEMVqFVmHiIA
Y/Zf1hJdDwqSYUYJA9KY2LhrhVo9bS2Fsy62i0EiqA69py0Lf6rpw8ba7kbaRS1B
G6y+5ENF5aO2KoGH+3fFfxKwKva6nVIq/hXO0F1yChxAmTbsEkLmCXF4NMBgvVa1
Mu1tptPq+GjtWBuCUmyz0z0t5a2DNgjs6dw5Z+kysh2ntou1FDQ008m8mOH9DO//
1crA97+gL5UYJ5GrI4akWD3WD+ZyXwD8VyI/EEB1ER1fQKmJizASbyO7JMojacOf
VAusAVEj5KEkzQOgeIFanmAA2w9MwO6JPstbdSEwj7+ZMIUL+4P6ZX/BMHxBauqg
QlxuXHzs7+uqHdn8GSNq4Znd5iKRZ/0seoxTGpd1Pl38BhPSk5bWyqw+3JZHuz6U
HIPjVH9Eqhq34gnsL6GYsFmZ14nNicgXcN6fX4eZsE+PWlD5YIGMSnNHB3+k244U
N1hc1vKyzBf4vxwX6nNjfU03bsLoH/LN5/hWC6iUk6c+N7Jw7rLVH3PDu1w4+oST
3hsgTK9RZGeh0rX23HWRJbsu20x3hnapnsyWQuoz4taZLfZHBFleIvGCd3U+VzEh
4gmoqCBwO4PGn1Sva+7VzPhM7FoIqAQezui22Rngt0vDYmy2pDCJk6TDZLEaSZkq
G5XXNOgHVr8fojTCT81y214w+LIhTd6RUJ1lUSzh8Ol6uCcB45L77pV78h0z9Z0o
ZOzVUJLy51BgsJTWjUIZakpRG26fN26YJSEzYBGC+0OdBEr1VA4JEio0kISy7uYx
O/oLT/XSLLZQmeqM8IEt944e76ZrN7ruopCLAbm3N0TYMwJyM7UrYmLh6h/ie/rX
dnU4kQEGgowpYj7nm7ZlVIgoh4trsh7h6t9dju9aNsVBOU/qstxZUT1JaCu0b6Sw
bbA1CApc0gt3ltNTjkXuvvjlEVqTPZrrJjjyT1a3H/wvpnIX1zLzoppyYJkcFTET
kFZvRdvKJp8XHXitIuBgrmiPmfy6eyNgQIcQwsT9jXgYkr9tp5ksKh2QEVxKh016
VNTofAzwbPkdz9ZQyLHoqancxaHad2Ra8eEnZQRGaX3bIMuLeJQGb4OYixS87V/B
WqpWS4ZYVK6DnclNrF7+RHAJMR4zB+VsRgSvIfmaIC+QtssAy+x2BGJQIhbNgVw0
Az7cg+6myvgegw+pFaivrk9eTrwhl8CYSz7RUOQE8fUiRuGxBYeYi0mI4ERo+Q4f
llUU0DXAtNIICblYDX3jrQAe3TAHUtlFd6lbatI5dYL5ty8nJ9GeHbI4rkSIFPiA
t6h5nmAuu8mH6BePpmGoXE5kgJQi4BTrp3N1ipXlwvdHsQ9IrzdGC9PxDbak8itQ
u3hPv1yX6aPJVt5i96SFa7/G5j7vpTQVgnf8pHBEeebsvGGs7Q4IDcKqP685oYt5
lqskBgzQ8a9IJUL7pSe0Bm/PWy1bqFXiPuWcsn2DwGrnQRUhor0cJ74E5+OVD1dv
d7bbJ9/wpbsVRfeq6e42q5DBQ3zJ59mEuIv2mE2xUZFe+j3w/HltHvKFvdfEZRVa
u1vCW8AdOOLKzJJ1jlxH3dpzpniZSbkNsiodkXN24+l4wm14mGXdH0sytF9fXkc/
0Bmpqocc78Rz/FTr6OKpDEpMoo35ALJn6zrlQp/euYBuA0q/sOz6GUlixdNRbhAW
H3Jxf1J3ekXcgUgrV15xFnnwiXh6sPmGMrn+725O1GRpfk6uuOaO1Ox32BUOz709
iVREna9UoXRkoNfLpAzyrD/wudgGk+1NiSXr42vW5Fiz93N109dkrLzBh1bUcbU7
8IiWG3O8IE0lyV5ky2O/+i+TBI7cr1oKRZXfaiNir7gvyjeY52vACO7VjH/8iztM
sGJBlg0M/Qf1Kh+LF+GJIwZ8yAleAMjKd0cHaJ2VtJOmD0TaRY+judlgp6pMpDzL
pPR2oNE4BU51kJMWPxj6Faj774TLjTAv2qCZlQEV7GIN7KFsrXMLQTAtiUzlIY9R
9/j45ihPP/ZXj3zjsPhY9yw2exdIijTsw7b9c/hDekExuTGF3ZysMjT8gF8hW+pt
SkM15cY8v4ZbxPwdN3/21aWTvaZTcs3ioLXQKlGsvYWAn9Z3zN1OEh5PU1DHPcD+
7pZekZebNb7VcrBwGpNkm/GIHJznLourF8c0I/vwwXkcYNyLkOcr9Dp5cZ9xrvbS
DwZdIRTOoM4X6p3qfQRetXQ+7Vb5EPrwV/Ri7o6PmrHvtPnVzOZ+mshKlREjoV2h
qSNfYL7NSVhtC1f/D08qvYhc2zI9Iamf7zqmYTswNhdH6iiZ3YQFNWFQWBRdDNno
y21OZ/4wUuPJgoLVY/1+nCeupDOLUlm0zTfj3oGszNVPj21hvFSyZHWdrOaYtSfM
RfVD64SfYJ9ou1wHHwBein8gLg24oSDOXOw4isBMMOpcGTK3U/KhYr4uro5VSLpq
FBgNaA6veAfua07nuTwD14U5Wi3JY6OEslP+CHiOEHcarpKWR/m3HRXPcaQmusLw
Pvqklq1x25/uDH0klZUUOlVVVS9wiGv+GCZ/BQsM1JbKPRlcR9gDUJpSx345p6cM
ldmSKk80/HkPD101dmu9Nd9+uNxUYDpx1rNBQFuXZdZKs9Ye9HSVA+Z+rHh1TCCl
6jKB8VIdQLgP7/zoIzhjFDYH0lQNgHMe5hKGWQ2AVBBz2FZi27UJv/bMTZ7UPgcg
wMWNk5xTeOBD5x+emCX/U372kQBp0EzDT1nrSfjtRoaevJpTpHqE6N4NZv1w32Zq
o1KA6SMZP8XsSU/sAZjTsjZ7k/obdg745TqqGFIwu2SUMITXtQveYiPiCyVFI76f
bgVJxsVsF8n8blYFLTNjthIxktIn7X/z262hUXusqQrSGG57PRagKgGdov5ya1JN
aphY1pP7j0uuaorInWPMWOxL4dZT+p2IPtOB7cNjPYdYtOCJYeq9iGuJDLxLS3u1
1sOYCsj/h7O3aqANHt2pnIlC+CGbEMyuRlsYHoiG6KM2xPKbpNd53+9H/PRxdraW
mrre2ItlDgoFvcDvM+yxt+Lk4+CDozNPvMzzPXQdTmcvJQXdTuAKS/TPV0sJFb+D
UgPZ+0h2hnyhfefe0n+I6Oy4WtVfdYsdU4STd5fWbbdFBcSahLw4YqK7x+jit7c1
VDrprmVagI0eJAqPYI1MbA8uo78y71VZDKsaqhgWin+DvguEpY/a+zWrYnsrh1sJ
+D1ucNgGBJ2geq738NjehQT+VeQF3QqjG4k8SDuJ6kEKzyjQDffx/g12bpKqzsUH
XAxKIFnrQwFdnlivFZbqJeO+BQu3vBCqwB/V8vPGmeY+vBBBwGpdysceqEFfnw90
xv/c2nV58rcYAfOzXX1VXrep+elZERwYPLLcRB/i5uJeHVssmQDkdrMSTm1znBTX
ha8D9qfkujmDnlie8/053e5uZk2YRjUSW0TYwylSUiK0mUxSnoevLSkudkEXxiii
9o7ieuUmqwYMHsfEzd8rYWu775A/g50HPWSMXxQi0tN0UWYnEbJMp1VyjrczFsI+
ppvrmLzoei5fw2R2q6AuI7IRlsd2KL4kYHUKo21UpFqH1vvgWVRgf1Ocem4XbSjG
2y00l/iAzDp4/vRKHnyTmZlyRpgBefCgNgu0jPv3rONn1e9YUZ7AWDD1E/qS3FkS
J9aU3OqP0ku3JUW90o9drbUjkMZqwXBvaJxmxTPzI/Log1/m+H5iv5ChvzZNpO8j
qctXQ5HL2iQnIp5oLRGue0Cm48b9QOxl14x9oty3fIQYEt4wPYSJnKpxnUMxjZRy
RMi6XUBbTjuv1zJi/T98jMTf/xrGdDpYXwxTKLETsSHiJxgstoB+rF/0DfivV8wy
AmPBSVjjr/18v18+k34Gcds2YXw+MmDsA+sobHvT4OdfBSW8/YbDZ9FjtOtKCmUe
CEj8eTIVfHFXbhsPTrcbgNtLqAqxzTyZ+YChboH8G9QZTXHWETaRzjcrgtNeK72Z
DcwxA+OK6588Yacx9vUwj1E3hGujp97xxmO44YUsjGp0sE6FJOujduqjcfKUczWC
6s54XjPr1PafXzT1Dm/5LHA1jWDrSdRHG5zvEqorQ3hQi9eiEVpYFiP7dPuJRJwF
+1/CXBrs8LgF+qh/Lzk8/DLiNrmnEYp5q+75meQS4Thtp17DUIIWlBaWpmq+T8U+
wY9oanxsV9TjYl/KwXicP7mvWxNMspF4xgevxuGbK3eRZcWUMlvK0PY24emIMKGt
LcO4LnEQIuC6q7rvfdolGW6KTFjClsumGShMq1CUN8MsyQl2YQimTx1b4IDAsuuI
yN7GXivNhpm3kU+OX9dwAxaf+HTHAFA9KKqmg3vIT8fnCUNmh3YnzhoDq0Yhaaea
7Q1X7PUxHH2eUN7NUEGLAdk98az/HfQMLR7yhRqHwYgD9WPEO1XHwbSYYUTMh1wg
rNmHVaczuRhEar/u2/wTnTu6rp77leNGzAgH7FQieluZHoeE0eJzc5YcKduSVedy
7fqebTt2tyAb91OYIkUdke63fmoA7AZpPURc/+rVpgXWuAK5AjfbpbJBMKVIRu+C
Divwt8l+LSA+9mkR8PTiZBAB98WcFwELv7Om9burLym2G/S9HfJgrDUQUjuVsKAR
ECycDE1EENjbt4ZagZdkQYodGvP1qpwMXJ2yZqO0GCxnUbBSUT3j+UjbVJaOlF6Y
vUVVnKMw/jA1MqWStGFvAvc2JCuLgfckQOk3wOOMmr2YjQtfBMx7O+vk+DVbc5IL
RORA6SECKjEZMrTpRj+xeajM40Jg9ZfkovXCzVgsTEoziITz7qss+2q2MOEHWI2R
6aObv20H7VxfaI4fdDpUi75r5/xmjjR5iH7kB1SISAHJyGIbu9zushYh8a1PS2al
ye9rFC2eDJT+oT9C9qc8B3DRMmUdraRmTsxiTpKRjfeDP0GY34hNsOWip76Q/O5Y
SHbR4wIyTI7cuj0KwnXE0S1gDENRgkPTVUzBahMZTDEtE5wWuVZELRuxeJobtS2W
3DGi52z+rakJDK+8KGWuswf2CaPyHMkD7HmTAkbh0of6M4Q/OQeNtfiFh1cfJGgU
o18u72u+x/XLB/vZJZWl2rsMCufN9/aKXbxPdgTbELzAdIf7RmljV8md/1CsGQKQ
/zE/3MF9zamVKSqKIcpdTs4tGnziKdWV/oFb+WASZhAX+bLQ1dIndLWp3rjnolOX
GqAXVdEHY1bx/wkmtS6R/W044imbCnttDc587MbjxdORq9jWeeUmckJbwvcU6PJY
DYWVDpQmUUxdNEW9OBS8gcbf1A6IAEFnkP1ipl5bn7blSxQ+4rYBySdPjJwAtKaD
ye54JPCxNSB+LBHHmgjfRPUT44hqvavCXewSXIJNK8gtHGBOnxLE4EDhtXhdSMXj
fNTbD3JfiobI5CqO9VuUqFw0NzjjljwbZspBOwMGXKXjS4RZnb0AW5+jnIBsIo3T
XrGAwLrL3aQLko/H+qhuMMP5RsvNNISjlXpyA5cAyKzhQFOrVuV9HFM28eJ3LJTB
ZXQ9HL+eNIkEf+dsZRR3waE0aLE764UbBhLWT3xuMfIk6KeVaPyUMMbtnN40vR65
y5oFf2v0ToGLUCsEKCoWODVe09cMh6IV0AH8tN7Vnehg+9cziAJ+i8YgEzfKGaq5
WXSSgkvzBbhBxh/fxgIW7HxDGizududbf5eIONFSzRihVVqYOKkYLHtQtflufrvD
w9fV1ieIGmG6061mpYIBuxitdh2pi2aZ6T1Zmr1x5POLfcGUrOL+xU0tZYyHariz
IsBoTiVE5fIkzNcOGFXUDCGkKP00pyPHrlfzMZ0ECB6QprgPD0kSMmlJXgQhiNb2
HC8Holk5GI5F8Dw5Fg+caDX8OuGCxY0sVZBuAz3fnHn6gKyeK0Mf/2pKi3/kOIRR
VevIU0c9s00nh8x7k7rnO4aj1DCOgD/i6zNRkR499tL+mpDq8Y9ktwnnKhokXUvI
mqL0KTxJ8c1w4SD2QYikl5Bg2wwy9D4405swtKJvWfIi2suVjuKbxTTpmksEsDHK
vv4hY4cNsO/maPzAhdQ2WWnnuSzOK9OT7xhxJ6Fk1eHDnDCzXlwAiJ13B6q5ZMj6
CMThibuILWbTDF6RmO5meJPDcoMrUAXpDFpwkU+JVUEXh+LXoyqMzOG2edmP13zf
xt/4h2I0wzNLox631n2CKQpM5VMete/KWYq7RImZagteXs2FPqmmDcT7zleV+MOI
5rb17arsvzqrmpAuvn5xwZ0Z23Jcmax7nXK56RzdEM0OX50Msi5MNtVsNqboJXfW
T0Njsa6TG5d3ZxodBct6dseuXWJ/oYxDJNeXULIAF3OjieyQYqsK38PU/PpW7LNw
S76sIjOcqQoNkJ8jbg62bn1D4vnqqsLDaZNAbT2rFbtZzgAdAUt7LYZMRWxDBUcA
58ciRaNpdN1jYVqAa0HgOVY0sggsFgFX59Qg3pYNMSuscS41dq60VQrSQtflHaD6
bxOWIkgyR0vmv4oFCZhiZI19m96FvhHNkcv5IKxfWn8EYEBBzS4Y9LH4HItRA76K
9K6bHfKFt/k6CB4NgSL/Jga0TW6eNvAypLmo6CENz3HFFAiT/iFc+1x5Rm2RT9Dr
0W7+z2dCCpP+nHZEHLUC3i9tx/hwH3c3jMIbNdGdKaLfx/UwJQrp2wV0EwQdRNlJ
FyhhLfVwrsoBazYmyUK1x8cDj4d+UswP/J8MuEff6gB3MssXH+NZx7VHghYG2GAi
Ld/Yjm9sWbpbLH0QFtSrbf9m6Ud1uJYgSVzeqh/4Mb8FS4w2eZ3gaB1LSZLz+63P
LfSC7yq4ndtv3vPTs5FSfR64jWu+nuB5aH6WwKgzumNLxtCSOCngacHXnmEYSyLP
hsvKQVfLllI8DBqJfZAw13Bfk/i0u9qIkhsJaIi76Y9n+J8qORMrub+j1zKY9Z/k
KJrL9ZBosu4rDraTCG0KOCQJcEgq+aJnexsgUXp5uj7q2ABdu76tMA6pePct/KWQ
Ue173lxioXkQVIrYtKL5UPRcZ08vFgJYvxvbykFOx2L+H6mC8W1kRVbsncfAEiEm
n0h4ByuFOk3rMDIj5QJUhWf+1ZhDMZTkGlOoM9kv2dDukHHM0nYGkxfiZGqRDUEW
MPiuuvmMII7q8MGfngjqZeVTPIPW2wCD7wmVf4Z+UMQoRu1U/XhuGDfRF3qO9qnD
JwxkTtPfAZCUTrjfNmhGpaQNR3Mn480aLrX4Kx418nCqxECVKj4bFpU5No6e0+y2
wpUL3XjE1xPDK12OmBKdcyEibXp7jIygAd6RucD82OYTOT057jImYocCmzVvljbZ
SMLRSG5oYaKOgPDaJTGG1UbmmyiA/ZDux5lfao+uzk/QxEJ+O8m0+sLi0DkroBzL
Lq2eCA2ReLbaV49aiOMfaQXKjxufRwrIAzz43ddIT5+/GRSGhJCsio6WBhZeLO+R
JjNEztl/02e6iUXklFQPpAAFW0cv6tmm1Ooxya9TU3sZ+xyAwFiDtX5OSmAkR0OR
KviaSZ9Khl2WIbZ1fkUAUfNNq5/VWILOKn3e2kJPkguxlSmddwuwzepJUBcS6lFL
auVDfIY+3oNsolrNsNEwaxSB6k8h3P3jGatkS7J5aBpb49CfZ5ffyoMK0pGkbqBd
VLI05ePs+9H4iJ0n/Y2VpPALjjMj76QX3MWjvTFD1xVMxRfQvWMEFyIewsXuPkQX
p7LFZ+yS7XtW1td4w2HAGeOFvRRiLYgiNExuWqHlgfckiiPRryG9sD+9QQR0zjDL
+dDg08t/rMlm4mWe2er5dvP3kIKzTTCdF3SXKnBOJF/kJyyASGhrPe1TvFMzI1BT
H9juyoDGPxIfXNORPqhgKflPRz3IfFAWot1ZrG/C5vvZ6UhEPerkgXh7wB6tUSRN
aDxZcXGO4TR9h/DX383qap0TgxvkuR7F3DcW4ZY55ZhWD9k7xr19bJyjNKrL1EYE
PCSt6Pi7DHtSM1YHM9lDwiFQCwWLA+jXZk77Hhr/g3mqvFAWDvFmhRKWSYeX8MaW
VMbm8eLw1D3SbwOS+O5UPsWbxzHlmNfwCxu+hsFWYHF3G9eTl5vH2RfulCUgL9NT
CajTSOxywVkbAvLWv/gsoCwc2tE9KqckoU5BH/8K7zAqUPjFoX2xCnFzmy6FlrRu
sNZY5XW46re3Jt8gOS8mcPpl39HjO9XWehFIPnPOfN0VeVobve0mgi00Bqz4yfNz
VQv9UVAixGYgucs8OA626W4jntgVI2NsJVSiYUtLcFb2KzividvK8PKVQ/a6CwFm
uPbzQi/j27MN+ayijggWuEv0ozUJNGuKlHsiCsp8lrrYXk9nTfGSDuVur0xtzcrm
VM7Ls4biVC+eNAwdLtSrLTy8KoL8cm/ReUp8oSAKKerhYoxZ6494F4l1GaWHY++G
wMRCGARgTSmjP2Q8/Hjs9q0WuYjWShfUpXERkVchClOPBk4oQ2mfRMj8qGa2sXqp
HGQRJ7+awOFjWFRHsxYnM0CeXVnM4FebUHE88LaKzMNVEkJGnc5bQSGK/5fgjuIS
UroQs81SLCHB+1Am01LMARnXhcE65XZfgODjftLa1udbPIN/OOKA9y8Yw+sAWk1D
wUezXNnnYKpasQIMiHl6fnW+d9s5m03V7dbxHwZZYW2lT9jhUv5qDKVE8W+uIE2r
/vTv5taY63rW+hgxBVaRoaUQGrfyGMPT8/2Dz/GBQQQSf6xFsKNf+GsLp9r1t+jc
n2AiMmUQfa5zjh1D7qMeTHhw7yjWk3NgwLvJBQfAS67lYR5jX+qewsRc/zjFdAFO
+zGZzNwurDIUrRLmuigfsWDQOqa/OL7wVyt9W+KQMpxI8E8x6WBrhRJK4f4l+tVh
jJ7wuBaNUBmhe50lGct82nsdefkUgQyxPysyQIyhcfrzaCcGmX+5Sps4qV0UXe/J
oh1VYaPhYmQWZnd2dQnwPeEHHss9h56MkpcrSl3vDb/M11S/KMW6L6L5c6Rh+5LO
+k+mRbaKsBrbpbLFLJvb0ZOFf8M6CF6U7AV1cnjqPXxatnUJWSLUSBu1A1V7UzBk
L0s6NsQdjF8edvB6Nxv2q4WI9oIPvfyWphXu/2yU6PoyCNLd3ittUmhJYZJ6kUSR
JAgrsgh7tWL2UEcLuToRVLm3gTnEgF2ayL7aAcg2dNmQ7rYlGRtmotVWlKSIM71D
PMLhqsMeGEeFzlyLb0Z6SCAhT8CUA3cMVEFXqn7geZ/zSwtmKyEd+vYfULlaLRgB
m0NJg0lMwhY6EYyA75yxIPG7e0d57jy/k9TjeDdUktd+Wjg+ADThDfkCpiwZv80L
QTkHif8ZqaTMrRRsAonJrNy7DbU9hnHJKm6NsSRyaTnLM9/FCoE9Lzswgn5KY3IB
3LVo31yfkplIm4CEL496jyXtljSxXY5oRpAO2R1a9VKU231RDfIpU5pg0l+7ISzq
p4dzFc1SJqbiSPHjjMfYQ8NDFHnEDTVihntZ/KCJoIRXvdX52aIx9eWddBTFOXCg
Ap7gNI/On3UyvLvd/tOADfo9xQPQGuSMWEQC4umjYxVXWvDCqN2mz2RdLHtFJ41S
9fQQZCvxI8veYOaepibceVbkJm4tAs6Dq16mPQ4n2z7fHXW3cyZWKw7blMiDg5o2
s/EE9IcZKpylgPZymhcCuy6y8kqsl6BFaQ1zaP4u1nPNPXL1QvjTKWU84J0PYEZc
GMpsdrypW6T6AE2S442ilggNq+J6ZBQc7okgTWs4elFl1qk6akBBxJEMEY+RjkxW
KDk/EA41U4othyMXvYgPmVKrX05QE7CItAyV2Cc9c2Tmr64VJ/C4maXsRR9PZ8ot
+n4pnhe/oUBDw7v9blkB1px7VWIfqdI3Mi4SxsrmixEth4m1K16ZPYKDSG21XT6m
EitWFbI2bzMwQW8kLsbF+mWlr+Fok/yv5habI5QqmvzDpEDjBDnuupLLYSoxR45T
bwz1bN0DIYbsyQt8s6t7CSCWo3JqKAqC8QAk7r14byUBgVQr0eTz3WRPmxe4EFaI
vrpRqUx1Cq26bDnr95VOsQRL03pAbc480YJsXf9QRpXg3aFO56r8riJW2ZZWc4E3
NkCznsyG5LS2sijqgAJX6zW70BhDwip0/o6UMPcRHoufK9T++FD4K1QmlmLegFNy
jqZcAHuwxkDpABAt04oRWGlxqZ9H910yMl/Vu7IaUijQrn9f0k1p+5hooYR9B1RQ
WgRelAoowRqzdM9apdRpPQqeAIp6sWm3rZiQgQpzdcxiXe4issclQ8yox4WwZy1M
M8J8Bu6JFj2QLEnknwxVWuyG9edKDw7GczmIbnamgZncfcvyrpT9hVwcnMbB4/TM
ioYcDvERnzTGYBdMTFUtDm5XooCkAG2HaY1hyh4AdDprTxAKTOZx//Sf86LsaoD9
K5PcU7+TJhXFYPH9CdExhkP5JXR6lGgA5xOFPAIvj2w/w4f5EofzhCnhwwyLoZ6k
2Yo+XrVfXEn5tH1Ah/96oC2NtmtswSU25bhHM5TF1stgqYZQTnJjlTWP94E01T/q
Umo/5vSfKngIpiQmRsFynDvf0laFoy4H4h3Wi3O43+I7hC4t6RTqvvBfJ7n5opCq
AjJWPReFdsl8ABeHGlnXstMD9nQVWx0hOq0VXa0b1IQaFg9QDm1Z3e+lWb7EghON
fmnH2YMMFzm5co4gRsTuUbQ1AiNAYkNYSv9UkEMR7WKrzQeLdyh4JsRoESv1Tdbs
gMubxUy/Hkl36ocTKAQn8H7glIgIQmH8kirptRWKtjdIHvmS8t3Lj9+L4POKCFSF
71l26ZZXFm/oaMOGYZe52rAerh1KkwYd0OB7z8sFLXTLoo9U4Q/RIbEICcqA1hiV
WTdbejuclzSlyWw+1HqPO7YyzNH4X9m3WoaMl+gjo12QCdpoOyFDqUxO+xrNvZVw
PnYGLx6m4DzXKpef5pQIW9nrUrnvbhyZtv9R5wOb2T5K6B1QjV5JyxhTv+XEJGXp
Iz5/1nr3ibny/4WxoAfIUvHQ+9vRps/yXVuJ93mVHCUPhmenyw89gnC0POY7USOO
iWwGtt5Au6PIEZiwgtfDNVVenGHpFOnxjSvkxAqbkIx8pcwJ5RLU81pQJeW/wNcK
S4hNeqirOHM/DacSFnWzrodZTpQjtqnx7jhBoNmeSWOab3vxxdKWUkderwIzNt5K
LNEcoYIyGIOqtYDNS5Cx0EOKN4WhrtixVGm5smyDvWzSb+gBu44E4+yAcjcpKqgU
G6Fv36WKihasbKFWQE/t5nt8f/n47YxL0A9qHuxuDBjVSMrwFavMgRwApC20OYyw
KJZjKnqHoA4b7Zdg+B6EFygfkMkmNDfs8gvpW4frRPBETWE2zG8776AWt8yIop/h
7twDcQubrUqEj7SnI2/8sX3CGnx9BO+7DthbC/dPRIkvJb8RmunKs95lb7MbmEI8
/mEyypDG0+fYI+Ep9zSz9a8ZH5CXN4WP7ptkgAkm9oW03gXb2ym8CogvvW8/Y6LK
VKdRUUyuLReUqqC6phzw927RGr4iDjDaXEknI1fngMWQ8vD4SBO02V9Xx862cRY5
/Sa7IHGUdR7eISAQmZ9shcI6DgP/GjGC9PEA1XdNwsn+kD29HaLVwbeiuelB98PH
AfQCPkheAfborfRvK2dmL3rB5KPFpnr4sHbbwYTkflNBPiqc4iC7j9ZE7FB770h3
ZV20AHlufc0mA8DFCjiOzUwhcaYF4zER70JFYfcQ2X81R1/oUQwqroG5BCgKV/mv
89U5IKPxkv7o0+vYCwZD4feg5u0RlctbBwL4J7ByH4RAS1jL6UNGKk1TOspNuoui
DoY1Rr29dznA+Pm675k6rQNN771Ivz3H0CMTSdEGnySlnsjEwr5+JhsO+CK5la03
8TJC5S6E6Ewg71mtq96gpvHS0BMO2TZsGaS3AII8q+47Uc3dVvf6YczBDsgPeFrN
9O+3UFogonvTicN4CtNrHr4rofrxNKMIlDLf5js6xEiNvdrsDN666jppjhQFUKSO
nbHhWuWbXE7Km8b6GfDOQp/WztkhmAm92vB93H/0M3z0IgUxC1lcEGg4ZFeh/TMu
mq5Xg9n1X7GF+zvmcOLticrljLCSJ/myno8tVIepI1jBxFCUu0Namzj2ow4XoLA7
xkwZ+d1EZmZWCnH5ko+dBRB3mRUqvfcTF2t7Y3K0vmP4Avk2SKpRLd5GDrPWyDFv
DW3vgRPTh2xW4nrmyrx913slFewq0wGn1v1DP6ZV0PKR1F6/J10A9PwX6drZIGdV
Qnbb9WGznKZoEHUAzZxae1kNYahklx6x59SGVftSvH/Ul/IMKaz59f9591k0ZpuQ
AHr8myt0JorYagI8FlSMdzX7HC8PcA+uPIaF+G4IwQ2Vht8jiOPLGSEgiqraRAjQ
4pQchIws6pldx5f/DvSzQy1Y5COnaJ86qJnNkzWf2DZHgnWwWg3h5Yx1xdpo8utk
51vVoAg463IAe4RsVKZHzvOdMSe0nrRKB1mZ51J9GvsKyiYB8Z85Z4IUqvMFkmpR
1o8JPxyC4+VqsqRPHwk8oYuNPEX/6YQrdvCBwJwLYOgQ5v2qlN72Z6k4M32VHkdv
sODf0P4jKy9k0WGjswz7Iu5WPOTcfww7yrMY9MLdz2u/ADeaphpbEUYu0hCnDuM2
W2jkr24X8qkWsK3R5MEnx1tHVJecvRy6wgpfD+Ds0bzNlqk/a8d/rjkpYs1Lf4dE
XpdIMo1uLzs9cAElsC09gYik7YKGt97n/eqPcgaIaPNV2qQEOwhUXeXYbb5GRkn/
JXpi3wiDOWkgsEnE/bAfKQV7b9Uva2KACnmX7jDld5T7ldQmfC0SHAPP/kKdbWzy
RXql0heGledPX2z5abJyokjDH5CL4ENPHG2prVwgqvXcxNAOdKw781qrPWfQazAX
Squ0bztWEhGBTUegw7dYiRmXRx/zSZqD44Ah8BD34frrr9/0Okz+mO7wz9XwDkC8
t9u6WWnSnyDKGbP5nCXQm5xaFKspT+sLv8+bgW/pUQOX5HJiczC75o2KrotvVMOJ
y9XIw9ooCWP6Zj7Ee0wQ+ySUNF/bDlXJ+e9MNqeziLXwQdu0x2ArfkoqFl3XNwD9
MphYCspQGgdxjOqwpbNKvt+LWBjDJouCpAFqTZWV9MoA8zo2q+l5bFN95IJPOyll
yP6jxQSgAKaLf3cRKNmfUAERfB5QKE+pDCbblCK0nZQeW5/Dn/fcQSS//0UhAHSG
slGjupFEBpGJJtf0s4TW52hJah2F5JT+iVhL33Nj4sQho8F2zLS8JxBFI/4Hb4QG
3Bs+DX2H8/9POq1F59tDEdhzUXLKjm1BwmoXy183F5V88OnqjzjIyK9O7XKbqA9A
KtyffWPISKH5tnUednolzF+6Kjcq+r/vvaDQ3hKptQ2ZwC4478QjrLrcQuUxZ6AL
alNZbmlakq+NjZlzF0bm3q5hnLI9JHKFAM5VMzxwDR3KlEFU0uyt1s4oajZP7AwW
77oJl6rp6woQYAIAnOWJMyZSKaw8rcVsF8Mn90+Lm3BvnEeGZqybD7/7oNquJkOj
j0bZMNDJE2ghM1BFOLwPuJ+lpRZBpBEL3vYgOOwDBNGOQIT7MI66A2Ce4KoMR7HI
g5SiwNH3ofrFEaiKj71j0Q/tRQ9csiWRdUIbgTKL/vfh6eKwmtc9FlFAZ3B7ipGt
HJuwCONNG7tzL/st2Fm/+dfogGZ1FrlnqzYPcOWDfCVbK+KuGuC8/o5u0RfmWPpr
moG1LlcIcVCaqtNghOX8x4ufL1ElcH2osyuJSaUJys9FS1tw8Dlhvx4k0XiQcnsG
45/HRNgHw2SinMGl2u1cAPH5yzFfJfV4LWXoNh5+kq/eIk7E/s9qnjHrUPpUnlSz
+WfZgA6PqxNq+BwIVjV22cn0iwoL9vah1n2/JMYEC5BFZ1Hmjvqgp+s2PT8+FVk/
CbhwvqM4XfhnzK4LgQ8/5NfXtpqoQABDlixkEgkOL+s3t3kAdADKUCTPOapPz7iE
Qccb6W/TLa32rJO/IPelcm2lZa057W79agkPJBNAEmsF5w64UCL4UV4f748QH0Cy
o5elvAz1/bpntvYjSD4N9kK8ntVlOwDRE9bly++xubW7l9VKic+D2HsZPzjbP4vX
iKuDiGBXCoPXeilzBEG3oC+X3rBR2mzChhrMwAWC0kn5i6cfDgtCvTTe6aPawyO0
st8gZW8261g/CTCSj9FjhziSjxGtxEilS7APttaok7Mtd5KLkqJKws03Al8RQ2va
vcCpyq6NU5yaY5kc/2oQ2jZeZGwN2pOAnkkL3zWmEx0FEIcpsOwsFvpHz3uNPbVZ
IcwcIESmZmudu1tWw+qoPXCfWghfD9rTB9uZGzE04H1BtMxMeeecp4UVVUDl7kIG
+JeSVoPW0vUqBtxtBeTXE6WDY2hXedlpSoAjTU93eVF/46NKzlSr3HrDzACTJxoC
7oi1HGuGW4BxaKLVXFRrOzhae7xfPiDt5tIu2bhAod9EwQvk566PAvTRnJx6rGg2
p6FBsICLwMRvO+Ks8TS3hBqlLOBOIJbUbNreMebLdubTEVvyl8KlZ3wKg4Zh2kze
FOzdfx964yFWrAXK1JFBI+4hJVueEHRY4qyAw48OygY5HQxm0db+r3uYqnyYe9bP
xiTT8WlL3FWaqlmy2yQ33oZEOrDxs0dnLofnGesz5iRsZC2GEUYXfPK7rzlHSg2E
WK5BK3X3cWA9fm1E7RBgisJoUtgrZ3RYy6sCRydpHilzu7gk1uzE1i1jpwT6jSrh
wbgaeqBtVla5hUTeDSxzsdTNZvG2ofqylqQRTWXHIqsJzcNZdocI2oxrED8AmYTc
XlcCALpvHpP0V7xHq9kXr4rHpB7BysB1VUU+3mOAnS/KqsSd08lofALiMUIBePsV
nI2oj15JSyob/enHaHjK2e0EC6ulJeN2eaMpMm6lHyXwgF28HjR0tj4dJrRcqQIJ
l9CXhe48/UVbHqajzbHOpA0/TcHST//w5RcGTgnW5IjwHztxobjRa7tq6LHt6htJ
Eomwe9u26VDrKX2nnLgyQCx3cF6RQHEWqSvSgPeoAEEVF48qqnnR3vUojhEPIn7U
X3RyZx7b4InDqj7ZFGXdq6Ykchy5oRtJjUPDE9N5Y2vhciKq2vKCIITxjVzDjL4w
W03fJ+0GGGMVjdusZP0ZZtTexPY7n9zkGQ8tCQtSv8JZ50tHcZ/vqv+qrDrYg2i2
4ZyPkTtCL6gJqnyAfOvTjnOF6i5O0KxAkee6N6yNiSabub4PO/LXOLoqrhx/x06f
bnG/rXoWEe8n8Vw245XhZ67TPkTGCYKr56KwIc1CZsLfmlL7wv02c6cQXN2wuUQA
yVavaXgwk+XccPhfTW67TieDnqZXdIBVsaYmZqg6X82OMOEko4mLCNoHv1Zg+Fy+
55OvcSbxmMTQgTMkMz3Xmpzgga8v3Dn5piiE2YPhSEZ7Onr6/YH0cuHMYSzaHw7k
NgUtguHql/Z48X2AVgvuj/ZzzZX2rtThpuyw7QdOlHwqiRP267d5IWKqWV7GpKS1
wGzBGrZUeDR/Fo8665+3uP3SY8RmRzkSzSf6fFSfJs2vRlRBb+K2om1DlPEyrKqw
/73pHCY4pFWYi0Rskh3CmVsiKU9GWXDob16LGcpD0+mWUb6LGBdENEsMWKWvmYtL
4gxOnrSQ933HSj5agwRHYiUuMdkeZkWEGHz6nzmnokQNPWa75AE5afpLz0+QHQeg
lGQ9vs20+3oYIgByjNjh2f5DehH8BJ67Zel2C0/AahZHgRdIIqrw2cmYIVLVNzOu
mnn6QPfJWSzSbc9Vp5lY2qwdjqeQvtXcC2ObegpZLAMUBDsJHRlVf0YP6n4LI0E6
E/yW0iynfKpCe0eo60FZX+cA1NnI+EOLjfI3WbmexXrFXGN+hVx9YAGTGVJeJzfN
ZSmC2gbRUz4vBMRImsGU0+a9E9EZHvDLnXlbxvpy0X5+97fWZOQqCvvIlQwc46f7
QFJltfoouuUXqKBaq92+tLttMPVoYYVRrTOAegN9EpVs+slQ5U5c0B2wb60EQ2wo
0yXMDBmg/czUdLfgP5kWofA+oxX3ZrHKU6YBQVw/k9jyp8UxBySiFCuYXRVPAZaX
opR8QRa2pdHl92Kl7LhY1FEqpH0D7LekPzSSIQkyJC2Y0POf0epCYNy4CLlcxhXv
VI3Gk0BgZ8/jjP58fGzGgTfOwvWoP2GswSVLWfVXSyM3A74FfRlNhuAXsX06YO3y
RrgoovT80PFr4nphziycpiQA/y2rZXgP5KrH0ZhiI9EcZGx1Sc02YiniU+W5sOh0
w7zN243UgCWcGeIRb/aqHJLZdGMIygcWCvGDDMsIm5v4nszv1XFdc4rYi978yUCr
JIsJw6opyFQEwQBnMUxU0plGhfw188ZFMWdMNDOcBVPBLMt4asNMqUX6HsGjKgH4
ZhkxEtDKK0Y9WadOYrPDm7YfEIxr8a3wMAS0sH/cSck27xkF6Gz3uQLkPZ32ppmG
8rcKCjrbdIyQSgNbFgHRDkYuCJuB+2s2+Pp7G02H06ZotWMIWV1jRYDDokNoZDgY
ZVnx9VTvMM+ks62scnyLp8FfTMZi9pAI0MMnpq1t23H1TScTCCOAzcsItElnlLIR
VCR34QURmAtXa4W/5IKjBfsIqicK4+fp2BVugZmmYjqGtXQaESLPHuk58UcyDXKl
ASVI/tmP8vfqINyZyGfQ865aBxaDx4zsijnfNEXwGvltlgoDRpB7ZAoeQnI9mlCt
z+OxPNEc2zZrdK4F3g2LH7OTivFQFM9by6WpDbAfLBShv0jHQScTvZnGcVm2YUdG
MjkbcJymenrjwTTb2rWiY1C9Pe4u3JZhqg3VdV6U8gnVw9MRQf9e+8dBcz9m0teq
50+0/LvOnjE3JXYHugjz007WnSMRTNDsnvrRLZ8T26XSS3/IGINqFV/yalOb4qox
ifeQ4D8lftP9I1F29pDpHN8ngwXUHvXXQwpONIRn5FwwDZvLps2+CZRP7k9YJU1R
XzIloyfFCt/JJ0M/fnrQ7lsAGQ4KO7qGASYxb/0HwvjC2wAJteD+pNvPRDKpa2yP
pb2ZwdQXO3i6kwgToqMw1MhdeFgb04pEnNNNBlIR4wyDe/4YHgbya9oHAYzy7nJR
47YKUhiIgSa/zeE9ZVxMIDhr4STWqyiiL0HW3DF4Vm+d1gGgL6/XxcG8oYen3Ltq
zFfHRxzcJcpyKV0rIoYopf62IgOhVJBCevXggOG1VLgDTMXptQrm2tdg2tT/mHh0
CZJuPFaobrCo13chFfxhy75ui+7fI+1VGuZajjbGUxLDf6H1OtzgxiwUW/CELRAm
v7Wf0+nWROrCwH/S9vW+GyRADydR9y4PpD4fPR58gKKlRWMNsIA+9dsSJHxaMbuM
GLsj8juDJITrbIE6hPFKPVQbrWiVLvaT0uSZwAAxrnE6pf9SKcSrLSiJrrQ2frZk
Y2R1/3cTMCAIwkgDZbdwm5CkcP0we46jLyiLxkTbP05Ri+KPqFFQoFll+raXITB5
DA0ZRITI5vtu6JGiWbDTpLswqUz07G0zNB/s2JyrH8j+GRrsQwfk02i0irse8X1C
mYjwK3GLS57CEiV2MKq6NGH9mgyHBQdEo3a9R8ACNDtT+KujTTU7RUIkfyAqG4KK
W+CxN7kB94DroRZONW8VwsiK3J3NRAStRfMr0/LECgImPUBAKKPXZhP1lFsBaEGs
4CR+pgzRT13kOxM4ZP7xxtMimPwaPAkbHAsF/VqPXl7juzQF5TItcFyzY32E4gSU
F6QCimioQkYWRA6B3Qgjp/RG3RvMcMvFzmOAQci4zUI+ZFvZYpNVV/nvz2o+1vIQ
itW5AVsvSqugkJgezoMjxqNOVS7tU5AOETZFPwzwfRMABRoQJfOo9H5xcE5O3OuE
7IhWX3pinTxNVYKnTqDeIPaxNlK9vgmXwzzCxNbvIaAKOHQWAWyZPZhgvh8032d6
kk32OH/qbf/yeyVUNNrsF2Vxj0/kO8rFSCBXNYN6P/yp5xaCgJVc5gp4LcP6n/e1
R2FT7xeikkx5jg0/IuFfei8FzNlychg7ippedc6/x2UfPRVgBuBgVLm7iD5Tcmc5
MUtexzVfQURDEE/FQPHLI7wVQVcGgvGDrchdRx8mLVrS7qetRocLUagvRr9vOq1L
JlI7A1bn6CeXICrCSnJMMKhIa/aP3FHDOWMn8h/GNEREe9KuBDsjtMfhrbXSjw2n
GV40BwFVazuWFWtbjflbLTkNDW7WGiUQ2sIPrTaQ0WzY7BGLg3m0SVt92KtS94+2
CtlFE5wgHjGEsJsUhVZ5WZFztcVLWOl3I601aViDdGRcYqBtsnMApBxRMgg3F3KY
8oPQfN8QYUQTG7kPG9LJdkO/mxdyn4qL03JyPwSIxfRjmC8ooNrU1Lyieo+Ehev2
RK7HgXpozoFI1N0f6WiKcXqUoh1uyBuAsIe1Fte18HPjqIdlZ7UVGMUSAKTvQZvU
sDuj4/zRrNbFgVfoL0Q1Uf6GfnfxCQYVV1eAQxp+88uzkI1/mS3GN0eYD11M+QNJ
k2WYdrKOOXJOMgGGGGy7eSzol1aZBYCVeqfEoRZZYkU47GBlPHpJxfyJgZPeG58L
XDIoNgfdcAhKH72wDJq9Q27CCRiB2PhBG/NVaP72y5eErMujzxntKyjdBpnsC6zX
P4dZzb6SvC4HFlAuF4MLrcGIatBEXmWdTlRuftPg3Wv3rUPARxpEz0Va+i44ExBR
ZJV0w8tsSfkQ5G3XEJiVzp0W0iO9aC9Zl2o3mCOzpWAm4W2ZMNu6aAf4sIgyw62j
CiaLtrQQ9PV7ee0xJh6yPn4ygt7DlbdByhoPQJo7DHkdMfM59PvZzThhkqgvDVLT
J70fAHPzj9fG6Pr8nICH0qX/KXkq0ybcMnrPDIZrRGe4CQH2B7UpnokI7IZ9pVC9
te0ob/mrQVMa+gKL8iimYBR/LepG/yvcwCT/XHmzLQKoT9JNb3hYtAzOtOeJS68L
nvzY0M4HQyXib/QR/UF4eTm7Po1DzBPKPLQVYdm4uP5IIAF/s0zR4ofR59byta4I
CFrIxprZd1AjGOC+lZhymb8QXPYJJG5Tj5fHk7h0n85nRej/XAkqBagBItVd9lZO
aAELbZxHO8HeRFuG7fe2jwFnref8NLpMAfjtyTyODJN8ffgZQNka4fzlhDdRMLKM
UTjF5A8EsHYtBi389ElxgCWs56LwTvcqbry6b3vTc802n99ngy/WMFOYAbO1G4Za
V096SGprLNTfNecyHKLabgVMWnrfRC9AWGHx6tjZ4sejvmsRGazCetlDuG9CEEJ+
if/Mctb1GF9iazxCBY6Xv/53XvnBcL0LVw6Cycx9uDaBgP67Ak0fXH8UNrOZrx1b
GbFQFTwkPyPWMLWXb/pnE0aIF1mCjHvlOxDOJYSECoMQhZz8vU9L9l7IAT+vRWCv
gfEhVPI78M/8Lqr9fSiCiaLWatp9V8u3cPsTdFyhZ7GLFdPKRerGstjIHtZLNwJQ
KZ7eVPz6n49dLMzzrTXIXfyu8G5OuG7ZwiVT6RWSjPWaffJQwmR2vG2rah+b/4oO
g6WIxraC+g4ZS61agOSvJmRQxMH7aJ8sno3hKBl+5YJl2sVWCtoY0S4h7q9up6wy
u5eQErhMFecM+aE2vDHrbmxxeOn1ATEKB/vBoNWZNpsw3FjoBxCC1aQvJ/FfSeu5
C7mKJZX/H5ITLcUPhIJWpiN89ufK9FxIvKvSM5ncfY/GDIRXjKF3gWbLysKuwxYp
4l4qu5YSy+BHjbMt7ZOAVFWjY7Pg1EULosgX2dyJb5f0Bu9IiolvphL+TycZPsd9
bi5yVlvdLuHNFZbNaySwhNgZs/ISslLa8tav1b9kh5ivoDs4KH25L6MmmtTNoFWn
C6u6eb/SUj8XjIHjDQMd3eEZpS3LQ9JiWxVyyLfnMmhoTqB/V/2B/KF91tb3s04e
+VXIH6Gx2pAkyIJsHSwsSyoSx1BzTlEF/iyQGrvS7fP+Mir7mM/rl/N0sO95Bg6f
E+sJT85ufQwsm7TDdvh8qhqzbk57kWtN805ZfhlqCurTtZWm5mkOs/UPv6+15Jnq
fpHgL0NEsEQxe07sUKCXAMTrpOH2RhKtUGV/n3mMKwLBsA0E3lz4o+A78a68PRBr
LO+UsMv/QwY9XKw4Dbks+mPJUMuvMkH3yPdfOvShq0+BZuRf7jrSbaexlevxi2Qv
zw6ax9axdQrCU4bO23/kxkJ7YPX3Wyp8RIveCHOgxeVv2rl5qJkUQeQRP4wAnHqt
eQLXZpu4GVOfIzJVsMlrLzCelmFyJAU85zIwCeijLgRHlW0XNm7NxXBrbn+5xS3B
009n4jKjIR7m8LOcwNytUa5E2KJBGwcjWU9ZxqHshSRRrEf5LN5SVw7ApPQsqh6w
OAnNKqj5higH4eI3RaVCb3asy3iU8Y3eEYIlTulIFpiv0BZYfcQ7H1XkgFl7s0Mw
9dIXWhGkSsFp/EAVdrCsm+00mAjJwXJkM5FzGYGXkjqOqHfWyQVe7BOoSN4BV7u/
eenzskwZl4aksgwbDS26BNoe3UmyS2TuaeiEOqLVJYthp9bG+EVCkc7SyNsQCmC/
CyTy6Xyn05sbcV6hiXjPgCXyW107rZ2EWbNfMlBZ2gSKuw8jxXO6edZ5MynGOUnN
Z+dqcf6L7gb2StkrbjbP0mUwIUuyZLyscmxPJXAj2vzmyN95Vku4y8yTXoNSRzyU
yWIplPBwvfxjT834ygBCg8bCk3vUyDaG+pAl/dM7R6n3W1d1hUPaur0dxrsmNlGi
uLHoGIAQvhznQHQvhTD9ijiY0XEDQlYxdygywzsSVc46Ilj/EYDqJgChy0Ei+36V
AmHizYyXDiZG6IOsgNfiTf974s+VL/PdWYto45Zlpstf31k8Dac0pgVbMyTKLs6D
sCCU0ssGQnz064MdxOgnkQub0ZAptgtUYPjh3KOcv6XE5/RyDiBCeJFP5AxLPEjR
PTItq/ffwBAR6DveK0qpZMuryO+4rDEHYfOrKY35UJ+UEPele78m/07VDz2gVUTG
Ra1yaJitmUeI38EmH8jhLeoBVi2T4SojpkP21NJ4IdAjvTi+GJctMVqjL8EyF8Bm
dgpuKmUTDKMrh9iLmvJF8n2beTjaHLF5uDFZkycLAPvMytQTNENX5F+bKMJR76OT
35u3JXjzco+JkSEHWq71ozRyrAfx0FAnB0lmy8ZisjUK0R7ayVZa7C/3y2lMKZUI
KtObkwc9blkuB7GqqFag8+O+5+WkZVcX/n11Mk+NF7Hkipgwx1pJzynbS2mb7dWX
EVtS8254RNFGFahz4TEeS+7WvFaA1jSxDHXUDpktrozr3Flfb5N6ovxfAV9N6j2A
BRtqtbXpHrSntJfPrQQfX/qpkUaVg8+SxSBDmS4k9axfmPoQ4HikfH8Dh6mM2Q9M
6z2cmIBNSB3IKJ23rTTXpiUn+9J9LXnNoAf54HxVQfHjoEAK+dPTMgAyVNO1+eJN
ivuy5SEKKNRs+DPSJdSojTQkwK9VJnvlhAEh7pqjjOJU2NRRFh4oJueksndMBp6X
f56xte0EXgZCfOcDfGk70k6BbaDwezqYYac8OTMua9wWL8tnXAHnLVN9+/8QsEHL
r64Xomkz2V9GVmD3MRQ9owFDsLPpn5Y3suqiSpJp5AxTcAp6541HVeF1P9s8AY4k
nchzOLLAI6/V1/TcVlbLjFi1BLNQDAfNj6XV4UV2UMWRJIeewaGlya892OijnOLU
uky1GieVkZd7MjEzMp/vUobOpjPcigxv5miXGLkwYtRoLyZ4tUQyRIl0/aWY4gOM
fsUXDEi8FJnact/ok1kketu1bp/dd60qCi6CnNJMf39qLrqSPpj/lPloFVF1nJtK
yJwam8K096Gb86q2sUnoGoLfA7HmyGjlVJ+juVIXbYV4niWIJV3/yRd162XJI/s6
7KgfplQ+54Zjr5qMf79WaN53SBhPuZEYGu6lzLIEYZF/+qoRzGZeYk8aUT6KXjYc
JrfLJoY2Mfl2bR7XyCpOxNWtWNMdOaOAubep0BDPvaxlG45A4LEb8gKCcSOw3qLu
cvlHOFHS49Cvg84xpNhAxDe0ca0mlCgUiAZmRtQXMKqHuimGSRCHI9xNHONFxwG2
mvI6JT/Xf+5DTGc1H2a7KA3T9qxJjFnv5Iffahnie88lPtZ8eANCM/dGQDXRveam
HZcO0Q949HcBM0CGxciZVVygtrfC6Aj+25IGOo6M3GqPjFe4V2c/b8nDA+fwdQdy
wyF9ilTDerCOMlocIlC9uvI26FgObmXw4RmkF7AaN4pNLwYvWbz66+9bfLTDIm2a
dBdP6FF6WIjMXSs6TpzoZJDOsUXFyaAAjcPRqKiLWjSeq65z4UbHjWJvtcCi/voG
BsLh8ELTSxuRThCFlYTOfh5fy1XPH2l9iy5aoYaMpCJbKOO10SaFjrl3BVw/ZLHN
ZKzJjmBvRjPNZkeNgOy6Cl4eg42OfwHP3Pt+Dtg8i9GIphqTnQmTBTUoVJh1Maf8
8K7KFDyW9BsBhnapsnGzy3eoVUy6nAfayAdXvzBP6gLFjVcZa8hCF+AHJ+WfXOLO
GFTJc8m7kYL0VEw7XBtFn4j9y71XOF2s8LBbyHKe8/HD/sf7RfrONj1GBRuVd3ZX
Q27TpSqLTd66Mud1DlA1R+66UjF6lkdDcALc734XG1YmO5/4iZBfMZGoJRrbY7BQ
tWPAhMyvVrqvrR9eyvzYIrgt2Gv88h+9kSXKl6xRPdZt35cUTRmpxruNqrNeKDFu
g1uEf0WZF2AfRsfiFJPIbSRDrBMBV0u4cd9O+j5mW8lsUncOKEQaT44f4TCKfIEy
5fgHT0xUTrWDoRIZCCDVa4VsSCUiW/wNMegyQLwIBk1OTFCCI2kFwyA2ZNwiVnJg
HT1vaumgd+iR/ma3uufMzdDZykkX8rPNz0rc4DyA7bj+fwUi8THo4U3Dwyt3urQe
/G2DPJfE5NQbclDkVw9mE/5jeUAWffc8347MsT4eVp8kO3Xk9QRTL9JyzOtWnSLW
1nwIsc9qTghEPvp4/99TaSE4Xf8faxnFKOqpsxMBR1E9uQdigZ+5NJNd36HE4qO7
pZCBFjMhnKbKn+sZOr1w5zEOBleJcYuyYAipmavIQdrNzaHysDmsXbiQLPq6ODED
iP8+LEJH0/vwFd+WoLVBr0U9/B7630bHKTO0ROfom+L86RhXZsCitkgIaND/bBkG
dl2jp73MlKJl28/QLZPr3DMLdbBB/S/yVAXaeZzaFXHte5w/1Z6nMp//spMlsqGo
Y7kW56gX+tF0CfnsWhTtLfS4gIJyfINMgNBCiZ2ttIGnwTNIevndr9yDxpeusxr0
vx4mpWq746ry/PwsMEARYsUQyN/JJfHd3VUrRBm//e/vSNf5nrOdk5NlEiHFzKjh
9B0sJtACLsTM5yktxHcgVgDTFkiu7TIisg9hpPMOf/S6XqmGs/pwJB9vXaFHRKyO
BBrbsGFa4+kkTea/FcjFGwlsrmO+D5LDXM+AC5DQpNxIXirBwa6Tg7bJC7Y1Ev/E
WEDJgeiMrw2wi+pT2IY20VjzRAeLZU8DueSEeivbeSQVs7arQCE5VIqbLtX5aiem
LpSstgwpxApNpdyyAiW9LnM40fXRo5qJf7cRnqJJIIiYoiWMlZwnLpTk5lfZWHtK
uMdtH67uDR3k9L/1/TmL0QDOExTrwHRpV0TyZCi00MRYMSMHQkNwdD5YUOnw7/8m
lTXAk/Uii3MMUIetSJ9NibMY3RfZSBqf2771LcCnhF6jc3BbEVOnyEBgI0phX2Sd
SElDrYj6r3ZQ8W9mg2w2RJW8AVz7depaUaDjTjXsd1wxZd9xdJ8X0pxSRKdHNOIr
KPNqxUVSGx7l6O2yT1NyLVR/jAYr2rUEDwWpUJUABYb26s31OtaSubDXGll98ouu
mf0Cw+EBWR7XmGSImxT1SzTgLhMqqAddWv1Meg2gckySCDRSsp/w4ofN7pDn0Qkv
IpBjKF9FF0pDD337KtX8MjUP5+MazDSKmVLlsnVGhIVeFb9ewDsSHJKvsD7uS0/P
r/dqF0/9EaGJPF18hA4LKhRKmjuCOm6w2qHzZ9NNfhdaZXUk+LGOspqLK3RlkMaO
4z2PKHfUMXqiMsKHXkduVaAP/ee2lJFnGM1Ii6pnO1ZyCTNnEegx1TnWf+EpKNRj
fMQFyyqzf/gHiyXKcrFRh6RP9hT+NXNQ/INKkqeVn6AQc/EX+iggmIwxOxdBZVXO
eqHUBbzSMBe3Ah3kQqur7w==
`protect END_PROTECTED