-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
hKXQahiE8c1uTn+gY9pidPwI7pQqUpPmgGVWuSajCWiS7oUSFDSSjGjisHGnU5mg
vfLQ2ky/bFuIpole/xYbMu7jU8CCKB7neBgqmtmBAul60RA2cylt6CSG2dabbdb5
dKRHr784x4Xb8jMvm/WveZJLhG5r668bD775d00ZrDw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 13027)

`protect DATA_BLOCK
ofdy1whf3sLNcNcEVfo/grv+ap/7QtlXa1AJedPxy1PoiBI1kYJLx9ynCrYuouB8
aoZ0OaR+TGUxEXDHag13ue9QZ1WQMManc1Z4bzIzGaBHesEzvVOZ2Yj9pwTfaD+d
6g/vhZtI4x0+fLRSk1Z5oxcaGFa0AgsR7OrEicHcNe64nMzro5uW2BaRe1qitZIA
FrVBmKn0C5/uH2cvNxUR59ML7XAkyf91YIvs95uj/bb47QOhO9wNzVjQBwzis7F7
h7mz8aDbU1jDlwXAnsISx+/uyDjHYDMHXhjj9BdmIa48tel3lVFtrrFVBa+/t2Lp
nRXxeN0Oy/KFeCIg4z8Q0VVV5/bRkBdvTIYTv1ckKuBkOYOcilnUOOwhdWwmlyQV
lyXXW8lmksekV0YVJ24dM5/cQ6idW09O63BRRN1n1A5SGq+JURA7X+p91Icuy8e1
BnKsq8kztf0Dg9Mpecr59FchPPaLn57y94vV4eix374G0I1USpgKpBHVfM4C0E1a
zhFP08k5LHXawrZ/P1ZGBIrUzdxiGm86xSWbJiLavrVQN6BZ9eMLxjcnkvqdFTCX
B7+WWuWluZNF+h5/OAXnuUH7UqfF7hLfdVoSStRYDbTAYmYZXNm5ittG6qvB1JQf
7MeuvINZLkITl6C+Ui6NkrPpJgQN+ogsehDQDN6bQESiiPWLAcmlwAskpS0ylCvo
CEOBN/LGmsgAmmL3OICGoY7ajFw8mntEuwD+LlCYh2E1yTehlnp+DleABkRxmrHL
rzD9CQw7bqmw45ZzQV3zWDZutuLdxnrXikRL9SZzXR50qmHTExC2zNo3Wtn9GiPn
QJWf1xpMve2n3b3Y1qZQW2ae1FqIJGoanNmwG2bRJGpHRsLRWAhUInHmXELWmrPk
rO0+Q/imjk8Oom9/Bo2xm9/b3KfrN9x47quPqx9QN0Am8iG46pLjGRJe9FoYy5db
2wJwIXTbVUVp07FFUmaMXfmgtfv5Evu3SlNrSQ+/V9itDXaGF3rvPbJBUfrjOQEZ
dimXYfdbdT8TyWquLGy0Fyw6Z1PdYH2nWSmbprE24eJABLdqmBkpSWtL54hlKwBS
GxRxPqabhMs1B0+X6O/QCZuwFVq2nuTtBAA/FQbRFUxWBSj79qU+upngxKiwnsPl
Prj+LCqM8enYWBwD5UnwJ4gR3KfZ4L2xOZlU3WkL1f+TIZS20780ejQOBYfkWZYm
m2LN5d37FQOOx8NNndeSzepguVsGLlhgikPtlRphS4oZm3Nz61hgdbkWfkSJRNXx
sjBukEDC8AAKDMZvNvC/W6rAhNuYCFcYSYoRn/U5RHmnPEsbvCQqg1Lo1NaBXBNh
kXxfpkkA4JI+NNo+0FWJOHjdpgIGvijAAoryc/EP+bfdN6YNBaEWktBK1rn/I9D5
loz2Ten//Lm7iUCB4JaTjXNduw9xGbn9macKrzuTD2YZKI6cPbBuwuHMlZEVFxsy
1OmeSlAiaN1RfcjjXx3RUf2WocVhgj1lB65VfLFt4sFV9gOs2V1+0RF9VMO/D/xt
uqiXSioT2LXJK3DMa7SCq1Y7phRAr7dAzggJdYoNQHO+HfQL2K+97MN9Ibc+m2UV
ChCIGKivxDvXRHQrN1znPpIdkSn3M+qV8P8Y9mO+bRtcxCvRaOFwHAxG5w7yKPal
7toTB0jYivQzkXIup0ZbwFgYFtW9UfS7hvkrqZRqL+liUF4nR89qu38fmII8GZRt
AnECfgsR3RJohUaXg3cNMPzMWWlrV5hf46/AumFdCRa6Soay1O8lfMSeNr/L1+rj
TVqs3GyzveH78p37Z3Ka8q6PRff90h5rX+hOwh1fprfpHhyBlWhJ6v2LkaNTWfhu
O5jVpQE2i3pKRHWaQHU7OMJBp4a6i7OV4WZk6agYNGR4BaNnGaTMJVQlFfQSPYbx
wF1c5VsI16PT9gkswwLA6ubnkr6vqBSS57YfKgnOmzftUsQ+IGnsxmcKtZmTB3vv
y+D/sP40hAf8QMn8cpuhHyyyxKoDRSqhPtRP874ucjDg7X+erZIa3wPS+zVLiYT7
sWsw7WCpMpmBJOTLzWN3BGhNZqOqk7iKd+iih1ZBwY51+udde3aF6oatHSs+jhyf
pka+BAA9MYeXQp82toQ1lBAOaV7Lnr7iDnmnxo/4jIrNWBuxOUHymvay6RlKAC9m
YREBLBbhS/b7RrfKZRF8v+uv81joSS4lV7hSv5F+6w79V8HXtEeTwaLpom8/YP4D
+cjrgtEDwzOBD4//HnyLyoQWq9JF8QZowXFzS2rTt7g7TZW1EA+cJCnvjbf6BrZJ
HDLLQTbWB8ZrwPWNoRIdTKVwjsQB/aFeqK9m24B7BewqelP45vGfLGwUNXZk24gC
JJKojBD4/1D18nFxdykUNYI41/NjA/Fd9Nturx/0FKerU65xY8mj8KR3YjEnwhba
rR7a7OzNEU9RrV/eM1lWcCQS5nWZA58kwC47YVJnaELQq22CgFBCHySihyZGEWYY
BVo6BvYN9SVbDdP33+rPdMxzQf9aGX49ztHCNCxnfY800fLdcM4lSHk/37Qb2bFE
dML1mMuE6s/7QkM3r6N5TzzEhiybnoV3Q+dbBRlnHpsInDoqrdYDyRZW9lYEETL2
iiBv4ebiG3cRA48fBVLHXVsFSgcxioPTQW8VUnfKh/Vz5/uJlitlSY0DJ7HFgfGe
z6Q/pWnIHvYC/zOwhGoXx8lphu8QeX6W8M7g/Ko0KUtEBSWFJEMgCp80Tg01Vu4D
2YY+sIKkNb23ecugtqWCDyxzXGJThFRR/MQdW1HmMXZHS0gez2vbveXqisb3UV5K
Y9QF1mXMa85j5E+ME4GX+NgGV1p1WuLz4PzfjoWoS7Idzxpifh6u9GqOJpSZCQL9
8b0L/4WZJOhD+N+yDRxtpn/3o3aXiqlSRopqa8NVzFJX4FG7UAFX0jDbKsQYm2c5
lyrEiyVSYrkDjgKkLQPl2GPYpRnwgbHklfW96aYRKzaUmqgjRegOAly2xYsQ4qXp
JZFhv8UQzgw08wkWtwhfNjmlPKwXq2R12FnPy27p1Xav9BOUPczZACHRtzcHTvgZ
G92b7ye4uoDdZLKurGyidl1EeBS10BaItkALnZbIuALGToRwS4DombcKHMJgAH0o
PsCoOVf1pAxFnKxKbm9PAGKIq4Z60D/8x23Y/dt6xNbhOXlx4UU6TZFYgxnUmF1N
miOzX0Vnbftj/EU0dfvMD1XKwHmQOuZNAto0wHL1VJCexqQ10z4lEEgtTrbLer5x
w7RND8eslx+pWtS9B94YxH86fA8gRIChwQmQvL1niUDn8m6jrpba4KHlcMzrW8K0
HPO2ul9vkNnLB43oAwhG7dppT+cajjb9Ey7/qF8es3vq6rbwIgojY097TkQed5OY
NALIJevIoYk+FFu/NbidKLkf/Oi2BmuCqpeSmUXpFSbE1tBoxr6pXQI9tI5+0IPQ
4KkxgdLS9Ch1Uk1cU0w1aBh+WyOGcMTvxfp72GGOeeoI/iT5aEf81/+61Y4Yesb2
kTPqvZ4GBbG5kLU9Srp6tlPMI9byYgAoQNmtGV8EnI+6ld9wBscvabsrKQmnAI2X
sduCzejN0GPGaZVIN6oGp7whmgeRnaqXikDO8CvtrDQre8yRfATi5wreQK3OBBfd
vWGa87D5NI9U2DlzQJ0bckb//mCBgYckhtQci9Yh/d9PJrqrHnucGW6VdNf2LX+C
yZjRug6A1rp11SLH37w0BlmEEqpvnoULpBanaOR8rLIaL9be3s3hZ06/8kEOfQej
huMmiax7jVGJWei6/OrWKDEHQ5empYedqiedIIhj0P6vJaaSjZdXEfw/EBId5iPI
R4lPo4yTT27s13EVj/e8O+KfqzeTJ7nmFYrZxF7hmkZcTulUVmNFzodIBVUOjFlu
b4sCEjIkPq/QQCaytdY6t0VSyODNuJgMDdvWtxHXZsO/RfyoeqLZahY3/y7nmaKD
1Fy5iR3vW1Yh+Cwkb08OjQwf0h0XqLv3pHaR0zSLhlR2shzfszPGEGLpHMjiDSXC
LZl8HtzNcw7xvSVQulBvzI4vudoaFO2AzGEa/BonJwCoUqZUnLYDVNx9nVIOHjdg
zvIZsTQESGmBdFHEebRKDIZDGAbtnsfJEEtqnfJGq3RV76C6yVgtDE4pfYRlnW4+
SlA5M29CaO3dMctpUY9ZSyZTunk/MYwapaXzMgrI/lfQ2qnYDM5Z61QGqMzFpMIh
umzUo+cdeFvbg0dlWf6O+j/M1s02SKuMvIQ6ty3lAhS5e8SfjzUG7PvEu3Qu9SyN
PnyP5LMC6mx+npyfbe0xOFOaOTQUd/IcZb4+fkopS4wHNsJgjOY2o/QSUSr4jdUB
6IuUB/1aXbL1jkj6sqymSsvTMuQLE7R1DLeHAdNfmu0OFACJJ6CeqSgv/gRL09Ml
86l8xGHurWL1agU5IYkCWP7FGtvbN+yw8X73y0qbrHshDmBKf3Ig+tgGEM/qkX8H
1mpZx5HHjHdA/X9SUXP+xHmFQoBH80GppKr1id+0wUf7rViUO+D2oN2b3qYKQ8XZ
6Nn4wkp7Kx6qm0FxlaS+HGo7NqD/DRtkHqDau/RDgegwa77T+9dlhbbzASJgM+YW
gORCYRn9SR1VysKJtO952tblRS5U9N2PE4zKFvsdr3L8WHfbFKg3qsugYJFMWGy3
lMf7dXKA9t0EkOJ/fLi5ZA4cjAnTT7wFrWbp1ooKIzyVu8qpnGwJJwVAaFyhUgQG
EI2RsJyxCDeukczGnQhtlkLrazJa/vxjsnLei1hLnaQ3+OhwryrmFi+M6f4sNOpP
WXzrzzMpRHYJrEcv/6dxo++tRry+ffJna39CUw437DQVuJs34Xp7lX4QZ3rHfCPq
JiNhQsphOBIFJeFhzxo+YC5gffOzYyODlh4NS4MaiA/Ihu54PZl/SO2S4ZaNZ6jd
BWUwYm51EQZhaSv0B62Y2T4ggX8uqRbnjklxmGhn1fJHSs73gBC4Vl2hzCx64i69
0+vACMeVhPLA6Aun81EDbg9N+yVMd/7Q95MwzgfJvpxrmZqz2E8KtviwC9M/1xmn
U/5MwA3pWs6NmoSkKk7uaGFQWLQ3BRf18xxW+F+LQ9jWCBR4jHLRzzS+kwsc05oa
5NDKFc9/+4WbckzoKYsaESGde5wehjJuEOepsVEWnwxWqlmqDFDgfO7KkOfbkOhv
Qn5UeKz36b9xyr9Td+Q818nixTWus+pMAZmbzmDYBUrFUm9BiJjOhsosOHuaBRds
arzoCi2Iigqx5/rPvhxeMZoHxfvEg3BxXP4H9/ozlWZciNc2hc/M/QZs3VwityAr
hjHU6HVulmsgzxIzDDACw9QkJKg35O4i1KTmVIORi66hzu9dlXBdqM9PSwwYQwxS
MS7gpODiO2+9+2f4UpYMlQhEWlKwIXSR6JYlq8Bkd/7KQD4XeCFK8FadTNvti+hL
uCfUhjCIWd3h0g6uNM3O4jz6MiaWdINkk98457NsiIZsKTjPKwU3LWJr/xnqQjgI
D2Y+vXUOBpAqyqVfajtjs8j0ndZvlrre1huSP/BqhvKUb0W3hUk6KDVGeKLNJNDm
v2HkDral4oJ3Q2NS/cT52guVT9DhFlSqRjU/bwA+ccmNfCe8c1OygUQzX0e1csvn
lSHKAwudgJoL/Z4y8MmxpewJFWA4nuVv9k7MafEsK4bd6nFbNUrPKQ2NPqL9n3SD
LVVhLR/H7JKoNKj7xK0Z1SKSiu2J9OwTXNIs6wlgC+1HWf9HF3MsdKVWSE5I9I3t
dWIIgtbFsvCJL4AbvpJIPJfLPiJEO+cAK73E7gTQ8pJHzuRoKnj9Kb5wqOKB9t3J
kp1K/XnS9BywPzgoTotE7TIkakdACRd3unmez2clLiUj+fOg3lIQtRclw0IDl6X9
yR9RNjEl2loDqqZ2izc536mMPBxAvrLwOFfckPckuaafShZrnB/ndc2+ge0OuLGy
F699Bq9EAFuQV1hlyK72c2dibjEWfwIKEFKw/v241IyAdiIeShr+/R/VVe49A6sj
ZLNU5PWoXePA+CKGY2w2lHzYyJF+ZO9CTKsAL+yeWqplzQZpW026UpZQ3beNRHod
KfxLWS/b9nY2k4aZl7oalO1iygAFzqrfFmLlD+/jdWpzJjA3drU1GRkm4pJbRFxo
Qw7RiUAoQ60bcCtGR4DKoM0zB9RL0mbToHOHGt1LCw/OLFKB8iltdry8w3P7LCg+
afrq1qoPy/GIACx1VQSL0s4dmzO9uPgOvzp7GsUZO8c0hJqyfl5Fx4aLU5gKFA6b
AM1knrX1qXYigCC1flcssS6S6HyGaU+KaX6VFdf9D4R33IRo47H3ABRVlzzkqtsd
uYu80I0pZQev5VmAmFsoo5yeangWAE+NYfMp9IJHQfDp5AuCAKTpagDLhaDpwGki
122iCClZLWjljHDWaBBWCX4ppojh+IYJfWJRNCjM5P3W57qZZjHmTNPjn8PfaaDQ
mPAfOt6k40FMr1ibusuaWtaFceeFB/j4Af+jhqD7PPVh2fFF3b5cDANrGjFWHsMx
u+O8E9kzQz+uxRPDkxrLvC3veUrZDOuZbcMV4G94r6y3ZbsOCk2NunLXXnzz67yW
z5VOQDmKnSUivwHHRnGQcEfEaJnz8PAX9fs3PF+TyCGTEI8apOQWNgsEmcwFrgIG
XuLGgotZmigMaJHXJV8B+4FyEa1TJb+IRkSsUlOJy4u1fm60h5UU5KRLBaxewe1Z
Tde8192/HMMaxGTFiVIKGg5RpyxO66uX/Gae+vdSJlkDS9VwjarbXuVrvaYQe1W/
b+Eyefsnv7jG8NJ14YEffR45g03mk4cBeusJCOMdLY0hABYubzRpDHBfsnwo36SE
sbJkjJiPf669EMvnRV4DIwEecaYJpYL7iB+WlFtdKUQPAlpxrYibMvAPsVnuGsba
44bmS8LZJvDM2sXYpskHYS+zHxHN2Z8oZEFnI/Rr0Bgr8QWQohENKJhY0JHMLbfg
hSCN9UmvHARoRniWN+8etzpDRib7JuGslzgVhfcVPALK8dIR38HpgP4Osbmvuh7Q
nA5YuRdkIrj5Vqa4gaqO8uwlEhIIPA1J9oJw2Cod52MSKWbch/DWtb3s23/1PLP0
ZmwKgqxklDGbv79GnVPEcxo4ww5C9NOCEK4xAKhR9XXgGozfAQuht4zgoWw8huyo
pyRTopALyTgRMR6dMxhgyycg9ABRUVUsdX3+A7anZ4ptXPVPDaaNjUGI17cSUlGp
cwInB0cfIO5Rlhj7gePuAaeF6qdujPFJaor319/b3gMVTAY3t2yqJ41KxCDMVoEJ
xTuC/1xRydBRCGZ2kBCBWqtZP+Xq7eMv7qV9VtOzWtGtCXs+yjj0pwJre8Vksmp3
mtZWStVqN5Ez5xEqNWOx9zYGKDjw1FgOQeI04+QgHAArc8fANX8V/f64Vasd8H+g
Dp3jT18k5Hivofnm9dSqcioDjzN46+L5S+ZuTPf1xJEp6beKCpdBGxVUrXtC93Mc
4dk/gUHd8Tf24B7gYv82T4Lwu0KWnkiy6yeV/mS6rDoOGbdt37qV0ekxe42mDa0E
R68Z2gr8he+aUbvuSMJwjHn6l6nhYz1YtrD9rGq88658TfVLJBjpHsOpbfq4Lf0S
yh/fXOzUu5W+ELcGu9n+aTNuyRUaXi/eCfez5isJUlNlDI99qKTneTs5FbFJw1sm
Jow9nCftMWJzm12jO++TjC2tkwcVO1rWMkLyj78i+ysCI6fVG7Nsj00cBFhRa5q2
L2/o3Yv9ICWd+8l0nt1bK3bJa93vsdVjt2z3GojgDYIISgzVPcBUfKKoJQhhAy8G
OhWmAY8OHRPHBWLo7lB3dN/BASP7D0jlyvHM7DyKc7boNqedP1XbcfnBTwOUqPsU
FYFfJPfWEUO71r5rEg8vdy2IDOgEMfLKMaReCIZk4OidrGyCG8vDNSyh3DZhu0wB
KXr83fz3ZEXq0gmQY7iQAiqhgc36IVUr4XeeicDYp4G1/KXKi1ALCbJoBzN7hshI
vduwfi07FcnajBL0v27k0+QWIUvtAH7eY3MMuVK6/4cyD5UBm/LK/DDTXOBFoVN/
VTsXKLYAtuZ4yG6yJSVSCKoMMhcAu7hOb1nm8bYNZVtiBSpuE6frDTojIMyZRG8y
vCpigkYlwKFgPkQXaK7O6TZM+NKf5Uf9oLcwnoRthTX3RZaBdnpechcLWu8OJTO1
VI36B2O52NZjgM9BZS1YvBdRhnnDD91/ftZ1if2XTqGmoUiOBlREYVyZBO0bilFW
u/SVBpKI41MbYZz0ugzxfQeN453kkCNKt7n0Mu7mXYXCFhgNYAKNSIXr0f0zkR3Z
2BDnI6aRgCcNy5gQJMRNXtvXrEXJb2WAzY04KYq01NMhR/ITcBAznNs7OZlGfbXb
OYM0KD1PxVw0x6sTZPNrc2sqatCrwo8P5NsXPVOD/oatEuf+bkOxzMPdwxN+hxvW
0MtojUv/tq5tMQD8bjxvMkJQBKFX8EW+45SANDtBH83qy2SPIyXMoyTkwBpVT0nY
qI7nt+Ha6HQmrPQ1Tpj/EpsuYpybDJFxhLytVngiWPyWqB+ifNRlo8fYmaL+cafE
0fkWsf45DknrSQuZ9chXttNWwXOvo6AXf0Yu7CuqFv6hSEv73UhoiKlqvZ2cMiPL
83twWqfkN4e2HAmm+NXFPsrlgndF3SbgGjVtAw5KtUpxyaqPR7gnhTTd4xRfzWtw
R27oEsCEG0qdeWruSZh+5HSUQtEKe6NAVbSep9Blw+q8alhlJkQaUsB01T3QrGhU
on1c9rM1lCSnK+hKrN9vQ2/OoSx/x27bJpejOJqxTylYO1ofkhb4K+HfyDFXf+Po
nJTmNaTpM1ZCln6czIznAFi/EL+myF5GbsthBNZH7FrZwsPtptWXxmFOEtRKkEnf
PIkLuVwRq3QWCn4txyiggDkywxg660jcnLLsxkehqkIZsYYiGyP0zlX8GWWvNdY9
0BZ9D6mwi9fIbNNKDpJHrKZCGXvvWKjZ89GYBjcvo1ERUIC63/QrEvai3vewkfMD
D+1dvet+4SdA+k+P/mt90gBB3AmS723CGYwX+atLj+4qG9C7k3xPnyM7eitHblBe
Ku+PY7Ly7vye/bKygJsxkSyL94waXT4dBV20kmMH74t1EIJiGH2oxK2rKqWF22K2
hjfN6EwBY/Cq9aG0vypiiNzaXv5BtAAxmZyNMdr1krw0zi9U7yqTgg89xwkGUUQ6
4IftIVuehFIoLWstJS5okRrLdzI1CZniIuYIOoeEn1NT2gZp3oJTYuItdA4WaQaZ
J9qgubZKwBHFmrv+IfpfgUlGsfJLk5eUzWO76U7pnHgRtJ/Pgwenh9S5tCm32WT7
WpVPJKEMHoHRB1bp9JO/+xPAqBvTZu5Q13DfUJ3HaAmN8Vl/zWdVOCYxJKcOGP68
VaFG2LDo1+7sEO/Zjd43aPQtgYgciFzWH5/TN3JrQ01zySKiZzqKv1Ti54GYyVUi
LXO1vntFYfzKZU14P1wvBZ8ZOF5PVYW9Wf+jbOYm3qbm2l4zWghfsfZZHys5vMbt
/gqhHswEhSfeT1prus0XLASrV2Nhz2C0LuEik99NRm5ITBwHtvNhbUoSGvrzlHby
jiRiy8cVpjiakxVoq2SBXr9u4wOyPRuEHblv8NCe/sCySe46vpQ7PSCMPnt/oPVb
XJNnDNgMBNxo0ev3117l5iZWaSiPCDFk2KJejEItGMc/q88VmA//wDilRetBYAMS
C3wPaG2qg5ym6bf9OyXCxMD38cj0+MyljYkWUhieU+D5ZbppJyljqJNH6WdJ7wAM
3uE9vwe5cgG+tNbrTCFO0wQo4ZKLXeCQsreETi01OGsYn1pDs41AsvEonDDd8ylX
AWPplY6WxTKyW6cuXzwJodIq+4rtIo7MLAqGg6vTO29UhegMlPRG1adZ96uKHAYR
BN60LeAy65k1j1e2emcx7fS23XhYdX3+P7DNIPDf8A0T7b++AIK5ZkooI95+YtHG
LTdcJeMHjdEpw6kaL7E+8t61xrkTcQzi8n5t52qqIjJj3TmW/fi1PzaXU7RmWzVm
ieXD1yNmSFrhrNFujs6FpErFtRquoDxyK9GTxJiKoz5dtF1TKH50XihNUVKHSLFM
otdEmhxD4YAHdqGBJ/9UAL7sxHwsJR7WI8L+zILgdzcf/8PyC4IDEpChppFGLKrw
GcO0uxfYG3kSizE6Fhf2U6ByXO9sHcFVh9n16hHALmmEKXXr9BIjnyMqdC8mEbNN
vKlA2aqCXPJ4tRFc++Iq53mwXrzJaCMW6fXFPP6JiL1b/I0yU+ar3qFxl15QcbZv
mdzEcyikZ6r+ZRijkLxPB10JcsGJEJiVjlYlpnroybAkGfecIDGU3A3pm39x+xlb
gM35OY228y2bnpXqQsZDv8tHnahRj0W403XWnDy/H7BprNA5H3S/+B9tIiCby/Nb
KV8h8CQodP/9gHi5as3y3h3X/4LYlMsKI96j+MgYZPrIopcG+qm4EmKkox37KG5C
IghtjcyzH/DCm9ZNgkA7c7v2OtZVxWMahbOGaC6WE72L3ZR2c3cgvFY56fDZSExH
gw7wr1SE7cvBV/We1Npt5cOWcePaQVZw/el/JWtobMbKGdEjF771/SnWygsKYF1I
7FZNhjlXDKdcGI1yU6MkNMEKrGslvLYFWa/D11wjXoF5R06eko9lDpJxLU5jxir0
yT4xLbkIqOMyLNDyTEKyVcqEPDoyAAAvCgf967DIyVjsRza91pOaF0cVAI2Fq2q/
HyY1dwqO2gox8QEr8k++uM+A1HrL3LBhBfMXwl3Y21jTijddztzjmPere2lRka3t
75C7sUUr8IOFoxlqJm6cLevgGJ4bnsY9nNFUMZdSTuii26wzv5AIjG88JWcuntjG
qnrk+zOZF01mtzCjhLJ9xfCLUAN70MT4almrTiPJ6/bsxDL0SdTfU9iRGDIGc3Gv
sGNfQ3kdjdqR8sqytQoCoxuJULPr1ZyR7JXrunneqeQ6pTq0pR1MeoRz8Xw69AmU
jHT1DtxPuvXm8y4F9QFcD1pG+SZfw2XxdvrJtab6hxgVkscXwMeH3wJjklaZ2keg
2rZQzOkyxuzm3YRqV6uWLLO46IpT89AGNPlwACfCNFktLqOOnUJLOoAtUSh6moHk
R/99xGJ6GgsbAB+RrDRjE39V3ChZHEfYZ1djLjKbpb7EW2QC5MYs7S1Fy9YqGT/G
OszQGfuy+x/RK2KaOtRoE2U5UrrcJnLwXpuKK5oUB827GaiwM4jtwcon845fH1wl
/6t5JjDoFdYGuF/h6Nd9e3DmuIRMqqMSwe0L2+J8LGI7ls14UXODvIjU4eYw5+My
mFWD0BDqOe6Ep4TIvyQRLIuRDZ3W3sfCAQRNpdbuEZOnT2fgSBkT8r2hasNgbD1m
UyHHFuSoIJ2d2iaEJunZ4A4zE1U1oaK/lBydM54WL0poJIX5Avoxe8wlZU8fnFjA
LTFlL0jaQ6otXG7wmhMTSLFpWxyXJm7/MuezEi6PcVFItcuUgB9CjZavevwyCR2J
1XI7cWPUIbOOzSsF79qdoXudHEnUamGplGOQk1gqFpDHi1Vh7K3MAIhbMUyTvqPe
airyDyNlT4ZPWjrn95NqKfkjqXRT37KTFaPRyhn/nl6TrxMpzy/5C9rm9uLNqS7d
EXmfxYG4LK1ZJb17T3FHBu2GE+FpRS5I9+WOGEkMCoLonyQdXlHOmyNQVj6r20mJ
XKgb3qI49CUsxGY9OPhTRciTrLwfmF8lYISXF6ChJBkye06RyWBb8wNVDJlOVJP7
VtLL259e/Ln2XBz5rT4r/hSaZADDYqpJm+IqQ0vUYSuvMDl6asus8SmGoIPK0jGQ
tnMDjjlmRCpaHkcg4S/kiz4Avyu/u2Wl57ERlOIrHXD8SZzZKMpEinJ9QO9j7hKt
H5kMKXYEROCe9H8os88s5m8WKvFv5GkOLowcGkErx01Yj1beKb2PEWrW6tbTjeww
QHkeWukBLfY9RcLFMSwgRn/RoCx1z64H05csbYDrCdHA2O+wdnIt9JKvefX3gXVJ
HRectCk9OfOZZBCh2Co9nHnmjlHF+MsNrkINraMLZOzEfD923vTX5NbUx8byxcaa
DfxnEFu2fUOXnBF9YT5gVGv7YRfWAhN9AztJJ1P4jh8m2zfDpNJAfeBCdJnuU2ju
PvkncVF3f5DKupOCAnpenbLcOezrdCFu8kBs/xfYqDlUbqmZw2G8d5MpwiexE3Kr
fBRen0WoqI0frMfe4BXYaGGC7jux83fF7XoVQMRUi3qkN8ucNliWH5L+19Z7QvNE
dJDz3uzWFyv8FuIVQxgVSFN/5RMlXfIJAs41ijOYxIwqefYgBAqw3rfJgsozjK6Y
Ngbjb/xEyc7jQmLFF7co0Okj5pchMR/hKhVyjyWUsu05u36/Oc7d0DOoxHS3MkwU
InuFPyvmTlU2Dli+IUKmj0riGC9sLUvjUhooIf2xxUdHYxxbHak89vliu242uBp/
xMOeD+XVwyN76H84SBGDOszxSbZafokdlroLciksfR0cfjC4W6wAOv2xUDOM2l27
b8ax9XypUuKqQYM/9BUwm5za4G/NAjGEAnBHPl+O/VM5h1ah6pTVVACfn+eNdOc6
a6yz16A33ly/tRpTn8HBy0RKts35fdyZJbB0lGnQ3DaUq1aoZaroMrTEUZO3OYh+
9XVtfCZwHYBYOazQJnWbS4VcUvG5GJPCUP0ewr82xC+Pb9lR3PRDJjfdCWb1h5um
0yYkBz4OI38HZBHFPRudcSpPzqxUXpnBzX/mmYtlHGI+wkC+r4TeGs4cVSXQ+iT/
aAMWrebiHQDsvizfZrRdNmus0L8w8CfGC/A7CGQLw95mvNPN02Ewp8MtCiZlfpbX
BHdXbpwvsZMRWms4dsXqzSCN7p96GXKcbfyZLM2nF8en4BD0MWJep4su0SS147od
hVr5kRrbPhOAxTdV5BQaKcMwXPVRydlHfwdEls6y5MczEypzw70mR0FwZ8VsQ7e/
fcPu32lq6njC0LWf7Wat4Tob58ntfd2JrV+42Zbp1sKj2UBI/fkzOw/2YzcY6eVZ
6MJUDdrn2uo97tSpjglbFJrZsGT0tduBRXWRKsHm7mSQNX++hXIYcT7nMrW5yXPS
69CYwZmiuHBuSN+CPeUDJHqpkXWYzzYo00wNQTKSJkxBFSxGr+a+SdgcVZz2LWKX
5A/S14/pIbdRQD+W8+JoN5Pz4PlvLS1ggtuGpnhDDTvb6H/FSi4G9IYMbA0pz3L+
kV0eeHneK5XvmluSMHZVdpKMKmsIP+OV5OZ6ioOzC/aSQOZPqpYVUZl4xT8dMKpg
vshIpU7YKMJkP/L2SKV5U8Q9dly13i/DzOntsasGXcpV+fAksUttgIfffnW8kkST
FpSvfYKnpn7T7KJgAIMUKGmZzVng5Tx35AYvSfDyqdEOftkmQvLek7wMNEKHdsl8
keoRQWZrbTWXVbC6xfOjrbzeOp1rJmk/5Gw3dHzU29T7Jb5FpIudNn5TsyTqyPY3
pNMQNc7ZbTtzBfNwrhuEdM9Dp2ansro350Dw+yqP1LRSNJSyKzTPZwoNzTpEdWdS
fbnWY0AZPX5fqvIBMsaH7lSG6cEuGYSfTD4GRDm1vRYshiXRVX7KNx6uUIr7PwcT
NxMbMvqwZur+8ENZtIUjtw8kLFKTm9fAEQree0JhmSDaQnx84w+DG5T5r3eqCbrQ
gPYTXADIb2NWXELvJhW7aLt7RS0RLwC3fYttdBasCl4NwjS3BHiqTmzuf9TlrgH/
bU3p7NfZslp9scdhiO69MCca291gN+TWWp1sBL2yyboOJFmDBtraCznAKlsH/AU8
E3mNG6kr6kds2SSKzRCVf4J0B6MA0M/yiX5+eN82XCio68/Epmr136fsrq83YNCt
2gTZMOCbGvu8mYh3RnshSAPGacQ87uD0LXPvU7yzNOP0w6/BAaItv+iXqMURjh7N
cVZDFrivJhgm1CxWy5Gws/fX5SocifLYSv1FIR5Ma7TVc3a5NjGWImu8QSiTrFHG
5JzysH9LLmfPNz06qJwDfXoN76Cqjc1t3EB2o3UBgDy3eCgfVQULF+bQARULva8E
LMz9lcmGKQMlIFD35NsQEaGZ+/oR1twq4l9SCqh/PHu5Xf+fRfrpM0lfXdiLabhU
WQtzHK+j3WDSu6AdBH7twbQ5PmxgUadLa/7L/HLe7mVP2YQOsPX8fw51mXn9DGy4
pb/Zto3zvhCuSJ8LKZ1e1kIrfW7D46wjxl2k7aAeiUWu7JvY0jXWhCQ7ofc5a40i
GV8d8mtLYnOudMsS1aLxIKm9TL5Fq4pXX8uTWB3nzuPyESbevI/QjXi6oIjXmtIf
L4pJfvim/BjPApmXUEEwZm7JCxLtwJklSMxljiXSEnjq9YGWQCOincoJn1i3vvN0
cYVRhbQtUU7Cee8STIoMKZzNdjEU2MYXwohCuCXWCZnWX2O0TRy7F+xVocy6G4wV
VpFz2HXgNnYb7qtVdl/UAPd5fnJolyiQ+hDWryya+LyFt2Wwu0d6drzRL6gcehMQ
fDOyJ5yTGxglER2rDMdZHoNsbzT8Q5qBJdn9B6MCZ/B2jHKSU6GtMRZlG2WCALY6
N0QRHGNhY1gFlGhiT5/l7zyO0obY+1Ymkro+hKW7EXiE5gpVqOptiCiKy5D7ULlA
hu0v/OJqT/rgCpCFykzLn9K9Qq3EhMlQyvDt4kgW9xZQ07r42Ds4JKNvs6L12jF+
tBtgDrtKmGw1k0UebChei0LvNBpQi+OCsiKLYNvrPPHhYLWh/pPvcx01Qk7SP31o
eX1eDqwB3yLfQx7HvYRSDXgqKtYW4XFAPpk7Gz14XCYQncuPsAwUzlMkejmz3hKI
o6aeJ/apL237GMnXTR2IIHofwPNd5kPdHOvtfBIuNDhz3K4ztgpKN7UcGmZAsWT0
fUbDWMUiID/SjlByBdoynIihP3KQVrcsBu6zteXisGyFsiEtE8/Szdg27KOyQkNo
k9f/werYYow0ErLA5geqhFEJxCcdPfyO4t1SJNqpVNVOVxSRI/HhjAyaycIGHGqK
anI2NdqWnRwNW/dnsR3+rkh16l3/ez0wLrKPd+yLWOqHvyI3LQo3a8eIq8q6/Ft3
IRKgRsO0uCd7X4prwoBiltanKXcGKn1JD61gh8bqvFo1J3ND3maDf9Eibbtxa3AO
/pKnyTY260IB+zZb9Yzl/bP0nKPKz5Y/k+M7Q15GBV+R+rKMXZuXTKZNkKSa18n4
PtHobWRixImsHMu540ziTJnPATyYtD7gOjGOVgBmlIGNZnDv6ODqK39PVs9w7rbe
QPXsLB0rLbdgpU45b/7KiNHbifLOm7Ns0rE7pIdOI7TTIlxUHYy8V3pvcf38VbJe
2DNzqdlmE9s0kQloLOMiQq/sb6w368rSfcz1pO89Lr0nZxxVeMe+8uvSv7L93A22
C74pXeiZ3+w69dc85D4Z+rTEXmaWViduWS2a2aq5p6J2gqkK3njWDnYMzY03oJua
UX6Q4nmrCiiMPsURf2ChlWywqBfjbptG1ZKHaetJsgGUb5h0bWh9yv7j78R5//St
PyPoUJFa9QNzAZ5r4G8RL7hOq+ItwCHxDZPed+Ssufjf0ybMekBCDq9xCXQGkogt
vfyazhT/IPSQUqALFWR8Q9uDz8dUWgv+0kEYgex+d8+lcz4xA4fWiNkjJKp0OI0r
mvlnQTHDn6LM4jkTHeIwstnLlCWpSZyE0xzyf/WPBspYPdJaLqje6w1+8VNphXdq
nEDFvj92revCqjM2KfYWrQcn125hc8rLEnvUFIK68Ttf2RCH3vnjWtBB+T+iEHVs
HGC6yosWI07amY0nOmCroC/H2RwtSlwNYj3+R8Gxh6Gwxs+zf5A9DIRA+UDIOJqY
curWupfKBO9AtrjgsrbxFixFNXD4BdG6VfdrQuYGzim0DemnFnnyq4tLPY6E4vZS
KToSLWHogBCZE0BKRAjnqAGEF68T7hzfZHq4awNm9++/9XLFO5uHOzCNs38AurCY
JrJnAoqaHMWFLRut9Yx9TM8OOu5cKp4J7e9fOrBZDKmszF4LAU/DmMaDLQyn21EF
A1nXZAC/7QM8uWmt7VjN4uCFAWTEaWog8KLdiRVdkXsieEEhyLUI2JWoX+axH+5a
3Pu87C4EfSMSmi/6a0P5J+OOg3rzQRf/XcptRPHngQ+wToJa0mi5zLnlOj2DYIIx
wCe9RacbvWMbaLfyjwmsm1T3ubn9TjwIR1kkRE59T0X1DcDS2pANs0l0idQLoABb
2G+x5fUz2sjJIzyo6NbpwkJzB6LUp6qPLIdPGOClWOry5vSZoUNx8NKU3flbfpSK
RrDAz0u6JY951FIN72s54GvREFvMX2cUmDGZbQppvZrME+w4nvc8tCLB930ADvw/
QlRL7tmELJUdifJH6rew6HiZCS9xfW4AcJYBOe643QATjyhcbSAVKzT4EKLWZJTZ
XKJVDUcu++rOMucmBExsfNwyFxCtwxHGqCaXi4ZLRIWWBlOg0ydkUq7Z14rnmxEI
3yTb9xRynCkNlVJlGxa0Q/jQg9E8PrVXrJRoWlNKEIdgde9fqgAsC9/D1ZPcgOig
EuP6LjOJiuQImvt1NWAJQALHGHEKysrfC62GOeqtpkvs1FF2YPALMSvME4lh4Rq/
A4S/W0Oli02XNIf6gWKharqZk7jP/ZQHpKYkv7OKeBauqgbYNapi8S67vB+v+0dw
mLksByjOzw8NQmsSnUQZL2b/C0hwUQ6nlPYlAlNxMGQzbaS5tXUU4vpCf4IhQ+FH
PJKdsnSjAy7q5InQDze8IKD/zoYWUF2HWWuR5EM0gR/SG2o9Yr7T4wsaEiARbIg9
zCyrqojqjnoR1Ko2QUgSoWog8SSpXnqOW9OxQIEWAc25AeEj6+Pm9spInmELvM7h
dFBNtW334+sj00280qjtmGePpltbw7IZMxlGiY0beHja1HMbN4fwfPRfc8+CGJXQ
cgCAbd38SQUQmz1Gw3feTtdo5+3qt4/lgJHXIqlkPs7fZ4BL0KOGzxomv1JVd45D
eikUXrszVff4J4SUWc/KOSWf+XdOhvByIk8Z1pAjGfW6niKeOOsA3WKM9fuZzUo9
lAYRu76mVhtSICHDbuc421SiLynQ6Ytf37clUPURSTrzeq+dXvs8mK29nGmfWVcp
o2HNwuBB4ehE81+EqFK96FMpvuI9IyqYU426IM61dwny7nIhD3DtDKG+tvAqecBV
Ds9+qQYmelKdWWbE/HgHTacvFGjkP0H/Gga/QAenQZOrth3tLj+rcTwqCMgrPNcy
s0yyefOLNGxsj5nANyF9OkL1EHGjCOsltuGiNAHbvyWOcRvLqH/E6wQzgKewBXyV
gu4L7ZRIrdt2VS6LKoQafaYxI+1vTEf7ReUAzrJEMwW+YDZ0kUUonzOyF2UHCY3L
`protect END_PROTECTED