-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
ZLtS+gMjKgcyACQLfqVskGJjWoFqgAiqU/fwxPdL6VVRN7LpUsIphDBnAfgW+X1u
VZ63inUf3VMWj1u0kh1iE8Maxk1PuVtbz1/JqqZYJA3Hl69RES1ZVfD/WWHwAupw
O0hwKpkZtVwSjzjbJJGfSExrIILpnidXWj0Xn4dNPTNORIrW0kxTCA==
--pragma protect end_key_block
--pragma protect digest_block
rpg3PDSxxrnPeZMFIQIVVO173qw=
--pragma protect end_digest_block
--pragma protect data_block
XhWT2SlH6NtzjuXnaBNRny6tXofUnpNgXA99QB3ERXHAVRsq1cLIieXHgjBAzAY0
RZ3fIRlq4OTlCmn2qEtYWFJ0Pi4wF6bI3p2cezU9xtI8WR+YzAizGOvBGfVUfxYs
MsxgWgPEB5LV0gaSDReQ4yZLbZf1ssRPWukkECfiN3qNV87eYy7tnd0o13ne9FC9
qYPdORD7WzAPRXe1PCDJoYocgxDzvv1IBHPimzfzlSKdkNfanGrduAoZ+47X34Bx
gYeVosoFJGiEjmZtqr3eGpyUct78D/YHKQXJd4rJoJVRBisW/Y2gs6L8Rj0/7xUz
bvwdIlsT+beuAQ1AWS4E0c7Lbz1w31n3sn+3rZoWFCSCQm+J3Riq0KS94vgoSeh7
zNMTH9m0oD149jxWflf3r5ClSPhIqAVbHp3r3KBoNlR58bNhELQxxrUKHaaY7lgC
jS6Hf6V2AAmTxQRSNA0fTTQRUwknWIDq+AulzoGvY74x7UCy+Eu4TE88RYw30Tbl
KHe+QdtaGFD8A2KBpppPcOqnZ9c9AOwf8kgN576JPtCASvNKMYQALmIteTlT1SeF
j/Rd+aWwoWwa1WQSujKh4MY7p05oN/7bSivXCoI/HGnZGR3pQCYhnKxbzjYJz/xR
RWlEDN42JIDsa4gKgwUQSDxM1f9dRvqqWCVSB8DEw+s7CE8Fvx/b2kCe8wPEHQDW
cEktcS3VnBVjp+xhCIQ74zGggtrhwxPP1N87vp58OjEqDU1qrlSizZ+ERIM1ublv
wUP4qB02bTLrr80IzHprIL7sCin+CPmTyEkoLCwDKW1HQ1fURxsGt9rsy8Vh9up9
2FxGCWCBfzERI5H/BG8LKDfQBovAeBHTq+LYN7KGeacLQbNVfs5bKjQfZKjj0Cyv
9shElq3roiAeki7ISNyl7iLPTVHk51rhuP1KxlJW3gtpUyD9tlat3DaZfgPD88GR
zl/a8mP3+vbmvQ4wqVoZ96vAQMaNvWbhYH1jDXzvKELfTk+pgjV9RonXclnht8Gc
QhfYUyeofcLm9KaVZP2/i50yW2Obep+3eZKzQUxxrS3FTEfb1jqlR+ifLnJJspBl
Zj4RCwQk6c8v1BmRldwszDjjGGU9jJcSUOa+8XTu/amCK3hSfhT9FWKCjb1kSIlD
n4ZOnX5LOO+6yB80qCD/isk+z8iUeFX1uKkGm3Pk4UMxTUD0w46Sfi1zgKdzdAv5
kMn2JuKc2YrMwMGhQnz/gwy2Qn7seudnp/gq2xpXAbUq5i7W5W/UQmagBqCZRZI6
2Y/YyNfORmu1eCdW5yNiVLir/fXjLBJsOIcS+rw6DywdiyzSHAa8DBD3PB5cJrPO
0F6A2+IJOZ2+fB7qIFUE2/5UVkrLlTT0XaR6zu3NwmRk82iNAN3VGJ5dqORHk2dE
iCsh3B94aMb+IZ0HWLWFmLnFemvNIwoAyntVYpCpzGuqSvJKc4/LqJpRtkLHoxBo
o28IO9TP1JfIPAQwhTq8Vwayk8cWlDR/BmO1p5irUvRAD+Ie/PqXbxBpPoDiPw81
XMSQqd2ceHfhJkcUhV4rcntt74rnEMmApHuN/XYNBFWaHOYcDULTjDmgWTLbFi7K
VidLUMr/bsKPUXU4ZrELk6zRXdZoH19H/KMniQHVZTXud/qkK1T8JSqkfNL7pAlT
9qzS8Fgi6K44n9KROWDSbdUOuCx6IfIRgYtLsLN834tWTa85Zan6Ow9mUgMpl1/3
OJYsE0ixs2eI7ND6lrbRDUR8Utks3Xkcw5N2sz3xRMOiTJAfyEbZxRKiykE/KrbB
QoPYjPiLmcSeFg3iXSviX7HtZQmF2GGgQbnQWPJ7cd0vXc2nJNhk1/Ztd5Ys05st
jkFpdUW3mbpq1dRQUioV1d86GtJX3rv8MNbIKPQDeY0rM9LCkoQvpiGvBJQE8HsB
5fejatx8/rsj0SH6FfgYCtCxV/CRBSW/zyN+hYHj83IVyQwMeju6CxM7yMXXvWq2
20mlFkdZ9ai7gZlh0VQ1s4LHZ7FplLx3DqU1Oi9ggWvX4D+4zTDTOqXoWyMlN+Rq
mVU5qGlh7gfw4vo3SHnCB4VtTK86fyNf+IJa+X5eWiHwkFnn8MBnAGty3gWf+rwJ
3sI24LC0sUcoIBVYnnMMWGHZbswi8+IorZGJGia36Km8ooswVn7BE9Yd5M47uHGs
UTZFebSuxM74AItCt1Z7tO1JKS3tsrNDlUav450kVWv1g5e7DqwTQlpYSbzqa7lh
QPWsAkjtjvP0XnbKfVvI7kq6O+BG/hkSJtZ79gsxVA+2R4cvHeR1phlEPPP+/3zg
apIMcZWFe0XKRLr7r4xTIZU3pcfEeuyqaujjhAx/mzDeHcpEfTgpyLc15a9+eo86
K1ufJGQI8178pIKMnWMkfhOXQmuRg3RQ1+9oDOMgUB/0EnicuIeZy/+1uQ9kw5cZ
Bh2LCcxj5NyWZdMfK6zK3W1hXmFcLm3BCmUBd1ME8Wub1qdtXrTBrNAe4qf+l+48
htpVjQDfCq0rrqz2bvYp4jmq1yL2WQa4dRweKDLYPTbvOMPnSBOAMTc/Hf5mwSM4
fOzMcmSdJKvWvaLA8I+b1L4zNfRcav+4dl62geujoPO5DxnQMAYDtJzgHEJyPWX/
y8hRxEtVrzK0yb8IBNhxuS3EuRlrppcwlf8CplwPevpgG3288ELUwDUL2y+525BI
YF2RU9Y/TayHDz6q0DhJnzJiPz+uUJGH5gY/GWFjFh37Rj457IqwQ9MPhJKb8eSL
BS2I1n9DvQt4mr39stt1z5pDy1XHutcOnVpM6Y+g4XdNDnsfDMOB2/FcRgYUrgPf
rMtxrlw2xrJvT/6oCYMYW6IT61aO4Z26yjPVbJUigppE8ed77g1Kfyh7kK4fynwg
zwQeZAHl4cVUJEJxEuHpBYn/VCHRCixGVKXqA3CHkWwmRV23c6+Jo6U4fARxmLgt
bedOszIzDWRl+CcqLRGLfGR9kT+oIT+gDCkXGs8cdYZxM1bCWmCBf4f4h95U84cM
V+H5sIBMnYtpnN6KXu08EHtRkh97tZVWMRTfHeQ5q/N2kgrP+drLOF7nAfuG4Hhs
UVsiPHQL4nSDcLDh6j584EQ8+q4iJM/YHqxol5WCWlTZyB7sHqMV/7K1cJej/55A
SQhjRuTmIiyPMqvyPxlCbB4rj0BtYqrLqmcB3YaQDL84I3xjWkZfAjzlh79lXcPP
L+7kxdQ2TW5u6MJWf7IBHx7fQWVmPZYRTbmNxeIBBRFrt+3R2a06wKqJSKiTLncU
6L0/qF2OmROs6REHcGCJ+yJVDPX8NeFw5kNwbXzEuoO9x0xUeTAwfCnRfJcgElLk
/+EqHTc1IzwL1FhJIzLGKUOmYtYgxSwcraihqrjFTelJPlznM6WqdQCY8TFhWHA6
VkkLuydtIHyu2sUG29lBKCOpcWCWzAUD2lsLPz8v/D03TNqGxnKcW8QwN3St4lP3
NDgvM9erTtO7JW/RAFXPMWlmv2pQzGhqaFUwod1rfvmJV522ABpPZziOpoPWHNSO
Tb9+QOwKXhAxHgvyMEd07JWkKNkH2uwdSiPg+A26yIi+s7EvgD9uNcz5BikFVsD1
C3GsXr33yQXtdtY4fwyvg2ZWVYyFivtfJPYpmxN9kXb/eimpAAT2aEH/mBamGCT4
8NNLTjQJ1PbqzizlTTP9fhXU1XxMbRCoNvti9479foiBQ7J+L218KCYxmo/Q4xXk
AW1Pvc37wavWPY8jv9HBhTaXkcXwgfnKH3jVH0E/EqspfY7IhMIghHMOzhxJNb/v
WSQcUtISgWRc3Uy5HCwP9a1gIgtPVFOziZ/MKqVPk/EIl/XEu3Eh5CEERYvpFeNk
Zkw4TBlkOa+7g2CTuT1Kvu7alWvJln9P5pqUhRNHmQx1pz+fQEFkuhyGD2uZpFiH
mLKPtPQPK4/pF8Gqv58yBkw/WrVMVJbiD88SbMCkVBYjoWRQGntozNYlBA9F8Yew
OwD2RqFqD/nrftVvaSvazg0N/Bmsp4zV6pJnnYhua3iz86ew3GJOstU0r/NC9iDH
gbMsUcRa12KGllN5Gp8wfo3J9Ob/lsvLEfyqCyh2npxj8LiM/iVvVdz9Eco2ty1I
o+Hk6LotKENNXtLVNu6xKp4+N4eF7OJfu/stYXXKSGFDQeaqMjL18nL8FrmKBS+Z
FK/OCHnYGCWrOpJ/VRL1ZqUqF+2Tkufg2LkINymZ63nFz+L2+nd0aHQgyImjcBc1
+El6kAVqLCnLL6eqcikoEAhWRAgbNcI6BPm25A22c65ki8ooBhQ8Kee2/2Xtl4pf
Z/jUTkW1oLEwC2NyuGNfA17CxTF+DD3q0MGqvLpXOUxhb/e56TWmA/xRE187sb9l
a/RPJLRFo42QtOTlE8dLkONr8YHIFoKwcVr3kbxFurqDWWVQvczrhh1N99K41Ejc
eML9JdGtrjafXIFKT/FfCUni7//se5MSxpmFdAeecdI1e3xqap62nzRj+IhkowqK
RdrBXj15vWSmh92YtPVvNQaELKDI3job4Wlw/eEBEVRDrNTipTAsUB/dqGscOSms
ZyJ1qFLD9tNeOsvr8HZCilcrq+3aK6P09cP8FBjWpTAFuBAtxGmpRFz0LMXQTr6O
qK8VKY9UNywXa6Whj5ts7p36t5IlO224edZByNBovJOQppfTft1KOC9mIfNbqN9Q
WX3G+ATJneHbkQKg+zKR6TtfJWyEZs62CMYL29gd1CYSXnye/6yFNhChc7PYvp5C
+7pq/t7U7KQYFBkbK2jYAEn8NPTYVaT9E8s2zAYEtwMZCuaNUJQXGgSNV2ntBXia
44TPGlG4nfL6Im/GVih+9r9rN65NXozV0i4XJvm4dq5s5HtnF10IOEfh67vYFDQB
sHThXVPlD2E6qTCqr14vboO3i3CFnZrR2bE/5X++K/PJi2MTeY9Rb+bHGG5Wtacf
mW1Cq26WQ3b76pg0M/FjLHdnrZs2ygLsnkyfRdm4HcBPzMLlx/X7JTNzKBk1+ge8
jlBLPAaqZdINQJgmr5vXOkBFVrYb6ZdgWt2xK4FaY3D/yemPOJT39CVQFjWPCno5
LRFXPPpvQWJCZMG9eXVP97UuTHchZprIJhsE1BmTpPVXhg9TDGIGRcvxWosal/p9
MZm0WuaEBeMF+jBbsg9l3hIlvlC9m/ngmzgQSMysNILjf3qSgdJJJRcl4OaZ/1gM
RgBIOzhD+fsrUC2x+Th8+qtm/LuM7gPAX4AerAyIw9v405fLSI9piKlP4UQEU713
q4JJOa8yFJXue4/7eVlYvAYB6kFrGV+NMgp9vPRDAT8E9iwvGRCPMUujY4FPQKmo
YPeP+V62dtiZO+jaMOiy9Who/6MEHY1NdydBxwNbhdSa6lWf1GZw4AA0S4WRssoW
OkiKYKhhuwxhQD14H2vK8JMmkrfyg49ztHt/t8EA28RP8T6/KPj2C147S5eBkyCr
IGLv9Jk17Ng9uMC0CHanUfB2RRbRwAATbx/uAAUg3pIogM8LXwNcjU2kqSH08omp
bST5u1SbjfOQ8Xka36qiXXdcMqhyGk/URt3AImjRUsdX0wgZjM7K8ziGdqQ+tRHL
JgFpeaemsF2UoStLOz/jWg5HbOvO4EcnZNFedgEgKpngrUoax0riTpLWhzc1rVnt
0DRiEjkrWtDmFwOZHEvIwY5yUlss3BvXVbfhJysBBGojPiSiP9oN/s0e3/wFZYxC
t8J0x4uLmnm4H2va9dWJ8hbidZeV33f9NBGVV+XYyRq2JkNhMDvPbU+Z6GeKRQEd
/Gfvol0lix13PWJDu+/JVYSfXCUFonoKmyO21c2LtgPQIM7oRyjfIAycerVpS0zp
bPO2SSbhWi/kiLqzf8lcsLKZr3FP8dMfyEQKaeLEeary360GBia8kD6CDpvm3g11
hOaJZGMtdJ34JcMcYgGm5LTyy81iLjm9JwnjNBFmhJk=
--pragma protect end_data_block
--pragma protect digest_block
f4L8TKyzlIsJYUvQnvkXnz4ROQ0=
--pragma protect end_digest_block
--pragma protect end_protected
