-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
ViUAzYi8nyZiIWgaecznzumxyPF68hul0gOyhOOVj4jsKuvLA1l92zxVP6Yialv0
EtOzl4TJMjIFOU7pGKJhzwupe1NP1megXFLZIdz/HiDlvsPdKP2A1vXH5foJigYv
tK0irCWk1oY4p53z4P9BuEWo5u5yWcCsATV1vhuq6vg=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5385)

`protect DATA_BLOCK
0IsEhPhohNkI3hOTGW3KcvQalzEkuCefpA6ZGnyJPD07CEY5egYkGvAj6jGV68+j
p4b1L8b3UsG+JsELJkUME+e09Nkr8mbIdfIII7F/Nme4bhuji2myqTcJdYymUC9I
X6FWUpcGGuGeyXzp/Qr3kEZOfkGpfuKDWeygPdLBQko/Nr1FcbGaBbFm414P8vS5
ZkKAc77PX/QKSdwIsYDjkCtLT2qRchpwm+d2aWNnOf5DUMPA7XKZKCakhZnyCEhL
pm4oF5Q9eEQUPNNWc3fOht+vcezWMfd+S9ROf3Vt3LBjcDKyQqAbRQ8Pfx2gfAuA
RjuD+IZb8tnkdxUrfad3h0Wc2bppP8+IjPUXmSGBqD6Lenh4gtHt+70J2p+eeOtO
xu9kefbdjQ5qrWLt9OGWNfLeh4Bds5Q4bfrh8gbngy9NM4vdV0EtZR2r/ShvOOs9
hQDLCMDiTRhoTejoSvFcTXMeDApqy5OnYZy2I/mXD9StTVo2avEQsBj9qs0Aq939
RYbWkPqu2377NYd5VbZPvbrSEYaGEgZbm2bwjn66OCJpmhRcYlvQvxNd8Vb8/QEN
u1oGtqBtcC+IvC58l1UmdbR54MVZH7dC5cEcRYEjUsFqU0k95CTjM9YtpHsJLjEe
eoJzrGgiP3g9UCRQGpnoI8iZ7kQOQMGAq6fDeiGIBPD6q3X23kKoDatErO1EnGmX
ldBuD2qwiZ6CcUvVxpF6zqGPcoeMF+WsPGXrsDMMolSxVK7vHnWRJNkmoSQeorBg
UkaDs2XRkiBVb3NcX9x+7GqtdjYJVI8pwgF/aMnhewbQSxQCMC0suCYtjDQDHIZC
e0hrCwvJggyN6+KXpSz7OVydx2QaTuOOmE3hd2Qqv8X9h0A/csBlOYF5xU9Fw9kw
tg94JoEWOqlWSMe4/UcWjKWhhr4hVDE5JJ1x+EYm2EL1PFu/KNgSnqiDbh1+hLFo
eSY2neiOCBO4Z7lW5FK4hju/Zg8Yeur3TBsKEDUXm6fSlRQluwStY/T9/PHwYg+l
gGscRKuQvPXksyK4/U6W0aXYPwJdRNhZMA/ztBc2aywlK4P8NrlfkgwlsaTjF7FP
UoFbip3VeeNSIhkGQ0tshLedvhFYplMgnMK7K7KrcMaqD9pnDCmc5gQ8Km9yhfx9
j/b/rAa4upFt91nrnkT6VFcmTzq9mIbArAkU6Oah+/QRUGgdRENDJAL5vwCI2Wfr
5gbHhHaNYDIoM3o9YMXlFAIC3vh2bzZorxLR4cgRORxzzuAVPByiJE94+fX04WmL
5LsmQHYiDqcjHeRpqnubW1yF8n/hc2JwyG7MHFbmOnYaVtsTjhr01Y/pkgwGaY9a
6cs92a47XmUXCDURHweavvNlo2ONJVs0sDUd94/MKq/0Q0a1fr8XRKmqAxk0IiYD
xkTRfCm0ULr7bofgGS82YJK9OEkJk0YFDNy64ck1KreTnpQovoOEdiMlxC42En1i
BzUZrTd4Wtja8gWi8Rs/zGJuqWnzWa9s2Jkc68zolHogmDrOvfrNIsd5b1ZyKLl0
rhMi/WVFjMH2ZdapA1HbHJeafPc750+msXvPoexV2OpjtWYFq0yy1GAnWlXpG0lm
hJMKdwQ6G9ce/ptDIhKeR9xQ7eay6ANEW3ugbNGxQsjVQIA+sSrM/qezYIU8e0gq
GQMx6FeoTa7VGQBF1Vt1uKBHS+O29DtMyXoHx49rxjh0uMqgR46TjlNFhr1H1PRN
XXfVIqmGZz8WGNwJNu89a8+czhXhFiFEd9vGuyS7FqzBxD6aD/+OzvFHOcMVG2oj
Lq5agcA3i6xJGRA9xjsdhpgtnnYyZmu1xxhikzIvWO9eaqmOWU2SvleoPL3FuE3Z
+zCnWh4jXeduYluAL+MLGNwtYtJGDIDhuiWZClFUOvTWOH2CXqHTqmE/auGPGxUB
KRQo+Um/G+vAiYYgzBGd0s9sOtOsa6oets9jniqTvfIB1Ku+dc40aZud+rv2CywY
NGXb+ilXX3zbnYb/70/3IT2BFZglUIgQClKBwS3mkD7+wZLRnaRS4xQnc/CMXpmu
+0elrkrT5tZk5XHXR83iulnerddk++qu+c2fbnBc47m6ENgoxpAn1v6FJx0Q7GWX
tfB8A2hR5jlUdN0Tps4d9e8UBHYcpmKySpe60SVLfho29cbtSgeVmLIZCbzPSjUF
/1Lx1JyhboAHY05aJwRTpqvJGhR9Umrvf0/E+1d6fTaqAdYIiKFE3sQg7H++97Nm
MKVV8oQFwNaboJaWkwXvKlCOXjHhVEf6m0jIrNJPxZTwRy0HIoQ1R+IRjGOznf9M
Bplenmz3o+5LnIBgFHo/+5LZ/eC1YEU2D0DwOfxsOgkP97xZ5xAaYfmcuqwig+sd
id6tnXYUEG+sm0euk2pyp+YO2cGf/FbmdNVz3uLshjO+ZlbWlhzsPGtNyaLNLoxL
TXfUcIBvXm/zClWceoZ0b48zeA22SAEVrc/+xgGnlSJ4ZsPKHcYW57jtH10ThTPl
WtwAinMNqJBD0Ef32VhttEbVkL2kPFcZg+YmSCjUsH27meFNS+z+RlXbrhwmIxki
UZDgC/8Jysf6+fNUhAbz6pMFPbkVcE3Pm8yBgJSozhiMuxqyBgC8YugkLYxc9SQY
L9rLp877K8/dtl1kcGXIK7GcNkOurrSINgnPBEluR9iRftRCDdxOoVbe7Wc2xd/d
0gbWxuu515jPHaWOVEmI0tKxsie8mCMn78MhSoPDKwnDUMrv3xmbD+5VDe4+wE5d
Cv36ywJoJqKTKd3BDqpfuitqyeaCvh+pEh43MsFflfq5d/ycIJjG/msSSAuJDITr
JZ4dfGpbq8xrFOzmEr0WAgRraAeoi+LIsoVNjmFSEtC3VV3XQgZjmrHUStnHebc7
1dFWXBbCDbmEpCUKlXV2JIQXUmQr/4IDnYxOZFNgAAJ6M5rDzzjzxOwGexsZN5wV
NUVQTkk6JVRyn80ljmNv73lYEX3xUS33X3YwiSriKpTq2pkvdJnEJHrJlM6hz0vH
ID7ceWSmWfDEfvNAfuSTKqVHJa3wi5HkBiELNpr+QSiPEkUD1DXXnIjM9CnuTfla
9p2Wi2Y+KzqKspXRnnQXdutG/T2w8B8mlyORsJNp3HejuK+xwisWBd07LeX8jxPX
b6AoB31OQ19CsoqzSoy44tlAtBMLfk0o2DRFIJKhENUO4WX8Sb24rwBKjYcbSGmd
V+qSwCg+RalrI9MhKEJbzppEYKMibnIp4vP4uX07Vcj7t+0JyD04FoddwW/4wQri
KACOZ0YeP93RvNZEi4BKW5jj9AjKs6zCwDNo/ACElhHvR0j3zp7pnS6rmSpKVCtE
FEGT6yq/Qz2y0UXGsKWdCGMMU9K02dQnn8v+zrjVkmT+TGi0l/CtQLaHqIfjjB60
4X+eSFrPKRKJbkaIuYqWUcv+4CVt4Vu0nyZtFe+ZTeopqcCbI+qdtLji9OdtbOUX
rAbC8YqZlcF1CWGLx6jZ+fIQ16nHtLq50U4T2Q1oeMO/H6oABj8/jMF7zyLFgPvO
6F/2bUs8dITS/UBo0ti2jmLjuKJVQOhiehDBB3Py/OUpty4dp7Aa/MtUd8LAVpCb
YjrU6LSAvtwbl2nU6jyR/ysV170/n8H1LBqigi0IeKtY2qZDmevwIPmJDH5JZsiy
QgiGOVaL4qSDZsLLtImxH/lgCVY9PwcaQexO3WvX0cJ+kVOvstZzw6fOiJKnbWHd
1GATmcD7Qj0hYnVus7hAjArPtb/nW+gGOToFaAOGn7+Dy3X8NFk+PwGFc2N9sLTR
/fmrsZ6QdyAKAPS5jjk+t2Q3KU9JcUWkmldSP/3fT+dpr1BlHAw0yG+G0vlK4uOQ
qQAi8PFjyT1MAMFgcQ4QFcGJQvhB9VxqmgrSaEEQM30PCpBECj+6Th9i53N6vIX0
ddjemfH6QOJVkkIcvopEaOf7VCfhgmfwICk037auZDGmb+TyM6lcHBdY/uf3r69+
6N6RnzOlXyZA+K+mbiBXlVk5fl6J3NhRxv+n0hiyDYnK1j+cchKoyrfMVPl2IVOk
4O0IsKf4Kb9zB0/IqAAFwslHRkiK0zYcJ4XLWBDGVpvq1xx7ABEFGu4ZSTs1z/tw
53fxIIoA7ZDazlC5LtT1TLhh5na0/wJ/s2qzfXXgS8Dx9LId2R409bOz0xgcE9Bd
EQUuO/dzaiX/gCtew/p94+yjdie5HG3PRWl/s90U7km61YilQCaNbNksvDss+LR1
5ZIcdEbAp+rBdVtXXKfNqoadWMGmwgIvZsBEIYj3rjfXQ1wosj8JA8M0+wdLotBc
h4rAd2kybFbFyiybOigvf7Gl9uLAL55FtgNM7XDtdAY/DGmFtJGKmNYnhuz5qMx9
JTZPvGwtfMlgFUpELOP6YyGCjsjvbXSOTWMc92VKuWfb2XkQC2qaY9Lrnh9Is/ct
e55Ik/KCeUU9ck0BT2pdm82xV1rOIB89TmHbHvXeX/0qCc4qfYo3+cAGtqs04Q8t
eyAMNbzPrVCnfCrfslWA43sZ4RGb66THFaPP/4k0iQhwt7YbSSojRtbY9Br6AnTE
UHv9yYPBCNMqxMNAt/7Ut5D+74aPHIO3swQfTXFSwHGJ9YbP472ZYQw+u34I5FRz
XxEcZhyJEvpUpsgkqprpn1iW7EpXfJyOVQTcpM+k9Ozmf8GTZ/WmFOhiMFK+ieC8
5rqXVD0bBnI1h7MpTck5Da9Loredk3S9qbT9gjNuilmZRWVpKGrSQvtC1WsUEuUD
NJpmYWcoF3VL0OleF/7qnwPtFTaRdMWRycMTP5mbPzsYTQ5zYyUovz8ZE4w7AZo6
0V/XsMOmIlq0jBPDdxB4mtUrQJ9jdEOQJoraneOFWpxwWahYZERNeTl1NOZF/TWo
EqJ5xtJpvNphgJjYmjHgRGvVnmaVYfe9DyyDcPBS7k9+zLDdZb3Fy2jaKXdaDo5j
NgTAxJdGyZ4FclatRxthrmbfsJA/WRP9M8IbOKWzRpMrg3ikCmo4W5bKx/Y/mj3+
Wp4yfXgyubMKQ9CrUqO3hIyfSr3ESpaQu0OzR4F4TdBfu69JI1E5fDnt094gtj7a
T1A99PVSo00xLTIS0AhKqgudQf1AfBn8Ymgw6ftdhzA++Fn5KCB56wmadRicIfWS
KCx2KqEgtbuxtXRixzVSjMWKOr6+nyLM7LHl+GA77etGfjXQ/5A17h/89XzNovD2
yOB31S2ex70+TNC/1frYmYz1pAXUBuZ22G3col2lopb3SSOfH6LTC9WSkBH8A6N0
2nd18xqLg8+Wbzjlld+JOw15b/FqeXy5gpupcVn0/bfTjbtbPVnb82SpueRpUBW3
962EqiF8qm5vSS5oxMa7hJXsQqUS6tf6xB+ot/xw7pz0sW57V/bAgH9WiK88fggn
A6PX4lZrkHxGpSCGDoPUbTwKERnh8B2q4yOOCxhOtGShqOD1eEC54TLnxt9SIVPp
XBtcA7oL5sEGQB5wGlj7QS6UOmltMCEa4Cux0PV70G/SKvlAJWPITDi3f61UNlYn
O1FwyYX0pXWkCXIGnRWfSPUzq8YjgDGyph1FQ0pazuuOSerTVuNB7eCL9DKLNixw
/FCFHW7WWwxnYpwkHzeJmHhqyehX/PmEwQdFqaVZ1am46dMMIwxJrB/QkoPhOgy8
1nBJouSrszMmT3JLd4Hi2UYR4dt0vaUZP8307rCur76067tQyYgqx/a1/Srm5Mz4
bTTaQOxnIM6sToetUXdMxXXuNq+zhC3a60ZdX5VcYNPGX4fpVppC0T+923314+Bp
wi+GkSRyE+qOdvxqxXL1OCivOsaOoK2fqYWUMnb4moXmEHjiRIqvxO1+CJqCLUtj
jClVDBS7wxQt6jdDJlq644C7ZBilugw7RszNbpDgg0+hZXhOnrtLlRgeIxJz8PD6
7BOHo82+mpsu0QH83hIrxOfp7CQQ/u4/zLYHOsX6vlm+cOMWfLdO0ErYDQArdl8W
u3jGuEMNMj38bFvfvtvHFQ/2RIl3qoacbD6nga6Hhit4+E8JStCt/5MojaYOljCt
4Ya/UUBgDGsShjr9be1T53uCVKFFCGcEqqg5VpUCFBxtGrwCGNSwEC8F2tf0lCFF
dJg9F0mzqxl0nRLEyLEeWSuH+GwlEEcCGu/b/hFtkSyOMhP/o+PJCI0d6Qy3be06
16xwf/YHiPDdpWua5NxEFgF7jtUgHo9GE0Kg27aqmK+v0fJVx9eoY05svFARZE8W
cYBooK8OJY5yHeRWBs3Ws9YorBoKgr7hpn8Nh41WD8ZbEm3YdUBKJMcHkf10V7J7
a47gSg02gKzgbCDgK8AqBpMK9ximKEzGAY6nDE3ccDaEejxIHj7PYmbJjoR4ZFWO
SOpupCKZ0BzcgoIi1GnXtvVw+s4hbENl2QA/Heu+vWgQ4n3H9a4zXNhx0wv11b2b
JjPfYsls72yeubVOAQkoEg2q9Z0NBWmIoQ2Gm2NU26W+1lPyv7AAnCQMp2pXBC0x
ogZH5tqj8KxS2LH6Y3eP08WJ3r+bcTkV2mK9Im7CObWqTLRIOuT9Q9BDGFv/KtyK
eScQ1bCZPKHQ5oMKHn3UJz0WZFLnrXP17KiZogTaBWkncUMYz8QL4PFYSRNjmVo2
KuSINI0ygJbtxHQq0baGueNf5wa27hjbPenjwMQ/BeU+WHtU2eFY46GXq5lLN33i
MT2fbkvlO67OV/xekeMQWKnlCLfn+RYKoK6QLyCgu8E9UnffMFTfbhISbsqbz4QH
FqOXnk8T3IuZKlNyJsCG7jvpwiFncSotLYAoE43HMoC+FjgIP2xDscaJln5Oi2dp
X30dt/zdH8pXceOgKNcXle9losajDj8fw81JENFhg1jZ8W8pOvmwRCWTLfy8x2jJ
Omew5EYKNRa81+ho/J7CAZoxRZbklTO0E4tKyOUdeM3xiRaCqz2khM46wY9HNNju
OpyDFpQLVMLHoAnr77Ovo0ArRazVTASHcw+YhFRsVTG83K7bKU4gs+jXZV2xRS8j
kOmPfsolJ2Lom2Q6HZH42rHFPP5R7iJLpZ/Fp3H8+OLYNkf2LU57/hM59IRlIv1w
w5Dwl+ewi2vNapYoPG5i6BPhYvbVWTcm6RXXWo5PjrRxOXoOVTD+Yqy0ZA4Z9Swo
YK52an6RgpjMJHATtSd1onv0pdceh3qDqPRLnPxr1t5t3mqFMFjUr/G7HVJXMgFY
070FTzM4s2sB+d9xi4RgYHI1hNd52Z22kCNLzIMPiJs=
`protect END_PROTECTED