-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
lFBRwxNe6kOviCO3z16uHglUbmexUkxH+I0QWOkPZ2Y9sRDqM6/JxG8lHVfdKwfO
b6waqQLb2DXdQhTqhzxWYAtgvY/gyVDCshZVzr3Fq9ToaQXnKz/pxy0Rrigos+Be
kgqyDs757c8Xa+hIs2mNgQI6IcP3pdTRTbc6fr0F2UYN903Er2SjOA==
--pragma protect end_key_block
--pragma protect digest_block
xq+WrrwlbtHCkbSvVP5GqpaSbSg=
--pragma protect end_digest_block
--pragma protect data_block
Iom3aRUTPkMafnZ8s5GaO2Qrhfd2bj+uIo+GYZL/YrTfcsttsECttO993Fm+xW3e
4U5ymfTf0MzjHV3mYYH8ZZsb7fOGHjywv4Bo223HQ0wgQpo51hyO9msv+b+kOc8d
oJiMOmmdedh28WLrVmwVZsDX3hZtlk23pCgOZyokKTgxr0A3QGjfw7JHQ+1oR2Ip
ZYgCS1+YvKvXPUf8aPi1iJWf0wlDdKdgLWS9ExvEeKuz0ou1fmaJBaNU9KsqcJtt
8KNANC/wGJeqP6nM2uVu8Qdnjhbj6NvqoH3wQp7lwIW23pBVAcNuypzyekU0TBfB
3yh/xGt4DDZttoqUwkuznTHWo3YJBXh+Ipp1rddzxgmbIhH6BaCEDQuAhNvG73eM
7VobNYFvRxQcMb645Q6oD3ZBXOhV4Aejvqc9OJjQsllG/isT9wDlPCPJVWqQyIM6
1jX5wOQ8uhGJqEh7OyLLTDRpGWFopymFWP3kHl0c/cUPAwbHgtxx5sme08Zb06o+
ltIvLXa1IyaCKv+DWNIXW/OZJLui6HVoQqCpjUQezrMIx57okW9PG8PRcJd/ej1N
555wsEiOuE6hADBkfj/KUBdYTLkFw8mdOWigYn7A2rZ0m/YnkFsPv6OCKeAZ/shT
gGd6L9QV2BF5AgW39TWEdIZvxU5OpouUmvjqkr+n6Opuzjxtyq1ULA0WV5bb+0+R
4NGLkh+a75+fJbWBjFRCbDFGrfMUZToK8IcFp+eoTm9PYpkoHM/Oc0SOZ0nmgo+I
Rhu06uQ207BNITs3pMGWGjQpmfQgvVahDvt+o4m1Lnfx2djebv/mI2E3KDMqzHZQ
45qC4MVtV4Y6qAb+PA1gCSBJ6ho4Z0KOpaqYSTJ3D6xYBStg54wy8jHFG9iG0Smf
thVWQT6u4ScS/n3vXReMnLuCgx81B/AhcEsQcj7iWwjepB8afZv5icub+mN06NGT
poz1SNClKTBgMxq5hH7mceFRn5kPViDhS2odu8ye6y7y/cxwhw7QAYTvSbT7ozwe
Qjzg0GMx7tUpB75B7iNgfZdnZA5TqHFs5N2llLfzExTvR5LBD5s01IJJrXxxRzXX
YjBTjY70oXinTQ6D1FoITzVZSVrlZRDrmFmPWIljXF2O8v7vvfnZiF0+4ZbAwFSH
d33aao9DaA+nLvNcd2GfiabqKBzn+QcEttQm8f+gqi/Dmt43Xr0v962f409dfSN7
WOBdqVLxzfyqJ2S497rZnGlc4Ks1ZtZtxmskiiF3fWhVfLUFKDywhn1CFZmYZMCU
INscOrgLl2yXdbTL5AyukoypQDE+DK9IUpPWB0EnwjDm7yJ+qu/sYUTJyn2kNqss
n7CTi3gHP+Y5OSrSvL/R/aKGBjZSL5WMK+NSeZlABomMLzM5oXcYyZ0IZ++8bEtF
iUncPZRiXQJOXR0De/9QQ4PyFT+vlZ0BEUvB4gG+ek9RUDTLZJnuWH9yZDePG9t4
0953H+QykcyzslMxx3JDyC98CR7tfz+Qm80kHT9KCCwEYN9T40O60JfWNLUphuXu
i819Gvwsc1z6vQmLIDzAdCZZ5XFvHOztcf88hWnA93w/lmqIysvaim/arxk083Hw
FWNwXKanASYyedShHqTc/Mw3/dCub1uzWlDN3DRxmxKBGgC+35kMl246IXtEi7At
geKh107KCMY86WQ0MhaE49gGQ78KfZYe6pfl14Y8rJAPN0uBLl9KY9c7nyoeuuUB
pmAD9oKhajfbqT6q6tdXInsob0v+41Pv+oscyy5fOzHWO/0jEWYdA51jS9Wg5VN5
04iNwxq7HVgs/KQoT8h5Me/9Ia0jv6IY78Mmj4IdJP5kD7wyvr4bT0RyP0g+NKib
qvuw8ufOrrHlScSznwIA+oHxulm67anS8Io6deT3J+ZyEsmkhcJ6fsgv5B5iQQkM
qpnaERzzeA7DB9D9CpZWfI/05hLl/dPYvDu6e4t/FjpHKU4vCRB+EFcwhJGURsm5
sxhQCucFljYu964Q6kOQqunrKfhBVC6gfQf6JDCV4UbZx6rdwvkx2y3ohntluo2R
cNeSFjCeQMAP129nxHIW4NcL4Uix13xuPe7R7wxNlLMK5IMIaXfYtjQF9StnW215
3+nYx/ymTiItraISvhHl3ubMyPld+DSpPyASa8vvPR4K1fehYcD7j/QXCyXCOXe2
yUvabeVRBMNQYAMRPgSRF8ev6tupUZ/N/QIKaNnNgkVPvZYkENcg4QnJUEDDD5v5
6O1aeX7OgSaG7LubZjc7483VPQxnpAN3VNDaS3uzXBjhC6E641eqDItiwb8+RhSk
s3zQW1MxQ+PGVkwcx3p5Q6TIaysoFCWr1NSI9EQ7+DCGX519orrU4j3tIaR258F+
kdxe1UGET7Yivsc54wxfFF25D8hE70+7+nxLD45xG49NSHTUbTEVqg80yqsReL5G
siG5JCrdBhr2pxJ7Gq70wMyAigZ+HfCC4pFshLXgCxkQE+CAalBmorrgcplJA11P
KG6YtFoFdjNPz7jYa7N2MRSoHjqLEyYPWK21na0zKumO22QxnCtMGAIC/bu2eCcp
kKB6hcXkB6SwWqIbeu5J2s1mCZzT9yYt0mNA+Vie7YASf4acihudBB29rFDi9ed7
rW7zMfSpbjQ4Q/HtIOE87luK7yVZbAtxYlirjanOCTTLfynCp1AKxvTN9Q2tisXC
sYNIce9t+eYUklzKliC9LIE9roHwtYCKtWfuU5kx3qlazCQseVmAoU6S+KrtlO8y
eQYEhYrsZY2FNe9muyPpfxwQk7Pczk8Es7Tu7v2E3ZkhfXEDh90iv7soYP8DjpId
BQ9+FvAU3kOM2+xxYUzW9NaMPIvNI7D/GLHaZEMv3ymXm729cO9yBd9hZvib5NJh
Izq9fCzpF1FNESGqSWkTPe2f1rj7Bczo0zAl1sIGDZ8idi839HZPK73P50AJYszz
vi2+UHySeK8tly5Oyy8oC85Vz9TUtBUpw9JUgE/dYAphiEbGRRMgTEdI4wWYEcLN
Kj6KGrCM7BCxROFFX+ndVXSSZjyTRfKRMydP/kP06XZBfjAhnZQAWJ4eGQfzQsC6
rcXx84lQg9C36mb7SbJ+PBGl9AnDaGAY4Ys7kWh3gPMP5RtPPiw1I8LBCZISCd5k
ZGTOF4noxioTKV8jlRlrGnmDyOrzN9NTNXAG6wHaIYjvmhBDG0Am9NXZ2D1o6K1U
bbGdVmCBvhfr3EYHWsQXPmAnhmDY1PL+LD4Ziar7SQoWR6veiw/Z/CrzpSj1Xk1W
ybQL6yFjVSkqa+YWacKa+zrSD3HQTIJpb7jAUZ4bXfBoRcBdDq/PJ2P9W1PpIn6D
5bieu05A5mnOMIMQhSIqNEf08qrM96wgb15UTLbmB05SJeB6d0o6Vq1uc6BkIuyZ
meFhi6jBoqH+q2KHZh/LB3vuE5kFPHE6zk7nfZKwlz1kemw6eOjoNFJ1LG2lL96B
/eAj7nBXAbGmE/ymIlbRb6CB/lN60MA6C4x1N4OxbkK5oi5GczLJEnDBY2zuLVIN
quoyy/lzKcc2VLTFymzk3ZBxkEczgVQkk6NJZQzHWf23Cm2s/lTExB5x+KbEcKNM
4EOxtzP96oy+iseQez31gvfluOcceVm8xM4bd8IlPGXnIYnBi9wguMpHe1QuEz1Z
ncstF3qp4W2eID0r2vxe6Aa6aIPcygc6aL2K51/cQydyKbx91p1De6sesbi169tH
djuXZW8U2eNOrVsSMSNeKbi5p5+4hRCFN2FHMz2Jtlxj3bpmOv/eNLQSZ875YaNO
kJ8unyPUjnVec/5Hizp7iAxCBaKe13gQEU71vuaEFqzvmyCv8VZbcwHTX3nBB2/B
m+9rsoWr+EPomC76XeTRYZT6rsjSVwE0kRr2FJq+orYZOQLSUClj//cLIF6vpKkd
MQ3omqRYuaZpQzmItuL2Als15BbBWzhyDPwGFYrmsVAXDO1r+Gy9W4f/SDgvyhYf
zeh0XoTugAX7Ix+BTP4SLQGqjMiBhrdEodurGZDlie5z62ooVrAFye/2m7R2D2PZ
rIPITsB5PabZjH2aemvpZ2LemjnNQH+8rgZYMBNwrwdceICO72KN7bLaJZfC7k3a
62Gea9FG64vHoSGL3CRS95FnMoBjQPOKD1qjhDazFYM39h4sBvwziOW3eVc6KnnC
7oFSXVvyV6AO//sqBEnW3TMoHOdRyObTBKvbAKM7LBnDlcQuocIBFTuOtF4Fs7z/
P0JfO1Tc0Ilcmv0zw3IcJ0z4x+AVMcvk+xNP/fQQaMXKvcg0Iba+83y26WaliZHX
DV8pPtUA3osG+bH0emvEPlAEpWGf8IHQTu7Hdu5jjgyFGI+xttR/rt9seVMckGAH
+PSzAuPywEcqFfH/M3+/04esYSn5ptJaCDbHO6KUOQfj6o75vTfQb9FtEOb0iGSe
ASy0F5dr92rQc9uo3dbXTcsS1nYXyZGbklEa6mUnCw5f4J/Awb5ZN+jFjceq0WAk
nksFui7XC1N4Ea+FYX0/4QfIiC6CPAJjcpMd56xUo+FCRWUg1I6AkNoEfzZAPtXZ
2jE9hC+aFqLSm/yzmUBwHZ7k6RcaguhRdrReiZZe7eA7ZRUAXyFikKZbq219WTTn
Jh875eLLpsdO6oH3lK5zLEkpYJ2QW7D3ZNM9boi6E9GK2DqOkev5PVfBs8i6/WwF
m3wXyxh5DP5cATQO2W1+rwgA4S68iEJ0kFQNB2Xrn5l/l+2qcd4gO4RhEnMBfN7S
BdlxO/BDG3FILHljM8jZevGgje4aTzXhsjjK6WSjjls=
--pragma protect end_data_block
--pragma protect digest_block
8BZfVjVBvU3GtLTziPz/gUiFZJ4=
--pragma protect end_digest_block
--pragma protect end_protected
