-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
HPR2Bn9/ZJR9ZgAFCPahiHngwDCgVxjBRz/GoTppMKMiwxB4jKMAoal5ocLqfuOGnbe86lRzG4zU
xbYYQ2ga1HRZY1qPsAhLlp6UD0kS5rVIPMjwNH2QP1ikKtJAZnB7/yGdp3D9QYIS8LA7j5Y8ttru
IIrzaD6Rx7fPscBRXBmq9Lanp7M0+YESxbtI6vrh2VkxQrLTAu/Iskl9/HkjVgt3ivWKtOr6+UO/
KcWff0yk26gs/rbKvzqpk+VrvGlYnaNsw9GM7iRnrZq+qSjNbcPWlSErAdqfpwFcxNgbkR+XGVA0
+U4LubLFT2NmMM2HSOF/1xBzA20/iNeKSzPLJQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17152)
`protect data_block
dwUZuMoeB17v9/qjUJOsaHNh8pvIi1LyItQKZNioX0x0I32EpGAk7ik14K9z9FK87Wl+yjGUFTGp
Gz8VD4KUu/8FZO9fcmOtepu+WGnQRrAukKgUu9FmADv9aukhOD5oax16qstApwPB7DwLmSXiqyNz
qmtJo3PP9jPL7pT5tIfZsDAgTHJYkEKfOlMicb6vzIX+XhQQk1Guw4h37JSYcDo+D7CDwGezp+45
duRq5B0iT2nCx71izTM2fG5ukpsPcQ6U7W3z3m37hhkQQ+s3xrrlNzvDO5QQX4RQTClKngj86l4X
10wKyDWy7SXYVlhlzRDe2NAJxqt5s5m+62YgmFXmHhZLYmMASLcnc/+8oBT5xv2wAhCtXeiNoeLl
EhBDXZej7LK9pzslPJjKRj/0lkiZ/157NqFd+Mz8/CcdsjIMMDleZePaumaob+wPxHjPXyapQLd2
LredDExKJN0oEtbHs3gYkeUpz4D3vC9ARx2EJy7HDThQimgjcKiDGtpoB19ZCezLLmRiYf9PYfKG
WfFN3xJgpQ5Jmb3QA+ARLoiXMAkKVEIoyfr+YwcFwlf+r+NEsi/78uuSepED2ItCjMnEBJ3XoOk+
suSObp+UnLRx5zwg143fc/o9kOJyAMjKLlUGvU80lv9iPyd99EADwYMniHCFPOW1tRZwDJRhsjR1
XbMCtkmO7PWaVXJLl8aLKkKfNtYgE4afqpc1/FX6Al3W13vISYM0oadNfIPBAwYbY8hEom3f7MG/
uzOCWUHs6Q71oURkMZv0aGqq4I0dDmfwruBDrbKOF1fElhtC6eHb7S24PXRSHDXbBd9y4TtN27kS
19sQxCTTPvj9clQiKrtc3QJpS7MfL1lDBt/UjQx14DrVpcSpiDLDXzu7is0JjdCn8WmRfgWb/kTT
fmrlTC1bra82eCiuhNYc95PeoVqBH2VTqhitqRNKkByB/s/YB7fIGq99gj3DgHYCCI1NLiskPrnC
spLpkI+iizaW7J8xoLPGWJOXAalfeeuG82lrSlwt/Xw5BnnJFirhLI1IM9Jfdf5KYvihT8/sh+ZR
TL+W+2ykfRL0vYm7AvhtHoDnEs3hfQ5bTWXHKgqIiZEIRFmibPIm0dnJu5HYPv7lL14fAB+sAEyE
Anwz6fBU3zhRHvcYaZveHXcDMsKFqBcVdWcuxFACyh0N6xKr1tTbKUO5VQc91Vy79KIjQh3Km+GY
zZDlNCb8jNUksGb4Rm+Y4AtNCNf/DQsuYdKPfFeQPSkMa+RoRB/Nhva6p+KAKhQQLeYt97kKP9+6
TYEZ9NKc0svzWPrLd+PKbaqJLAAKZ0ziz4L2zrJ5ACe5lZiqDOngWbokzsGqZmDojTQVx2ThpFPF
63hS5RZBNJ1FFKuBykkEjzxev39u9nmiznhJBtHDqkd7Y1B8c7k+jADyB+lcikDrweGpYFA2KeQj
CoquvOPVLqNN+ffKdJ5LQQNo3ybvX01pyZ7EWz2GySWYPC89lJfYoRqz74xLIi/DKrhjmVhDeJyP
ovjJCOJhgH8F9Wqe39/JkQCllEfgPKOmPF15oVjbxCVO0Mqzd50O6X1EW88+5lSqhJrgXwOXcKck
/km41h+UJn5vYK8YWNcL92u0OI1mpCqZ+quGwFOjjCWL/yo8cvZx2JepHFveuzXG1hPEwMCuKS0B
9UxZ8n/poBt/Wghi3mzubp/McBuc0r9HSCKjuuUi9GwrPI80WYH+4yiqpIASg05ER7ocm+88aPIg
yRIVZzT0po5hM5mlNRnmw4KwQqWLCkplhgavWhMkPP8Y4zfYe7irZz3j/vQruhvrIxz0RPdzkSq/
9e87SdCqQTlV5mtbc18fRlZg3rY9n7tXZhqVPEooV4F52yfkT4GQna/FS0Ui/R8h9r8F/Yth3eY8
A1ubrGPBNIYw7FlMmpRumGwsMbJYbgwOE+T1YSNvR6OC43qj8mj7l4+zxJ4F5lc6tjPQ5EysWOIr
1vp6eZmy9F1dnedvIgZ50vQcA/AxITHcnBwFGwe8iTFxSUUIn15juyVcBX4FKwEC8Ahkx4YJ8oDA
TNN1G+dbQsjLjE6cJD+LRX34qeFOW7gkgAABs9AUHRdT6KRZQbfknnBrYQnlO9OM9Pv9mcEV9Od9
XkVzQ+Gn1k6G1gfBr1494g6Ulw4Q1DEwsEuiMZ6dmQAdhBmOdFzJbN1jbq10xtAbVN0LpFAQtSHa
A04HP1H/GY6dlF4Ad/WRcG+i9WV6zrxZv3vnSEHHjPHBFQUZID0A3JTpDL+QYKX1dHciG5JRnYCG
mWgR+97XVDQoYjBgg2HCUF40pT/S9CTDyM/v0bFC2BGzv0Rq/jzU5qXHjrjgwqt2RafCljasvpd2
lJg4QA/Vobk6HFlooj6ZL9qP2WwpDP0vaoIJz88Flhovqj4gSpsorr3VoVSAvkzSAAZOV+9qoJmL
KxfIKkU6J60bmXsrnwRdfEWb6nEbEv2cSE/WXwFfu3KB4eWs1yLrGKDRq/Nzch/wJTo3XnHJEJIv
e/DtIoRJfGRypo+XvIkMAntkfntxEkkWPH9b8Va/k/BhKZO0/zz7bjThhhZWfjy9g1LfqEyG9qNj
IQaqFR8lXwE39FQBUnKffHrxzyzOoErzK8ondCpQYPYc539rWGKeIssz+ohlqjnJO6NQX7iGePfm
nDEUwDfWu2+/WBajasNbi/gR1UIIOXIN7UycvNeeqWg5/3yQWJPoPRvSCAGs4p9tBGnrKGSQ2fUS
0O3+ABt6l/6hF+Ho9PHqKKzYDvXZoa77T41W4hSVuqE5zExUSVKNTATqq1iofqOd/m0YfMOTch4v
rV/5RRb7cHAzKKV0pOafyytRxEl08WxINgpvcYAj+JlyILhgJME7QV7VkRW13SGK6OrspmRljQsY
NDcAswgJj6gkUJ6Vwd48C8s4xc/xKELnos9LVBdBoPDhzVqttu5ZP0S/3AVzEpG92EDZUt67XyJY
02X67aSbHXHAUe8ZSBUa+rBYBtfFnezpY8pTM3BAJhpx6kUWHa3x87hLa0Jsv4xeeZSLoWE/HiW7
iJTZPs/tAmSGHiSfS+VF+u5cH+WwYQ/Xgsua5sIIGCeEdQoeCQKAkdoPGhx0rBQGOvs7pV6kbUBV
BActQBcRP6ma1kYsDJb/McoRPyBWVghmouIRS3JZ3W8EUGUTGL3oeGwyUc+NnDwLefoPSfJysYyZ
qpcsogkAUiacxUSykSDwh8iTrVW7YxeaW3g2Uj5YnUlvR1B/EPJKYtQcYF8aex2tSTRhsR+oj/E8
+FJg35hQyJteC+Zz4s4wP37sbIPGEa0KT1XPNtb4p2/Rfa94VZXx2Mg2nfRXOMxz9+ZaVgytrjJ3
JDBfLzJp4/dl2FgoJa+jrAWSgDdZkjpraPXSdcOH9cWGRZuPcMiGbhVnIwZ941g6jmTwjh7XtHEg
0ncVgWus4DP3k7UoH3gqbLZcd7Z6VGikqYBX/7qjXkvSXWq7vfadHk8qTH6WZHI9WCkofvrehxcx
U1SlKA4lGyMlMOzfkup0rJlMs/NtHTC0Lsmr5LyKcUDF/ZTusquPuHw4VGUapVImobegQvT1nqHw
hk2d3h5qHqPd4KczZzPEw9OMvuRqXOAYU6mE4BdyeZ/vsdOLQyT5dTpu+1cUaL8utgXUFaxQiYZn
3X3fTuPn7t64T4pYhM9MPtX4d4fpo1fAOdXlhVbiWmnwxueaiMlm9xv6mAGR5BFRDF9x3jEWhqqS
6aiZWuLTVhCInQbi/t5WE8qF8MBDQLiMR1zs8SkJHP0zODOiCIdjNP27COkwTTVK900NlWVs1zaE
mBiHpV7QDf7LgzpeSSdJY0WbtoGogR2zB4a4LMHIB/VaW4HHELVLpcHRGEgiHchcSAL9PZuqvHhV
PDWdJCBRifVbekG8BtzV2n7sjJHOhPgXv0S6VlkjDfIJQPcMOGbJiDTlzspYpLlxtCxMh094v/zm
+t1cIfrSHsfaVDMGty1/5JZ0CrzwRq7mBP5RGmhcT5kaJcrEQsBMWfnCvtbTyivzB3qn5kMF/wEb
STbMn+tiESQkIwGIupEUoo982JOOmGSCJGa28Vh+cx9eyXm9Rk+wujDvs8EgMqzLQ0EGIvaNFnQD
+CAz27DQ5znpbORJG92B+SBsbCbH7HE+RM82KKQVdPN1VEXFPDF3OT1ingjd34J0CVDFsOtfSjQB
WK9w7ljBbGKBmm8606OG0s3dgMkF5t0JqcDOESdNuV6zm/nC8w03sKeytnngzXzswtN0nMNji+2z
UjVFuD/pNZFtz1bHVi8t/j4lhF/ZNRrXa6ltzf/Wjnt1NtQWFjLSEIzg3gqaPLPwOssihPuoeb34
NKETfijvzhlKlrQX5DD21YudNZawtIi/2b7Xkwo/Ydbf0imDlVli53Yxk6xi6YejgfJ85+5/mmy9
okGCpJfSAS9YsZJ17VSDbGRoovAJ0LYLIaRCcutnGemXU/JfQjeOluvBrRnKdn3UZf3pY5o63pvI
8rKmZMAt6IDsn3qBxsWIEXtJm65BoHT0xV3KJ6jZYcH5ACdvV47TFz9VVrTwn82Dsa3eQYNtl6DS
4NsP9VCGKA/IAN7GMGPtFhXNCMaR106+boSZJmVEyD8XfxZMtCx9LqWdmxpj2v6Job81IetXRGnz
5RULkb8tqYAnX8/dyWUDJ7BF7xVUVQyIWs7R8K+/XACn7pEvRGeD9eMEQ92mG/NE9NWNiCrxtbC/
F5luV0B6rQMRClh6UV32t9cccJLQv2Y/S0mcHZdUq2xRbFnLJ+vsp0GBdK1FVVtRPGScWUVW6+Lt
VIxwQYiwKVwS+2hS4gUaG7mgv41fKEiKRacrZ8zT2tZqNFPDW0Xa+4liOLwID9tSb1uj5ej/Ew3I
tcDLZxXU+tk7aWbkCLLf1wyrY46xt+1y0csLZhJeHrQk+1FGqJ1jxiiWiZInY7q+X++kT8idCT1I
0riZ63zliDdy/SeLYBxwF0eQvMfd8gNNqrv9vKOhXGshYdZLo0zDPbD949k6HFiEjj9zu+lnX/9F
bL+Q3HiCDNmTl78baBeVvaHjBWWg1AMHe0ZVic7/YopXy5Y/po/0BiLtwzMyphXRz7IYQSd+6ras
cca8pEA75MS5S1bacbO0r/qClxd61ppVlxuyZsW5eMK/jrz3gwp+WQn6hHrrEHYYk5StLvM2Pcp7
E2eTJznx8shHB+6D+bVVrtf3i2mOhCxAAHtzPZ2AAaAySKRc5R5j4Ft8Ad9JNjOdvdKGowHP2sDC
T/fvrl6WFn9ms/16QqOcbcel5uxCHIW6hDMZ3nlPGvCkeMUjuZtUuBv6pOaj/ne+7+q5B5AdNiEq
jw+8bsq3bBxu7n5vSmd21iy2rju1lBHe+ku37CAMx6uR30vahIERG9bwuQyQnLzLyEH8453Hvs5i
wWA/1WsBNi9gHDztz58h7n4YYETmA14mhtJCqQs6TBVLNGh21OeC5e9pZd+/qnkTk76CnrbMWJ9c
TxdJ3YUhnDPxeP+I1B1Oq1hDWsFdb9/c1zQPseGVkgzdpcps2q/X4oEiweJ/Zyky9TCvisltdmKq
dOOSwqRJKNsrbJGP4nz7LrRWB08EVT4ag9Ryb8QIuj6KAjgCK8Im/VZ9fBVqsSkvhd5Gzj/Uan9A
V0z7bQ2/xTHIgNp3keG9l4hX/bGyGH9FhC8mZg8R2AXynLHjAKEVYxGrRylK9ISqNtrvJgtwjgKS
9KvkW/M318PDv+zQxLRnB/Wd5uvCaXd1IZ3ZCGJqssSQ2TBeOSncgCJYsthqinfhFIg4hUmKSzz9
kc0JoSO1N19VjuehDigtE/L0lrh0Rn3BmPhREJHf2Qe80WHF0PiDiHwApQwGVS4G73ILmaNpCUGq
rO7o40QFZl2FMav/NA1K0Y5VEew8jEojZWs42MtYvFO9d/jbsX6FYKXmsALz4qhi53sB939v2bGz
XDZNY/Zlc5KCz6buFaYdKEPDDZj+Ut424LrquzR1lSPX/4ffT41hAI8bhKLzixB+0/SSXrgonpQE
cH+V0rU9LQWjNyTWUYGh2sAnMYbTRaDetYRxhrLVXjqiAkooPmqpGZ5Ds5ED0Q18SgpqWkdbEsHe
uOFUUjphYmYRdyflMuFZ8tbXVfBL+2yohEVWDkeVzk/7EX1TxnRmuyrdkY44o2DGVNsJuXc1NXfo
S9vfoCNM2AQ+1enVlvH7KqUXr0D3Z9gZnq24J4RqIfclMLAdSGxxIbYFwDK6XuamoKw3HKpkOVTu
BNAAIIKOlVaZholsm7SW27+F7lzjDeHSjepBxnHYzvoH7ejsCcPRlwecKsRgqT4iHwHBqQgYTSjl
FrGgYBDzRTyz2bH9PAMysbdfnZoHv0UIYTWNDAsNUZLGN9xysj8Fkh35D4VJ+bRMYEXIcONOROyg
vfo6PWl8GPh5he5IKDPz8nqZDyWZY8eJUO1uUQEgFlXtr7YBYG3417T76l2p3NwvpuvOPRWzRezb
8HWSSp57Gx0CAosvBfI8Ix78fWyzmRTeXZdc8CHbSFPWwW+wR+oWK7vusj14OIVeiqnTVM1dIkcB
LrDibMAtUWHYyhZzJ5Kl0v+zXBn90LwgctOEgqRmgCmygSVvLtLhu0561QmwNhMKne0uKYr7I/AF
bt44NVeoPxInFgbvrbc/hkteLPHCEnuvdqXSvEgBBQFfAeTkx/WHuTt6ch0XAWtyF0z/plUBV8KJ
xpK9clPb1Qv0UmkOJx9SloXbF4mNihqN7Eo+2yp+gpI/V6S9CTm8nwQQAPYel/mq3UJhH8U131Gx
Wl0FcVMLn/v/IHqCyLOnhegf0WtpT+lBKwAHZ3SzzVrdVhIHUTCaxZlDcRuE1Praw/HIZroP0/hZ
Lo8s8J8dd5H/9extwrQWCdRmbBI/m4DcZ5E7Eg1t49hqvxiZPwNb0f6Bhlft97Tr8ESg3HhXr2V2
iCu100vl3+3MfsKleB1VDpfwhe0MTxOOd2OL2sxBHS2BUyoGwVpQtTB8iWwl/3mUUNKtk6xBcqwq
tBuw4+Qq76DPgKgF2WeaRxmb/1QGMhNFPhF17SmIjtfdty31fygS+p2gpC/MsQDFNWKA4Uk4vU4c
yRRYxuJnR1hlJn0spQCSQeG9z3xVEGbeGcAsCJZtj+0RrLuQSI6CWEn4PX6ojOoj+H4O3/yu1Sjj
Sa8XUOWU+iJ4gKOkERvbfd0TvMaoqx2zIywj6IyRwPd5ai2ASP0Ssm3TNVFudWklGO8VhuhzXicX
+DqQMZ2tmAe5jPFpKq+sIx4p0DD/7OPQRiyDLfQ53kXYyY5YJz9s/VvqyaCCK/DXxyR3Phh4weik
h7XpJIoPLrIKsRqZ9qAmVaB3AQoBm+3RNpy0KVd0Tv0YosyNcSiosvMP9Zd1oebX/4ZRzMdbEngR
HEuTReJyqIqh86WXnpoW+yw4DVVcaeVqHRaSdK+XnDmovZhuZv4ZYTq5I9jNHFTmRUr8rAS0KEPf
SdzmB4Dc5oRk71lVhKfvEiTNst15GIR19J45/yfyioct5NK3JVOJOXs88CCN8hqGSi+l5KQ1p2Ku
j99z9gBx9lrW7uPyNAR5dXWNqzkdl8mKhaoO1gEGuibRT7LZJWgWAn2l1VbFu80ryQiqFt3vuYTr
wuFFNS5REtg0ZaOReMoKg+I2BdkiqvTaDw7SLtZO2leTp6+P6GdcycbP67X5H64UVxxYnUsEhpkM
uzrytgSTa0twalLBJOmOcyS199V98vKyIon0kJcXvxoXHR+tTEkvt0RLcdHid3KqA4cA8RCBacvm
R0TAuTAr0caW/DGedgakVdYm1IEdyqeeGHcpDvc9nAHT4ZEDVJOPqTSc+ITeSaVdIAOrRd/gVOMv
NtFNW8E1iiNQUlQfuwC42pvXUXX31IkwEtd1xLnUGUUuPaoyv0jOSOzAWAnWNglq4qE/0PS507hz
3pf3xdlPXXY9sO+cjfVmDdFfkgdHKsL+q0wE38JMw4bDQEH6uqzRZJVcM39KGfZZVGedEFmI4WQ5
ClMOccmVUeXk+NjPGyCm4z3tCoaySRdSwHTWokGN3VZAc26EKu2oS4kHoYrk35DMw+e9P8jzketF
5qITRV+lhLq4ezTGmjAbh7Hvvo7F8ALMPB0TtD0/E9094f+RQhutitO14E45OHHkDn30bMde4DsP
N1qzNmRNC5qozCYjnJPlxpj3MO0yJ3/7t2mILqbTQN1Ah9YyaVEq2Z0wc1SVT6yEzdKXps/g41iK
sO00FDmvDUb03SXyfuCVuvV40V9S0LvX8hGdmpBZfjVJaYmLk2ruLvFc/9OpTYnrpuC/zK82KjxW
S6wkcvNr7khU6cTDfDUtOewEC5gW4OSInQoQsTsVzbUGEnpAVQ+0DiUeSeKyZe9jhQ070oSKNjym
MIxpW6QV2KIgmDe97HZ94kzy3pdi6m1q3AWsl5MnO+JEKQb3kBW0XtMo32Rf29KGlpX2/mj/DunJ
STGsG4JUYKG1H1Qhgy1OD3lNxglCI5IchXWggZkw76flOXAin86Ax71gcphKm/tG4YvXL5+LspAZ
gmKxz5w8fixNbPDoLBvkryETlZLSpmAuHsfulvcW3JCQjBaY+YaRaUl0T1byOvYnz4WfEHFiP0P+
QyAfdvM0uHUjxtwUDq9pM3Z1ILQ4K+8CnyF/GpODu/20+QOW+xDBebdYRlXU/EPNM0Xlilvl4U9T
4LmL3RSHML9MsYsWa70x37mSEMGDee1qrwSvZyLHpsAE4BlTLBQtOOYCeJxZoYPGIfoljoFS1fW+
lxzFtq1oO11LHtgx/HK9I+biHq1a1cqQkMAgSlVGMsYPbntS8N8QAR1+PxVrJCuOav4KKM1lNqC2
Bp0cVzZERk500+XA8RB4x+4KdJRbI/So4AiW+GxYvbbFfbtO4KYPxrPRZRuudbkyuVqkagN3aaGT
pmtQg5LFZPaEforWSqM5KzCWX42cANvRVpjfA98FPT4yByxsc/FNn0XGsF2/98+0Pp2TOhiHgLSD
Lt4SdHYrkZubt9VgIOfZZ5y1F79TcXyUCHzk3i5oxtT6ij5Yyxo251mvAJAvLfghWjsUXBFaFp5u
dCpUY2EP9kwYDn0NfdHi7G4RzL4zND3o2OCKs3fFYZJEK3zbAWwbASc+cz+y5MDzfasS6Wwm44GJ
rgJfUGoyN3wqgKX/jlaPBxA9NQQoxrCBFe4WCvJnkpYi/SL8opz4H5lOS5oAM9sQTDBAwlfJ0tY/
pt+uc0gum8rhAHseBDvJmeFK/CcbX/BJ7/iMGomahiRMGM3v8pVopFGGbAGVFPsA3BgZlvvDGClo
zuPvhsjqKMSioHj3Lhv6+EI4wt3kaMFButrD0wyX+mnzATmzfI1iw3q0aLSDHGdbHx51mBjOyuPE
OSFxsDDpTuqd4LeXe7/+9HUE0izjk2B2yHRtBTw7Oat+X/pXu23TZF79aheMPlF1vmGaQPxOTkIB
9YPd7+0bUb1nqkpepKt2pfWAADcOdk6bqPrNQ8AJyazXjQX87sidgPCSdq4O4yYjiXFBP1l2TumT
yTr4ggYpCLjN2vawMB5OmkslcjuCnsrXqTu4m+0pNco4ODiUfq3UKCB6Tqs6cshiM9zbwBxcjj5v
65bVFNOnun80yo92jHF1VwuXrcB2FbvSGRX+eeDAC9sE8RGVDdwRK7A6CQfnBbyFpMJutpy6vrTD
SMm7xY49YufqudQjLoFZD7mnMkUCiP7+mee2JP6/kfsGn3ch8VlKCrG6ZK+sDZLovhhxftSd12lG
9JL1jLw0uKIuFdhdIvmNupTPLUr5GDYHZPuZcVrBySh9qM/EVS7mcNrRWKe5WcR7Kp36D1Jtnh6P
ygSO9zsPx5WQ4OvkPckGF/vFRG1wKuSh8BqqRoVddpUA/Zjpd+Bmow9BCBaJYDfMSezcXtT7JysR
onX7NAFIJ9J8XlEiNYHd+ZLW0DApoJLuhQkV4CuPilJCo9gDuQyvr+cKrJRmad3yv2+VnmJYuEIy
FG29gDzd4UhfP0gLqyXYhxG+GzxIuoShFLtIrO5uCGKTPOQYCbRJLTxI/zkfHUudod/EoqriUy5T
BGwHfuTAfhV2HI61Lqo66TNPQyHLQAoOL8qT1wGrwXwwYhZhRcvy4Ptc2Qqy9WWdhzkvFR4ckUCP
3zbVCDAkC3vD8FDnxHp9sA61fNkeeH90IrkMsB9UrqFc05jrj3db05wtuted036y4Aa73HByispU
F/4puAWobQcjaoZVRUfjqEvuOrE47M7tf5D2BRD+9YcRSU6dFXtcMw9jXSyOvF+HX7+3o9wPbqTD
oDsXPcGH2T39SFaccH1AuGJZJrYz9GDueyj+gDpV1/b+gJhMm0kexYC8xvzD8qifmyded5/Evhin
CnjZKDvQ57UDPjFsNWQrcZGLcL9cLGjXC4b8DcLFzYJM1l5yf1gfhGtfChTZCMJhWxa7U7B/wf43
UIMt8OjttKuYZ5+Iw+sMdp9h3yGihBIhbzCOIfrswk7O7ZONg6Rpexgk2YUr9Jenq+TkSwGWqOZ2
SLR3v4Xwd4nHgk9+uniSeL42kdOO40K5hdRXG/mfi+IxSv16V2aWNeTPqw/M3hj3d5IkiEoG8Vy3
CSrPYujlA/Qhatlb2RINoePyXQDoCLUzH/lSC54OgCuGro5PHLuJfdynd7sLNgYiJqtYrVVu/t59
GDNKzSP5l6EcKoBILe88/Kua2f3mIiCHHs7cKZ/tjihMOBsrI7NrgpWdVR50f8O/PxvT3ii/Elq1
UUT2udl2Bw1qWEWFuGatX13gbsgRb87m6RlhhMNAxjlBHbtXrSZyeM6Gi41YN4cVsCmGh3nME49x
kbofObqbPIfhSLdJiOJBh/CvO0DyYMuch8Vr+6qML/Ki0/zx1TRW5Y3Ss6K8HvPpcvDKXxw8H3nz
8OadN3sF/J+7R6EYDw2G1FwCUIxWtVnIJeJrXr72ZWpLw2RFWJIpTQn1wL7dCXq3caDybUtrfuXO
6cR+1kGLo0ni2S5CWorDZc2kmPC2j7xcrMfAOBZhY5W9rQrg+PmDc/pejH8eXIUc9pXGSJIxvtMw
cW/TjEBGRMn3++mmacVW2uquiUcl3WER0QvLDfyVgS2DbGwq7G2AHiAj5/jNA5Oa/gL6gEGlnzPT
ts05/+7OV8e7XGRu8ADWfxZ3yPBv5Sh9Ttb1GXB6xhSExT8ODX9aGUc1ueNNVKcZ0boebobFzstM
wRnox2OL8tQzuSx34nch1psHFCyFWY0XlsYUrt9UAqkQVkiD+gnsr0RaHiJeKpq4HxWk/wVhmg8S
Dh6KS/LUGREm4HbcNXzYSlz7AjsxQ51ElnQlShgMkreM4J4EeJR0Nc+U8OI5PcFasp7JhGGb9yKl
hKDLEFq9YJWhPSHhrowsCkG4VTWHTDI5/kWR9IMqT3uup4WH99bWOSC9xPSm/22BwtMos6FOqwub
BbvjXqcYIGnf16kxveZCRxdogF1i9zVQ29+W6nU0wKX6+ajt6n+vx8EIAjZQ5g3Pm1dtgnjKhRad
VcTGIc1ZXnqqNj/ZnTG3aI+IW8y/acciet4qqhLcCtwA3zKzQDNzrI19f7UfwZD3bzwyR/TkgySb
WlKBgqsq6+GoXy6A/MG07H9C2mL0LPO+GOCeIvPKLHJo/Y/4DXUC+aLCEmRJBUw47Xv0Aj4ZlPhm
NOvceZKIgRrOghXvR46D4tWMZSLBzo6KgLDGG3sWraDr1lg3GQQ5v//Iya4OOvprDQz0e0/0PxXw
CxbCa6EqIcDNUxtLy6stAF3nNc+/3tXgIbMuIG/+v/uVGc5cyUfHLtVhLwOvgq7nkoj8jsQD7iGi
tsTabhPiSlBH0BbBo8gGYEJImd/RClI09swQ9+jV9YWs0xMhU9WKRHJVprNjbgT5/FfIFWbEPUA+
aveMhbnPW23VPMsdSlpOQjTUOu0zLxhjmWItCXXIEe1obp3TylqoS9ozjKe/TD3h+6vtm7PAkc3I
slUf7A/JUJah36RNsgPKIlV9lNo9rJ4JAn6D5HiBslLxGPeOqtNEEwr8XELr/cxtdiOUjXYNpbsX
1XTjbJKa5tt/MGLSK2msaL11P1qt2tHuNk1mBmm7zNQSQZoTeqoSllTYBhEnkf027IAuSlDEwCcY
8wKE8j/P7rzvtXwPxpM/mFtM5Hk8kttOeaK6jr7bne7qe0xoWTN+ro2aNuFs2UrRpByZ+9hNiQQp
P9oXzpCuWUaJOJ10pTmxG7K6y9aAgaigJWAYSR/BA2OmlEd0VqvjGwSZDVdcad3SpbI9Kkjiv4DP
F4lJw47WiptvcAusUPxb8FdZp6n0no0vYTYH7YX5gOjJlWxj3Vo/pz7/mC6VaOvrXVyqAVjs83ep
unAtGtM/LOTbW6RU0OLJggbdpCG642wOZfrkL1ciOEkWOIAVNHjAh0eHSJwDHnwvAK6vmj0OO47Z
aois5go/3hF5f2KaQByh6+D0hKpS5Hp73x2/D3iVYYc2TruSQs9/2i4zCbhrEit5n2FUbcDAY78z
sS76725btXdzirwnCWtMKyxze59+ixVN8xyXs+Sx/o+CmLq/rb4Z/cFnwmzJB/pAFyUEGuw4tQz7
aeSRIDjghmI72+zOhFHozsCW3cXKhm88tVlU++xzZR7gaLYLXxN7rsvI82FJnyGJDfWRwNE6MpDQ
UuHJO9kbiLMwdunY59aaTcINfoC3DHYkSAgB+ydeMIP8nefDubXHoPXJC6wbQ3qccEruoAwXZXP6
Wg4HRLOp3lXOrn7C+754bfiKPFo8Sb2qBoo9pBZghSVkDYfzum+GMBlnflW0dZMcuw2Geaiep9p/
UAPd85cUYwG1HV9Q5hBWjed7jidvFhAD0F6P6A1//4IPkAN2YUKHFzfnTT7JmEFZl7amYDLqd2+u
K/9+AdmHJ+GCFpBidgd7X8f2ttQdeB0imAGAOuGp98OsIA0aB+nsCxJ7Fm1CVPjNovI1dOgUDqbm
exaD2TKMX9BiCbpxkM6U7Yu6elZatEolJV7yJQdwWl6eORNgpgZ2h/xroyYdvlCjq4mPmYYU8k37
xCulDf2ye1hT4jR5joa2ovMZ3nEIa45Dcxc+zutBIVKeiDJv3O7X15oGJsrS7f3NM2K+2iamknRt
7OjP94roWfRyDO/HdXsUQWXLY24qWYR9c0L34WH51J4+EOp/0chZzjZR8XZzMRux4HUHeecvB+bP
lOVzl/PID9mLeApmIAqBqhS+LpotPEJPXFMobvwcNDYxB4BxFYRidFq1NtZHqEnJyjTiXYpFYZUO
dDwutvCyWb2EHjDiLI6UCFUrLnfGuDa36DgRW/w8MpB0KvxXbuwtVcYQD968WAVIOUMTVy9wmreW
OxwoVApU5tO+SU9GzyFzG/eFIbcg4SHyWQ/JzhxER6vg7cDNeHEg/jLQSHgi/jx0LgaRuozkD143
Fwda5yuLFqU9aWWMg3n9VctvcRlt3T64zwKWV332sVFMqlbT723yd8ndH1avSfgYzKcV7DoyOhsu
r0aG8CIXGOs7GcUNKe3HjKl6XPtsFatONP7xNuJkO/E1NKjvs63jZFBtv5N69AqW0i+HblUQYEhV
pnupWmn8YUDPo/OBDW0qN/YyVulR7y8AuQjhQTDJSvYGMHnO85segUG5Y+nXSPxttxlUw++byOIy
VJnx8rvKPUR1iouEw0jCTs7rq1XJ7hOR9r6SZp4UcTHM6IwmQCkSC4utcQXgVh2J7/kl7VRipCRG
UYTGeQsWGz14GMwPCkpi9W92fNysVXBDAlCkKUrLsoV+Z+wbHdWpHqVWtjlueMAfYIq9kwkK6Jo3
H1eLKIwDpllRLCEungxNhHJUVZvMSD4xCBX7jlCgXoSdFUTapPv+Dihjths37PPIyMWxdLZMpS/v
fjLsl33w+R09CQJulgqJfheqvCEkka5zewUZ7VszRf06HumIYHIUfnub4SEvbcdzwDT9topzwscD
WneOJd7f3Fg/0CMB4xlpp26iuH5qm8AEFszrG5EG+uVifDuE28/jRgWvHJDGDCzNySqTtoNYseS1
wJSfCEzU/W+Zna7JDOKYvim81s4pA6jtflR6KKMlQDuly1WcQcYQuNmJpbAB0TQdnIUPWyclzR8k
LNBWvXRp84gU1CxxGFE1FJQdT85Bm2DGqy7impxX3ZwMFEJN+wHX1rc6uotTAvZ6TJakvPt3hgSu
z5NULdYSSYN6TYVxTUUjd4yNsi7WryVaSYZbPAuq9H73F9HVLUxasWxHo6gHslzYntZWX5R0om5I
dGPZsl9HXaz2SRz1VGpL5FVMWttlwoTfFEE9NMJjJJJ252Jw3fKxDV1kZnhN1YpG5WQ+M6RWXADz
UibQNsYJCbKTq/wYdLsV9olSxwfSVwJg4XinX8RIY56OlQte9RH3t6uguXSRSSpIQlJWEstKMuh9
9/icfKR/C0J5S8t6KkE/ddFuNuD/BPl6xcw2FM2LWre0R4iWoMn/z8vVHAnxp9Zhj4BSj1ulen0B
qymxqXMo02zpTvRHJqrZYU3YzPJtzEO6FsW0sPorDFxySRZNyRX8MFLbooPlWaGkX7mfJeeox9up
lG1Et00D/btWmLicYCsNIDj2EonEi4QzEUq1yl/QiK16LzlA9XPnvcya9dsPQ0PZWXhTuBH0eS1q
VmQwazyxLh+AzwYAMUUnghNulnNmSYoDWaqPorAfopSDTimEDiHTxE8QUCnJ+4b3poPROWWC4Kgi
6ZtHvpI0xU2B4NS21TFWU2QqLNk2Oy6Lp4xPvTbE9TGDXtQ51zZhzNBMhfyBG6SWGpT5xpQE2v9f
MPGgSvQ86O4g8B/bySTaTdz7l43tFy4cDgnHLla8FVw6EqyflSW4n3fzgI7L6zgicNpdKlPLjWXa
6hDjZ7tJ5EHAjwA+VIMa9/mQVpRPj8J4pbQMRtCbDPOooEq3F5uMXBGsfC+hzQoI82QZs0J8k2MC
2xG1gIafkogYkl+gvf1RCo8+tNKajdvq983Toa3Cl6CWeXr+L/Gi5yke+6A/5Nzq1klPCTFoUoEX
79GigjnFcFRwfNriqty0ScIqZbGle5zIggvXyUj1ME2x+inkWVFQB2Imdq05+PgXAIwI9VpJb+MW
z+ess3RQF++EVBIZksg1vQlo1Hdu5hOTTNeDy2ePbAf1BE3mP85PG5dftoOEp5IjeoE7wJeOj6ry
Aoum8QcPzlsqX+qhKeWih1U8UTUCJ7SAn8kUA1Z+zG+ZpzNJHVz+F2Dr+Qei+2l6bskufVYJ204a
men4fbxIaGiNp1L7lkM/CCPn02iZIoPkRQIim7AdBEkaZbTow7iPvLVQ3fgMbnSz9qsX/IQIPGGI
uIZV1vE4vZAmhWT6FilipTN7T6sBCu41uDKz3KHUI/QE+C9axUX5+SxxIhEG12TLViIc3LSF01Nx
Ox1JIuLRDTjvY5LLCL69AKnsVbPK9SsiPNB6VeiAgXxh7nOe8SYwC6w3Vxt7NZdRo7oG6SR4ThNx
roqCDG5A4k6hksSlFuaaJQbk1f0n4IDKU8tsrQakZdUGlx1Twi16FynmSUZN7tbgrLRkIEsIWNyY
xQfpfZha6btWEpj9ZGU2U44JE3blDgljtnD2Me+iVEpbMeeAo78ZD7icWuzF9FIOt83SMwr0WoEq
GsOOMfV5Rl4GV0bXu99QOshBdSQ7cAgmoEy0abMfznPH1ltQt/i+NQw9KbruSfxo1INKKMPkb09Q
6LmJA8b//pGNJ/8seJEnksR42GOPPUWk861x2/9ibizg12Jp16P3rVYk/hjk+P4OssdQVXFBlpkx
stNx736aOU3+it6HT3T094Y65DidNs7ggHuGY1MlNpBYhMivLsP7xvI9oGk5WmnQmeAYKyhGD46n
+j8jYRN8FPI8B/Mmr5W3on7kp+KKWy+J/ibUYi1F827861XCDDQOcBACJnmmUWN1RaiwaN851CsW
p5PAya9vDa7PDZ/KzTGBGq5gXPPC7GJG8sqy7sy6A/WLfseJ3XKB6TuE+YeYqq+WtF8IOrVqWYXH
TkhzdOMGmb4UOi5stCRu+eJm92bf+V4+LUbxpVxa/3OnMsbJwK6X4kUOdVxGoGC1xt0avpu2vgSo
0RTbIYFZlErQn6Qn4kBZqEE5IXvWDJUk115jtJ6emH0ITUdOwFokpM2xSBO2bBt5HjmUekAJStDW
2bb8xXUzxiMIAtievERdo+iNmR3WS0evg8X4tA+RE4iNWA4ANpPqe3/rjtia8C6MmqrOXL38h8Dd
DDUNF0z4Y6aqomrCXH3xP2TtDUf+DjUmpKYd80h8YraQf82lGMNJcBxPvrPrDCZm7NoINiiHZ34Q
IihaTE5pk8V9Z4KcfJMIZeGEW+sCsop5M0Ezhirlu9CRLQBXaAlXPjPbfh+ONqDICUr/VxHO4CLh
GCqdHPqfxNyd+ZZMdiF+mNcSIuhH30c7xKC3EhHDBkFj09gaWHxnUDZlBtSI1EyhkfLBTqYBilcz
6a8JgubVDtph2i/VQTB2PIx6NJsiLcfMz30qS5s0oppP9cSc/X6vw3xtf/WKZhG9TQYOaCM9TVA1
tTPeCN3KwD5QOH0mlD33bBz42I3/G8Hmu/kCsuqHfVkr5MiHIdWn9nr4FAUEaN2JR8b5NzkaP0mo
uitiuOXdXRhboW4X77p7lJRPwAWRbtWkszFYhtpvWdqsGSqck39dwvbecEwOQ1Wm/ukHhvjJojCS
7ruqx1ST5FkFJ4zDXYvBpoSAXDQiecmn77CHN+tuBjuAkKtiy6sulDYwbbx9E3FdrFAA/AXLnuhU
u5aPtSC/jfZG52Oy1SnWTcPDHh7auJGj+T/wDNG3AFe68HcPJh8QanMJev8PHdCEapyvzcuSHkZa
eBn1BLDkyx/vsPXxUzB1RosQG/Whqeehj42TaTqCCWUSe47ilLZkb14UXDimvUkQ6Dbj8mWu4rj0
P/sU5w1syq+WEHZRoSSJnh9wYcMlazGuuoc7NfckPBhSPNpNIRT8O0wkbgSREN3vHEWGqVSl9fHF
m0B7kY/JValaXCZ5f0isbncviC7BybV6kq/AZx9Tu1u3RElTWzJ4i9MpOpTGtoRwH2TiXmazubFw
JOaJ/StC3903nX8TdS473jpw63z/VlqL+gllOBZiJbvk9LT4qjoWKN1rIAsCvO4fvuecWkdfDCnA
WZr0zfTaoOPaKFhQvqm17ZVROLGzoodLxUri9LMkScbtJpyXq/c3dotB6p1YjShuvtPBgKVeJ9Uu
9MQ7rcgi8Nlgb7hunjPTIfmjTmd4XSDI4aQIwxp44d/jLT3d0ubgdhTf3lz6W+9FGMv6dDCykuyJ
LxhHBjqpDRCTfEU6cdpVAHQRCQQiDDC7fOoS/DxN7YOgVAYamFw1pFwYY/vi2/4hk47QuLTl2Gu1
fgCkifbnOqNh1VPG5XOveJy0Eo3g0FbGrfnBue7HpTlPd4pUje7GG6gjh2WECbxKUxBZd/KGTsiy
V9RH9FP7IxWA2Aj4sBsrxKb4GV3bBGX8zCD3R91An2Z+oC9/7kO2UiNqQgZksYWntuTaJtj7XKrD
TK6Vuhdxa68W5VD4ZNrVraxhYFxVvGTT4zqQQ9PfMO3EEtBR+qUZ5g7XOSDYyoEfqdw888trh6AJ
LvTxcUgnYrSDOadk3Ti522b/ePcUWNG7puRffl3m+yq+FPchqUrOv08pXVE0hSvZ5qNV7L9krNjD
zzegynfB4P/Uih55o3EaTXg1snJxE1UQDKSY0whAN/vX0nm0ABSvvSvMJ7c6FKBPwz/oJxajaQAx
85am/kxzaw+lz+ATjmG5PR0CaPDfyr3AYDPxFBvtWGhvrkkBcFJ95pdL5WUzgjRlaPWwMkwSpt8J
bmLO6arVlH0N0VW+ks57JkL1JM2OGc6o8AH53iHsnYdUR0p2N82ZC6VSrPxy+IyunTiXSaMhboIm
yYe+rhM3gjBCv5Y2PnFV6FiXeDh1GywpP98YkZ+wL6NOOj01i2dq9KQvUXYOcnDs3hQChE+C/5cZ
f0b60bZmaTh58tTGPej3KdL3mD7YIkdhLZjOYoGd2IS8R049xIwC9a7HRdW9GtOXJZYwzDb1Il8R
k1Mkrqo/s3u2J0RhnIKffBR/khh2IUjc8a1uXDo3wRerXrzhr9jQmcefkCOkcwZrga8OPaHcOD+F
m/LboTJE+hqR+ECImIrdAwq25ES2JHVUYE9QPzMrCLqyl0Un3pxqSVps+tFNvGj78J5yVR3vGp8T
T8Dsae3JRwRT/v0IKcvO0vg8UKsmz/ftONYd08edYPcxSj4xAozBcafF9SCrNhtTKQBjlUdW6dRb
fEdAnOaM+Mn4qDVrSjCBkpJOuOGBKwgUcZXatPgfJmBlam4gsG3E3H8VC/mqNjfq7lsgt31PLMi7
eez1+b0WrYGlxVc+a6v5MZjI8zDeqtDTsQuZV0wfQAz2aldmbet2b+IJjdEQpOg4zVs2SWnq8vSJ
7T+PB1AG0GSvq8sHwQp7xo1TCOcbVs2LEoDNeBgcdPiaBUtc/WXiAjSW0JDwcbamnEoB2nj6SURV
zlys2MrSffa+xumFsFYNSRbTLjjT81QpDLl9keGzhoe4DVF49WmPqOvLZamiPybqr3mrgSYgfSSp
yQNW7pJWnp+xQtLJ4+bFfQZgWHlMpuuhypj4B2h5yEKz9s4w1Dl38SDHrkJZiNqUKYKuY1ZZMDj8
xJuZz4hP54da+mkJsws0m0t+5OlVyqK0euleNkp9pAVZlEZYcByJbSbt202rzmqAaEYOOP+DVrap
we8DpsxNSwXoS/59PDH0EpfiApuTafyoKqN0UQDSs6Hxq1gFxfO9Po8fYQ/FpCUpD/ob0gbBUZ/8
0wDEpZY9DeQWjpUnDdacbz4Uyd/okLWki1NB1o2L8LF0vgFBkQJj7TnDYnr4XBWeoDmmiS29HbMx
kGyqt9uUvv4iWVaM7TSBGx6qvD0SCRtP9v9XgER7iGWydin8Oq54NSoFdb6YINthLblNT4ZD16bm
PC0vgTuxo4wxgHW5AkukEMmphCufBvbo3GvK3gB49W3QimMjOQ1g5dSiUHI4kxt8q3naGAl5vpFQ
L1H7x6+F/7ugg+XOXzf+yecTO3yr+wjbDhnVwSBVg0tWuVaOyZdvzyoJ+KSA+55m1Juidxln4c65
OiBZQQXlx2vsYsASS1t33b7xTPTSACjdg9h7xbZNIWDYaUO1EYvhj+MNHw/OXT84cdD3tQfajnZe
ZCScHXB8LOzNL9JXiynWXsHI7J9TN6yefnvvJ1+XfMBTi/ZPd+0nLUVP4JsOFLRJDdCjuqaCjvx8
QbolP8MXT92wP7P/ZqPIDzK5nSh8EkWgObumrk3MivlWQya+zqurFgxk7zqe4FwQztJN/LtSth6k
9Kl73NvjbwV2WTroMyTo0sqWjC0KpDSQW5VtNEXtjck6XZc6pGQVNHlaoFUIANMmgySdnHTd/qZl
pxbbTlbCwD6hAYPTXVxHgZ6w8Aqxk+jFrwhd9vYydtqln7A7HZUPkqa4e5ZPUWOZJpVGuOZv9pwm
8fUhbW6dcQYnhxZjdLsOaC/tb5nhjIBNp7tfkWvTvZP1dga9Jt1b9hK0MDqsV9AWUOV+q9KWFldJ
YjpWx8raroNi1H1ifoaSi3p01Gn1n4SagGe2mBiscaW5h6fuXQ4TyEEnaLB0/mg9bPl/gLPubs0w
uYlszDI7iFHHEvbGXjo9Ch8lMuwRB/iRhhsvGyu1Q0OX4jjyrabMDFl4kVFzrq+MIzwhsKNEYaeY
5F3bZ8z9WDO6T2ZGj2EcBK6TSUc+ylASuv+7y0DjjRjSA1+3H5jA2ow28E5Kbwx1iEwV2J+/BODp
XJREGRxXUHwD7H1SsIhqUpQxQZBtUmFZHhlniskZZq12b7Ps7Y7Sx8ESJO2cLpXJ+p3HHi0foYlV
BPHpB4s5RkCAwNWmgmt8oL0hxDGBhWAKYZku8MWP2ymkZT5N+KuhUA9mYXr//J4texYpfoV0VysN
g+BAq1JlnDso7Wa8qf00OIKsx7nul0ocfDWSSzu4N1F+U+OSezDJ+IQcP6GQfTtYYJMQvrXcjqH/
RVURhvX2wMWpiKVWy6wzTz+mKTgbMVfKHmz+LHsSSlErJ+07KbeHu1ocyqY7OWu4eLuSmnbTy8dv
ygNTW/1OlcG/xRJ+BllzmxuOXpno21qoGNC17Ha04qAi7dOV42ekG8ykIudytzYyD78qMqXV8pkb
+g1Bkf2bOvB0xtNJIhk2n2SXbylCizGd5h97dZDYuuDB4DEz0vver+zfdoVZKAn5VSnL+uKXcXKa
yBY2XfLSgKm/AHSVuQ9c0jyJNPO/XvZrmloYp4PwB+66P7kZ9OgNgEq6PKFG9R+7gr1I/s+qKNZz
G+rw61cebuHYDt4rBpUt9hmD38hUh1wZGEBTH8UHUekDZ3ha+pRsOJtkBW2xpFOq0wzLWWzCLtr5
JQf34WUhjJHkoctjSsetkS0ElwSoddx6dlwtPhnCNmUbVP1kG5aF57c0kDxMeM2lNXRi2+x3POdG
rXZjabJIQeFHye4T+RE7Rjt8UI+QVYvm1j583oDxxzCigIglK8F8i2RmFOfUKLRIFUPquYXhYHVF
uG43+HBc7G1YLwUELoP0Q6OWTr4Aq0czGnKjZgJfvRawMqgEO7t3JC4S8FD7HyZKbo8N6wyoH2MJ
Qe0LHvvXjwL9aZBv5PlV3ZR236nDM3gYCaD+QluNkOJZeYmYZ47c3F/lJu3zsqHLMU03RDrlIRsP
z4S2yMwRtULNrWwuV/FOpn44SGKfLFAvmOP9kky8iaKtD4wiq6CBCGZCG2U8PKySCTiRy5XvDuDy
7qZXGkbCS4mxIEKL6ZIlxlqFr1g9RJ544qSd9E6S/QvktV9XNCNX0rFyMHJHcSCL29lCgcHlokFl
HZPgo78BHIv+igF25gWqTd+hTR7HWVbQBvp12bBy1NxJaVSP5QNSTEK+QNW0RgO/5gNrU1vmOL+A
s6cQRJrI/DC4IKMjbKrXkfKQAJiM2P6Fy6thVBw8/ALzRb7AhOBpLWQFNy54NVp3ETZQmV+tIm+K
KRhpyHPoHKe4AR2DkNW6mO2CCl7lnR116SPlJU0wqz2I2EpXtGBO1+S+v7Ct8U2H+OAJr9piJRPR
CB0QxU/P1JkTaZAyoHGKKKapYR9ARkthUu9fYTEUCaxvfI3bARgR3Vlo/2bD8J/hmzdLTGSx4ri2
Rxt9YOZg/v3xlX+4Bsq6HgRSluEx33wY1dJ3b+V5an+A0OPLoyvkvuKmcSLDnhvASWat53FgmAYU
/oM8gd3P+zjuVqOh2cDD9TtrOEdmDzPLzKEacx+oGbfBOpcxNUhF2VpuPbuDdxoxjNFm2hAuqupf
YHv758Q0HSmalEXfkS5dj+d3hS500spk6lvMR7MiSSiXLDTEu8PI+ifLPpcTWKeZjO39Cxxs38AM
Wdt52R0F2jWfl3SXNnnN/hGxZObxaYRmEa7AJA+ivPE+0g72TuDp4E5Mp7k9tBWRMHYJ/5lnFiZr
HMRcZu4lVeB3hYILkSONEuGZ2HXqBz7yrKl4ryUiMPgzt3ZxNUQEwpefH1mDXBOJ+GqSVu1SUtQo
T80SCaYmIfhBF8J7KydlS3D4h7EGrgTP2aq1VxdiBrRTT6aRwuTNw2E+c+CZd2nkBXtJFN9eKov5
vlYq5UEW+57ODHZLz+SMb+siQomJvCmTktYjfI0/E8iOt9ltqKqZw4a/ZG84xZO33jGtv3SBgecT
0OQJyXCIGcmQVShoPjVfxLHtAqxDiWEDVPn4NTD6IFlCP6zwY97C1y5npIjybEWx2C2tVuRSogow
Qk7pHoi/6pAszU2UeeDkkqSzsFcHYi8rLq4zVtanl+7+79pY5c42qh8FhjvKGq1e2rD2mNOb1Q6u
MHAkU6pVwk3UyUPlK2Nt+0NcSMDrud5S31IMf0+eNhV+JhB6bL2ft1lFjYBLE3muFe8zRaSVTR19
BO3dfzPaSDgpQg3234WtxvHTPVGw0+aiRg2ezAEunP7mdooLM87CT0BVV7Dq9dnFByGrtD80GIQQ
NPCR7OXneiFFZAax+L7r1fe2deidHvki9qzId3ATsJ9DSyO41wyJwTeMvoHBy/vSRwgBdBZW4lRg
HNS8zKXCUtziUsQoavDbIMLVZqLsrwYszh/3SzLUao6Jax5eMniDZp105O7+LBj99B+hiew8GjxR
fyOyMXuEbhtS9ggcY7qcJ6rF/dgvXKRGGPgoSHJDd6Na9rbI4M8v3O4FuQS2xyvKMH/0dGf94TGF
m9xKHrhpxfLBgkLjncqkTZ4DM1ru7LIm74MwjgEO7g+6TT5db/1SLfeHx2zV9JzxUgWePKEQl0ny
TagbqGn0lzkPW64bcPwyuV7o6Z5AegQ0fKnBr1ioKwyP0Cirswk/TkP6a88aWTGFL65zWZFa/Wzb
wtPIDVe4MYUGYkUi8HwgCj0YaxlBK1r2Ii9SV3dChFEI0U/0RplG0EZQzx/vvn5Ddd2nZWj68LbD
aeJ2QtGcoguedPbVk6phYA6340GLiePcAjMHwjguf8643GNUBfUViwNwIEOVDcALbLSIMunt/Qlt
4t+41z1dfrwZip7V/46RKMfJfjpxZjyBLf2LwE8MuB/LLxQ18l3qDtr8njYsPIJPD7Kv3JEC0qYG
gSZYgujcihmhdBLOQVA9iYMPryyxjjr/4xf6pAbdcqV55+Jg5z2qCUcOM0IjVRBiVqX9qnumFZny
nhIytYhvZYlQlNhXcvg160MwEkBc+SU7yG6wIyon462+Ee3mC5NImG07fbQD74PGVJ1Yd3zGdB4G
L0WEupfvAQ2S7SGgYTkHt5t2iaBbNOTWkGT3fQf0vrl7JsVn+nAF/NlKx3Ej20+3RWEF5v4RjiJq
z4QlySt0VPtSRRpYIhxqQSd5wtG7nMXSRhSZ1hQtSSMCLhXPqf9q4HfUZ4tOswp9EUuCzA==
`protect end_protected
