-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
oqXNBTnwS7aNTGYV9V68BvKxMPCqgGf1J801jG51tL0l16Q3SyLOIwO8GpsGubbM
YGZfk4eV0ySRY3n9oIceUQYrxtwZpRNWP+LwpKahSIpvrBSQasvB8gtS/9GGlMPa
QFRXCB51GAU8FcU92ZDMHQAE32bu5VK1hf5dClk6yz4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 19698)

`protect DATA_BLOCK
jWYXJgwLeQlvY5hA35J5HdFd6Ljutc3ljzUo1TMQV1aeymVOt71uWc/LjpAG0hJ8
OTrDoVX/eOK4+TRmxACSmVedanSv34Yk500sQGBcW20f4RUxF5pyXUyKJBIOpG/w
F6hVUpiSRrik3NWLqL4r/iUw56LcTxQfVLPS9HCwLWwY9Ud3BG1EkIcTTgncZHwW
/Xr9Nx7Sjzb7sJVNeyjuQeR+hAxQaEJYLwps8nffVYZthOivtq1fjKk5B9NmGgHd
l/i7j6HY8ybH8iUCJa5tV3Vx7oFfWCAMTeGbs1ABnyYuLCtdmDrfdXmvyGg1vuAo
dj4YMh+YhqGkC9G8EwSFRJZWqwPMWu91lqbHXRhV3jmB04qzyl0b6eqJ6CC7PKcV
8WW1OGDERrQxRrxu11EwkZpZnYh+DV3zXtJ84EuxX4Dk6pvw9J56ErANXg4Cv5m4
2Rll/oXyv1EEdfhaxLNV0wXW1PZlXXbOtvi50TaBuahP3PpCcRWyxJAnVbcF5Afi
IRnpJHlFRRqhcnclBjBNpFCPloXQlNv8Gf/odu02RGNTnzJyx4qWjaLY89aRkDDu
zGnk/+XfsjtTtBff3oCQsmQV2JgrxgM3nyQMnajBbeEZverZ5i6aAiEIMFQ4ASQ2
UrXWQ90E3PVfnm1M49gOKtv1E8XFrYE7x7rQvs5jUy4e1c2+kBI7DXcOcIfWEGgR
wvtO/1UvOE6bTZMyWotLQDxxB8NN72LfIvvot8sMOpmw243TRB2qOhAHzp5lW/qW
O0gorNrQyKm7YQ2j56pHloCh380OC0OaDwmfOJDxen+LuML1U0cjNsBDnvjlOmSn
xUJ2ShH85+puZEsBX6kLz0Jb44sN9OYWsrEuCUqH/d8bnjn4gDWM0vl5rTOOxMxF
HddhBIY9OSIdkr+nP0gTVLazJ1D2CDvo3wNRhItt4p5jInxjLDQ6xmMNY2Y9A52x
zPqHSj7Z0KZdRpzk4wp0TOfg0/0NQc4V1TuhzrUOtTr59dxDv427qd1MlG9d5KUv
z6goMPgluyh890Piq4IbVCuG4r4iu+mpgGzq7Edoj+KwAGEtNUe88M22nwcTys/P
oX9XDfyaokj8AkprW33xPtHAnuTdGTd4hK28o+mcLjQgaA3C96nA7T4WyxzQfy8p
I2ChESnLJ7lkEHxsvREEm2AgSI4SoZ/rUQoM2CV1qU1JNnHfA74dC6YEQ5B46fH9
JM6R23V3nfrrs3avi5VdGAQw2BnSrdg0fi+7yq0eqeNN9DuueZcJGzOvhh/iLLf/
hxqwxBweJldJineB1oIa9pgTZARbcdTFeEfTudAndgVUAsAOdjOyp0/E/bQt4w0z
0DonqnOiS6LkwNWmR3EMIDYJ5XG9e30DVqwpaQW4jJpwYRvMdd1yz6n/MrH88000
9y1VKe9RB0b5vihNp0dGuTCm15TvifNLnqqHYAxiKPlc/bhN3fhWFMlpvg+yoh36
rrV7gnsow1DW5Aie6ynLrnbvKa0/KTWZbN/gXFKxIzFjxl6ExdxWvN6B2O15TryX
knduOZw0tPtchUUHid5R6z/iOa06u4838nvIjESpBRBpBIfNls14opLmcn681Px6
DX4FdmHiZRWegZDRZo+A82eU88eVoV1K7/kTVibHMoBquL31XhZC0sTtBjLC6zvr
RPgCtcMSCeUlGsmMsT2xReIGTL89TAxEpjvZ2s4G0+6DqSvexWolGKAgFtVeXLh0
b6WCA2RqyuWppSakW6uqK8OvVwWg6/4dty7hCG9C55VJp8TyyU15YdjODy7n3qlU
moGpcx0IUCsjJSDq2WsK5WDVRLuNqKkG/9wNCn6Pyj7AROi/vdMgJtQQyVWlp6wO
NLiHwSaT9XdZf4h0u2EGE2KzMXtVBzVnkcH6Vv5tIetT+voWdfDRvekeWSblTiyt
i3sDALsYBhWBAW3z5Afwuk96VwA7YMk/W9wGDOo2yQXQRJzDsPNwMmEm9vcKxpJU
y9dGgkh+84mcTRXn4qQDL42ohKOT4tD0Scsr48436jAVfwV8dQws9Od+BnGuOY0k
D7LoxcBtmYKqyPzigc/eXFwRCXWGPjf90pdCCIKA6MSRGUBRbEtQ7m+so5I0kQsi
7lcWOaDRW8k8bhurT/80jKRJn2u6nW5JOp52uomGHV6alT+rf+OtjsaAWChnRPTZ
ob7vPF05o7O6B9VCViYaRCI1j17Q5ucp9cUein2yerKstE4PzvO9tPnvsqmG4Ku5
KypA2WmCd93OOBfZEE4gZa4uLUIAPfTfHdIbE/PdpbNJ+sUEJGlHNqA8Oq8ZyAdo
BbsMWMcKyZ6a19PwHxS1kw/3PZVue/sd8r5c/QIs1d5md+8//W/gjUOo7ymVIFYR
LGfhcwaqhFzbNvwvqImyFbQxfMmsKy3dhdHWKZ8fwhyvWYz0sXeOCQGN57EsV95J
5VeXgSSR82M/7El12R0Js7DnAmPG5man05boZSsgauvYNp++rl/hNpahYbKKRTq2
rI85VFhno9538TEEiGFTvmbQqMkSk6ZoZmvZ+GjJIC3T8RzHTKxGUhe5zgzwf40g
BtB1irLPKuibT9Ciof2ftQLiODB+zq7Co0yIFrgBkPDOYZvTsxsdMsMJDyB+Yr4S
Z/Tx7xr+V1GpPTQmNfhBXN0Z37HUoPHOc3E7vb/66Io+JYWd69i2lbm0+R4su/3D
FFB1O+SH+uBM6EEzcejfz7agw6bfaCQu8MhivxhEI95qgcIO6yrbx3wT8aCuI8Yy
IJp0TpNOWwjjHZamH9dXJdiknrrrvgNohBC8tg+uDDAsW3wYlvZq3dEj+lfW7tHm
gfJfwzbu5E3CjWzkfddmr67W0hMJP3O6bVUt58k1HapBZbqbTZ/UAzWAiooYGFko
jb3rXcfLDL9VjE7BKbV6em6KSLhcWeU52k/L5eOsg57DdHOlkbRdCXYEvwUGdLNS
q6ZjwJtBiIZnG2eUOfrXa2WBbZriD1O3msv+6g9ZGbbQAf5V3FgJ63rD/ckzcyvh
46eROC9uKrunokUx+VbpK3YWH0XN9t39PhV1JjDk0GcEOcT3XyIkuViDi1IUNbDF
FVZxG0HD3dmgMiRECelriKvgL7+ZAgBcFyY1s1Qhc2IGmLcjpYWK1Am9H+Pt0Pkq
Lq/HK5DqxuXOS6AxgIa4wLbReDP5qjf8wtRB/3BOZ2K7jJ6rydLd+3ltf4PsdckJ
aALHT076DTldypRgrkx1bSyrTds1bMikT8bHA44kaFZBmZ1WNVNyLwCdfbFYdiUa
CEmzOgory9/98QCpHhppsoERqNlFMCOOWzf2PxzFOpJb8bAShDjgAZ0xyrFuWcc+
lhLY8r7OJzj5Za4YXCIWTFE0eNzWWB0WG2gl+l0c8L85biW8/9TBvwygBa6ab1BD
DgWHKYcvU2Ve9yW/MrfIg+YqmjxSC0/NDVxVzjl8wUJSiZh3E2EMH9jz2iyS8lie
1ztdcPaPSPCy6v4Myh+9uY1g+AOH3nur10DgIGoK/E09xtl7ri/BSSHnttAR87w5
tL3TChDtzGakDybn2Z47sp3cgTP1ILDlOVbYV+RUkwg4T+lv221p6LxfufdLkuSx
cZnlWO846S0bbjaed/h4eP9+RbkCDbFgBSqnvio1P+UVRCCN3blxUAIyX5/H/fiD
tfd5hSt08EbrEllPh+L1tDB2zX0vOtew5D/NUcgr6Q+yW8uzq7MpO8em241ocrv9
lzT64TdRaCb1qnoynQTX9wDLlzHuowZpGYT3VUw/8v/K1HcYhHq/kDvWxE0mgKUG
Coer2b6ZhEbxwk+2r5cWE9MaM+wufkuqz0s0XzFisfVpzQPHjVMLRrdVYQgRF5T1
gBH8124V2j2hKlt+hO8AB9Xl2Agtr3QCzAHGdIw/ug2wEXyjcaPJH5fkMyEJlr4m
B6FINMfJ62Sfy2Ihec2dmBQyzewHczphhHykIBKyPqTMg30urNEhRmjwtcnTBpPh
vGAggxpPlHZ+oS2UBAo9VuSu+UWCORfpS6OvDRFnxHMBJUr+qnwDVFUFKYXtz8/B
Kj4TfYFfGnzuT5AGPMMjWuuqjgBvuzoS1BVOsua8UrPw+xcwSuGDV30fm1nuusZ1
GpWaq+kiN+ntqhwzKyOuNJTXurFnJpWRQSROwQ48YTuquA/hw3QzAE7dwpGClNxV
fm1P0hsYYdDIWqWzTJ5SljoPero0IyW+4gvWjHsVCO+v7gW5ARWvTiQJQL93r8YH
JK0LPyMDiuDTBPiwkea3QWUJTVav6SIca/DXPyMcKIqdTGuMNVXqY5Nt/BU0s3fX
anZTowP/j3GBzB2E14hq5GKkQoTUjzJjSItotm4kmMEpi7qgctBsQ3lf/3nc1OwZ
8qLPEZlwVO8ieUtrzBTSmvx0K0XfSrjRmLK0zGOCPRcjoOLU6UwmiFhm6pDda/H0
B1ojYv2RLRsoZ63Aa7evL/jtt0yEWW7GYK9FIMp1PloeISsiRZaonSg8bX6Ts0O2
1L/sQBOtjkLnN1G4MWdMI+EnYaFIol+FScYrB/uiRu6tWbpDjOAEyoRAPP3NBcAT
Y6bWqe5/hIfVftAVqdGQJsq9MnHOo5OWqSxVttGSw3+nNRrMdEPvYb/oSgWLuHV1
9z2pFVqalEek4lAuj7CddTxNBluVmRagOeAFYYYVDX0hHl4ldPFsIU2RoYGJJCes
IlOh/O6z+Jp4BstFlLXcf1e8x+O6r5FzORZ/MzKs8BeEgCWGIeu4/MeD3HtsrcmA
NN70MOQRolocumfiMedg5Jt8d2m9DgOzIfbTYw1tTjpRhEq7LAyg0YXU6wkG7AKz
zqF/o7ayiWWw3vsPW9idL2bnku/FnQWvbhLoQgKAi15eLMNyHzLI9epR8GLeGTJB
WSBgCUTkTuopngXb+qGKi7WNVy8GloscfZp9wny85Nh8QuvUFO2JrnJfDGOtQ88l
MaAdu0ZsvFmmgWoY9KL/RB1BUoKRVXs5POxpuuAhMQvume0pp69L/rlcOg9OD7Sm
u5338C3NhPXELVpZj7u25XY+F+SYlpXE2roVbZcx1Ht0G6DOVdNqjkPa4CNFkyxo
luO0O37FcNHEKdgcmx7SKsLve6/l/fujhP2DGbdXUd5NkP5Xw5Przh2rccndw4c8
PtbTkzBbLkmEqWPITh72ujA6mcW0H00cfFL+DGNvUMt3kZmVfUDZkHxJPeI2mXKz
tvnI87sVjSGRcNqBKo2ih3xmZBr88LBl1yU3s3D7qnPdTndtveK75IQvFvjCaOzY
ypIS62BKFA697hddzZ+SzxeAtXtkAvBoYv6Z+ikJNfHLfyJ6GhRB9PNNssm38+b7
PXdoGmEvQSvxWTiado1NmMqJxlucFs1ewD0IoTMRbd860SeapPfFm/nWW/aERzTE
kv7tXliupmx1VXP3BEt4fPrkyQINtB78c4aHBs9ZeZMeI0Ld3hSewHSo4+uEe3ob
5hT+6gCjiITCBM45oousRzzpGvqka5XZAHDBgPq0cvcOvX4n8nuGwqqWt8NNDo74
GEGrJ9yJu93l/9Mh88GtGlLBS6Kjb9qqPoVjvBFxHujDDBvskQb/BjtDuotwqB3A
0nLiQCpQPCEaBPh2Msd1rymjaA34A54cg5vQz8gsUWUXzdrTJtI9zwiCy6QHg2Ek
slKxZunF+ii2J/jdJeUtuvdCwJKAt/ya+Mk8ZfhlvRUWb8W3Rekn+6pxXEwIhfxB
mJoxYvoUxQEQEM3g2G/grhg/EXi52w3RGESsZQI3JGy7olF5Nm6i+ge9FI9Aa52o
u2s8i425FMaewtw9j+pggzt1IO6YR2W/EYmeZBx1upLW3lwln3rl8AfphSOR4bWU
LmmVkrD7jbhDNmuuvoD1D2ti4InjUzHz32himpRvn57g2WtBWqZYOyWNnS1BL9hS
8L7UBWRdbRzzmf1q+XPRmO3aTMV0gzOCCw4vkMMIBS5ob/0ssRp6sGgozg333ztY
AlW/i+lTA712QTIo4VyO8HAtyIXFOdC2NNBMI4vST/Q/dgwLMmQMjNIvkkzcw4ZK
jxiuJPyibMf8awJlbJ+or7c+P0kvV5qrMHxZcxPWXuCyOmty9fV4avHHTi+ZizmR
7twPXHd/LWazghl/ZZgAtjIJKE1ZSEk3jOpF7n+Eh2CxXIqhlhZ1KgYg2RaUMZIC
vGiua7ZbQsNG9gQsBzlQeEarqLXaIXqP0CQcyD2mpGO1cua5FfFu2nqHvcG4QFbY
rFwSmmPjybrBgzCAeISuLmZZtydgZ2QUPHinNcpytmME639r6XwKK0S4peJdpMu/
vxHbJtDJjErQD+x8+5DxQznxejCI0RJWHCuo/7LyY3ETaSfuQBHXRewcuUenPImE
v+OtAzhknFaASND+MmNc0GNESAwWwtAIeLaS72cNuflMLaeuFtahA20vMYQcWshj
a1D60jKNymr7ZlkzT5Tn7qLt2pI1+g2ReWCjy3Aqw5/aACI3Pcgd8yT5ecVXYGuf
zdkRpZSpgVO/VcVSmwDlK8dHz/lNysg6xp3twJkj4V2l/ZnaeJyAEsX/s5OVmGhf
glsoWFGta2rgCVVXlvCJs/khM1KdRhMvkJ93Vn5lhhu20IqqUT6NDQ6hhTvWYfPB
fvrAxrUd0dbQbq10qi0wqkYFsj3SOOIQ/LA3d89W3UklWfzonmK46aNGIcqSoA/A
rPrjniNFaDBeAIBz/NxTRZF4vNPiXLUFOmkFXdr3WxxYGkUyvX7TCt2u2KYzj25d
hCzz/hP6lL4unJW7JwLHqrN/hJ9Tt6SGW1jqHW46+txUS0JZs4kXi4Rb7fGI8Yzt
e978s3UtpNpCmcDI7VDxyoRQdnTus89LjzctbiHSNXOmTWSOgUnDAIfKyO2BsiJP
spEF/6tPYtb8UcnYgbam1TVeBZUPPS2IYn8ywl5jofw7zqqTwG1YMd5M1GdIVTHh
XRDdr7YG2zorFAl94II2gBw+RT0v4QaUNhZCfYr08qJJ605fCxoJCriM3LepmLaD
kMtIIW3MMUcEcSefHaaqjZaXHxNJ/6kMBLMZz1byaeOU56ZZ/DKdPrRvaVX64t8g
wZNd6T7wY9iXVFvoXnE60vOSug+NX5VNObaGhGLOZNHPlD2kPs4lbwky8LPdMfhS
DoCv1YplKj5dmMIbQjEiF6SiQfBd7i8LqET//9p21Aye9ecAfi2ti1fcpwtzWa8p
WI3ew8woT49/UjOkLRznvYl1W3EmVxn1ZJnCNHWhVLPKfPLXv+6/EyYUcgUmAyxm
LfZWMao6mWtgcO3XTqSReeYp+UmzWbY8zTYE+yjtojLIhzcUYHkB7OpfoPTpWyWe
i476r0kyPBkiIFVkIC+qArtf3Bx4EdL/Pp7TaeETv7pK1tFZzgmzU5mj18avh7pW
cMPPDzQsRjtwGl/eOhmPUwKAjJxNKiMs8MXQ8Wfr85VoVkKepDmWckTx3L+oNL2O
lzAvcGFfNv+rTaaIlCnad5Cw7w/P8GU4GD/SPXRjGYYBueRmoCjPQmESlhowlr7Y
YyQwG6w0t+s3t7NdRPKJN9gXNb+4+YyzvhghyF4gFDK662ibMuLNbdijZpYLPi+w
XIdYnxBsY1DVNC63htW9/71EceqVL+q5AuUquo7IyZ4pg1anaIJ9elAWxTW3LrFC
W8ceBY3saVo/NrLENhM2RKzaPY1/LaP/RIMixv1+5LOEqh8NO4Fq9xClDCvtewpd
yi2juFlYy42mMFGgNDAzQflhbINz5ZQcfwcPU/mzYs7W3IB4g7WF6c+lljLI3I6z
mMPQ1DeIAK95HJNSJQAxpa7FtLtakgJ8BBQ7te4VuMRwD3Glm9DyIQlEjauprIFd
i+qF+dVStvW6dptUWU9tPtU0J61iRD7NDzFBBbhzua56tSVJQfXxmZ0VhsHcHmk8
RT1N80wIgp7Jra2IN1onqtGX3CHZaq4joSHC/A/2V9pPpwAbkX07jl3/sSCysvyA
DA+VLx2aPQhGRbfTenfURfvAU+Kutrlldd+T40BOSRlLZDOMS+bsiy/mT2mvn4In
eROcPPdUAZKJJkzZGSau4+BiZ5Mr+t4TCGp/JJtrIeFNHk/179vsKkyVRkG8jr1w
B/EVV0y/ewf1C3dOTjeJrihQSgUcDhGE6fBcoHMe+DP6Kst7PurHNWSPJk6efy8J
8Qmf7l8PSKb12tMqGLHY/si+l8L9Hv78mf8racuGoWBpxngLCu6uoeU0233wlVmS
75zLeiDHbWqDT12qqcppJs/pr+f6ORVbGGLDZMLqVRaayGx+rt5XQyzTAckrpYnI
FZlvVg9r8EI0rVatRX3eDhRhXESTNeD/fhmlAY06mEAtry8P3Atuspc8Bv5eIV+T
L6kDjQ8h3GTQ2U9nINIht3WyETI3+BJmkPmDMLIilyO6s4QT1a/LBMHaXwYkYKUn
SR4x3CH9Xx98O5f+dTKGzNPeqrKsl6MxW4wr52oJTh8sKV6yShWCkunkHvlrzo9X
tC/hlWzYwSnBxWFfuOiz4HBWl5jPaFxL069UI+Dcq6n73hUp/AtAY/ZcXH2gP7wr
BpONl16JTRuUJ7wNZq9NXnSFJ2FDGxEoXi25pHVjfyK6rJZf6Prt5+XLtgsGhgHq
hmMYzMeOVjcSIJm79FkGfPNPB/AzvwN9dG2oqvQZXotaffOLqJKMVJeJifus8K0N
Jsq8a9Xg/f+rsGZEZftGZh0n7Jyie2fguMbKLjU9fZG/bjVTEZyqLVTxFgWbM+0O
8G+YQBx382zeO61v4klsst6Rc98KuCbjEG93nqT8I/8IBn6aVHuv0teCFyqo3Wle
d8Cwd87MY9FYjD1bbYbhucr/3zyCn29ioClhVqgYrR1P5EzyEjfKXGBpvrPySrq7
lzawqyjY6U7x/5aymwXDgYs7ixiEkitFER93ejBQzrKVaV4z+Se7I03RdhAshSZT
gDPl0ozctbhbrQW12aB8DpsRYv112Nxi63vWT/c7M1cTjAoeFvntEGhP4fMckt2G
G2ODBSulsdRpJtf2ZUjV40oP4+WeQDhofB84XPd0TDLJcXWobrY9gtFRmOQexutT
x1gyFa4FjevxLc8P3I2IhjjM0+aOhxT0CBIorBKBBTxDZcF0S9ntN/i8lwZ3toVs
7ZGg8nFXM9eJYBBlGlDvK1zb/eE5PYrk6idpK4Axpbmynx29uqNVjVJsENdKQ3Z7
MTLSDKiL666ECLJ+BfyMcr629sw+JJYC1BsryXWxEybhJWZJBdAy0fBLiXMq3C6Y
UUSnih2IkWojHwqggA9MenC2Cze2v03WNl6lhWxs7/SqcrP3vLkNhVGVIykLQ6xI
hRuaNh/k/c5hKd5Dn6mCQ0vC5zQyioq8D+qJyCuasyPyfJeLYulVUmBRR+3aAMzh
HfbDw+KVlD0kKsZsjQiigtKeLhRuo0urDpbtZ0CE+7EExNkyzSJ9JGh7WEEWMNsD
sA7uiEWHESPAdQQ9HFPPPLua8o4dtBEb/z3p5E8B9PfnJPI+16qomOiqdsUFpf+8
ebLCFOCxTii5tDWT3xGLZQHitBIn9p10nVPLaa4+x1yFNT2e2trgGsZiHaAaqBwK
iJYXuD/Y+8u5Y+T6WOqrjQ9j4V1HokP3yo9P14c2iTwiUK/tb2epjD8ENZwhzQeA
50GinEmoT+dFbIk4SWePVDNx7HvnP6P0TCIeSs3AdSlNOkMoEXX7VRyBxtVlgUOS
iD00Q68bld/E7JPfk0dEwBZsvJ61srKj+gEg7dtl83fm+B21+PD289HJVHGpxLjs
UxFPITIXd/bUya3hz0dlbPqGZSgPKUYZYnpzVZ7NME/y1cxbtUiHEvJNxcwCqoT5
Hes/gS5Elre3bHMO9nWz7o4zMebEO/NjDJCkDzWUSoCXtJTP8zXHsRWZfiAc9aEo
LwomrUL3tuF2t9M2jg4RobGCDZ4zEJq45N5wvY7bv9Gm+3t7jw6nl2yKFHZaVehj
i6Vo9WbiWkat4r7W6f5GApwhe5YZlFGUOoTzryFdTuoAfma8cOvKgKNx1lpFo9r4
2SRKyKE9KHIJR9qFrZDwq/HZHeu1p2FdZYCPH++FS2dimSIlMhTBpkRDOoFMw0c0
/lTUnwwOFNohL6fIwMj9p5o9w5mixJJu9zgwDJkBxXHrsccAfX2hMlbicvQzanPa
RWzMtcMyPtF2A+bVmRpMj/Rd/eatODBx/Bw850cnFzpPlnATZBXVIZUUmAxZaoBW
UPplnt6ZXCgzeQvNTJanGwbMXdhRm6G4HJ4x5xVqV0n3kkS71H7679Yy+XEEFXgW
/FuXhHsjl1mDezGPlwqKq/hXQX8Hrank2vjKo5uUUgDqAcOlhsxWP4EDhCDK4l8g
9QS9C29msBhMM8QK4kySxi5l/RF0X3yePofsP7jERrYhm2EHjRVpnx7nH5djLgbR
eMzmswpO9D1D/HAD52vXLmZ+TmWYL2WNsz6WvHXoD2CsUlEXrkYZ0NnJgdKuHIHb
oL5kgRpHp9o1YkjD6F5BRabxLkLlf+sjdYq6azFPnR0CkAEPzj2Adbuv6Cvm0EER
Q6JnAqylFu3pPF5U8Q90K1Sn2/6aaJz3edAlGr/GGG2BoYjTMWahlFBDl9FCMTWM
e2cPZF6/gwWM3DjFSSGqdIPFMzwR5bD45bLDbHMaWA+onAJhKx00AuY4iPsLho62
5r+83iAynlWiH5z4twQCR40xAn/iLZOTWW6DvrYHWWRcFfatjKIfU5U64rW7pnkr
G+l4BuhdAzxbkhJv5ihrnGgMssyKwu06zHmwHycjzAgcdfTN5MlvF1V6DruNaOdh
c5DnZswI3GJRwBnaSLGyXGV16AAyg/bo3sLcp3vWOTOczXZ+lNv7RT+2qTDHLJ9p
0N7qd6WJD4GVUpYt3ghvAzlvdE+VmydKLe+6CsnmRe0PKBN8BaC36nzEgluELaK6
o8d8lhgaLKwW6U1icrZjd0i6IMU+lpruVO5aoN+heehRG4XpfF0a3DuWxdMPXV7J
paxdYzX/0dy8xcNW4OH79/j3TzC+IM4fI+fmnCsqs4of0hcv9s09XkU90ISdR9j7
39nJ8mjwxL2oxn1h7iCjiXP5fdO8guHT0dLiE7NcVFmZh6E7BOPmzruBJudIolLH
6XHLIQ37Dq6j8LKuGyW8T8xqSxIOhEs5nqvMSCxRCh4u1Pxd2gLqyfCOZXo+8n3N
xwB/9vvzwuLe53PKlqMNPtJ70oj2iKuyPTVgEiRac4qdgUWYdzGdKoU3fTlCVyaR
FqHN0MckLtTdc4vfy7T7FZHSJybGO/P7/YwvS53FfD3JwpeY/aBToZgANlGup/1F
QEpgomRcIEROBIm1poC9X8dRC9PpH9KcWVwmt+okedg6JuE5Sx/3iBbYHxVVh0qi
8GWyioLVvZnhowHaPXIopD/dHoyCihj3VaxTSXLYeSBqJCHa2v9NJsXvdSLzrrX5
nheGtpcMwk9kRyFqaaeiK4Y0DrEZzH1YmqKHkuFr99fb63tgqHkVlYaoyZnGXmGU
zNgaMxamK67pLN6Ov/H1N2r8ZLvcxm3Lm65J8annlHM41zZbn+77sZNb18NGw9vR
8Gx6Wd9j8KjdVkFHHIgSWFWLS6Vf4lyIKnKcGXpbHQu7YIVZPmZD9q12itXMpmFv
1Etvvorxfb7GqhcWv1DfO+ZbvQjIbab8ENrPHVylfC1wT8E/gl87zZxRfudYXpY1
cO6NoUhyPpHiw4Qat7oJV98Nr7gxJYF2VRyaXlblppYTcnU4CaBZ5DG7acMip449
oZKoOZmVkt5m72/m2kvVSo9BBMRVJhHerRK0qo/N0ClD8gibwm0FMktmN6erYmTy
IRsBxzNB4iBLJN6oPIzI9yZbBqSJnkUtR/lIInNeQo8czuv1VWZLTYFDPh3UtUZt
Bfxq+sLuwxZBsLjSEyz3UpNYBps0ahGzXB36oFuFn3Molk+X3mlwPLT6VjY2wBpU
U6Qu6MGX6lMQonX7YSpYVmBGS74RZnCmnBVqPXv8OKN+F1XQ9EeFocg7PVzS0P+U
s7YtBtodFFqJWmFe01EJP6WXdDQeDr9BaUH73OcaWJoOBzs158aI049W9XeXeN77
2et7+nzh43B/T2N5iJNp+f1KG3CXgrULFugupmVdQRekfqfn3JJVE5vwY0Iwcq8f
4x/O/gltkS44ehHVjmPFjgBW9XiCE1VeQwq4P6CZY5XJCwXoqIvF+LnA6yxGCsaB
p2JGD4RwviBQtptVcnUmZdZ4+jjDYjr5AofNKo7ZFDKHniEnFqtBqUq6YUdW+3s8
ipzIzmy64A2b16JjrgYZqjHpr3evsGaAQMvRP8G179LJHq+qZhkRdKi9Q8zyTekQ
pGfqnfSASYLucdewm2SuUulBAC/gJmeIhoTb4Vwez4KlTJ+N/jJdgDe/EKuKhAra
AtX38RRcRErShmOzI0aJzfIHbopsl3ilcYu4T6SyoLv7nDPh0EItMmGL8co4HaCo
TW4FWb/VebM/b4QMrvNWgO1N1KVPKxgJJAVJhnCp/hCeaKqhXMQBocNfPTrP8pEc
iQneMjxb8mfGKrMW6rMTc2YlsQrhl24/5aGE4yBrwU42KcWB5pv2jgvYtPQxwRkj
LsLxQAcPSCB3bSB5MU+bOmIcliyl17tCRuV6lqLyJkhmtkPSKGYD16C8VmTxAbTt
np5YKYFh2vNQNerjc6HdAqxkpBMoirts9ZSD6Y3OZ122M0NZH7m9SXMHBa2Xws6o
ZGxA1Ze7D8rEwDDzuE8njzS2vHKBN1XgYYljR3I0tk2wmq5+jZkx6K2ODh3DR7h6
7vCHNgUMKItn/8qlk2bU0E4BBgDO5G7iMiuL1jXFq3PKpFM0OgVBQKZU8wv9oyw0
IetbXQmMzV9N22/EKBZV29Mi9fP2w70d+DN/rPVT/coY1vl9xD5heYGZCnnJAIni
7pWaRF6AZ0HxVDrN1pqWVXUt7R7/AMbnHC8hoQruo4Dv80A5XH7UUMNlH9QQHNp/
QOr1jgZg1ghgBCwb1HKPbw+qWfKd0QwsW8DfSJUX9YurOXEIMXbbaIFr8vs/jh61
M8YtnonUgBydedAR5NARvt9UA74F+POOGr6CPDAeeRoRsocf7Ux4a5yslNUyDXyn
hcqVyKmn5P7K6kuPGUaXGAXUZTlKv3Lr3WW4OYSaKgefhH1KXk9et8WgiGsxSj9P
s+b+Nm6y0XTp/Gyo/0b8NEkG2bIkcBfFWII9hx0VjNXaDY2jxjC1zTFFlkbi2Rtf
F6TIdRXhQm9Jq7ZKMWu3l1qxgSJ9F7ol5OMQjnU4gyDPG6ZN1JlAKPWmaOOQqQsx
t5/5v2/AZcxvx5BN/uhPAFEuMixLesE3FU2ENiEzBXcWdU+gcg7MzVf+uzQoWdcB
TmB3DjNvoGed0DjH96et8ZJBuBoGus5Xzx+brYs+8WZ42IRR0rhxt0sAPz8MmpMi
n/M4wtwhfeOmck1abXuV+0urEMhnEeIyIOdTc9aoZityHH0uGavXwyyf5ZiQFdSI
uQwxIxJmUYu7TwZTagMC/OKGEP4srBaZm0NzhASZlyjYtMKJiZlsHHvblqqE6oGt
Yfc0Br/Dols+uUq0UE0zU6e0xLIJaARr5yChzVAUxAkgNHBDrnDW0BrNLTk8osVV
SMunGkJHXlab6AC3pA8GlR8R3MvFsv/2gwVUk7jT9D9Fe6qHebJaSimzS7J9cxGR
CY20o8IbFaO3F0OrFg38l1zZVHKt9AxYBRZBMy2ADmx9z3yMgknRXOJxwn+ft/Hh
I3Ne9fsSUnnNkzRvcst5WzE1VLdGfn6OxHdvEqqzrAW5CxRq2u8Ta4qoYNuW2K1j
Ui9X/PN94UpHqhHmCkG8UFPH3JYoxIzUePCTlL2xrc5hnhmu+sCDzUKVqHzaXeN4
yW7GJVnGGIZH2SnukkkSht+ZKiClR1r95OOCgWeaDUkx/rapwloYbNPkN5nUrAMp
ATolViQo/rEV2C7G4w2uZluoULiLTIt9Y7DnN0dFuljAC2PrPm0TWCfMexnG5bpl
nSxM369BQlpgNqbu5huPgp9wnBWenbWps9l3obMdqEFc9uOVQ6F6JKFxE1F78GHj
WYp4/bDBu2j4BRE4ybfHtK0+Pwdg/ePKyfBO9HxtG4ChWzUAcd0fprBozEOH0Mj+
7phLt6eynyFei1eXLFXm0kuHLP0nAmr9AAMW2bAli7XkOxxQoY76/fhUx+/0iLop
grA4RjuVm5E1G3BvQ70kYk2e7APsil6EcLHN7KAL14niqrKktET5Tp/0gTZ4LH6N
v5jR85e8bLOtEMZjOO7sFxqlcpjLNXOEN720s4JiNktGJniKNFmmsiirc89+4FtX
nNKhU6/0n2/+GtKztGJnf4+fmUh2dRCaV6krzYvYEi7Bs027ifTsFmVwv3YkrmUJ
YPlBZYe7aTbbDyXcW9UCLYPnfbWkuQvHF1y58Tv2/5Xpre9Gfoyi4iCZQPMFrrz4
2zks4/UblYgbJyT0xEOjJ3CLXur0uTvN+pzW8uyvk+jy5BFzQLxoxlm0nLA8CTY/
YClZE1RjidGOIPSAZpZnKEzwxt8INlbCPRqMWTIOV3aPfX7DDBZ5N7xpz89QuyOd
a0f233wNuu6HjDPovpS1hXgtMKkEEucZkiCYZm/nYW4KaCzIuGJmmDjSF0vJvV2d
+DRlb5+yrUVG4E2SngcfRTWWDnTjuVJaRZt8w7xgXDA/dys+8am/j3I8t0NgAUR+
Jh0oztJak9cJtbXElbB4sNqzQVmzD6WA3RtVdRH2hKEUojjyOVn5JlbzuFTvQ5QW
E3t3Oawu9kTMTEeU6nxrpRJF/7Nct2DOqATXAAECLbe+8Wo8v2Wq441Vafb+GW/U
qESRPgeB8cJIiTTgMLNGWy12GpdL3iI80LmlspB+EnDF5von/2JmxJqcykYk/TKD
P8WeX1RgPPdrXyTSqZENCDGVjD/pIce+GmfA3/qkX1OE+Ox7kyx0cRwdiKpdWosN
knBXBu8Rpu0jUDS78djj5LG1sANF7pp+UHZS95o9rb+tdFAKTXJm8euhTQ418imm
IdEQZV90EuXy1RPxLCIBIuppPHrZ9fSuHbgYUAMG1HacQ9Wj+aTBCXjQDgN5wUOc
WNPsd7bmKq1uz3M8BAlj7KK6adPvUlPzzGJieKYScdWyazJa92VzBXV3BOtCTWJ2
+SHH1VtEhYnww4wCSAxpzZZ1/8svIvIwugCwfLsTvlrO76pa3V4hlv7thWQLYoRR
GZvPSSKqd5+ZFAOfXdeSG+nu6lyRwwKDR5FfkMFVYVk2ns2rus2e7q9zvxRx+Oz3
eqvLk23agoA1UpbYrFKqB5vuXftjPP+ZtyD/ayC+nuPNiKbWQlokyIvn7FTIYGSz
fvUwFokKQ+hggM1eRJstHaJcDQzsdu4psVTalX78FPSpFruFNuxMfClB3NhTubld
iADanqako8CsW/32Q1XOGW2gFQv+9SG1ScklM7ncrjHaLWj0xEOTvb0OcQPih0gw
EPyDpPy01oo1GsrMKpNWkRgv9a3rvc+PcHx+Y2jAm8rDdkskAx0qsJ1TqoEJIrEn
+RExbfRJ0yN6n1OwhZwBXf+EhkxF7l6Fj56RQtfc+nlDskY8mIt86xX/10vl1JfP
kRiXdvo0mOPCOIw39oZLhiC6ikaju7+TGi0tyMH5XtOv+VpddqaosdqtVLDjD5ob
2oCOrZ5aCp5XDtawdV30Ry94XIf1x8Ni4r7PJHX1ZRfxrAIL2elm2LCKvBxV+7jb
imHwm+6MotHfcMxiV/olFJqVXReVotS6vx+hACWhOX1T/WK2iu5oR/KBQJHpneZN
shmZDNzKzArPvUHJFsqRqna9r8r+bU8v3efkDGVMC0JPU8VvXLNd1dVyKopY2HDD
OsNjnHZPMMuYkkwk1qDBRHV90OXJeG2b/3kQRUjWbs/O0RkcxvI6wH43TDnnTtMs
yqxZfxVNT23rxHIoOYoOEL1CXkyXo8ladCe0Mmyi8Swa3BZp5SQAG5UuREX4tP8F
EhMOTnI2WJ58q7mqxY2/6QRSxxQB8OZFT2iBh+0HfDy+TgxKT+j9uhR6fftHl3Pc
ezg7KHEQ7kumv157tjKWFqDsdTfEmCVRf7/HdegnBZMLI3VlmW26350KO+ryQoQs
5UU0WrCi1lLhmfb4Ge6mh8WE92Vy3QQHw2+lsPKpeVujfyaleD2kZXmEN9A/3WL5
THbvR4cMmCHIhJp92pjNhh/bvtjpjUs7uRld4c6rQled2zExyfyfEfK2eWPw27q7
Chjwx9RS3H2DHQio3Iw0DcE8t2HUGP6evL0+F4aDOnmIDaqm2A30JyyI6FGst2fs
SCZD06SsCFMgGsxU24rXIHJLN76+heHIdzhJ+eADrz8k5LISVjFWFMmeF/uPrd4U
yM8VRMc9J0hVQKhBw32WnJC+hkpg98rnuMylFVCEpHobLU+iVhQ9BqJJVTUr0ZtE
wWsXI3n6ENlhnoUUn0YbHoZkQqH/WUOp+F0xZ0CryeiPbM8q+txqMauojKnUm8d0
2KIV+s4ar41Bnf057jI5CMdAwJ/p+KPnUhC1Oi79vKpLOhjYbQMuJnc1+S7GQQ5y
fVZkHZ7sEg/dZ3dXf7wgtdN9Ij5hg3RJt9KLAFca950FwQWRk21WFfLLutpAOd8u
uTTugqD+AWP+q+kh6vbyDfzBPLBWJvTf8Gn/Dz9fQPyREbVqPAhTjX87S0S9ofgB
3qyEORQWOQkKVedK5K+9rJ1Cew1fhc9tWr1eSe0x3IZgzxz89dyxviuKGJyddt3r
ZbzdM//vnLY0eB6Sbo3OqBiHwJQkC+WIUGBEtFbdT+QmDvcnmaPMedkl2hwcbnxZ
9TmveW3DlXBzeE6Atz0WeZhxuqwfDsL5XD7usBWCgvqdGPo4/qz5iVovZBNQADqI
1IYYT2yoDpH9XR3Q4fEwqCuHjGovGi6gbdrbv+/5DumhiknPhBFG6KTC7/oFIvQZ
i/t/h11uN/CpbMC4NPO8E8Prp/e/c57NMrLK9qYLcKj7C9OQrzgykLJmWyl6da6s
QUUuHi2YF6JkI/vR20k9uM/31/GMYJORA3ond+eduOOWVsafOcYpzQ0+T/USSfnE
f0WUqvQn4+9QKGbeu53H38+FUYyWZUybNzepKT5GPkScBvq3gphZMkrktHddspgu
e2ZkZ6K9qelRnWu3eluMh/rqPWGkJs3LnsVcX+5dPiEa9gfXLIyEsAQz+twDFt24
jtnLSviG7R889woUQYfX5vWvp7pVg+F48Qn7d865eIz1ihiWBsq6oV/tB0ilPTqn
ewJVF7I/gqHMc6tcLJQEGjjGHv+m5Fa+pNAMzJcktKw2Pp6EqoCpl8Y8M86HElfH
gGZvi5Ejl/rS1xIVFsZ+g8g1Vm7HYZXYX6nv6NnRZr0ckyceNjbUewv/f/HLz0gC
c0Xe4f6YE7nKjih9PdwvqNpKblgglLk8YKE6mch19gqoDemMUi7GkUTorRI0eRjx
g6R1jepEfn5fmFVpF6H6jJwjOu6OKdyilNwG6o+vH+IqLt/8WyJOI2+z7USPCgc0
LwfcFhav8+sO7MPJbYQqCDWFbkr0IG0MiT/AjpPzB7W/ohjEvgkUAPHin+kwRLY4
mvRZ1+OTIfo7pCq6HcLR8BvqH7Aty3YiVQs5wWmgE6plpfSLxe3YZtfIxEuKZCwU
FCWpQQNfaIjY7urKQmLrUzAtzy9KeAbNoYRN8H8FZOE8uvGNwq+ggUkr2uGXjnee
VbUjoBhvxwZtHPuESEMDKXTNk+FYiQOEzDy2CW+mgkWuS5hiKA/DJkCRYhHXnemk
utY6s/QYxS8lGUSRhj2yp1LX1vmqzrCQoZs8tKDI7q0rpBcE81yGDmDrfdZ1LFr4
Y4C6SCeSkLHlYK+Aq9H6umFqsblCJh73v7cjdZxRff6hPJ/l1aUDr5ms7bK1gr0w
hzU5n5W86HlyPIig9FdgkdXnh3GSaHTQE7p/peHk05WhijuREXjQeUNhFp0KkbaX
KRNIk/LN+jOZq2yz7dT5rghHs6liD0ZHs6lGUqLQQoHmyUKbHxZcLEibWcurMteV
rqZi8zadL4r0t7vP+t82JwgT4kINBgHB4lm4Y7tQrSWQhHON2xXKK2h/z2O2qGMp
jjcYn2sOxJN2FSpGy7EMqelz+71iUhdJ5sB73G4HZx2IG6RW3bSg3s+oVsdbyFFG
hcQZp6ZKQLImmT41UTOdURyTA+oEadFWLan7jrJxVLmIhgVDuPPMjXha40pMoEqN
8MZ15QE6B+CrCCslRGegW7JMkUQajTWyxHyZSA/E3wJxI2DeWMev8a9cyx0p/Lxr
NXg+AF8Up9DlNPqUdOFQYmskca4pDWtldg0XHXLrWnS1SLW5U7ZkAdp8jA3QbWqN
M2r7aA1+x93Rdv0GGpkzcwsCOoDo3PMYNUNuifTY0pKOu/d+Sdo1NQar1S6QGcK5
XB8kptTXgdIS8fbvJM3DCiSIdTRpysjPKLum7Kp+mIJWGJ5Ar8kwQj48l2zBYHhH
DzeQNy4BYtchh0xbe0Oyd5ylgRr0FnzdqG5DsEkPWnLmkP8VKFIiBaj5BwiQ85c+
BZHyZuQnV3O0IznXrIEJOQ+6WiZPRQ02FBTYzmAa3JsEMDgEY4CAiFGA61h8NfzG
1+fu+VO7i966q1zsVlGR2K2cDNCE/3Kt4CgJ9h3ET2/Ejp+tsswJRgcfrG570qWi
ZcfgpDPOAKlKfW7AzXYG62VHyUgLJloOCf8G9dM96hYgWa76WG151w/DbhRCouBs
gNwMQb2+3lmCLSA3TJnhWw5AQJayiVBR91dzYg+iLW0UWldMzTPpmzIYW2orS0sz
mAmSLmWpAqWzy4pkZj6Td0TP4N46NtewcB3/QTMsjnUqn6FOMhc5qf8Mzn8JktCV
sTmsQJSxGIzpcSws37FCE96PjSpeLR4cwpudD1Qm3BXvm1W0pr0PxIHD5XhACflI
93daGHCSkhps1wMDu46U6YUzNOZvGyF50A9olhZTVaeOcGRpVvOVOzUIqTYL98wr
8vke/PBTqm84ubNEebrPq5jpLVubKh+m8xivVMk5BylRB+7aEuwLy2Tr0Xo90J4C
CIZfTV5Zoo6LpECnYSZo+LBMwVi5kv4R0iJk5BPP65Sb+Egy1ScvxFQoE7FhEDTZ
Yrf01gyXIqsrsTESQb4h9GGjbg6zWJXtcKdp+PtF60kYFyfmbUsIWvSm1ScnSTha
toY+mm/C4sLKl4ECY9eX7xgfDzjRBXvWSK505PDontNADSQS1bbHRGi36H7vLiSf
HhA01yZoNOpgBl5C+KwnyMgWbH73m5idM1IpN2Ls5u+yTnlQYJlL0bFwFTI1J5w0
Pry/pqu9dtxs1WeXdVLB5zA2M6RwRHeU9o4gcDN28uBZlHqP4WuPpjXc759WWUxB
Zik2y5FxTB/R1tcUJ9kkSfeIR6ho+1QaKbiqpWjQnADZmDTBvfP7JmVdeivBqmlI
08Pa4M/7adTpM+5q110Tb3ZsY6uqXEK69JP0of8siiZnESYSqJKn5Wh2Hs4hKjKu
hdjR1Q/y2oYb4GVUrxd1fvFju5xybvoWOcTZaaZRUfeO+aeIIzRnMu6AZAGGF7ue
O4Uw+kWqLMCwC21JLgffz33qhDljQK3Fa5XZ3GjvZ/BWK3d1qgG+yHSY0zvYy3CM
nBci2+5F+zqtc2TUzwkszQJKuonuMRbPldIxBf67V5jQloY+VB3noyU905bqnPWV
quBD0sDw4EfMOOPsECNFP0sjcv8Yor+tFFEQaGnSTd1pXmUnkEAdt3WrcqgXzo5z
PtvHjlZKC3EP+yyEney55BYjWq3ieYE3T9dy1e7EF/A2bC8CXNdq0Zc2+E+3jX0Z
hJbLlu5/rdhcF3HQROfkh+0iv2FJf1iPP4VYdIFAYCGpSCjR2/8atvxCpwBOCNEo
3HIPkYWtmYH4A1CkIvL/agrFVbp3C0ydY+UATyVbX406VhDIS4UxEFHkfD1EoVWL
4stHBeCYrgsk4186g+LyDUa2psjJK0cZIMBpIe5l5bRQc7hvYUM99tTIPt4bNqTW
ajOuMpWGuuOR1qADC8DVMvhOaqqgm6hy7qaBqIe2OwXI/q3gyP9FjmxEXMsaVnP1
bP7FOx0IaOl1W9V9TRxVYkvKCCFSIV7+Bj6ES8d4q5SN8aRGkViA5sO6n3zqBGQb
Y0HS2nWgeiRkWlAMFruvAvrR98QitzUdL0ntymDfNWXF7IrhLj8ozf+OyEvisdX6
9MoiIViGfSqB8DvCOVDnrL2Psy0XLM6Udeq5ttUwWSmwhv1o6R78Gzls0M2xBXnn
1qA2TAtvjJ6iJzua2KnKxAe3dam+5cmmuoK53qiLJgNZk/isHc5z9WHahWAI9ZKs
+qsyzaxs5lRfPRBexYvLQshNUy7/WQklVq2YDzPY4ygmvQeVtVYaLbL2pDYKCsk6
iQFtytAhbyvgdU1YNiHI2XbAMUxH0b7arNpdsQlO/wB/reupPGRcM0SMbbXE7gkS
2lBRQB+q3N3sg+YGTh/17P3DgpfPSYadQO3dtL/0BalHJF5IWQYN1T/sl4KAJDF9
J0iZkLoL/vQJoDj76dXoWXD4s4KpP9YJS2I+u7573/D2ycS82dyJsBkk0sHrZ1Og
0Ay77GDEWI+G+KcUODXTX9EkmNFOw545YTeUqwCXIkrWWk7dIeyQWMlhy8G+2BwM
L1enPe3v9kw85D3oOZ8JbQruVQwMH8G8PxktaLcnsDmYfhQcjTM2q9NmhUli9WMB
WuVS4OhckKmAWDlN394HFDUgaoeUpSfPGyWQ/ih+HlX6rTbVkoUJr+XmjIzdMDiq
vVDy00jDTECmkpuSjk4kNlMPFGoMh8G9YYR5bmloiCgUbBeTQmkg+4yoe3fc4EWJ
7SM6J44P2D7pTL4NSfjdJtLXoP6e57b40yuMuNvBWUGNzWAXfa+F8WlXlvPaBJ/+
F2OkpPLAqlTa9UOdI8FdjmIifTR/s7W40S3YCBKxBvFU0BvUsdrGvsSUvr+kO/7i
7gxA9XnLZ2UstxmGpthRz4qaEH6rfOSYXQDfgVnqRrcQea5uKE3E/oHati6XCZj7
Pb+5MBmVQXZ6ZnptInk/6ekq8xUZBHNupq314LowuRYXKB/wYBB8bcBTaGhOLHcM
fTL8PmcdR2gs1oAVEiSPtrXZvLBEFMhC1k3ek8tPeBAhTMHb2VnO9O17HGG9EEdp
5nUVQMX5rblvqtpZ2dsfTgLzXryqi5SpSsLboE9ufXiDVqdt1T2JX6G6wAt0QUcm
ttEMSBtK09nfsJKrnvLrLqgCSuxvZlISwRMfiXrP66k0lD43NmKM7UXvkVrX6z0g
wr9iExsILd3f4H9mjFuiwNaSCZUJOtiawFvHG6GT32h4Nr14nh6kxEuiR/HUmUY9
uocw/u/1KzzinTv7n96azK3ZYnI5SRLZeJJ7sU+hbAYcyoxUA9sPKqY4wZ3eV7qT
VtenKG/h9BNiGwNtzfnyUpfBOmFGMPDZ2VuaSeEk1T0QCqlTwChkPeeIwLGW0Sp3
dcnLNq+aQJlw7tTvT9hah4s1AXuJNdbYxhlFfeI/2p5eAMXVTm6yi4Egj08VsN5D
nwmUDFpoRIuCFv3WtSRXVwQQtBKCpyaoaa2rZ9cM3BrwCgNdm8P/KQNTfFNGLvwr
4Ek0O76mwQKtPGPi9UF33386sBzyAghZSI/pzUqLIZXY8xXktttloGb2nqnuAn2E
1zyuoIiIgHARQUCi1c01qzGdh6vcTzYYqgViIg1a7cCZwksjXAc/9G80T2ax4RE3
NgzU7sXJGRaOCRLyyA1DGJUrEGKQ4s1RzsoqjOGIEy1e1Kk6cB2S6gcxGpapyIUN
kfsBqw/pPYxSafAIGPJtdfwKcItXocqI7y0Z+sTzTBw9mG4A3N0c30Y3s2704YP0
RVvORVUmYiniWjWDHUNJbJQAPvaBWi+CAQ2VoR/CelXRU9D/lrl0LZzwa3OEMH5T
mcafoejpt3Q9BquHQwrdwXyfAsJlQczXsD0aQMeWXONDmExfit9GLucotua8ZL4J
2LA17J8hxAeL25TgplegEbCq24aDamPa2Uox4cw1ILt/1INm3k8AE6d8mma/ZIHz
CYF6fFwjkR5HYwcuOuZdAvO3sQM5z3vUkZ6gQ3Flp4Nly2GYbhF9wh+nmT4668E5
UhpLp1u3cduZTm6dRTwaQxatwwveDPwPfznZ9doT3p9zaiMKeXtOm8tnyORtOSuw
Z1yUimLmHwdhI76tRK0usOR7YPW+V/Mu0xPaY4mYclZHHZBiwT/atCJKutxxgWux
qG8D82IHP0/7REhgc2NctFnvnhoIeH+9ebPeWC2CqYVJ+rBfJd4T/roVD7i5nnC2
rJRcCnyaTC1w/Z7c+8HyfKWs5OLherV1j++cojLHpS0WzPjEvOl7+JMYgpLuHTWD
4EI92O/3uXszRPp6i+u7f/RO7HXTXCXcsmalxQFdsHhA3UvQnYJNlp02J+xXBfkf
qJY6Pzg+IT4UG50IyXPp5X1ySD7/RDBMcp47HAmxVsHuMVYtmOwTrKTOWK2HWym/
UMWAF9a2aGo+6THz8IXYLgD/8/HCZZZ1OzPReVp/6Q31dNNyb1ZtwW6CNnSnmzH8
MgEZYa5eLqV+LR20TUY5NxkqKs7+StrGbhI2XVHeC22Siommm6lVyadF/vEmmeGT
b8K0lTABsnVUSxm8IqDF1cH9w9a7+F8Zc/NfwtpeReZJg1RdHPCpOTj3n89/7dOj
iGwp0KOkQhSTdqS3JIEBtU+7qxsxjA1t4VFjoXcnw/Bi1yFrFMoLP2+o1XaeCDJU
3Nb9lhrRmovTVCoH6Wxr7tY8LIPbs3tz7r8/0cI4TpUa1U/xYzTaWVof1PfoFph+
W0qqg/5uPcE6XidrqhrCZXLSsBm2G3tCvckXAsiPY2l0wjrBSnHEcndA89n7y5gJ
9L7iK4uSWNK7o6JYeXvxTdIoE3qpCCyXy48l87ebElnk3kfE5EQS8K0XvBPDMl+q
fB1EChBKC7sXQD7PURvU4+A6uKtlunUstQjw4ekeNXACS1kPlw8cOQmbFguWRQMj
hVyBejlkZuC4/ZYdIDi1NC8uzG2j6bxsm1eiA/aWbZ/FcvzbF3y+SPa112D+gM39
cvW9Ayjhqak5H91DcJGRWtezk5++1oRaosFUkEBYVpxM7GpkLuFewDbVxMT4KD79
GfJrzFwQL8xK2d76sjsZNKmT/oznro16Ixp0aNWKiKibSkdkeW+f4Ta7k5CrrOMu
gNySu1A5BfuUtV4pIzKeGRE/tqeshIIObOoedCSqIwTTi1k4Xq/Jb4p04NFKD+x1
WBT2A4KhLVo/yIW93/zd6DlMJyKpEeb1o2afYAt+9wojSUCCnNy/p3KtYtTvHrVA
Ci8VBKUfq6zKCYx3pTrdOn4x2BSg8kvRMDY2ooF+XCd/pZp9WaFQdYE3ohnfkbFM
PLB7trVTef7vUcytozbjBfG87ci1eyCv3j9BwDS4u1Tq42Mfr/6ze/+Ti+4aOwh/
7eGz/Cqlv/oBZWaTM9v1P/VFYHCHiLXFD+dcU4uiFFymrAEy1mIndHP04ujkn65t
9DfOo8rr9LQdG9LrFlx+IjkEyRNmtEXM1E4AvgvYtDrqs6o/Mm0BpGIFqsEQxZsl
7sagVVXbPx3X2fo9kZmiwV81+X/6lMMN/fRX6GIUPH2a4/hWvdL7JzM1H82CX6bw
ygUAAKMM3g+oA2UQR22NNbCrlg3fIEYXVTf8W/motLDAR3yr5XBFA7vWUn2eNNtM
97qRBLSk3Jaj9xXt/b3r2NraCmoiTPn5cAGVNz+bUzX6ieX2aCAAQcYwuM5xu3+k
WGi2NsUnfYyuf8LJpYYEKWoi3kWCWMidqWbvgF/7cacVKZrJB8y8TylLOR2QnVAc
cuGf9CfAHsZhn5CwIAhSn6NmLvfgPVU6G0rXUqgiiLFhEtCmra89TJSGwT/zoOyU
m+o1UZCAJ1rIQu64zNv8c4qCDIP/0DFRz3JEcOXux409Q/t+TWA2a28EHXnw2vaK
kRQNIIq3Hyhm7yOBwNA3bpPd/ejx6EExqNKxp8P3Lkt3Mty9PI8EqvCb3kci9Czw
WALNnwzrahh/9ReZjGj1p8nc1FhJZKhnfjJUstfM/gLtGH0WU5vUofJ1fMCiwmQq
p+a6/KnhqneEpcAJZ+YLGiFKVIn/30PC5O1UJaHNUXLg9RlbmQJyvq3JvrNr+EC9
jTbPunaw+lR33tEczNM5GFXUZoq7E15/gnJknQvDGdfSvnxUoYTU5jXkErYkY0eG
0bRBet9co5X8j4kycpIustU38hJnvgXHWCnwBV8nH/8TM++tF7cy98b5KUcSTi0T
TACmD6mbh/pB6q/N1WdWfaWjavNzXUb7K/8asdhzz1uagjvJCOia2DPV0LIIccya
dQgZGHTi5y3l+vtXl2RP1kzeq5e0ANiMI/Y9p4dwPpPBdcFVd4rcfCWXHYoPjsDn
xcdZYz+5V87DtwdEKa7lkeCG5nT8d86Oa0hbvJ0IBtZNPliZKWF2XEbF6KRQS/v+
SVBB+6ZXjM3HtNNh9TqBmkCrmdECiF+ay8KSq4fqnooQdnHHixRatfKKcEsSkEqf
0X4LnU8G4scALN25A2U51jeDnLtvAM0YXHRl0XOm/BTGlYs+7LuoD3OEssa9RwGg
G/IlZeVlJPnvuKp0xUnJslYpm+HvwyIoyf/mPMXISqNM7e7rXP09pHysjBrUTT65
NZLGIqSKNvhYns8oo1YS3EoaTWevnoE3uPUrDd4DgE8Wd7ddCalN1uwW3qU9qgJL
hhO/zDlggwouabO75jHaOiiFEQ1YQeYC7BbMGBO7xCJFBQQKVLaiyuxOuPJWeq4c
wjnzbzZTF9aKEnhPF4/WkZ9MggHJTPxQQv6/4GyLJ480498DSS2x7JW+Eg1qhbdX
zE7wnUDwiy+rmL+qOelJTBRKlw8wSpUVtiWwDXRhuZDor9hlMBtG3bRXIWbSVqal
UHZqDXqGCDwun7YHTNBF/xf4HRQ8WbLwygR+AhGYorXtCWkfJ+rF4qb9Zzrquhms
ewfQg+8stDF5zCZW42CAkTB6mKeFgSLe+YfKHqHjapA159l3rxorBLqdnqPna9dT
Mw4eNYslBpiGqXopEtfwSrIA1DDT+hqbd1N/lxJUFyRzQNQNtjYI9HN9RAPheNiE
4Zd1YcWp7iwWgOmYJT6o1xURxqQfpG5BgHGafij+R3GHIsrGYFaMcHtB+O1wrL4I
twHDjLyNZI8m2bdx0XjrH5t7/oOIoWFsdYZ17scj6k5mCVC5vEJHurFwBJlE4ZSH
lok6Xok/RN6+N9S/KsECAfbzesiEM9aRGAjAIoVNb2gJIT5Pe3bjnA1xsuNUyy4K
B68VDky6N1uRinQIzgPIzM/LRyzUPU/ynLrx1GBQJRpdKA6Rk7AUp6QIwdLZHcO2
aQUs2V1jsgmtWehOZKlUrxfYsKkSCyIPpCNj1EqndmCkB4Orb0UbPVUsaJs+wQAF
KOcirJ8ABZBReR9u9ZXnZbmxkiYA9rcnocknll4IvGWDDUg1tJw4vcGi64Mvmr9p
9imPJzfbXa4sVWBbKwUUDRuOauk00h6tveVxBf8yT6EdR023VJGRr9VDBFFUEGlm
NwstycRdnss5GN8hvoa+CZfmW7IAX7OzAiOOGy1zTfO6IOI/+B8aimnpCe1ZAuEx
otzfsR8NOBEmCsCgHiAzxRtJdc4SQumfUNAF2JozoE/9qEwB3hXz2ubd+rkKhmYf
6VPqA1O2bwhNim98O2bU+v649fKO7dM+prHcrOFCOapuTmbHRk0lhiwRiVHDlkYp
6Sig7HBun0Mmsefttbo2UI3vh/k7bbGv5z/zuDWspj6COR32rOrzizAWcaYuAY7B
ViXP85x++/MOQajlDr97VgnKXiq0xEV0OnvRZv2nQYkd2zxMTK/vpJKH9D4h3YL9
zWSz6dNIyscsgtxn2WC4DmLWWe+c/wAgOax02tXFgR1yDstJd4JHyyXaBGIL5+NW
ndH+KiNAwg+aNZW9wLSG3+AGmRXk1hByhsexlnFMrfy97H1G2Oln+IEYej2yxRMN
3R2u15GnjZ84dbUFIUQpC/AeSacyk7vpyun5Q7nQ9eAhe7J2d9QivanKHVyMgv8j
7Suyv48cNaW+eIouPY3XURP7uecZftVI1WMhLZD6e2auaIhKHWsIzenvELkylmt2
j79paZNNpmaFv31bVWMxVF7I8DAaIMM2fHWl/vM6chnYZ5L210PJ1Ve71dywO8bA
38i5kPbMJ3XBhj7OjITyXc892tUIZQgXwNkci0VrEwj5+gaOAt1cjz4VmpmVgg2x
sgfb8t5Was9k2QgHEw3YuhbqPKpVdrKjhnVrmWmiqJwemupuaLSaoQ+2qe68CUUh
`protect END_PROTECTED