-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
ubPSqmFMZKZ+pr2KPtpsw/9/ZkE1yyABcJgvp3pCYYF9WHGs7lT6rdamoNHAh0pS
vkjkTXOvFFMMB1Z2ojla6lIUdWBf45u2meDNr5zmUA4k41VIGRnVemQaF6liWYgi
pa7LTy2Gcxj6MUziQRSXv1LCGNDxsozYsN2L6jMu6JM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6000)
`protect data_block
s7REMmmsFZvbK8v2CrOwtVPKlALCQxrvkJ/TZ1nKQq+bBCPVsag7TWJ0jhArcmy+
gzTOqdHsVv3reFz9ofhXThkpIa+TEdj5CLq3KRAoeKK9xcEVolM+1ADedYdZtvpO
GYGJT83Xusl/zWoXj+DoBKZHdJQlELJPypcfOUbNIymt3wV9pomdjPEbbpLLwXLk
0OjS18p6SMSszFDiCox1fLQ2Ke5cved5YEyRJEmAPwmVKwbWIvlbwt/hQNjnQDh/
7axhY4pqdswm6b/LmWnZC5Z6gH9uXrmDKKXAXHpeAGEesi3IRwPXIkfdFNB4vbNS
bkxwseLeWmVIF7yY72HFkcyk2t6pb7SgRXLB3orPgleNPyt7GFae6rc+SAvfpppL
kBfmihg57+VflyhE6NEwpuSsSHYv/Uu+vOH4JYJsx82d3i+kWQZDZFFs0niRCIQg
8mb8gCr9YUtRfi4Mc1I6icWPKtJc2TjRg7gCt8vkKhY6Tlc8OLCPtA9zKi/MHw1g
gOnJRfzW/2qiK8TU00HdLCGi9mCowDyyJfBIBRD5NrnzRVbAQER6zTdTCwB4merb
2aItP2smV8LG1DGCmLNQvkD+VLSwwQ39Ffl0V84g+QG2VkWeSbfowPW7Ll8NRek5
8ViTyBlyD2xqB67hAd1TneLU+vI5pRWGT6DdiF4ArSozPwvCDMlS+qdjvGwNCipq
g33Oww+Q+WFaEQ0NxBEUG/XuMOe/Fbj2r+qdKgfV46E87kp5M2SBpksljwXya1n8
Scqen9rcrkbDcF/CCSZgaemXJPrJgvTCmpIt+Mr1MnzKdyPRoMg2xoMFOp+xTUZq
QGg5G9A0864YhrTsRKn2Un/jEVhrBMisUiMGdDsK7clkgoRsmoYQ+sxQniUpae9u
KfgQS3mZzCDlucfXv8QIjB6EcU4pR+Ri5kgtnE3AWDBSvJ+NDs0ObCKhUAh9wVz4
ZXALZPQsIsOf62pISgtfucXvjso0K5BrtUVETp98z8UmgA76jGukVH94zCZJGNEP
fDWCO48+Bu1MPBTQbt6y4ht5aHqT1vCQUjGj79v/0mPnwXBtaEb2eUxJE7DASeWb
d1oIfjJ2f/MEENCenmXRB+5jxxy4RxOkrd6LZQ0h7uF2lJSIGhhqhBzM6MBZyr0t
vFd/DicxpuB2q2YP6Zewb8xgtzRC1Tk8QVyxP+42eeSaoOeYiMMBsRz3ENjQRb6F
xsBAKAX51AIN3xnd38JaJcH7pLKIf6BogDpzmlj9GbZCtN3tdG4zt8aAhKrpgNuu
BfS/WDd218X4TV/S03aooabIEPuUrzzY25X5auwsAAD/vaKHA6DHQmNNWk26Nl/4
T8C2wEyChlTwFL2zwFddkIhIr9Dui6zPQqV+C+fCfdmGzivYzLqBfKv/ITEJIdYF
OPoYeicF8Uj8vKcgpzY8QKf3CPD0rmZk4c7oOacDLHN5nyEUJ71n8kcWwU9eSAGa
lV79AXar2htwLvTV/Qrm76ZRXbV5cB6f9Zy1R/LK8bWwXksTQTvsnMPlqq0DpG3J
2nWBS+bpOG2YoUFEK2o7XK+qFqZSjlGWOLEmHeCuKaes+knyb8/s3ZkuY3nNwsOy
yvkbIc6x9iX1HI4Fsio5CTGrIQCoeMnzBpbUlQ8ofGlMUsa2zEcbEqkESwkl424X
4yyY9WWzGJ024VDaemwAwdZ7hvbAlO3KgaPOFcmHkkX9/6LhmtxD/tQliByoDaxv
nqXlhIEd3ehOchG/DkuBxTcRDrC9t2fhabUxmFLNyFq8aAjZIvMm8Hl3cLvCTzzk
TwEnhcxH87GOR3mELjq3vQ+9wyno3lDUQ9CXj7PCtlykx2UHPv93QfiMM3pylpKa
X/Qo3IZwcJxb8SdBq5fH9kY62PjeRP2CUTcOvI5ZRakrdlJ3NSn2U6yjxg8TNRCL
j+bHRI6ytR9omHyCwy6/RxcUovsyBu4IP2IzwtggssQcd2CTXsBDP4ocb5hRdYsA
+Rof1iTfuKI6aixgRJ4oPyw7NMXRGO9J5DwcyrOPxWFIY+8cKEyxrDVyBy2Ou+Db
lS23VS+72L6hoYZZRv/x7T8nVOtkrxKvXvY4ATsxRMsTXMQQiMwjG18AKjMFUQV9
sduIYjl1i19l5gJIloqXNZzLq713CZggwtFmwmXGQhPyF841hV80CdfRojUh0Sgf
g2UhJgD2HaOQMNPXYB8HALJEmyVDclvKXi8cEITT6VIXM2rHXvRDAg3nNrN7qTwd
4JpZnoZJ2qfGilWUx8uKFuy+KWBq/Bm3JgQPqh0F+9Ml8QrGYdujoIeulVwORiXu
UJjSMLQr37a19jf/MZDPuuaIQwxubFyXP5JW4ymlRZldMJC3jXad8RVq5tIzIknv
rLXyATwsVd8R5IxoXdRGyGa+W+6SdG+oUOi/nTOXHmqBnW/dn3B/UuBXnHEoqFcB
9TqRbqnV/nf0Yh3wqViqIjyhBirIvPIM97WAhbi5Udd3vmXJ57BwF564T02DfDfK
YqueJ1gUeHIj35t3Gsql3MYHlGilsmcV0C4nqbcAN1jP4VJ5Fjn/12HMUVy8TxpS
MNXiX8n0kQ2J8Iq5HE8qxJquJEGd/XEfntMiaYOnJqJ9FT8MVrIClkX/N+7akrXS
QvAqcpVDrN0VIHpsPLA516StvkbD/ulY3KnNtZ3HyvBWVElhHTHO3L/LQje7nGPt
QahBYDH0xkS3dXkNatQUJhFxmULnGP3ZR8CdU7W9gGPc9RA1GYBAJ4sqXSJoKJRX
5T5lZrSCNUaSzJ8uZnIl4Ax67W3DlRxNGP0w4r4H4PNUgwVJwOOliqrwGa24CISD
UcAqvxn7IrXnfsSZ24NbCGxBbjkZMyW3u0LXiMpdzVab3Ntc2ePMvTjl4gtJ/Z57
fN+yXxpdgmRqJ6BsYKoUaomwIWcI6yzMjQl3918+oXZ9zWe3xfZRqaz+aGAg3CT8
Gmd7qdEjMOeXOIPKfHpxRdFGfe4Sgpuuvp5jWRBXwLqJNsAXC7MgC+Ctre2fZeBT
yOQhXj81sjCFcC7ICeRZhrU2qfgr/BI3aS6tLGfDtVMKj5+AKcm89aduIGG8PT5s
qI/8QH2RHrDHHJHxI4d1bRcnloHi5EH0xSOjSP3vgrXZTSbi9sacWnFLyEQZzrBJ
yPgPHGBrKjrAR6xP4SxgTURQi8/iwkoWs5PSxof5QQqyjMOqEZIC9RH9dHFAF2iL
skTm1eMs0HrGLA8WX3GLBiQ/XCCxsqLVbHZeEuSXDyEmZ3aKRyVrUXTDic7+0CD5
iio7Jc0u7w+raMx2afE5dIYSbEStpsEjTiPBpcSgpdIUTBsIfjHYwmZCFjTdcFRw
/H5Y1kYNVL7KYVnChHGODWIB13RNsFrEC4tNWc1gHjN+F8IXZ9y7BSLVxdL3YVT5
bz+LtRsdDn65Il73FGvAjRKOEeTbZniKSrOfKX190nu1Ggi2JgrK6WS4g1BaJnur
TggxY7ajGpZyr2NOmvacwMQV+IxTI9pZkHDMD3r1j1uiR3yQOF43L5J6CWhYBUEg
z6GZvLSRqKToeDjp7rOsLbKdrdti8siLB1FYV1FHyu0fuIuQfUjayQENeWFv9tLn
8lCWOIztbNyTOr4kX/JIHSPOFfm9cNP98rnbmVCmEu5Ej3v/ekTZ8Z7OxYV97gbk
+cosFhBz/HdxcFirg1ikPNDZrnKYhK9Wx0Vjt98xvsBs7cKqpyyFWnfGiczyyjcU
PkeyteUp/yo1Gt4eATqxdDgLk+Eqcw1AzouTZZv5a1zspTKZjKMekB5mUkluSsU6
pfztmTlvKHb65cvIGc+5BqtJOKrPVBpCrw1naEBEdXH6HSXVjJRWPMnrC/uz/b4C
TqkBf9g6BPYbuOYZC9QfgxTntjqr0XJpU0PjHdPK0Ok7NI9d86GoGZOJdCZp/SYc
gS+yXkbryF+VnbPf3iKSM79UMbNgx4DzrQjIcpUyzV4CEJZfyokd9qjI46XA1jzt
+aJfl1iuEaIv9Q5a9u5ja3OcV8yTIBCITx0Ici67xrzizFF0b1z+h94GEL0PuD4j
FMCgKG3BHh4Nfw91z8mo+vJ+kQ+jPpSp7NSOQ2y6BOCILRcdP0sxDXQ8k2o/5Dp7
CtYKjYCTNh/+4+d/Fqx+K27PJmKbP9wj6rkrU/m+qpKzpyGypQbkXVJA6aCTNlqZ
3KG+NHWln0xDP4rXjv+OFN59q6PnZxo7jyidnyoKkiP+TxUkci0fab6FPgXIX/pC
/3okRsiUmAGiMxsgbjSLGAgKV9tUJ5Bd2cf9m0FmkZJzoLQZyqRJNw3F9dV6usGp
01vSgY6fSLTwC8zqOj4DjU1opk64/PGBeHJQaSX3I8H4lGFKRe8sa2RkoSGeuo4V
jvuf8eRLybmCUUgMtlfKgTrHQWgGdDF8wg/+N6YOBv7PrZxnraGPGbz34L29zeu9
v1QZLsdsbIS4KZSOUHPnxRT0yZBLvi8avx6v1CJYJWOK4FxEBbBvW01uaiqYa61D
to75PAd+hU0t+1cLqG2+7Dl522d+UiWzE2Aw9ALCUrGcTb1aj0kOveYF+oIPJaOm
t2XIF3TIgpAvgcyX/xO64rzySpsB7lfEGqkpNtT3g1KoGktyNgqw9ksk2iK9Ihdq
pbSOVvYyYgCOep01ya3XlbFgnvBEJhIN6KEAwitH2J+PrqkGy+ezCJQMD5SUvrfF
PpM9gx21TdA8UwtTa8V+DIZNucVVg4D+xtIl3FQANIN3ZdJo31rQD9Oq0EsreJYS
lwuW08OhfPR9wW+2bxDitwtsuGSNPotmrYt16g2LQM47AivFTEcUDcutfRotgTYu
g6zfa5FZ0cblAm44h43KGm7KGhlPzckFc9rj2UZu/5dQmMDCDBh7OspeYeldy/Ov
fljHNPKnrI/7l0JFj+yQ6hhrBAwY8/HcTjbnGQhvB8b+CIl47zlIsKmyY8omM810
F5kRq2U/4XUvRTmNDI/+Q+NhUjYCuO1R++m0Hr625ytNozDEFoa4zMKNUnEaNZIb
LZHSUzukho4KtFECW/2iLKP98EH7eRWvFfJLNeBDfJFIvgD4tgA/TFM/DB2hWtHZ
IERbkpu/7Uh6HaT74QBECkquHONt87ErPjd7+74Cbnip3AhuFN0L+ZzmqOzEUYlU
PDBcYo/lWgnyBapHx5rh4JLWRdAFHiUFLiJ0mBL1dEppKKMoiqzcO18mxyYwfx6Y
eqX4glNF5V3gbOW1oa+tNdpY8bEIAvF51ofpr3CEdq+MOKjKkEVOPCoPyKYYHHRW
bW9O8rLXauzXL2CMvRlPblHVe36L7XkRTHR0GBmDfdAkrjyuW29YJaQsrExCcUQt
vBUaGxcgRo4NjQrZXS8nldP0beN7Ogh3BxEkNojsnDp3AKjgS9KATbZ7CZVEmCaC
7Iy7LzopMvR3kbSxNJTo3z0KDd43tI5oskeMd8GcbftFQkxH1jJnuUySn/F/O6zW
MxEwz7qej5WiqO7zet5jSSu2G1BfZxHzfAhJnZYrC0riJMBMwRMBJbwZ4XDmLvA4
yfyFhgu+K1m2TYDuCKBbFohb+Wg8Ws5PAb9p0cHu5ilkMI/J+I+XFt+NApSp0ivg
noC2KQDyTFfMnM/nJJj9otWCFrshNHw0VNdyK1CZjhYChaMZmWXZLD862j7WxMkg
nWwZSj1Mn5mKy1wG3c8qEe9kCc7brYCFKlYnpwS05HRlJtq5iyj9GViNGa1AV4o1
yxjmxVta2FaLiXDTMCV0jYT1hfK2aejEVy+GSduGOtVpOdUMYog4CtsUghnyqZfb
Gwlep85DD1rtjFj9ZxUommBjq4ub6rea0JhKDV6in/jQFalTrxbPmLi3ueHYFKLl
ma6jcAq5rfUvxPrxSwAXoyHAjRUyXSWHHdpKY2Jasl2xyu9IMuv7CR2eQQeDuL+Z
8IOoLr8eAnivyS+1BCnB7T/uvzYplyMRG1tM1r0mhx8sLlbRukvux1GKVfywOcA7
HrBoLNA70D3Ic9CaUz0+ONp8dbvi4Sm1gSaZ2t/uUrR8JuikQ2JctqHohs1H6sZc
XF6xSZf/6on4pbbYIkdpt5fRi8YTrAH0L/88jYjQ4DCqhqLU0GKCHaNDux+tEqo9
dVWs27D74ijy+bcBMhOmjL9Rbuo3R/sCwna260GUUeqRxoeZ0F3xbrXuOr37BneP
eDNYmqERN9J9KAiepg215j83F74LQqlR1H7Nk+Y1NdXnm29ftFS0dHt5+f3HaM8l
oTJAvz5jvo6mQjDazybrkTjwM6obFAbpLf/pIBEE6n7LaiB/tjBE9IZRjprcMF5l
1Vm9po1j+/j+69eTSl/J/tEQckPKBbnchr5YIXTY6AsgPyzljYSW/r3fwhyjnFS6
gG/2GF8R5kxkvQgKEzjJYcegFcqgIEhIOvvYid4X5QODP4wTKlfjasaHdkPyeNXK
SVV5ZJnE5KL+XF5ye/o+van+WzDekt7Cll5+B1eTrqO+oBdIkTrrL7afksfUY2Km
aRz1fpEvZec7ioZ8XeRQYw7RhRlQWa+W7rgsHQkDYUUwSjlwTv/1CDJ9tzQp42IQ
EHqllzHoUogOzFhCqiEuBblWr1zpI6P7wGyVlFqTs1LUUrx7dyAbXSfSDBWqwu/b
i6wt/t00g+4i14AMh91UJaKu38zUUN2We33VijS3gRntpVz+fQhZve+kUz2j2V9R
i8ylgUj1dpl3X4+UlBFmZLiP85PJPOqwLsXc67/TFmmgxDcGoEscYJfYrk+iAIbp
Qm70GEnBsTis+VYQ7+3SEEqj0c8YiT11/abC5INoyRvqvMXOWm9tEVOvSxcC10oi
nWZZIIg6oakqOO7ib1CASIfPmoOQHuSWhg8Dcm3WGzQhBd1eGFu1BxQchPRw2AFX
yQezA5U4r6NBka82MfisXTg/u5lNf/xROWiCbwGG6DLn1kvpn4lJzMdxGdo22iXo
iJqcoKVsLwmEIcLSqszvw4jszE5/bnmaaoEwWjqYSPzTBoxzkrON9jZPIesOGHQ+
FKTQtEv/Q1k+ZityWcfF4e7awpLxh6H6k+sywrz+aH523vceQL5LmiQlveitMhX2
51xprx3WAwu+GS6G8HLnPWLOuFqdRfVu9vphH/hIgdfHEvQPD2DVOwKl3bCCHQEh
lr2cGsSJYlQqPRMrZ4oCZ5pERqOm3LumunSA6EKdRq1t+dc3p1NXkSCW/X0xLi4M
aSm9368BvNFqHPq59B0Ngm5GyUcJ3CjTdgWG+QeARjy+HUYsTO9ckIENluBY5mV4
T5Xl5tXupjFM0w1LTb70bDjmwICLm5XbyfsYtvttMUL/EGafLjH0oMcAcgY3J3rr
cCEdVc20ng40f76SILYV6ni+njuRRvGw0ATUvjW2w1sMDPxa8ND//r2d1A6+86kD
lM+UsXI3sRtNS+9CYKz8tMA2SN84Sg8O5XHXpcTlWt4+jQ65HHHKy8liSgYXMS3o
TN42sKvdWZZVlQUYZkYJfERNiIiD6qWjRFQXP+TbrYYfl87m4zWFdpOCgwYLN9yD
jBUXlpKgD1zpRwCSfFZaxgrexs0ZO1g5VHi+mZcYxj6Dv0ZmQO2kWzJJvif9lNGp
iXiX3JS4rlXjhU7Ug2vsI6k74/wPGjGBcdwQ3jgxwafENxALms7/g0012N0mM34S
H5MT2dMrU9ExAEingTPMR1UiuABJTGfcIPfrZbNKq/g1gldQXJWlJSv8iTo129q1
SDxkyKNQ+i2DJDbS/z24iWqFNhxeWkJOMJH4HwNu16tAVl5H4HK0ZPeEdzTpPcb5
162+AHBQRuAKQDw7H71rgE6aShyEnT1SqAjBdNkEBHPEbmnCmOPSar1Z0GuI2JF0
m51ZbrM94tBKrsxwAk5boLlQkb8w4rpGBTvG+xMCQ0JlaL+qxMtsN+n6mCbH0ftH
2PMNGG+cEhIqzfcpYkqaBVaZZ9f5yAcO7kqFVcK2RgdKLylzOd+ulSB/+GRZlk9T
xCxbKil0Xxpf/5O5ZXtNuYiPSGsnIVLrYtorX5+eRgAwZc6NiWZHWa7/oRBRQbGs
`protect end_protected
