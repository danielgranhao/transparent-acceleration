-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
PHNBvtyxVEZuvIWLWjN8Q9jWTVuVVE5XoR/yDVXsvUwm24tR1ZPR1mfFg8A4rHXY
Kv+Ha008IXLcJ2j+R23I8+S1zWaC7RUmAeHqymYaFChUt2pL3mvsIlrQ4zgeOurN
IxnGnNyA2DDGkJRKRsB0CR1Qqy02bucTjt/IFFKcg9A=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5488)
`protect data_block
LUDScxWzgESWZPwMgqEO1xuC933NNSUKQY/Z++7alKf2bsSnHhfZEpuMfFzgd+vI
QB+G/kmhWcfJv2HKUdT6CtIS/lTg39Zv5Gtx+r+BBbWMTMUec8I/R7fg0aZ2ez//
2GFgEDE38jKdQGLZFOJBl3r2YnbYZZelHbkzGkyBB9Xa4+05iGMGcwGxbzQ1npeS
oVO56b5mrDNkQHPs2mojx/uIZodBler6qhuk39LegB24p3AAkhIBchX32L+9AHe1
cP/SeNnQD5O2UF9xPLGtCm8hvfsXQ/8pZaknwLlhL9jErpevFlnEbRPUOpYyFZ+u
zfsnOKD8/5x6xXqJvkiTSfaOAsxUr+G2wlrF2qMqDsz3faJs/wo4qaZYHrUEDoBv
BloQKEfrH8aF/ePgx26XcJA7o4bzIO7vObjoqVzh9hXeDxkykZ7DP9fj+Ib46lQD
sWbhvF7T+f87eHDP9Etm1Efb+R1toHXz6kJC8gp3HZNgMIO2RZQFKCeuFIBGdZ8X
/8CAAqYceednmDVhSJFt2cVz1Zc3aAYFS4WVRxoiLy0/sJ2M0TF3K1t2KfwAozzt
5/j48T6YJ2LjsuIbj3aoLwMmUoFwEQrMhAk1IFtchdkS8B6Eq2Kse8bgZb+QB1x9
r4ShHzGhJ2POGf8DKd3ieRAyVnhxRIFcSKbsUeQe4GcOrO8sO1FJjrev+KDzV96m
prdQAtCbiJsOuf/jARRv7kDj+4bm3X4kmVqeoefcf66afijiMR129wKKDmki3SyM
BbDsjZ60HrqtDf+06ozZH08OJBDiiimxYCPD0ceXPSV5D1oVzPBHGEJko1ZAW3TY
GsxXNaRdvLKsbjVZHGWViJlOAzQWs05gAgdveKen/AIFbQuYo3hsh4VhGjZbMlFC
LfvN6FWweFf7WEYP0JXK2Eh8a+V1IveIBV9MvylxrJbSL7NzV+dyBbfE3LLCQ+Iu
ROLqdhcI/jt6IWndhXoVOnhpBDBDvrSlIQn4izcWzMCxs8UdSWP8L4I2e9/9dHW7
kSVK7G1Z9GpqLQKAEDgSsyrp3B11SebZgaCv4MvlKx0G2RR+le3tFFrzZ8FfTppg
OV2FggLIf3xUo0VSscG6e5tJLlTfAU2j6mXU53pc7dmxWnU3aqW0TVlkbsHnZiUm
yZvT4ny/Zuvihi9iJJAf8ArB7X9OcmEXBrBd4q2t+ZUzZti8qp1lG1JH49f3q+5E
WOEeFLRc6hnnXWLDZD+xjcYrcoIxPcArJ3V5SmkclyUqH18GqXj7dYyhGX6A6aDI
Gfnr++Pv/emdSF22jppiLwKHksTbj2Roj9u799ItnvQrJLbLqtyIQvdYE6kCgXt+
tV0YYXoMq5Lto9U+YZhgKMyrOc9ib8z5XzM3Zwjj7UAfhlQljZgci37fcuRyNp9i
URAsuAutCBORVEoTHpgYFWrm+q43Le3OUwKyWDt45kh46vhWiWQ/Hy1hVrjDXzn6
grR4OQaISD6hpOp5jTAE9TXIJFXNGCRfFh7hI0aegzFY2XABayYmwpvv6Ex7/gTh
js1FWRa6oNO2Xgk0P78HT6a+QLr9Gb2ToODHdccFWfeYFKJqwb406fvYxX2mXRoR
RW/b5bF3xMW+PkGWow2hamAQ+X0J3dQV/U/IVVtKyU5FUVLnSvJYpCqESoD1r4cn
VfLMDwPe1iFxBXz9/Yhmxj4+eIyVwl84HeY5W5xAtA7c7HXOdki5DwBAqq9c8UE4
6BoTnX21F1KykNABokgkUuPU4dVON5kAiUHOsOUgy2iaDYVyqZWI2xshnlrA6d1n
gPIY/NgWvFtCd5BWfLZ+HlUtRTOBXASJYeOfEf1uB4Cg+ZbooXbZ8rvU7ftb1jGi
Z70Q30uo9fC1/kIR1FPKAGApI5oGkM+OA019rPVPcdIvoCeEQF1FQrlITDHsa1Ng
lS88GDK/T6jgdrcDeSz+UWx9tAkTkLAH2qPuGmuaBmTxKH8+cAV+dZa+5yTFx5aD
9Mu003ZJQQZUrtmHLWoS85zzLeWZZbPM0KFG2sQ0MunIkWHemsmEpB72r6bo+p6q
yuRYhgZ/jAFEA187b0lavFHz67YwC/pXBpAsHs6CbxWizx6R2DPneNj0atKiyqmF
7G5GRzKSLZhZBq2whVXqwmeXcPw2+kPkmEElvn5oy3wDCesjMOaNlB/WmMUIIR6D
ndP80p8LxO/pqY2oSvjJkIxl5FE25YePUofOv+TgPWR9r/VT3bf12jDF9XCWGA2o
mfYLUJUPWUtGUiyAv0qEf0HjLW8iItINSVlIDrNSGHYRnHxlTf0AOVr+rujC2QDN
QLQl/6PtLaaM8TorSV6RkSvohVCLBue/WLDzD2Hu6muk7qz2reCdmCmCHxTZ6ank
Ohczkjvh23UwudahePolThATxifj79PsRZU5s1RyHX8smtf48g4SYHfmqjgLLFMV
lI1N2LIS+gUsmzDZnOl4+afKJfSmgp6Dl+APhss/f0xRi6yh9ryYIew1V4CfS062
A7cmohr0U1F1skJ1E8BgqlzW29eLzt6+00EBmZCSuEEkXEf9U69IZT0kuJTGPuSy
MGZAhSjJRNG9t6yF1wFmXzRgkiSp76lDQ3iepQ0Y45+yVNjrDjzMUS7v4AE2nIKY
dE9bHCbgQnBjzSVSqIFHqwaUpiixtuzRfvFI9aVrjfOIb8I8V1CBdVDxIXd8a5DN
OYPnyNy7AoVCwsSIT1wrZcnUkgHJ9mc0N5JRMzHcBcwxrmuk7+6y7f89SgjpRsXb
83ZY3jNEDwWZ0iQSSZXAP4gtC61UZjkfoEBHwoJSsQWPT8xhL0TM+2LSRicy0RM6
4xnGBujFyjKuNDN0QJnhqiG2TakCxexCvDHxbN0reRSTHlaHJjKvqFGFvzXA9aGH
1Xa4Tv24U74Zy6/6qW2YAZqgxQBqo1G51aiiu6d5+Etd116rIihufsR5SCboAKdy
NvF0PrhDE4jYt67boaY9oYAM7BeFSvVyNC5p6g38Ytq8nhBH/FK5+68dy+aR0n0P
690x0TC31uFhRhS+vqfqv3WRBgMWZZkJ6Fruu7MN83rik7UK1mK2lLQbUns3gWJ5
0V83+pE9MQKTvxLw7+KHYq17NN/4h9gKo1VmW5g8pyU8Jow/dH5U5JQz/Dw6G8P+
sYzANo7akIRQ6eNqckLkmMkfjR8v7c+JkFaNPY8Rv2joxUKdmdAxykPTjgw1WVf+
JKyyzOxcD+3vUxwuExoGICQolEctuk9byH7R4FImw7T+cEvhtDnBZpmmBmV373qN
WD0AjvXLcqS3LvH8w16Ix6tdlouzMeviGTz4bZf4RadbpIyH0wcwD2Fym3Tkosek
ganqn860QLuqZuY5+T/8wbuu/t35vihuKQrn9iuJaxZ2+MTnpQRwf1jBAbZCWHpN
XXZEVzUZNbXzxhDtnYcHZMjbdw/zEUxyztD9riS9lcR+At130n391pWlV43GDC9G
9GZkPqx8W2oUQA/ZCFifcFeyR0mnydoiQAvpmtGyIzfDT38+yL9Hqv+GS5ksCGrf
iIJQLawJiRN5VFMwQ48KITMlcmbJxAHES+k3YItzF/0G1dR3YgczrVxkGKXGFh1y
blMgDBEbH0m6MGnaapIWvfpuMGAT7Unwgoj8WeuJqin+L4PB/6cdn6g+y3Q0gekH
CCacQeHSFmv5rGwgMb72R3O1Xtf9byFS6K2OrnZP0J0dokKYPW7D4og6IFk9AU99
A8vW3zTyIvtlwPg+tY/Ow4jhWRTdjwRNF2w+UZpsmTJbiJWE5Oaht9jMr04adt3t
ZetpE++jSo9z+rM6FOAtElPFJqDK04qaeo5k5ZQqODQejr6hyTt3nqVg2GUymJ6I
t7/uXyFSFUX5fU6RDP9DpoedIXnAmf2gbprLQzsuPzVwW21Z6ByNi0kMTV8eIqwn
Hmlo5xiLZNG3Bbavxn6T10cq6gYvYQPseez6OoyNQM/mxlmTFR3QhxMzbXYRf5cW
XQ0GbFOob9ize1cD7r3/SsKhdfHMkakqpbiKbo325dCVbd0oOOdeYZqpikTriZrd
tY6kBPXGKT2bD2ipzbXtKOTQwm24rHxsQugQwIUgzsG1RMEkJwilONQXfCrV3E1f
Zj+RZFF+GUxwevHL+/896t339H3aRJe3xCxT+7BZf2T8dE0ts3BmxylC7Ct33oQ2
WIo5f2yltY2mlxLmLCIhVEWNbpmCOIVhpRVaXfPssHj3rLopryMPE03NEvzaZQ9b
RcJSo+TEHEmwifKmf5deIyaFjIOf/D3LNuX9p6lLvn74SAhY1Vm/5GjatYWKPqeW
514jAe3aW0r19959Kbe+mHn4Jx36IkMQtqb7F0baNb8QIqZ+/KkNbU8PzMiUfuST
VWXJ+DCA6YW7i3tlu6aS7jnUSFnBVqGuFnw+5J52qOTsp4HzrQaOHvlRvTb3VAJP
COeEYThqBgLGnbcSBi0V+t8uQyKd8g0y5aRX6QDJETJ9qzqPT4Lpnyy1ABgPN+vc
DRdTVBNXFiw0wXaMJ0rMMr/G1de0eML0onuWCDy+rumVpGHlxw22QjQccFIBVV/J
BaQAqoGbVk9AlNbvDFMnevbPbNEq8Q6SB7bdJKqwIrYN4EKAkDuFuAQg7vvN1zye
A7h2WKddUZCzhEkTf83W+hVVGxjAb6tnDwFK1sIcfj4mhZvXFRP5Ov5Im/bMGN4W
Bq7VfZ2RoEhF9LdFyIrCyQMnAZDWV4/eQ2b5LGHrFcnydfCaz0CQPIHz8M8T4YxQ
/k2e8E4wdWSCme3+3a9QbQMSA7FrJQ92xFPa5fsUYLS03olTQSDIzFviJwcgLhOw
s1DAT9ydy8tGy63FbuHIATKB3QiZugnQV3lzTsrwG3rUNmYYcSOhTYuQBmb1o9DJ
jw1yMowUTXhIaoNcPIWEu2eGouOSNRqsx7jCgdglLGKJGh84WVlbc8vRtfi0OXIv
nR3EXQO5HZ9vZy9cM6oXl0G/OYy86E59Ad/0ePGi7JPzaSZozIT6mdfz+vOHtNe0
Qztj4sJMgc68M7ZOYsQ0Rf+htQ6DuB4lbkrah/UjwIGn9IuhqvH39XgI7qqgMy4F
L8yvLZEog39vuU0fvCWW+yOiiaTB1U7po1tHUPZUY+H9iPOC1/fOR7TkWZSRzMMz
ATacymVh45ZIUdCTVoof8xeB8MjiVWq7AMFfh8tYjEDGXg5OnboELbwewkrYTE2O
BMiwe8AUwccKWN6Ele3q3ujlrCvyeUvcTu0rmeAq6omDv6xlGIFPp2isJBh4Nx9g
nXveQGgGbpYE2drYkNQysm/cf1QLSD7SYN8Juq33PxFnFzJZhZf9ylvYg9n3k7Mw
90OSyt3qVVS35m1Oden7gAwlYmLelD1bsCBwn1zpXscUo99+mfthBMHmgd2VjdIn
tIe5LvMeaP06o4HgH75WnpjJUwuo+Mbac9hlUXIzo7FjwtMmi/OsxoCfLHqwvjz8
7HE10gnQu2y74NpYuCDeUmABlBfVzLyaiYHbYZJwgYXOPj8Saeh9HjZ0oqYxHpc9
1OQcANU2DKydR71O4K7+2ne9bqyw/DDxMIGVn0uX+04MCwKEjbVVvZJsH20eotDl
fBl0AtP6D9VmhM4KDNBifbs+eTlLc+M4QWl8d6M9zh7ckcO+42uVhApIjDPo/IVH
G8CEESmGPeSp3Rc2EYi7pykjNShQGPxuIzDfdt8OiB9ektc4QHWFKmHeUWgGKdoA
0l5RPlWwQ55tjK8NJP9Ru1RWFglWuQq0Cda6EzmxCHeMkOEZkZmaGbywCioPPaJD
enTzL7y5boz8r9WVfnxs0uAaxIQ5x4QyAYWoNmwyphR4s5B9DyoxMd0KYnJC/wyb
77JXLZpZvJvetQJHw0HBIhRZdmk6mOb3kQG/h4rzKfzanjXvQAF5T0d7WTXhcwP3
Xje5sfX7GIzZMU3FX/oibLQAT23RtcafGskXY0XRf8BJAOIh3+TXwS6p5DjRT40Y
KyUSeQ5oFK4jZN+AxrE5pawFbUu+lYlAuPaBaEd7vRAMp31mEb6lIxeiyM6/N7hg
KjoV71y/F8cgKRHi3Uo44nAVsKaC0lS1lvC+fm/wX0KF3a/KEUMOMIj5K5sHNVBG
eodwXbVCfjsW6t56QnEsSChXB6VImSaQJheTw9lwnMWRmiWfmgg0C2OhVlOLWTsy
Ij+6CrO9yMAcrzKhgrcQn+tjCpN/vb5GlMp4orQkD71q9GZKxGUeg9jbzXkUiRDt
GfzbyjpvflLEwbsRFeHUBQVJtBzP9cs2at9bHBuYv1ZJAsG41b/AtXNP6y909n0L
gq8qv4aZ+AvIkQ7FDPPO+Jrj/5lGPX1FqPJQ3abDgk61L4bzCl22ZeQLUU7IBmUN
DJi27tLgp9WDcnSbxum26W+sRrzANHo61Q+UQtt+V+cXjRf1HCAodP4fYFcV7Uf9
WQ0RgR1rS8RVIOkcJ7WoZeSS0+DoI2gHzqkx5r6ItKhIGyolr7QD0h4viO/ilHLr
Ue8qezCGqyhLAofF/wlDxPbrelfeZ2/4gmv819MLlD6lNJENkrXOsk7/Z2Le+OUe
mka0QBZb66RcurLGjfighyyK3RQi3HOvN5CKdtqDS1e6iH9jurdG5nKNOYN5mczg
lu33rU1Yq6RywOtawFS9Zq/66vJv14hfULQNCHkeOm6FAy8HDS1Rr9t17STF/kMQ
LlK4QSxArnIeURPvhBZ5l/j7pIVAx5yYpnI7tvudNxeMqSo3bBOxPa2A1Uy9hcFL
42btsJrfRZuAwxfGt5TC4EfmMM8Tr33iOkg4KoE7pApblEB6nEd/Wq0IIHwS8M5i
6T0oHYMOK6nwnBHrf2OO6MwaTc8129VAbCCk/1ji2Wm7xlVVTXhKzSvIOkXyGP4p
ivq/f+9HCFuNcME4Gbh2asS7UcifIpU3w5yhD2HyTVWELPrbTOxnSomR1MSoMBml
Ka5jWSp480SVkCIsrBUakGBcygIuQztcjugzgOaXl8tPhl82FlkNwiDJshC72Ni8
WtbW0n/dE45JfFUm0hYlHAM3ZXilxw8FWZEdhWVUa5jyresR7ujOqdWGXNkiLP4C
qFPOdaQpCn6m9xZct0+TOCxl8+tPTp8iPcn/rj+m/J2hpKEg6GPm5rwFIxzNqrNE
eWf35VhGaRiB4M4B7x7F2DEdfXegMJH/w3vL8EUE7p9zSTsNv2hIQtAElRZQiCIl
Ekdl1hQ0dUz5Hie5jeBxsfl20SKWXOvVg+gEZ464coBE+wi+Nj010N7/XBRRKuuk
aNFtQg/YDFuDGmZILtrTm/THHtUtyQ4yJEGoSKmn2ci1PfdhWh1dLQWHSl2upEbM
ax4d7gDGiabRKXN6Q+e0KQ==
`protect end_protected
