-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Lxfbmb63aU7oPeamflVNmbUY8+HEcAr37nzGYqYoapO+v6f1Zs4mISOocNn3elUg
jaV5hTzqEBRPh+Duk9RLb+lAsKj0RC2pLIP8qhaj3hZvZhIGiLWqvTofS2CPXa2q
RsK5BEMEAUWLXkpbA6rbX0T3gbnbgeLaGYM475Ma7qU=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 23328)
`protect data_block
6faYUF1RUhLwkm6cYW08JNbBDsIdke8cF3a1Ob6MbanhWIMGGeHqhluBhWxiPYtJ
NWzuRI3SP1vjRehsqL3fxglOv727nSzIbhKj35bPKg29PjExoZKgbTrFAiNTLYri
qP5I5Pt341x33UV8fwBWOdJHxyUZNRNNDlDMXaV3ol0zP3da4spTAGZuPY81HJs1
A6ahpIOIaJ1AJQoQh9dkw27yaia0B3IUFbgOG+AlXTuHBVjO1E2oL3RMEQWRYOEG
jfEE+1y7rhZM5qrqnIhjiGU/kcKHO8/7MsNF+PoIko1ZrvCQXzUmJerlEK9S3+Mp
J19C+8Hc8rEjSNxISbCzm/RGfO9Q4f5uM/ZUqlZKFQNQBB5sdn7nLtNZ8RrSd2ph
RPrdkngymW6KjEFRyHeNTuHZprqnYoIIKcT9zEltncr86o/hgJZLyKP5fk0xv+3B
o3QwRWTkG53EGxpaSbDIBSrn+eyEqjhB+kJ2XvKTH5sN0UasN/I1tIN4ZY1h+mGl
thSCIC+HD2418M8RRm0B3H0Eh140reAYkbmabFA+audpvXd1YhC5PD+Z+8IiYSs3
I23+gosOTZjSdnyjVYog3vEKUYxE+cIVBgZ0HO9MW6TTa/iuoUOB0ROH5GdDCnVD
3g+k8uPAPQzei3gjHkzLvciRmn9P/ndjJasmzbpBAvWPrpLzBoqBNEskSUv5cVtJ
ouRV34FULP1MGXQncvjDr88gepMZxaFkllTPPYizq0Um0mjDBR+j24CDSWe6RfhR
mbVXXKYQFGtpdxdbZPDm5CXogSPty6rmP4eHB4X+iiboGK1UuP3ePB0miH2g+w3m
NvHZbE2SYPH208HNJGB4ouzZ84qO0FV2rVKCwHnYFmhzxdZsmuwBDG8u88oAlgIV
0FkljJapO57RrfFCoVM4QQALYK4kolcc8bIJOmYFLqOdpVrU8IzFU/Mmr0CyMNiQ
nAL3ay3nw0MbtqJsJiQ3aMqHfJWRi0I6QddiWGhCg1oEvhXdJwJBGbsVO7hbUy08
LiHIwQukSF9rOicgu+RJo2LdOiH6tHa0VDf/jE4ZNKBgpqPxIWl3Lb3FwNFgZYBq
XF+DXCNKgVaIMc69CjQGa5THY5UePBjh9FhcneS8w8+V+PCChA/yPHy1H/jCePHz
gxPWp2YETh+Z7uwoWYd5g5UUFP5qtaFxBaqdVq7x8zG9WMeIW6An3PvwcfcU48Ti
DSJh7PdE+VTiSCt8W5HyHFCnTy2UMg1cxkf9Qyeb/tG8f9bB/p4wEH/aFaHIbdnp
4FEyKYIyYD7a6Az5G04mIYhbjgJp388ShzPHStEAdH8yTfgGwQDzdzt68YP/fKRN
5Pc/dFzbBbbXpEGLGzwXqsbeT8udKFQoNDS22Laf8FIUlnVv8M7CqJ0eUVKM/9yf
D/c05TROHCY1+8FyQoKgvoMaofzydhdgJqUHdOBhkzjgsbN07bl9/PHTio0goFFx
J8Rc2/0LK6I/97nxeNcQd9pZslk2rMAiPwb0OiZqiAi3GTPA4JcJNCs67zmGdaFK
dXSJXudQLuDtdBfUuzdIbLl4aYEWwctcmuLLSIeN58cDGkpJYkNKNnQuUv/MoDgX
wj8hqBy6rULUjgLvXD4CGXkLAskcuigQ1YhCfOPhhh1hiXsWfEnAjq8iO5lGm/p6
f9ojh0FIJEy+m4vXBPozZUOjlNOCNThVds5AMhk99FpV/xZ5mYFGj2a1wnCVVG7R
orDKhAkWinHtFtUwmeN8wCWj7ASPm59S9VofYNYDyhfDqHfcW1acypkFoNOCwmN6
LVXJzBnPvJfnza0IR9UNExN/ClFMLH5CkyHzKO7vrmbkwC46HnSeqW4W8APLxSl+
wXXtcQNtFt6BYqqbX7dTQ0wzcQsML/FVL7Y2cjoimUdOEvKGwjzFaf0XpQ/6lFbW
JS8JAnOnFQTQ7fnjkwtmNJx52s2GzRBAFWe7XfSISxVR73V3vto7qO6dKoSpm109
+w7/Umwy4w/TcEhoW1s0QzILR/x8QAuI5idNi6GupigR6/BNNKHvzUe0svWlv3d7
3GRLodLff3QwANZQbYxgPnPaqJSJ0rfEOTt5XxutZZX4V0E95Lk2kipwRnhLWncp
Ii/736PhpSMFfLQ2aYOJKMKHcaF/y+nIxspVFeIQWJM5XYP5U0FNw9zfbNfGyptN
tInnloBxtSMdsjBFTjH9PS7XZ9SNUHzeaWoSaKg+tfASLUiFav3f/Oycn5/enZzi
JtlIdS/7vv+pMTQ5aNMpY4j6Vm1YB+ku0ZQHzAzUteqw6OSkniEzwrdfyvpJByjd
u5WUppoUvst3+pcsUkmp0xjWn3qIq2gPYYhJsFXiJpso7u/AxTqxTF0fO6Wj31kS
t5io+8JUlynlIXZN1m9fl6UviNBJ7NEdrGrHNndJbIPOfka1OajTb14yK31VEEq+
YdOwsd/RaYZSUG8z7Ka6w3iYVdpJi66yz+waaSWWIYik049C+J5kB00a9w4alRCL
U//RHCRvJsh+/f6q1oSZgrXaFktSDDiERzUDBH2Br6K8xqKR6GGidgctAsKIMJ+Z
pRlli3zIan6lWjxSpTCJgwOtRjXzWastMfNSH9BTPORTHEvtvXnprEzSGQJQJkcQ
FySfz6ktXua/gxDSGVbvdt6NFZw42y+jrS+TSDoIodIbVFUfDdiUM9oEcOerKRtq
tM0rfy7znzxpvGJ6io7oDI4UYWJj65GHAhRVu+j+1lUPewm4G0Iqb/Y4L53s3yZw
EFzXoEMD7NDsnGXW1EoAq6rHRlZILetM4bH1FM4ZDlGaN27dKZAs7QZ8pDki2t1S
5FATRfZGZC0bPMG8Pzvuf5o2AkicGnjoq/aQGnMNv38N8FUyff8h3hnWet7Xfn5Z
bN+1DMT6KQ/JKAJULJS+B8H2LCtVccLdov8BoEAUhZ8tXAfCvhE5VW/UzIw5Lzib
U2xbwZLT6H7KW7qBrTuT353M7HvtEjqZoZe6T68MpKC1BWML2nxnU4wM2UJyaDxE
5sxQ56n/ArUY9YXMzJeo3FyV3Qn2UbbjuH3wuUI5fjQbQWche2munj6UTAOmbdnn
NyCEm+9sVaeMAXyrRivQVaYXSTT9PPefrLOdtsddxHFLWXF1f1ylXv6pubnThaVw
uKdYiNnJ59LAKAemEuRnQUpbgotbovT5UIEsqk+/POxu3eG9dIjUwoBE3ovAM8P1
e7e8CeBf7HUdZmOznyc0eMPPm1DCx58MaAXtq4S4xccmTEfe3Sn22o0iFQpE5zuq
XVt42a+pLxuKphrbNRvEsBiZnG6rYhAFAkGSKpCijw996ETFfyBr+gC+JlYMpIz/
zNA74if+pzgG4klOSK/LWq0ag8LNootB1ywXF0UOTGkY7FLjmZLHBvkUXMG0s4FE
fGncAkRBWfYddFeY1F+H+3NE8fWcX1xrvDCssSofgM3sxy9lCiMrS9fLiSj7YE6a
xeAVb4qkpYnV9cvww1sweSqzd350l9b9QqY/2PWoAa+ZkPWS334Y/k9rmSyal8LZ
2tMuIMyp6hd2mUF2DK7IqguxqHUZ8JmT1q2pgiu+A5XZ1HUU2KuYxiwBtMbDTHg0
+ya+Q4rK5T4U7Boe73yCgVKT2877Xu4s4fHkaCT3sLYCyXpqy/EAjopxLScxstlY
0HiNgu7ifCM+tgkBNbqbgPXtA70KEqeTjO2USA8G3xQ1CPVf9uv0YIvOigqjJvbE
GM2tQ2oHd2AetoqmIRWgHOMOQQETn8VNSscNLW7u+Un8AhQPzHs6nJ7AjDLpSrCM
YUbebQJcDUOq0K5wnykmmGTLF73g2C21p1P8pa5lKBkTHgNykKOXvoIa1GjoL6Gf
plZK+yhNezRuvOFeTBMCZ09f6nrX6/zZ1bk8dLNXqUKqeZjOdk8qKOfiSaW4Ky8u
pM2par/0cpFNryzbDS7XpjX/3HneoNhn87ub3ZWZo+GwQbpnT7VitQTUQ7j6cI3w
Bt617ukNUyz3DFqMmLkwIG+QTLRPdOKbv4xNa0LFQlg2o1blYlwCTkW51ek0BEXL
9QC/wiErdLfqSZRYqJrNty3xquhYcBmOzlLK680MUn49HD379JPt4O7j08Ge1UW0
fNoGoaU74HkLXNZfToKeT2jUsxXCOWrZMkf6pMJx5nhBD4GnWcBTiD0+wOkwN2Oi
RCCPb5I7lun/cuuymk6M2W35Dra+qjca5zrey/sT/psoKQbmS+eZcJlw4aVhM7ej
m3IasbFVVrOGm7Rg8USpGiUrRXxrcZ9hl/OVXsMVeIlOLLZM4UqJOl86YEETmvNL
JMrovubvKFiZnj9AKnYQBn6cGeECDNtO7mywJJ9Dc/T/Jh7wVProProo2B2ahG0q
kRsnvNI2iMJC+LTRpqEqb4StF+Joan/8o2HdejuEX3Ebdf/EDwe8NPnEdemDyr2E
ytMTkdrn/arAIXe/OmmIXYdnum8HvSnsi0ZnELxXh3mgM/VDk1Y2mnG2TyjpilAv
5JgSQjW/yyu620lNYbHImVw3R8QrfjWDvdNzzBQFf2KYGqL+owb2uD0S8vAzIZ3C
MX0D2+6Q6IB+DEQlNXx7c6ygWEXZPZikoYrucVfJzZsejAmpFaCxvqkNAu6XzU0h
2XjE78+bw7maa+C3FJjJ4Ndy0WszVV05P5MNQ9fTb0pMYt6AGYN97FqhuQvEXsc1
McIBX3oJ8hQrY8tJD8F0bRFIb5cZAza4yTz+fmcT5jnHv+U9nc9ShNnGId68xsBM
QdQ3Piw8IWyhOzPAHx0UHMu6GoPyqyKlmR9g0IPH0wur5Zt1+NVwUX8PqwbNUVxp
TDFX2trClWr0UvO10SdFKkYZ7HfgbKsBuZsjixSD88KCUvwXyaNzhFIMsrRe6dO+
eotE9J8kexmETmVp73KLlCl6G3r+xU2OYqeEgD3IeS0Fz+PWLq11q0L6NTYqq0Rh
xjhmYTXIm74xzurZqeznuttL1H7o0+ENmJs21Fz+r5C/0LOCM9cWM0JKKryotiHF
wLEN0ZDFEXVB3F6dDHcpg/sLndHxDqyqOPqIPPPPkCxYScIcebUwmT275XGMsEgD
WbLh32TQATKNwfSUkMT3JacPS5YRZ51ldOu9hm/lKBKnJmMG3yqTTEbcLKz0k/uB
BZL7+UGJa6CgC/MzddG8wptKYKlsabXLu1A3MoWRZ9RtPW1bcE+vekoAmly8Lrv/
X/mSjWrNo9ZCu8PA4Hw/fU4To8h8KX/U+70Z1pOxzy8mVyukRphA4hoNtTdnGruz
0Kv8/0XtNZPyIDmn6YT+3enuwa7HI7Pg6I4txJxNxdNDm9Q1S/SwitJ8fXAzqggy
dCmFzjCz1oGxTkwNBHJJsNDpOhhXJBPb1UB+nxiVYAkkaFr8oZQg9D6S/IM5ZCUZ
wVXFYnNaVtFBTlyLcj2eDT4geX3O8xOUSW3z+MZb69l5PWRZFhWEjoWGXmkqm89L
fPVFq2cG3yG3TpSZjUfGLnMBUkWVu6mCEsm40mMmi9d/7SGIuoCA6vTAqsqOS+K8
GVdd0I0pbasikPXee+Nl/d9QUHfTGptxrEujuLDJl94M6UbHQ+YTt+kfVCzPITdp
7zwfmlNeto+x1jIOrngL0JPqUqRPBgwcdN17vb4J4GtqwhoHkSPYEhAOucQ/fmAY
jjgkhQyl9mrojNrPfTTbSGBNjO1qtj/jkqW7u8zS9nvQCn0RBk0U8pR9qIsys0w1
fmppboZGpooMF+bKk9mkLefypSywmBD/HwLvgGPCHFLYd4Xzil5GfKO/BpYlx/2D
mSYJwWjAD28GkrzspHC5zZk1FNSG0mGxl9DL3JAA21Evd9YKl32VUYdQP+zjQkLK
dGg3p1vgSAjvllvBIhBI4xo8xty4pmCOPKgFs9q/oEyjtjZE6nxvybxOr52yzGnD
WmN7s+t72tmVy7Klesg0E9C+yPeGemoj0motSGsfVc7ER6KW+pdmU3LtCEZZlrzT
S5avXMyWQAmsno4Q785ZBc0RfXp9zd+d8Nf2Y16uC7lPUzAbTPoIbScGzfhWMU2H
u0rS24svsgBSh7MpS9A7IUm+F/0ykvrEV4UAuBkY/IJbvwQCED3zvOpkBjMO2Cyq
topDXfCDKbO8H/JYg844Kb8xMnCBymwMsrFYETUtNdmO55fOH2gXXuV/XtmhA0x/
yD8j/e07gge0Wo2FmL5iB1eQoeXlzk2WB878lHO4O31y+voVlhpfi97UUqpEyNYZ
3FbNhcD7/FbbgJMRLORRaSg71vmMGqXNc0We+GJcvb8AS0CzQ2DlFJFYWYJ2B7ii
dOKiL5lJ+MoOyCY8FARnzDck0zSAN39tSCrKrnPqBVhMo3RulmeqNUHOnKE8wi92
qfEkwSa/RkvJUaFonw5wP89Fq19yyPuqYWoByLDS5rIuwpQ6eIk7A6Z99gQxmBoY
dWmn2FKZSCqu8sY+XGF8NHBiNBytgVhEG7lcckkAfWta7dI+N/KR418+6M5x0KX/
8SkoZzy8rgiqJJ6JMItTwzgCu5UGtbHz3blQaXft/yYBCded/4Sq4OPSfd7rwHPP
/TQ+RQCBButfkTWgpxJKZ+i6M7ZkMyGqEMYMCLhHz73KgNoZNlwDH0ORnxK8L1Uw
qIs88ylIBRZcRNROJe/QpEDslsOoYdbuUd5HXgkWTzUhvS9Bjkv6Rrjw1ADYXgi7
26zTBdlAXpJt3z7K86BL85e1PQVsyIAE7RHuH4wK/mfHNB8W7D3jU493FYxW48f4
tpB2x+KuUJH+rY+fPk+m53ECzN2VGEegePpvnmNOY81X64tT9iYiwt6BdX8oRhvL
uiWYyAPJ5aOy8U4cov7J3V1zf+ucWlqgSmz8+VtJ5enmQDUH0IiEP3n2uuxglUtD
jF489MUE2si+Q3kRUReZRQKZJ+rNx7gWi4y7pOQN2ZUKh7puorGIH6Vcdfgyakic
/IMO5EmAECbx0Ke/ITRvrN2AlQHRcDLwcTFc77tumfAnrVti3eW8NWgFFUZhqAbM
so4ZkJFwoGjZsNqw8TLzs8AOYaBdXPYTBIUxkrWaj6uk92m9xvvNQIc4BjGWdmgZ
d4boXuKmcnJxnWgeFtBXKS4vY9bcB807pAMxdH2E687U1iL0rOciw+gMQLDgFisP
Gf0xbe1tvmbkkyRxc38rWXC/Vt1bUD6jBfpen2uP45RVaOwTw3eElNL9c9sU4Dtg
V0tPzPFzEu/3F1BgXbsiL+Z4qvT82g+PRcO9mx+4LvSGj0TrFUN1yGMJ2vbGz+S2
6Ja8faiT5YhZH+30cQ9Yd8Jm56I4Dez7CktexwoPLRGKVdXtvL6Rj0yM70jJfVWq
y0p5kDF0asaGF8Ob0g5X+hVasfxxwy6QujyJzTuUbs9zXXUw2LXPfyoaX1oTucvI
PAbrtUTEpuCD/t0CsZKtyBGKbrQZiiGewByWbNKHTscpGnb6f6T3orAaGj353S8U
HV6F8gx/gp6F+BzXngGG4MSpeevpME17uefamL1+MmRVHlnxWY0ZVl6w994Vyd8X
TMUzYrE7Q8xbXerKJxh8CFjWO0IiJ+vZuA19BJ12N9Kq+3VIhHJqaSCm72oypM1W
KcHV3zLY78GPCEMgVDNteAf+FXNgYrDcOCyBz/MZMYOYrr0WCVZJLhW5+WaSTrVJ
bweFbg0hbWgoR8l2Hscep+9gGoCWwHvJRk0gJaOKPMVm15+TtRyvlhQV8pzuCn7s
HAY/hIk76VCVXbYLjjd+cLUpkB4PWyBlfk4DfGK9GmuLtUHhH7gQio/B2V4r7LXA
/eUx6ArVCfDmbob05R8KLKV8knAtYfgEgF5rC06zvcbuRk7Kjy8Ei3HuAywFC3Y6
nosFJriEgPDTQMsfc2FyQLyR9btEIs5pO4riXdOTVdQIJxd2bEmt2zsSOlGvEK6a
B1WJ1fZJrFfb6oqn7vWDVce168I5eAnsO/iOMTPKCDZV6u5VDMH6oI4MHym2Tc9z
gv6jAKhoQuBQUiHmj6DMfUYotPb8Rkt2MiO/O5Za5GMgfVLVOH1A+GCVBbtQCfP/
sZeiKoFa77MSJpR0BozuIECTj7fxqDf0uyK1+gM/4Z5kE4zz70/Rp2VupQODeHVq
UG9GtH4+nQpHNfJjtnDSyuqXNeuGengboeF6AtNoAsTZcAP5wwuGj8gwkFF5hwsv
DXjcSxZBV2YAKe9rr7TTWWBdNIr/FbTI4WHUOYSGFwOSY1h81L5hzWNRymY9rYhV
GI1vCvL1kdbAvZH0kIMVW2gZupVps5GcsOlyLtnuLmRgw9wBPc2hds7+LFfmecIB
MKqBj70O3v5nIPG3Wro3MpwVZWxAqm+YaVSkPZNkI+Alc7LYOgAnEYjVbOchiyWI
xad+XRmFK1UqCcfUqGaQaQ+DfV7uh/P3PlRgQxtOVXvmdJTe0mCCd0DmkkVvnRjU
LzdAumwnoEU8Lo3vJry2o4tSSLPghLB+7nxi78TY648UL7nNl81CtRR14h7Z0182
huaPekbzEHhJUPPefFhTqu7nFOmScy8tuc/hFbogrSnkR6VvYuVKZBDWzxvqw2D8
Pl1e1mr0TVlj3aHT29r764hfGNaKKQ5an7vNjS90zgoIr/uRumY4AQQUvcLAPPWl
q8P244FQN/0615VgrFQFtNhhjj6GCL+F5MaXdn3nojGMeRGVKIhbn5S7rbMMFuhL
ET/O6s2qBa3pl4CRW+cf3C9cvqRCdGwibV0hbrtVRB4L0jsRgnszqrCUuqVgwxAe
gCr1ezRjcT/8PJPIlWfjacB2JxWlZ9BYe/56uInLJ7WiDH1nZy6VvqrGNadbcUqk
A231eZ55wegOKiAKZZ21G47NoGsG5LPFlwOQ41YTWDXLAHoJYD2GU2mELZcsiFwU
IHCZKxuC5XwKVaU95ipBqNDIgJfoHwc8j4P7FSe4B5+heBJCdvIla3ucNi8p5civ
V4KajwWRYjNLkNhGxcmJC89E9q6bqXMOgZQ3L5EJNizt4IsNHqDUrk05S4SPuMNZ
/UFsMtsjY6PG9mPx9kLFlsBQ67fTVojoPgVRcGTioCoJ9FihP+Nf17RoZGUso1Xv
qXoW3LUEyjFdTITEke9QbW4sJPYUQjBjrBetMVPFNAMX05BS4mUHRj3caeaZ6vNV
wVWSKqdoRU1lbAmJycTnXecxP2BM04jAcEmaUtOU7ISo+tCWMIyGuIRgo2Zblaqu
8e16nq3CxN7uUOxabkKYYieyshmf+wRPa3CPHWBZFhYb3mectagwMDDCJAl8fo1/
CKUYl0QL6IeGJYBTGxdTR2XbX7A5SIbe6lsJYkhonY3xyOu7U4OMtZsA8A2QMYjW
uRhsNrMlJQb1fpuRx3tE2cdN8yrJIqyHnUr3qKXDG2XQISVMVg2D2mJfz3glCOU4
l8E0kqLsy+wC+MvCrQSG7NXUh4r0p1c+ndLBLS+FOwMtpzNEBO2jg+EmQL4N4+UH
V+lfIzth8qxm37O7w/dn9AXDrF6fyav2VEZrwQr4WFY+uHzMKDGVwquXeTvYC/tH
ewiOXbafAbKuohZhC2TVDruDThmJe8ytadALGwS8bmwFV0g3/XhUirEnPCwJnE36
TJOthTVHWBaI75MM3ldeVEYAIRRciqfpgndTdT3EuuL/NrsxGf3CnGzRiKdo/HES
TehFQO5IjT8gQnB21bUVl9l618nwrrcRTKUPWEvz1VjWYKOs8pdSvPLH0qUmds6d
EEourxkCabvxyKBu5rkHXiuvgxcRtw3gz/uLQ/aW76jwERz8NjFw+6dvatoTFFLG
dmhwqqeIFCYUG2t/Ef1xTQOUf/CbAAkCKZSMF/y2OOZqegWLc8MjYasG//eBqK/D
db8vdH06yma+5jr/8KHSqzN+KTKPtP9gGd+oszIg7yn5WJMOX/mKtExiJY5zcWsH
N2RnBE/ssJXy1Rq0lnR62N8e+OYX/m0hIQK7Ab1BkWE+3UtBiSgjgJHbZ0Z1uhmY
/tbdBKUJDirlQQ87Mn5EjPsgaeh7W8jhz8hC6+ArBqaJ908I2Htywzuw3V/gz9QI
AV9rlwkLqQiMPPfc/HJNoDLDCSYacRdmYoXgPe6T9imGvePuoalgeDxrB/KSrKhI
nwfpVGiiUHQ5QzNHvRXEdPRCwN1a3F8cVj6qVxgz4UV/MYnZ8tikw3MOisvVxfv5
0gZsd1IuZyqBf/asi7LVRIknFrfrIMGouaw4rACZLjFnoRMvso39bKph8RCIazpv
zXRzsZ6aLWLBwC7uce1r5C3os2louFLdvcUk/soh+fLFZPZ1f8c3gdKj9MDEPI/0
0Yq/F5bvsQpJC7UozfzIeVCpOKglceYxLStEBt+/acAUTI7vWvS/Ei0wAzCXVTyW
ES5km4yj8zCRH7S6BBAGFIt54MNO7LFJ6SL8hjIeTV7JP5nN16JcJUztp6XA40xH
8Bz3Zji50r9A3xY++x5FLUn65crWwA59I2DPqM7bnzuOH6YkNCrhVEo48JnsWvVH
rFhTH+DagMNzHTs/mqDRI0wPHsX6DY6o93wkIc4cQAWhKtEKPrh7OU5HXKmpQ2Vp
5MIGvG5awlXfvG/vdEvevP6B7qG2k3UHws9vvpQT+Op9N0LeHSD+ySAWfqDeSg0v
6JTR4JgB2sVqBxEMSja9e0SNQkpzzBRlIPTQAE9zem+WqxwKxXXtOvDxP+JNUQYc
X0m68TLlg0d4ZnGxc875c+fJorkeDrDjUJJkh2CNwgI1+U8F0sswAzTOWf2YsQpo
AWvFOJHC/rusmZP7FlUoD/9K8tVZqy2lmU4skKY2k2OHEtny/bdeBxjA4EqiaTLn
2e0Sbk8nEYwKleONjUEy5PDGPAhDPX1JdF8G3TY4/qNUp3mbIDp2lxneD+MAw1UT
Giz0c0dHBBJQYLn9pknQWxRClSNZ8xZZs5AUz4o+Z4WKiqSpjgPH5+bvWf3DJKz3
w1wHzJmmjERCARAZP7SJZbp6bxvVvLAh87VTaKhH+TVLZ49h9GkupegXsOomeXXx
lxd3wyv5wDre3ZuvB9k8R1GZWcxhTvn3BMmF+DIJv72vwrezxdQ3pz7I0n4CFqTW
k9QygO3mVmeQ9EuYifnHzv5fqq1JpWW/TBOmMxNi8GYk+VHtmwibD3A7zPaMsJnH
LYRXv48YUyyf6fWQmtc6UqEjXq/7kJDhLVu4koZ1u3wlcipacBiSNFl43JrX7qKW
6QDaKyQbElMJbakAc0yLCv0lewf9RvT/qtruWVr7ggu/dFxOlgdiigq0/ro4yAIv
DaR85rbrykzd9oCbQ7MyFpLyXGB2lOPUz+edfqU3vGXf7johTSYUhZafCrkxa8Sq
zVMX//YJWL2d/R+raFGZbeBuZ14ZEoF9lf72CTVHweEeQRQe4ZsSIlUpUNehVb5G
hOFYU1gqCkCk6n45O0CtBlyhTT8W8V6RaZvXSxS3SOrCyJMCGDb8ehOa5k2WKh3b
Wjvet9b1mZhKOTKCkhRft6AZ+qvFfYFmMR767gQ8m2/Lccrj1SkdABGS2cTwfRez
FGRAQDr85Yd99Ywl6ccgkQzfUZqNJZyCuRWVeIcRpi0dtkv3gIvr1+DAMtXE66zO
DiVevxyBAUimw4X61VyZRy+Ry8w3xK2/FgPHtEfW5otoDQCVFWClGOrXSbrkZu4L
lN2QuBIlGrbTt2iyxeP5jR+VAhz3qbGhwR4CV6IqBpEckfPGoEC0KfNJOVSQdIRY
nyQR+KY5dyE0qy2JjkekpgUnaU5mdaaxJLeT272vOgS5kGgJT1cQhrExIMgclOfN
M6aqdn2jo7RSqx43NNgTp+jnp+RfRj9OTlPhK5GeRUqfrPlJK8vxWUCbgyxq6xQW
lAd322y/tomDfvp/vl7tLEC0ZVvZKf81NzuHD58Vvls12BtHn1qDAkBWOFeYFjJx
laG6lVwyNKppTKQAc7nRDmHP2jqDIkAbN/NNJEd5q6+gSDfEJCHbzlh9Dfihscd+
fu9NI9AWtdUlmukP3xhr5C6F777B13cMAeP32guNvpzS2RsUIHjiJcM5OiMrMWVi
DsyT56nrzO5vJ9DEM9EEUC9oHoVQ5/GuXbsTZ6hitQQzLgeYGPWviMIAV66EKVRp
wrzuKCGDYnfPyKAuSMSSQ+ghWujVVRyFfG3lANX808+u8kUxgVa5XiecVskWTkQA
bWBixmFm7XN48CdS1Xhr+tJOBH3CPS1MOKZ7Sb3YjNqPNWtAE0KBCqYKlxPLreXi
FMi2Mji5FAMRM4WzWNt8toep9A6XSQM8L+X/o2+x1prQA3GNbBh6W5h9XA7KwpTv
gu5Ta/8FvmyxNEeE/HTVQYcOXjlZ4MIiX68s8aIFyoKmjqKeOF+5bmLM4Lmxir2G
DBLGADZ57ZHRGKQtwx7CazibublrMdmjFoIhicYSgbLu5qhR7hbkF3ufXz3gjh2T
vULYmJIgzZKtjdg+3Mn60vaAQuYxGEjvgmWWkEZryDZoVoXLOCbyLG1KP9+fADPS
+ogaqlmrL4QW5qNOrdSPzvDF5hhpa1GaQC4mCtlQpNlzToCoIGk1JjuhM2WyeNUM
bWISnKxBQL9lIJYVQTdMqhsKSsarPa/Vr3fasBRT3rYs1bLVLcbO7Cb51sqvSnb1
sx+NMWM7rn3Ne3EuxE0NCJo4FatKe5txreVGdFuU1TUPcEOHXYyaY089iJf4jj8z
HW6B30HGgN5WJXI5CuFU/b8nLC4S3J+fOlAPk8/Q1AH4Xw2ZkgiGVu8rTG4zpjvF
+Y9S9sZdxZuhw/S+PHPJuZDIPh7PyymautssrUU26xpTX3CSF6w4Y31U+udJxNDR
nG3SAhHOySNh9j64Q+Bg3Ah697zxam5Y3Fcbs+pdxcZCh6dUVrGNXEuFwSD9NDXZ
H7venigsrgW0DoKdWHG+vCJUj8RmptsmdfiVvM200DMNAlz5WOa9K3/BBu3pbFGc
0bJMmCngHCIMh/tVXpbxjr4qqbOIwUEGs1sgQo+qkgWJg8uEbazuvm5ldyB1QFox
6cKy/g92px6tBrNrOPwSZYs3v4nxriqVGYhC/LOPQh6+b21OCc9oMOrVK79JSvB8
gpOX81x+5+ZHR/DC/vVRTZNYmFo6862SfaTVjvH0TEgrp2p7R4ikX+U0G8cHj178
sfLIHUiQpRljUV+gHacSkmKzTyEVeAbRRZINbVEJ03rFjbxNJAdhPzQj9OB2VbfC
qL0ZJqSboZjPVkln30RZLfIwfUUJL49DxhQRgtMRsBq31CmM5z4VIp0CrfYQaJEO
UxM3tQJga1TQr1UZn6XFCY/rkp5zB/elNq3hkQGxOqN3HPdfP1WfXdCDxfjlneQL
pzcKOS5WuaB4IJcAtQqXWQr4KD1ryX3cdmE35t2xtCCUHiXQkbFMXvsjZNnY7mD6
roLGNrj0FHZmff/W4eIJoNiz//XVW17H2c6BDuY6Fr57a3Ec/vjHncJr7txA58jF
aQgoB0mG8chpyMMAjKc7GJ1gFbR8cSZC6wyS5m75lSYrlRhyRejCqYRHKm9d4Cbo
S8CcbdkKkCIiHl8dVE1frKUDyX0/IgB5bgehVtOqWBw5CKlgla/4BgL2cjJJV5yt
LqWPtnQZRKS26SE1Kgf3MRY977mqKLFvsfiQ/V2e2J65RVDTzhBA3NlmjxiDZGOG
6+bMjahIJOPd90i32cXx5TlEyzwL5G1Xxo7toGn5XYal4V9sj215SspaOt2iidfT
HVE+6uqyeL2ApPAevk7x5jeSaxnsgstHk0L4ngWD+3IR4tt3L1NB44VKy6tEqtPw
tehKFZFDDY5+im/H9t1RCI80pEdUOGBktjKFN8pIEfg8NCT7QpnABovrkVAOl3vx
px7Fv3MHKPyNvPtVZ8v9t0d/PHez6f+J8CKvwrlktwh1VL0nK0Nw+X3XUKCldTfX
EyuxZ9rq3kvptohoQGmQHwbLj/uF6Qu7cYmTPaUbjNHOgLXsxKX5OX+ipZ6DCBmW
G+cf2qM3m2wax0XwzNfbJLeCqaIHOIsR8tDXEipc57Id96jGc52TahFRcEls4QuV
FVZuBpzZAf0gQOP1ohXswPm3cYvvL51ca2bkX1rCJdZXfiNBWE9XiBUgSmDgGd7F
GaSFSbanUAwP25Ujt5Hf+3W7cFwNPdXXliiH2v/kxPd7+S1140UDwXayBVoICO+S
tOtckSeGqei7bHEfW89tOWEkaRXXRu3zLzZJiaK2wiQGXRFLRObprl0ooNpu1uku
BQq1Xk5cAWRBjHVnVef1Otc8QYurWu5vsk1218GluPilNzvS+TAedAivILol2lil
FjpYVMRZzXM7wwjsULZkqMmPF+AD9nScee9xI5p/gQZh07nCdQn56xr8+VDJq/RU
oK1NnHJpOqOFkQITaiHaWIuQ5TtNLR4WO68+FiIh9xDCePJpE1I6Wa1rKNBsNAPa
Ka0ZT3jciJvTF3w7eRXrXFRQJ7MW8K/RI8j/jayUDmKtVk0VRTLPXimsa4yOQwg+
9MgQYuGoIrC8MqyVgzvlFrOqnE40EIsiwD4UA1Zn/Q5JNwCed9A3pM9JNcGui47y
oZW9voO0smZNE4vyfmd8plJZgNGlOGtTh34+ek53A1SbVNNuw51PMp28f9FRawz2
DN20EZemWGLtAlcrfWg0cE9nw2LXv+fZSvCzoH+J/ptcYHgxkD5scvL1U2AuSJ2z
xz5M1Mm5cB0LpaW0jHccNF/+LKRIyeuj98IyIlQwldbdHhQYJXcPInAfJQsWAj5i
wMB3eS/tXhj9WdrqKXuC2teoiBFhOKeHUdnyiO687FruB/Zvl/CJ87A3yg81P9n8
A6mLF/2oadm1q/xGv0Bd4N5zraabVT3COKwQetEzkiub5E38xt+D/AfQHQunO8ko
gJFTP9iuX81CSUwEbOP8yc9iK1U/v6GV73T+uUe4JeConFDzksYDH0uo74oKxDAJ
jM5+57Y1Kd1TuapNCzCp2zVThv18u4m7ICdWjXmJ6GowqDd4CmNozF09z6S0SiSH
FB8UBhSo3+EEHUkBpi1n2pVu+ELqIYrPXDZ2esa61ZnnfyHWYb7zPK2S1nkcmnZe
r9z0G2JR7pnH0iUd+Xs92FCm2fvMFmrBZZmSbwR5w6R+QZGvKtGMOWG5zkru3XDQ
xuByQCUFqeZsjSUzxafpR54QRTUK8p/9JCc2RkFhlkOTcGoi5p/caEdgTpxEKbXg
2ZZTGOun7O2ocpBQGFXtjkc8E2MRrFq8pgt7wallmluKVFWZn1RZVWirdKALqDVy
5TpDrVU/RTgsNscI2XStkTHidfDez9OB1EDCLPYeZdturJwBmF9lup+zOflVU//6
nteLBxNY4USu2yng40P8WBT47KYZTKho/GrlEVBONSltqVxRcpW8HdPUyL9WjK5a
6URMlr3jtNthlZEDspKgdQRusB1zhoUzGZYr/PgSvwlzxOgBFC9ckeG38GldD5rk
h57NIxSBGDgYniDuZsFcdJlapwnmFkO3tH5MwjUvtXtVHnBvyk+c4BmQ4+QS/YNy
aEnGD/1VV5AcHyYjcBcyp2DtL3JyzTNzIbXzCoPqxHZ/QAbj4SPTRHunTEg/NEar
T7WP1NMSCCw9+0EGA0YXqpWHpLJyOndWWoldC2kiDxvS8B2ZfK4SRT7B99xlxZqs
5Z/54DlsPDIjkkPLYcf2m4QN8J8M5D8sNpSl0vVUgHOEJC27R3IcPhNM4dJRkTSD
2TDRLhXZnDXbHm35zn8sCPicmfgF6RpXFK+qtORgmjJPQo/7ovHLZbhQr1w+OV4U
/jMPz4jaEii09JIqGhS7M+cMD7IBLv8fUtzRBvkuEp7yOgalOc6JYl+gn3wNacsO
4Q3XB4+x8x/CKOrVSVn5hOnRgW/K3DMqNDueELj1xDHPbormEder8MhNUPpVi4GF
IvoYW28fDkzW+jp9s41Nmo12MePHQRSJvAEedhDwp4Ipv5WqMO2HNo3uKm/0ugXP
/z6jUgovSgxmu8Jva/Sb4imjwR3amkdgSX+qEFC96XRfx2wR1t6zgTf6H4QsDyND
3iXTNCFlNBPE59dVKuw2wstRdBzJjZFhrgfwHB/yw4hTVT9wFyzlIvsxkCIH3Xi/
9bFxy3VVmihBA0ftcTOqQgExQzJJ+KMQmKAVuS8wtfJWpdVak576g89Dp5IEO0nU
8xRb6QISKtgxYGk2UAYQkHqR75XaLp+TlcC5m6tdUEOMTqKTeQugdIr0qnH6fJzh
fN3FGhMH4Ik9G8Qk1AfjNnO2R+dfoEJCiNWLOLzfeTs9QaZyKEVqnLyaTDq9krEa
NFa3KZS1lixYet+TMnPFaOEEdfCfOrApfMqsCcxbQgkTuubU1HSv0yV2tJ/RwzTR
vCN5dAB19nzOHjjJu1s4pgvsdxhbX6/Gpl8zAU+yozlw9fgiGr6JHmi3Z9e/jbo8
2WgMNU/XDu/1xyP/0LMtdQ3PVAMyDV2AXUI+a7ZAT18/see6vlh+kUGcOeTrxy1l
YjLAVFHG43fEmuQ5oLU7Wo3UXIFOzAqAdvFKzthjtU/gvqtfHQleDVkBCt77k2z2
pj3zOyPfn+Rg+y00wHJhvreVlbDSoOCkbkT19izoBDTImbkWbiq5dFAPfrykINXR
OrG859hrQcC70JpaAkKcuaWEoVeIrmta64jDuyyHTUx59HUeYXErJNMw0wkMwyOs
4HXs8wzyvTd5xaA9eny6t2at1K9Ebq/6Oft78sxxpoJ4laqLC5Cq1FUF1FHHhnLv
L+yl9f4X47/wwwp4Ch7lYcagKF7vE81jV7FUJYWpy7/Bm4yzEHNgm38wOxInjQUK
hAZ8rtn0X3fpS2PJcM2MFLG5enISpo3XEv2atSBXPjlnxYUSLUQJcFBCdiAWaz2s
+VP0tQ8xvEQdEWbu2hKn7K9Ly8I8+AFIRVLDyPv2/9IFrd5krKXtntZwardPzpGC
Xc0UIiMH6GaM0OZBOuuWZg2LR1WPonMp2CwzSuIgkTEY6O8sNiLd1v1jbS+QBwXJ
YTp9PAYw+Lo2TX9oaf5MWX0NnmnpXAwxJntDLU2ydE/lIPSDDbZFjPJrqLoRM1QF
0O5RxE8eCp5u0rj52UyR4J0MbgEGgd8OMFU32Ymbb23rsO4Sv1vPqsC/vx2xLwVd
Sq8NzAD7cYzOmvOg4yabp4t3MYqfkSi8xo6YeOOpeomqHHabsP1JqvcWjimq/JgR
VI0j4HkPnWUQ/eMhAI/OV7r4eot42k7afvmGy/6X+yUQtSprMS4xK5viJzZJmxoa
CkbGHdFmuNseqM7RUC6seyK+YnZZkx5V3axtK6fUj8BPWkH3xTJwE7LR7KYOaZKd
0nDBInbu/oiXECqYTLpstwFlIRgtE4TL5KmRTslcybIzj0DNORTKBNgkbeZ4SWUJ
b7vmiHQRmGpAi4qXfC735LQ9nh+bdpf8G3/6F01A35a4kD3OlAzTgfqfSr/GvyU4
fNDObeWR+fKtP0/QxdY19beBxWhZP+uNtCFxLlKIRo/rH5zLF1Kg+Elz+cAACO7m
d0oAtmw3Drv6knQ4Ymg0LLzNhLUJECBxSjx1bqdmfBVX5ew0tbaNdwdofvM3/DKD
nL83GxyIaPdE6Q9GPsywpPdc6sO1Z2I0YpZl9ImQOOqJ9RN/TQXjci4o4nvYqEqq
hdT4Ipr5EbEjIYzrWsVelT1xL1SDvHmLznNWnKk0EciAPsSpACm20D9gfddoK4I8
s0eT87EpML4TV0SfADt03+z190g8nKKEfSurHT6AEWYBU2CFfgvyvFo1c0WwUGTR
vsciWRGJ1nINfCpuULiLruGbTkuWZwxFCZPUfQFGO2qRD28BsUXUstA3C7aJWs1l
gtpGuub/eePxqsZW72du3v66FCS50WCMhXFTq4Julvl4JpCQ0OnqL6bte8lICSOZ
oVG0ornkTnGxYRmYVr8A+qRg9Mk91g62ONT8icGlJvJrVn2rHRtBSUlwEluZWaSW
mFSi6zTP1+shCtnQaiGRJIBzdM46xuQHh9c6I+2G7B3xfLMpuu7VrEeUhj9u16ro
MDidvwmmF08lzc9eBOe8kNHqupCxaUrpeD0sf7ZkxL+Rl6r3obhuMI4whb6vsZiZ
Smlrx2NE1oi32X01s/ePUISJclKYkwJHW4uJpvxrHi4mlldzPNQ3AxYnMP/QrjEX
jLT+zleg8INS/37lmSq3pMrvFK0/XNbTciOpMd6C6l5aN3SY7diFfHxSn3jqQk/q
mlbDAPS1g87qIpF3I7s5leANif329lcGcLbKmwqokiGqyIK9fXi/VyVWFoflSR4d
nOeI7eFNEv378BdziN/7obr/mGa/rnwvN08TSpzDfbNR47+NxPzwHepFaFY+H+KR
1RsyjZUEPGepWpt9VqwkYmV840nffxg0JcRkZkVRMkd0NOrOXUls4r44DFlKUYvW
+jCN34XF8uNb0+JfNvtjt/rABu8DZjlZ952Mpk2LasXThK7JeIk1CFmyraHOsk43
4f12y+g9KrPR54AzKNWLr/yMZjn1VpM5jPZQemvhMpe2CRukRwsYkf41N8jEtjIJ
G7HlvhT6AS1ec30DD+gypof7LqHqcFSHmEM3++2t5WWIYzKAJ4430XS4loNCg0K7
6fPjjzuDQhhdyydzMDLa0GC4aXau0WF+m6eFA/s4ymYjVb8aVJHXVcpIkaob9Fnk
GDyTuWe5cWMtHDFJb+OR05lFqb8eBFV+uk4cYt0y32+d+0WBwCjn4Fwc0cHDHNRq
VDDg0ahWzTN2CP0HwSZTrwUQlpcih7VDjr3rxSVKh6x/OVTSi8Zw8zY1sTEMEw+i
FmT5YtlcCGpT8sqgFND2V8G85w4OONq2lQFuKRT7TtRWluldKQrtuXtNwXa+ABPe
Gc/tySb22e7lzTOih1o26CK1s9VENcnBx1TihigQMqjXWBulTyBrpMACwEekbMam
R0KLTWJwZzeqtjw81AoPtbyvSmV8Cj55icez/l5nGrfdJroE2XLCXCEQ5uvbxlKa
0roTt8tUpE8b5uCbHvHpwG/g+9LzuO66VHrrwRn85eqdeOJq4FbSTL2G0+FAIABJ
FGrarTnZQLGtyWr3zVieLra5wbhG+e7bcRxbIxI6J5mp95JfyAEG9oRnycZJBNTO
RFub6yHatTgUjCgrIGkOwZ5/FOPZb1FmU5ORmbGb4n8VVzyxB/fZ9AxlgCZMkn9Y
4wWqWGmxDSnhAHThSqpD+TBxXn6cB7IoVpEFFrQvdn9bjgTfh+WJ4aXTjdyXEAx+
HsAO6ucS15Ow+MyE6iyiwxAG5Ds7TAbE6485a+fSm9ouKS+tmQ9f4P51rcE5Ta7i
ou1DZxhs/GWuM5CRvofYUm81x6Q8ET62OuQjygnLAfI17QCk2n9++bRj3emmSnpn
of84RIA9i1nDne+DjlmWDC1QXidZey7s/4RlJjO0Ij9ys0vnWltlEGMbDyk5NZQe
qk+l8ZsrcyZmC/3rcU68I9cdzwy3jd2QuIO4nYw6elhj53BYQuGs94RXEvFGP6aL
9ltkfT6KjKridleYheUcvVk+ZcAmsH5EhtO3/qP+JkzqFlsDj2lHO68/+EqVeOyh
mh6Jd9uV3iMAu5feSaLZL8No42h1OyZiZrMBtAJWDADTs4YCKjMDGy7kWzOK2cFB
xSD4XSCcfi0N/fUyx3upu7p/WrdmC0PL+Sh0uRcKY6uvn3Ow8dQUAcaGkp9KBrzH
qArTuuxhNC1G9U9qP+U6ZHQMKc4VPW7/HefBLYo4FtGjbc5xJYc6rkzcx4mw0vKR
QORMGEOl9QffFLEdDwk+wYt/DWwMvphLJ0RUPodPqD/YH+Le+yaRxKQS3KdzQYxG
BlsmHKealugdVrfwvIuTTSbbVW9+6ZgurSU2PHiKmRFRCHCyUqbFi1D7lQbcpaRp
ePu4Ii7XDbeFOxV4SXHm8vuemCqqxPrx9Pr6idpMOuqWQgYYwvC8PIYCQLZJIpCf
lKsm2E0QyX+YD8aYpKNRhpZdg1kFyDsfPdrE+bKXdmdwnIu1KGrIFRKVYHKlpgmw
RNt+7+pFmH+lHTL1uEJSZcWnZvkDUmQmBhp3Z0pcSS3g9lv4gNh9EDKsd+JEIQ1S
F+wl+CB8wuScR7eAPPEaVf3GiIanAIyxphBNLmncDwCRWpNhQy5wJkyvlP8jq4pX
JA5kjR4YEhjzHEAzTwZgj/sx6TBM5/C7k0V/mM6uXhi8IU0xpxsamvkh+uo/W7cn
0s04m9Mm4IEWkhg3yulgGTy8lUVmm0wchKT1rGO7I5HYDElAfGOZQd8bEaGuLTtF
AZeryukz7yZUZRmqTLEZum2zI9LR+oHHkMDq1jZTPq7vqljnsJ32bkYz2KUDPly1
znjRihoXv2/2ztwYzQn6fwffchUxw0BJRZZdxByvP3rNHmqMWqeQWsmkSWnBczCP
q+WrBergIq46JBpxUtq4XYO51ICBeSTE4AjaN6K+51/CVBAIeiRDO+/M/42n5uDc
Fi5RZL/0V0EWS26t1H7HuOtgqkgFPjtFOQAjz5KwHTiDqPpwAF1TLBW7mN3eq6ug
5Uqip81zr5C2eQxrrDCVeRwrbAX8CXORMTlaqpXLSyjbF1/10FuX4zoVcNIYia3X
EUZb08LUPGNW3KmQaIdoVVNrjslYIG25yxoOHiAj1Fuib9fVqMim+nMSd7Vjo7ZS
GyvT2hFY7fJnN5/ppffrmNBw5NZ3BikQq///GPddXxTkqhunPVGcYhWo9roAKpwB
fYb52pI6ZJEX24geAxC+W6+zO83iWrk8UnU7CKfQv0RGaSTKfhsGqJAj+/FQbmL7
kTAXspSc29bYh3GDwB9R/QmVhr5rByMXxsxJ7RHVqERJQCDIwUwgS1zdTWW199qb
2zeyWtevC5m6klg/zd260UKdJcLiJOOcMc8mj1eAZ8u5KwvvHf/i2QQybHQQu9cO
GjJxeXMHO7fRnODyIjlARhazQQZ9oL9bd7OGnTp3ODntG37naSjIbsxk0ChKy7Xa
qBPmIagiEhGoEfRtypPg7ynHbHW9vT1NCKXc3m942g4+hs3ywQ+pDZyUyKFvT+j1
W6v9FgNEafa9a+obsiBGk0pjlc/6RmIE6v+9dZ1v70KYG1xUkCm/S/JvqCfG0pC+
aabEx/DPavifBg83Y2gH/AZTbQwOBm8w6Ax0ir/aoMqV2lsGel0Nbajz1XASWjR2
yqeWQ40O+PoQP9+QgvNpujO6ydwKS3H2Qde+u0RW4i57oyJoeuGLKGlM+iKex4W1
p4GEOB1FukW+bhJ6O4CZI75KNGBl2GGGFLLS3jAx3bpA8/ORiQHOw1Z4Hapbcs9N
aa3yN7XUmNgxOURsHtm92FsbY4uIViOCnsm3GllBWqKjJkDO/v12cZsJDwUhVUQz
MZ/3AKhrI0jSosPfa8Drc6ZDB0B1qiH+EJBKjBRwJ0AiFJ/htF1AP0RNPQiVVdNo
lkjTCuXa0fcJyO/uiBQ9oBLG3HoOzT57mWstBKQdY94cs4z3GoYbz/hTk7TPQSeW
EuP6TJ77ZZyGNrBw8opIRd/L9OvMQMBwRODVXrizwxTvCWtt+24oINcgRV02DoYc
epYt1LhfnJjOwBFzZ6CcmB4XuyvBhIluoUCcSqzd4hlTLSxrIkhOkEOfm1StmEFv
j/0efj2eYx7ZBhTSYwAschXnV9mown3TGyb+KVUAJ3hXD5HUiS3qpJ6QFPsAiYmK
0Pl33sF9kzjurxxyPY4RBsb2jSkK12aixby/7PXEi53v8JC+VRFavLgPJZcLi4Lc
FZ7zIUWdtw7JFIAT8jpxf6RZiF2IkqBUCY9WUbxuWP6dG4aVf6bjIHJgqxop2zHz
gQQ5Y9/6eroHgD2gbMrJlIwzPE+lZsOMB7255W8rMhSfvVG99YE7DLH4kBMM7N8T
3N0cCaq+cc6AhJ8xBK6wvJqEBOZSif0/N/vFypD5EGd9j6FvjPxMlYZhBLsW1af4
WpBhQYJR7RKIC3cvoj3FOhENDm2k+NgN799Lq6nXOtHi3Kgt43mk2974D6B9vaAQ
tvtOWzcrGbE/dlDl3GLhr4Mtk3ePoYYCh2ekVVSbtfcYHAgDi/64CghEKFznmmIJ
sLLoo8iRRQFCcV6t3SXFBNX7hWCskBZnZVl5PwGgxcruugiB2NFKZz1jdsNnaCfn
1C4wRWTlvbzSVfHTM/jFxJkVUh1XCEmfHTRIMUbw4KvChxjQ6iqBZlNt22BLQy8r
hE1ObeuT6HHlCRCsneaOz9ANzA70pK3I1W1xSw0DBwaRyIqF7J891S2I8h9RLtyG
ZugOQB9uUMHHSHBtfur3tX2tc6DcWgvdpaSrX11QDjDyp0XyoTkJyaTXTlkwoU+L
jPc7T444x4pjR/HckcgICo6MphKxIq1zVxPVZlh5Q+6YjPanhJjrKIHyIZTyGErC
0WCIhBnB7gI2OGvNPDI952aTU9p5YPyDWSS6pvr9lSqoewf4gWxGKBYzLdfGNFgT
CTLbdlORub86HebOtlw+9dXm4r0W8wWX/0T/R7lhja05U3bxNaLerXieQ80zhfIW
XR46qD0pCbqgMeKEmY+q1UB3wAsPP9YjGr/iHKIPx2sdXrjqgqpjq9o88EYEX1p2
+Vvci30ahlWF+6sbL38uojcarUKKYYv72mIF5jyy6m4KiQF62ko8hpNfGIcya0NF
TSj3iNDWrBm7G9knAvjCESqcTtlfmUhlDY3fz3v852foLjKpClWV6dbXPLahdaiW
uM4Efu2Eh+9JAgqqHEWc46Sm6XBqLSTNYmLaTBKp+e+8/SyL8dZTJ9/U4+nMsRrT
Wpm5Zi60yZY4fFWzoHVgwHFQSBmWbDic9qJYuYQ4orQvhDyqX65yUqak4y62yGYS
+M7HGxsSQJ5CB59xwnliDnR7dOYMcLV+aVYyQzJEo04+bFpF+If0EwHyiNwci4NA
pvJ1/VqAG+1RvW8Hw7PpSHedT8vAULKQU1qBjXHsMllHczpIyH9weRoYRTEJKoh3
m+d5ehT6c0DMmNrZzEa6N6ziRtqzYZWo3qu7WtXboBiYw+UAg5Y0aK36Otsc6om2
uboqD6bAq+sWUUE3CEjZuzV5S0YWwleWnsZtUcm3FkdKeokE9aEf/l81hN3cTO7t
gELl0ifZQR+JEvaEmkxPPi8TetENrPSXXWW20RKh/Mo0s9qnKBUD51vWV9G0+Hf4
sKBYSX5knrwkddNIFOcu9E/SAlO1J++USrnoq2HXUaGjTE0oVe87llwo3P1Mwzh4
G959mTLo3YqXiv7T+jLZQa12CQ6lZAiQXnglotaclbZ0kIYt+U4UP5K5/izglVIq
LEWV8lZzU/0qR3thPJO4+rZ6fdYdhLNWMflHQwQlCyyhnD4+9elt+Lar88X/R8G8
r4H6Pam3SzPfjiP/gqZcVGUBNDETIwSRk87sEyAtjK9cy1lLbF4DXMIVu3TE18Lm
lamEz56Djrmj6MdxQbh3xuGMUDa6sDauVOGoLOFz58JO45XoFed4q97pMOSvYDW2
NcjCYsxiXR40EyEVc3SN0h/Oil8JqfBTzNq+isBKCuZR211K1CpuaapyXkIiuzia
AhGtYzLGaXpNqG2YcDdvPSee6SkPnWEFkSUqdadieKSyZVtJhcpSSrT3x0dBR1BA
N/oztOJ1GwvDUtW9vg3M62ckib5Gu17WYlYXHoiDw0zLogX6wxzWLx6v4d+UuPjO
9DB5SufvYdb7nF1EfhBpEhmVRU3fpt6YxmwaX7ALiSvZEWaCVV5EHNRnuno0jBmQ
MgviHQ5sYRGIBki4p/qhse+ls1Dg7pTA552DR9OWpCQR5wyTfIk/zCp/xwo8fYK8
omTVTGIhl0ck7I2TPTUPll7ThQuLEe09A5BhJGsoSCxEX7a9m6/Ceyw2PWg0R1CD
iGh/rgthYjR84qWVkwRHvGr72EUmlwPVZfOGRJ1xxTqQPdn40uwk2ol9E3O+zvDW
Sj4h9mMxxMjmD9XN4nOuLqAlBF11sebzpeoG4M8nrIeevPyWuI2zotvmZ0d9ZE/6
2xr//Ld83kC+re23tnroDHWBb11yrwp/8nQK78gDRgaK5OgJK6MBt5KEJuc82d9u
yxggr5PTyHVT2Gc/TpMKon5eyoXFj/MaBrFXVOJ/Xb2sWqDrHWEt+6O2dwLdZ7PQ
19jV2OZny3eiHjDDmFWsfLGYOhiMohy/5v+AAjOFm7g8HKRcr4qhcu/7g1y+uEMH
TWC3mtRH3sauFF2lgw4qrSpAeNGHD/dktzkPljFqxPpuGi+xFReedVaxFp9LFxEm
yUZ1zgTco2GLnxG0Uddu9sRVVgm0KfXFmaL8XOb+jiEVFt7MgSPLRg1Z8VWny/4t
PiKZdorvjwTHVYB5B0RCnRtd0CNK663BgliFHHTvNEKvWu5tydEkgiGxaqTja2dD
l838kZyte4rIVUNnuYnqzroReVlyMq/XVwNPz/xncvsJx70tB9pbd2U2/2fKzL7/
PjtA6v/RZhlhWuYkFX1NE3m0g9qf7w23U1NVY97lERgAjBBh0aYuR+j/ZgsaR6vP
9BiiyPv0/RSaXhmzzeU7j7GsfJuvS0rEstvHGq6ZiqrYD3O9iLkfmFm2Bqa2eqEw
iD9Qe3a7RZpIBHF1XD1PqwovsDr8S+HYsj3zXn7raVHKtkgreRbZG95ZSgNJKQET
I/TRPTFIlDfs8KtfOsGc0TZGmiRLBiW32u3djB8mHIo8733lu0QzT/7KSUsJpMJN
6XHcUULNyqlEJhKRrkuppQUIAQubh7ZMuuRZah4NJWV87EEpF6qxF73I4YOAM2BB
du7moFCqQVl87Imal7xJDrx2gPpd6sV7LIcKCX9ED9spCAVuWGyn9116Jc9OB8B8
ZlIdZHr95zGcMi2cBIee3kTKa7hLHV2/WSssnAd+XMDK+ljk+24mjiy3XKiKvSgn
4HO1JDJKOl5Erj9YWQHDZQC5Ye4DSUVJiJpkNGzXpA8vj+EWmYxJ4N3sPUSi0ML4
swYkN3Y7UbN8m1s0cYXoMCA7R8rJlN/M1/cx/jZS0vsWdBAfqD3DoUxVs6CVVkut
oOGXzTeeIN0mFXzWrCdv4Nta6d/iQrZxDK5qq+2L4EUd8b9iF5SYHIWFogtLtZ6T
n2nzApRXE/uF/xOnUlhCSaR717AKnh+lPzYfN1oziXuPefrzJbbvs7zqK4zZsVyl
E+QeG5LZhvz3Oq1096FbobUkyIJnaxfo8skvpOPf0gWs8g74GhcYtZoSoVGx9wXM
Du3sfFXfPBkW/sLF986UTsWaEYr0MUtnMgku1qWjuD1EVJf/PcfjpiduBrtQgpfn
iW3M/qAwKtvGrrQOLWI7BjpVjbDY25xv6nxQ8D3sJjET+LlyOwZJK0nl6af1MRAF
JmKK0F4zFUyVXEzMtuMtu5ZCXP5budjbYqv/eaurAGi9JMbN13Ua+6qnWNitB/Gr
ggG2/sln86cci9MFEkBlhTH7qGQDFGbYEjg9agnZkpqQPPp+fHH5mGGJ37x+nRc7
H0eV7+61qa/hSutsIEaLdOfFrKxbLtUliHOthk1K0Q1yTc5lN/NlhCeeAWVZ3ais
rcCkHZsNJDyKNSgKZYU2R2n7TlSlCxLcQOzSCQvsYVt7uZngwU2u5V5uNRytro8+
uGlFvMFcJlGR6X8ed9hxcLrRVCJ03lqrb0mHsWaVujwakopP9Bx9dIR58wliZnuE
6aZ9qTRH9zY8eRqeYrE5dK29FM5LNAbHqDgP2YuOk5vuS7JYwHb81CJQfQHiJEZN
REF1wikrGjH0dru+32AgVgU6o+k9bP5eACCdpPnw3fPu6dCH8EFdpWI08o6bGW8g
uvcI60PM99gp8mub3ZsIz3C5DfS4jm04e64xBBUOOzVZpZ0RNR2TKZ+EOSx5rTo6
uNcXuaOK21pIwSIQwwSzwjEJZRKT/ovWd7JjEOTno1u4azvt+K/WWV0TN4CvmnQK
1Fr8J6c7qLwdCeN6JPaJksHC5GiVWqAhukLtN9SDLhOj8RZCeuRXcdnm3IPX7hu6
JdkQORZ6Bhx9ZwlDXnJ1iW2MY1hwyab+vWrEwe8znxd6CFw7ifdU4pY6wL4O+bEE
CYN6Q8GBAE8g0sDqUAazXB5Fhngy+liqBPlrDTAwrsJnLxOzrWghdnIHmOrW6f1J
JKWsQwqGp4mVk+Tf/alwwaOvG/2lxoHTQRmRy2oG9Dz3sARogzoPLtyus5CV/yrU
SCtUJ2+oywBnua08bT27ZSbezJehGO5BGRk4JUtTK1vPBjU8lN1Q+CQ5ptkI5VXZ
4PZhbYMYPIQg66v1DaosPsW0m5oCHUMdH6gebQ6vj1+poKd3pSRBa4+u3dBb/2YM
nMn8rjUHHukzzwZ/e4XugRKZXM15/oycsoB6/dPl1g5AlKQMwq+dSv1e+JI08td6
0lsd1EbMorm0DkzQF8scacyMhekonqtP8XhFDUYElx4z6q9vjFbOmjU+2TMeaxcP
+B/aWl7O5k8lkp7YKpR/KWzZnWNkOXrw6pN/7tgEqllShXgRsCZT6p24brBgWMMQ
8TsQP8KhfUPK2OEDnjz3H+b/xTvTrkxZQslNJTtrr6bq7xoZx9L/yt4iRAIqKuN+
w322TOei+CvqodjM7Rreq6R88NKvddkhUU1hmBeK/JHgehS6fP/4M2b9pSUozwLw
2EEubwEdPVBG1y+m3OJsnFHQKl4iuW6PrzDPKtVb4DqzE1PZml2sCCDwoaiwGReq
IshJVDBvfxO+Tn6NU+Sd5SBtmX3WPVFgFOKGAYvOyHt+FOLYLuxoTfEmFPkgXZSe
a3Z/IL6ayzCGNxjQUaNwmXjkB8dZnwhzCA0yEKeGyZBn/2SCqftrK2S7UrvAQ0LA
25rQgVOLjwNfC+Mdl2+uxDmIyiL2FmStNyGfU+CYVpIeawYsEPRT1FtrWDtyxTvV
XXfqXFiw9C2iIhsizacr3bpyRGYXwu3gOdJyvJPSGyf/6OXd5rEzlJi/4M9zjLGS
fZLpGy1xQYf9zWnEy2sIelfgPtDRNnslC8ZZVKji1S/AIpxS9OkA5IZPDuEaIui2
1+hVWlsC0H4tlfYV1giZXzHZwSnASlQVAauZgEhjAdohPFVxjsFAqusANKMSXLRz
QhkcooGh550iqC/xuf1ne+5UbVBnKd4TwSURlc3+XimnlSj92ZDKAkzHPtcgzjQ3
pNld3bN7dX9KuTboEImmP1yip1jNTnK4Rin9r8Sh31t77rSwYSh85jYaF6kPu0wX
kBLV+gkWFO95GsHPjCTUZ4fZZS5xyKGbXynf5UoqNfpwM2tyFehqKFTyYCePPafd
/qjVBWT+x8r7vumQnT6Qqu9Xzgtm2l5JJQ65cPjxocvfzT8rQlcsYiP0y+Tx73He
YAmPmS8g1ozmtOxpz14XcswI3D0di44cNueTIbXqtY/cMzCqSb72WxuPkTANIG2R
CjNRWB0Y/0jPAaUPHkk/CTyIhRC31nCxtwBs+ZF0WNqru+ZC1w0pX8xfaueJZSlV
yuQDkYaiK/8drWH7xyTcZyPBxE3bcK0CLakkthyAa+rzxJU7ESuyo6mjf+H8WBwm
Nqf4Npcnw3Kerb5PAwx9nn/CV0KpUcq81CiPHbPR+06t92xN8f9EqQxmyA1sxYqT
TnffYZNuRbkrcJ0qxAacLsZCC6Zbr48OCTmCT9fMqUmCvY88KTaZ2HVbivluUNBb
bjE87QeblwVGmx928qXr9wfSukaDKbWNmNrdKswo9LJ0EpKANUGR1gOvr4corVsZ
7YBXl43M8ghaHh+YoiEC4TndWG9eahaO90mp7vr5HpJEpxbo0TQJe0BkmUjTVwwb
8XzMY6WJYZuPGqQM8JhC05Lt0h2fNka3oFQhtedEVEze42/8Uz68fIdP25Lgf20N
neNVaQx5CqyctXpis4ELTliWBEE1DLGEzFDybIomSEeIj/e9DappzIyQWNPKfaMO
BkNIw7kTchvBKI5pn/IaMjGG1AVP81NWJxJi3Icp+RQQYz/I8eDVLFJej3jLBB2M
HIlNyiu+bCfZYajUqe4OvxDxr2Sqa9iNds7o5vrghp3YA9VVDDu2xui3cuqZs7ix
Hjb8FBzjBMEiLUIr1l5sL1c5jgppoGeH9pMC06BI9rHd1wsokbjARerq1x7e9xSn
K/cSqT4Er2o3ZYy6ZnCwx01QfpPm2M0OQE58E2izEoS8Acq1e+54MPUEZPbWX10L
TWF0Mo44J5Fz1cDVqfHKI78qqyMvq/k76urkglyjYi4i/krsc7/pM2yaOo6DHe/b
PyCt89q72t59FOM62bbO6TU2zFj8YHsLHpwr4sKU85nKsJO4rgUxESkzRyoAbUQr
xlfJHI+j0tjRE+7cCDloDA1ZbZboVvJaPDNBCY6TDeKBdPpLVvIwNA1KFWmd6fOs
2Pgiifd9mX0KFkmC8yqsY627/f7mQxCGCf+NfPQSnLWDOszZeQ0lHPKlOXh0Dc6k
2i8LRo2ckXk/3RYNqqY09Hdk4GjsOpUwkU8fhpsNZZrsW76WyKJCwidCqmGqOCWj
pzbjaJuxQFC2kRyrMhLuvGwpFbL8cbkqEwm4SsCupI3IlvPBynoMP+wAhMuLJs7B
GCQ8SxGW5esuGGDZLPVdfC7FIni6sYw2lndPaiEDv2+2oWxAkwd6FIot5Uj7A6vs
nQAmr6IUO7JCpZO0BGdgKMY5eHFBRWYsOPSxEmdVUnIE/8Bid/Y9E/8n7wNd3T7N
2epH/tyuL6UFTZS9rrI89gTB8mFcOXJz97mhRMBbEenEvfokUy9mqqeWYeLYyZ+F
mNbKPPO2aIxM+KkjUwBvXUEbirbwTCGeN96PmSIU+KU2iblUU/CtSfIzpFax1gpu
rD5BJfdlwfZfiVSPa+Q+YhQJdSBNhJrXzOsf0TM5sUR6pSdpsPCGkcCcgw66/pGP
Xml45UhO4Snw0PJ2rSMXQFttkkeUfz8RLupfv7EPzRr3r6HEFDOFp36UHlZ3aIsV
MWoXSy3214a0aRt0PZ7akHP3rLxkqtS8Lxht0B5PB/1YVT5KBsbSOrZBiVeVB5Gh
UnRSqQwiZXsGRwPUXK3OOUIOh7OLtG8xbZ23GOzP1/Fs6HjCbNoEtVAw82CtWF3N
JYWSHChzq9+K2n3gY188lOEhg2ujRizygNIs+IugxG/Xua0Af1fBd0zSyuXK5n2U
d0Jg/3m3pISMAP3rANCj4t1GJ8ki5YO2KWD/p+W6n+UptQNIUqmmEDfp//QPBTRK
zw8o+mqRu7FuDQetwkNSIgFq263L5sOMyrv9Tobshd/7aA95bBMe5F7qB9ya4XBu
3i+gIusYx6ITuviNUBZr2CsPYI7HlGy52y4EnhP2q6O4erasH7DF1CttmPF9Y9uz
ddI1fSvhRFyLD6BKOB0vfBGGtn4JwkBCv36i71Na+R1tzkMF9NgItgC7KkG+LXp2
n0k08HcrSuIO8Vrh8gDmJ5CE0Ogyafd9Vk0RZhT37szOlI0Zoi++WQ8+ctxQmyh+
juM6pUEgNSNxDGFYp7EsbDyBL+Tq2kK8eshBVWarXbRdjyCasUs1x/V+ZwDA0FdM
bXGnFWuhtSFSUbMbLC1e0UZNorPRwBq6+MW4k99SU8VvNhqEYvtQKtXrVLaQoR2f
4qcALHuMcNZYI+DWbeCVzcIQb/xxtEm2cFZJiV51J5CZFLZ+0GPneOAa0iVpZohv
8GoSHEmK2x1CMUiNMnZVHsxcOz5+W0JjYoe5Qs9DuwU72twNttzhup16Hf2/elTN
LYQVYjg1/WHe435OJGqypnU98BaIYET3xSNe4I6odKCMLIh8mgoB0/EsT+IJ77YS
Cv8bKUyfIo5TtxOECcuULxNJlthNKkQ83tPEHW/L/vUZKb7kJsE7mpu9N5c+JlaY
UoZ4+N+igtAPUMNXX33m8ijTKO18Ax4H/otn465iQhsu1AFPnHTGsFRTNO9l8v1F
yf8S6mtanOgh+x8ZFZJO85T8cHi4V1yXwk3uv8HEKbVHMX+gYI/N7WFFU+XY5ScW
ZPHnWGsSaDPG3fhr2gtohQmEtEU1oPbJSbNPv+0RHtVjOJ2iL/hnbOhFOvMpFpBD
ZaM+v4dL2z3Q4O60uvZfr/bW0Kv986meTUAAcqWZ3nhbj2p5Z1yd1BZuB/vhQlQX
XZpXf5NoHSAZJYIlKOBj1l8Xl0RwAlUDSrixrYkPg1YsEzKMvDADmzaJya71w2SA
09n7CluTWEM+YSw+aVEbcW+R995F8KXk7a1W3vpkBvlLOfjY9CLS3ZzBuZ7Tx1ak
vVF3MgGQo0umNKU6RCYRecKKjJQeiLafW+pQ+con3dTHUiea+9gU0hCSFUCKs8a2
mxfwpH99Gaz+mt6RtfX4qE5W2z+87zkLg7wQncFDb6x7DWyNmfvezpI+xX2UIOX/
GC9x+TsKo/6vdIdy5z6wPIRRj0X+UnYgCBtFs56s/Le9yNQtxXC/ky2Rky4bLtfF
gorgAVICXZLCy/A5LOjcxzEf9WT9WwiTt2aeflLLI7i9YmayjsBLYz0re2/lf5oV
84/6ErXfSZvYPnXHhq99IP48r98eWZ4aqpgW9gqVhGZanPAozI3Hun3GdhA8x6uL
x1Qg3jWg8b11kky7ZL+vb37ipYsnADWsf4UDZCRV84ARu2wv02Hc3nxVXnvRP4Bk
99kA6deNaElf7ZYOzlCMoD1FIAnEgxzCSXUxGQyXM7gHjmqQmI8GZBKK4uZhjQc7
5Ir6iYtc/RhH5FoHosZ4WfJIMGN2jSQT6JRZF9/b6DKf6GjtjHu72jNxEvgydRIT
PswXe8DQGm/FPqNHTp+1MadQNZNsKfC8vwwZou5EXuPqyhZYakXc2605Dp6bjwuA
ysDaU6hz/iuoU4syfw7BcyGqqZLTjqAuBAvi5cgQ+5qsVPr9JWdHYOslR3/oR2pN
f3GX/Y7/NzTINjsQrFmQGZ+BBqgGF/vDkzVXSFqbfs+/TwLz9NRngQGY4ZwqXFkr
iQjmy9PzsFDUmy7UlA/AZ16tMXky3xbqMOxlBBul9EXb1MxzKIiz7Vf8ZEyiKLbF
+Wjz4aMWm4MhR8fonjYjfqQXOl8WhAeEpO50hRx/co8qfb2WPUvuQSjf5HKYUbY2
buoACHM5xM/hB/bXxv5n8s0TjViKHTeScYdJVeZPuZIXyKE9BkK35K6PXZmrBs7l
/v12ajUYCGnTujVf0c6vR+EExXngaRt7XVCpuahhsGcVFAKKCR1s8rGRMeIx72JU
liQzMIPl0HIhc3KS5U+RfrpUwpurMq4EWeeewahC6HTh76opYoOCcF48rXOvXHDk
`protect end_protected
