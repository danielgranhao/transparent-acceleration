-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
c9Tt5oTqpFmcAegSpFuOgvqg7dFpgcEkBxRMTBoBLDcXPM2jXV69hXD+xzxHyTWE
Sf7fKavblEuJXHOWTFwcWEgXf2xmaNnyT5wujZmxVF6dFOfGfVP1I6RJzC7F0F1p
pX7p1uLnZVwatLuKVv6PcuI1Pz4n8lZoRaLDiLczatw=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 24912)

`protect DATA_BLOCK
0ct+slUPxZ+6eUR3YRIC+8wihh/9jMiWw3Ci5qbwFnrhkROLnb/vgcRr8XPxjCyn
wfRGd152W6aYH64FPV1mzQ17ketCTMhXw6uP01mU/3Rthx5rugKs4dKM3xe2caTc
UJnW97+MvGmG8gbZbQIietSZ+WQ5nym7MIOaqW1xQLxIUVl956M85UGbJrnnWhzd
xCYCdBnDpiwOHfpCaOEQtXzUeeX2FtZKBLBSQYB28OeqAE+g5mR5eJQlzWR70fh2
fLXebTEWzKBxfahMVQIjDZ3cqgEhYOaiUu/w2gquLhnhGtkTkJzadfOQKzKN0JiA
Ua7xJO6X6d8NkyHdnBCOUdJC0mF7By9qyYOIF707ZglkjErqMEQw7yqd2z6WFM6y
M0aiMSsmfQSa+ZRq/iQk4mXiX4HeTAewOtHC0MM3LpZQL/ULYFvsmJYQjwVvar+4
EYTlZJekabNBfPwIlLyKNHzpsc+HrAPeb+OB8Mo/8qZo11kZvATJMsxN/7lSHT+X
4cZvM3YVoUbigwzOYWpnqbiYosMZQ9Xt8cMjR17Z9K+dvihL8rqM0SZn0ctwZ7uu
l5QZnge0IQ3Y1sdbvgJP2ONl5MnauV0lNeZNbFEco1EzfsMSzB4XoBZvKdiEYjtI
1Km7/hjAT+gFz91nfYy6d5NKct7GY2l8dG6FjRKWOchbi0v1cJUnchvuPpASwL//
A2zuw7LEPIYrJN77P2ieNfCJoOPxAy3FGYd98/dNd+/DbKeZJqV3hXidk/4NrXuT
/FujGolZl8jYBCyGXkYf/WpacN37hgUPUmRWTsoZ8cGog3ztlEE0Uu7iSLkYc10h
MjlDuu55lqFBIXsIZVRgCntkTqTvIeux0vb8zBzZouIxgLdUCz1C8yZRCpYNMdmr
ga9zJyx5LZM0gxsF/ARTh2gP2YWr6GyPeP9mSQa0BoLg3z5cAcKkUURKvVk7cGnp
+wyu2I7i8kowEpr2Vc9lt9BCf6Zv3RdWG1RzWzS25842PX6q8PlwxhLiCjDIn0J8
w4poiWBjgqCosHRuNqEC3/gwzl/g3OYUmFBF0Dg3HakloJgnYl+DgZYREb5hRyOb
mng6sAfGc4qqoSe+q1hClaSO8dzv2RprdJGmQ7+ffh9NAO265puL6ZpYa/BcCKmi
FS448xRfafyJQ+NHwduUQ40kJSUcxO2NUO7GLcId7Xdq2M2RBOt29BXmPpjZYl5z
0BtIy9+dpoKPXRxQM/3MSDYHsUh2G3ecb8JVwLK1FSvlfJZnH1xVinvEXdnjuW2n
EHFYDGgDlGN7gnLZnJYlmcPhCIsY8ki2vmP36MoNuu7+RsUnF7vBqvoZ4gNhiOYH
RecNMeNFdQgeulsvqCvAMDooV73Q2FVAZY6Xd191SqyMtLMcxkRXLJ2v/a6kaLTT
Qlx+zzCDBcS8iwC+qrBAHg5ioJOHqgVr2UJuqijyHh6A1s7WtA5Y+Ro2G8J+NnxY
Q1NDeaUQ8JhfbUkeIVQtNxOL7k12Sp5gdTTd71yFtTqH9nkzsi0sV0USBJpZO+Nk
yjOWPxyOI6ITCBU/uzxaGdKpRJK8LqbYJhqEjsXWy1K1+pbQ0SSm7w9KSDN7CgFT
zcLZhqCbx3XBHSw7NlIgV08kenL9dzMS4dAuBsdUG3BfsBjcLUBbxYBFc91M/Pqb
BZFGLgftYYy6ivenYpyi4RAXbZ1fOyPPUw+0H+MzrPn9ELcc7uAttaUe9/yogHw7
FcRtq1Imyd1a3mvhWQYZZkql0V2hozYzB0NaIs/zVfXxe1yu6KqGCbtOBfvrDqki
1Anx8oLbOVbqWarffxP2foRkO58J0UZJjd44jf/WxebEb1EAJGJ173JdPCtoXQLU
BD6lq5QUOlIrRhhpMLFXLMP/ZiECw7XVIEaXBY1CEL7MTyjb3jHO3y4aXdp6bWx+
Lq9I5RrYPPthD5RLz6nz6FJ2eq9x1xUCdAitEstRn8iycoGTr6LjRHLkr4kgEbxO
ID4Jfe4WSVB1/NjKknnY/fSMEKhXaOXF1bEys+afdCEqYcwzCQAJOSTBTiXOaOfz
Lq6EUmvdfFLLRTh0khLnbgQIFdE/MdwyiPduY9rBit6ev7RxtKoSLgk6wgDd4y1u
uQqXtVREXqWBLXDJMWv7QrAU4jD64ZHd6ePzXgw57p9KKcMNGUGxeY5YbPvvs4N5
4onA1TmzxLhxY8RtcHyPPHQcNTS3+NYD4PARoq9c0e7fO/UlUSlUEpF5hC4g8wm6
YTnPrs26FvEDtHtFn72KgxwL853pU1JLMhftNEhy7bkQ/8TdfOH4kvHDA3N59LiC
WfBiqD8ArIQFUALjif6Nq+BgEdABkKFsYIb0hySmyv/ZQnii+G9I63T4Cf8lxfaD
oPSSMWG9zy+YuRPZxs9OkbDcy0By8yWYaxevS6ib6eegciOzkIpX1RAbbmWYIbao
Ccv91O/yqMFYrBQka2zaTHh5ymirn9QnxwQj32u1CwL+7E222+0Hjv0qeuLJCeq9
jIHQPM4O7HYLciBK57+wiAnLkPCv1A5eMuy9jKpr8qXVmmQk5+K2eUyh/KD0dKHH
0KXFvQfFx+NYuuQzAWPvWKsK7G+hDKRx7ParwUgy+nw4cGEUDMKW1YkcdyRUcot8
3VjGOu/CQbupW6HZ6NAjUlBmDjUmMtGkMOErVEt6cI6OK0hE4O+yYfIPlGqrPpJ5
hB9AGo35STdb7IE9lVMkLTJXF/0swPcLC6zeJsaM9XODadIsyLdYuqLk8xk93WmW
eWRcTEDr56u8Yku3/hL2HzGMwD39ebTyFXUBR1dnYRNLDga7J6rae4jH/OeA6nin
5n+ViTeqdt/GYbuUIijOGdKJGyxeZ0B8u2rZkfb12oXWKFIqfxScws/goCAynot4
snQRKNkZUVhLbprMXsHfxu7iYmD+Z7uGZNm4NBPfp72jw7Eb6JTlIKBirW6v3alR
O1+cx7pAodwrVJ6aXv6h6WgOAeKOsyWItNoBcPo2xCiqMHzeHUH4Mck9ptI+Rh57
nyDzk82Ds/wyT8w0h+aXYEVQ9UO6sNdc8jMy1E7wp3rFQKehB+Yr/9BYG0ADj4fY
/D58nTEqsmEBFvt+x7PtX0SlKwMO2kk4PpZRuVlaADWzqZdovj9eJqAhrycg/hFV
x5JbRqD7PYbA22GGXr7jIj2UX4RckLCPb9QH+DVPxWlgiBABzNNUgxCWL9a0ziaQ
cgTmBXjCF4KwrfYlhsoEgaUjQnWbR6XQrVKedhz3wdcG7bHOSZbSopexboKpTvvR
9VHD2951YwpodKsdsxb+KgRQ4gSLazs3AA8Q/+FrsXBsSDsuklqn6mNADFGOBZH0
ksxcTv+/OH3iUQY4HtWufd1EweCRXYmnypniDK9ueyviHLCCe1D3zPus4ozTmshQ
Pk3p80b71COSqDE31mmeeqYGny2s8J6uaceVZYPpYE6WIBjD1RVn+p+hkm1YgSKV
Ahpg1IpeYjYjdBOAqaEmTlhdFhE31tgA9U9lUFr1ShnAVuvxCNpVKHwczwOOOJe4
BdH8PeMxTjCCrUZaozGmfipqMP5mDXvO4QDhSjENy1zjinEfrqRfEnwkAxNkSmHp
z5HBPQZHsWKXenMmCDRYH77vDiAKRvOTU+B2rh/rSDv/GANXyx58X9rRkOx41B2q
5jlADXBpKun76AM0DAAH3H73qdii/eh570FqofDV2BQsJqY6rZwmLH4b3Xdon0JM
oS93uGoLO9wF8uWsGfw1Jdy4g3/qyoQOM8IPiT1GvL8abMU7s0nLRTZNTS5oVbhY
6fR4kGaJYn4o0HXM+JRTPJlcPj5M1NjBMCDxBxVFUUeJRiX+20u/Nh/fMLw55Unh
sipb6yfIbYqhcuVm/3MVwXZkXpKmBXLjHquKALrbju4jQjALmapBQ349CypcEBnE
Rfwl7tQVsfupneNil8pz5kDLO8z40szfdgl+Q/775VPjpVkHG8siAAA7GLuxaFjy
j3Wkmb+LhqwDqSmtD5LP5p4t3LzxR3ZOGYIvYQUBk1c57hPmugPRa78gWDPbMUlW
7ws63qz7nK+tJ+362N2Fu8zuLydrYC7td9KIV9OhHwQldBNOeRZ0va2PQooz8I5U
09yP+RGorU2hmvmVrZjGKJgnwIzTvH+Hl2jWHTe7Qd6cckQ6A3rlmN04OVn9XM+R
YlVk2laUVP08FhEUMjEA9rm/TCnigqjsF8ankbjZts4TnAMGnEl/dKvJtC8fOzXw
d7CkY/sqFuGqYFnevVagwdfTptXdmLPTEhFkGzSPj/XKiTd9qaC9aphsS6uW6DE5
pacEUTQQOC6CbexSqNZeLjWz3NcrseXAz+iCwAMfV1r8J6bTUH2L17IarPY1W/ka
Dz2+hnUykb3tqfxP02aTiqffjPemKrIjxxymLzmGaeRa3uyP6iWB8yqO31116LL0
AzrBSOUVpNesq54SZEF2LuWZkLK7roYkini6xoBl5T09ltRflfm984mvha/c9Um3
M7eLLJAe3qToZtSYvZwlSsNFoBQZ9g9VW0Osu4jX5Wv2Kuftn8reSqQqhqEamw7W
e8oXFKL/La5olqCDIULYB733XAuGosrqWmyf4SzDVmSsTb3Wz9Osbb/j2CqVEGQ1
DtsLISUwVo+ALu0WhZ0lq0TyoHgCn3cYaWKgAruFLRnkOp+bbNNdtV4xt0wWMASX
X1aKOX7u/yM1d96ZJ/jIzebKpnASEdIqU9sfoNTH2JdwhAQq4B2nZu6s5svVQUGx
cC5PzbyoBOJSoN5vvzrI1uOhZ8T4kwWqpd/niICac7zbjMTEiIZsYID+ZrUHbcDf
GNScz3BneDaCLX0ST/IaKrdubnG2WNtJglLFaPkCg3Q/RSbhngdqfajtMPHLTFd7
V/ofMaUIhZ/5oTIAwPcg+QWmJaCf0UoRnxBYiDECur6tqdTAT3EQi16T924R4xDY
MPx8xjblpdlliTDaNcqbRq9OuyPdXYEYmVRDhZHSDThsPB67juhphFfMktBpu9uP
VSLlGHDJU6Jko+oyIl4p8vtOVXWVOX1zKww7XT+B2bhYgtzWCFvbZXSF/FDxS20S
B9Wn1RQ481zS7/d7/ejvosBZtogwbhWQ19bp/sKzPOr2XqSB6L+XBzXAa5H08zUh
8MfozAmUn5fa6kf7O4mEJKORjuaT9uIy9VWeuAPz/7QB8bcLQAjBTyXxPNpJgbmC
AYmoI4D6N0aqm0szyS+vnP53nHJAkpQyKHR5RO576dBzpVgHLZ9OP7G78Yg1Lj0M
PwiLvqi9Qk+5iLQ6/1YowfuysIE94JF12Fb2KKPs7O38uUBsoEx7PhOc9Q+9PpqX
3kNHUY+/kxVtpZYTrBIzmiB/YjDreqG1ntHnAYquzDijFvZCjYw4B7v7G1372T0R
m9E/5D21UytLPpF0EjYaVsZjk32M8J0bicpWgwdyCya+xr10L89AY0/M/lawiGK/
IDxnneJXe5ISiUM2E2EUQ4HvH+JaMm/uUB1wA2mMXLtItR0RdPOpiVcRWvWLfiPB
lLKt087OlgX4XlQWw8Cf87NKu/lR91SD8PW5DsrXuCn872FSsAglLzKB6DAVLLDD
AKdJ18soPGlQsQxa2iH+GofzRb5nOfnwggn1ENKCfI2AE9glqAyFcH8bUmzPNuIP
oThW3ag61swSbXLUvs/r931RU7TGU2trQj7Il8Kkcf5T2+Vzy8UhAlqRgbNSoPSH
eZdcu05xtx8wGBkT1Xo+fvj+XLTR0JySIk/yHyYHyBQvCYDwSIAKI65RJvXl2ohL
kPYbvkaOXspYbPrptzwu/5OiIydn8TJUeDnUI85kA6wR5mzKQxSHpxQCsJpqwf2u
61vvScyf0S3M07iiZ5y1k5FhtyyDFadZP4F521RJXso/5z7OMdSMtkWzvBe5Rtu3
f11Ge7DFMy0QuPR8c2+oNeS0xqngmn56GeRGDznqTk8r0opKlloxj3cps5LSSuPC
pHAi4x86o2X6HXjX7IkHRJ+Kib/tmlEMwnT9PMqlGTyOXAjqpn0PJGzW5rj+n6kA
OCk2w2+GqJkhL/ZKY//CykDiALyubNjMHwWXrLr9g7OhKWZPiineow+9gOGzqYo7
9FRm2VRVqLws7d0s5NMpqEzNbXEhcR2m55AqwsDeev5HrJkJRmaHH7n4kgmuoCjN
/r5z3z7a/0/rueRxoxSX2PNOCr/EEKSoRESSvbVqY1cNADmDrW0tzOPJfJ5djXHK
8ybLgi4689piFLdpRzqRXKeMGdVQvShSEDUdGuf898uT/ur16tGDZ8Lv/qhr381y
c/rniGiPEnr6sorlkeFQ7zF4+5PbvXsx3t+p5UKHDwI6V+R3qqVz3Ytvx+UHOthD
fWBpIJr13Pv+FbBwF/yqz7tcZbfT82ZKXEQwMP56AN7Zu5L4sKz57ziF4lRBczzC
Nc56/QeS6+mKGEi6iKnw9jvdNw0+RS2Q48IBqTFzoVoPgmQyMewWKsqUNZnrwV85
8/8gitEhgAAcSyXe8xteOILSv8gHn7fK3zT0B0pDZUXUCVum2xFhe0NOTYL4Zy8D
gRR5iS0QZ+8BMlG9mQqcIqL1XpTg9N0MAffcSEDBW5Ewu+R5WOZ85HKr5B2Zren5
8vclHxeLNPRyNArCsEx90d1yaHYUoad9v6oWbPoo0JtZhR42QV/UTMsbvuAHDiBO
fDbdc6YDzKFak7tMTB44PG6TRw6DSC1T7sKp8JvyE72PKuj9xYmrA4UUUJEroZiD
DjS1L/DdH7jC9s+vdgKP/Hy7E4EkEgcWe9haj1m6S6PWPqu/rzlCjHFzteVtvGj0
+fa3tn92VUlYcACgWYyOzGyMVeFyDaxdX7w7jRra2psOrVG170xsxhzJGUmo+phb
y22UFqnag4GoWgNkdIFTF7K5f+zAJ2gKMzmwrYdg2SeesK8XbZ5J/WBcGUy3QURR
JD6mlv7yBX9HHAVoxzB0lWckgN4dgrBMcoQf5KmcN/gRGBLe4zTHL8vwoRQcW/Rz
g4uM4Ku8q2/r9xVLL2aVDU9VGjGlmA0UGvp1E5jIyldhPy+RnRKphV+9RuRL5TlE
QRboDjs1mrCe/eaWP+/p+zvjWKJkW6BO+hZJy6T87bBc1tiME4yIK/JNfqykAT4I
iJFcNLOjNYu+pRc51hRUra3Eiety2jchXFy+ntZgDhgFSK97T3fdsA6bOeMcz63x
JKaKTynrVHL9WC/XWm4xK9dDR1wEtbOS4UrrdoDK2ir5DW1Lo4kciqhUsBAvk4G8
lNTd72iVg9yt+XZXOzD3HgtBIqdLRtBU2wqk5hEpbRw5kA1ADQB2mHpusbrjYdh1
TZn73RC1+rTQaTIr1rTnVdkko7iXOuOfOGxEUpWPmjptQ7GLUgecAhP/cgZkxogY
1Zsu8rsiIbyqeMgqWUsXN0/RFEDFaZGFll9Ho9aF32JsaUs/vXFcpjtpAUga7oWo
ikpCz6XKZLr72rtsbgIRnLMq10NEGfwROg44W/L0akM14J54RbffL1hY4YEh49Ax
4bxiLjFDbZOkcfbPbjQXnIOvEZRs8JfmdiVeJTf+ZeNYxO9Yz2A/hc0jP4Efb/wm
Y1nW248Y5IyQo4JBockL14a5P1BoRzfzeQlWWUcGoHK9OCXTQba9Q7zCHmo9lVM1
EytxtMerAd+hNZYfbiN4lZT/KA3PUEssBzytRymvgeyPy08ows33imjEOqNMaCTw
y9H9/XS3Vsl8zNqpjn4eeZy6WO/JZv7X/+aB+Jn3YwzHc1/MKphj0l19xSXgmVCS
kAgMEdgprF0wluS1ZYaLCm5mQyr0UxmS50SMD6D0+n6QUfuyQyXjvU3Kq3H/vxcd
jQ9scsB+PGYCJGwgTkG3H0+Iz09p6M85a28mjRwwxrU+I6Ck8DUjaWNCTG8nF4sx
+zQJExftQyvC6bCDIIZquH38s0nW5WPxkn6VO5fNQcV2qTWRM3kDP8HwTaFe5VQj
4fy09f+FdO/oz0UQgKhN977HnRRYuVIjoobkh3Tl9LuSMM0ern1QDtX9COIdrzz4
NPRaBsT2Uljmeds1ieRnKbmxB+XVy25WYmVza4hSqHAUsX8fuDEJhRYY60TPVILa
W9W+rnX0ex1qXqaqWWXqLGphO90o+Eq9ScIBmQwO68YL4IfcMVNPory189V9EJEg
XTjmWTPbGaACMG7UQxDm7YFNFcEhonMD3BI3DEX1Ti0PXs55MkbXHTcX9Fm++WV6
1KIUbdsbYA7pwO1iaKuBSGJdC/184f8A6kAxqY2gLCTevSRXzSnhVRCP33CZPfaD
6PMlHRo6U9W6dR0mltHMRitwl9AhYNDDeroDf7jMVT5DTNoXJ5nTRK1tnD39QPpN
LslRKXU8/YlEdwBweaiVLiyreCHnNQJnVJx0tEz3qfcAZfkD2Qs9O4tIIUk+IWOG
09nbC62WJeCRR0l1i9Ydz7B18PKGTSAoU2vbyM1hs2uGGFhCvLlEOu+Y2+uCFudl
/PHnOKPcJl/acVYlw3csc6jxFVaIq/2RA9y30ehF36YwBHk6lFHqWRY74tqSgBB4
S9sm7GEWpkN+oer/j+fepdcJDUL1NWhKZse/oz49d3rqkdYu8FMGf5L3qoSToL/9
6wBSE3koCKHK/290MmUwM1Xqi3UpX0WOiHCeurscTvnGOUhopTamMcGWPgfkQLO/
OAJ1QSdpLIoXCw04pxbh4thg7T5RWOK+MyGcNKngxNY3AvJ/AIKcpCBLUqlb31Qz
XUzFK49wLUMv15K3ihRGxZVPRAriiJ3cl7XKlhfje/w6qJ8WLWUTFskp7koeyC9V
G9Qn7lDE3eBVe+kTxfdXVKQDoN5llN46y4W3Gj3pnRuFfqZwe3LIZP542Vjh+A0O
xL9l+JJuY+aPV2xhUHmhZPOyZCx6Ee3W0NQu6zGMwa7KW6jn4s1+nxR6Wg+MxACS
m737nRPOF7rI8aFW1DGMH99YTXnzPwOJSyLqr/RNv13+jrBUuKZcSYca+Tz0NuXt
c4R+cENJbmYFWUgdJ60Pt6jqBKFR5paAWoekujW+ZsQITn99FJOXV7YrxnpoCKpp
6OcT88B52ykQDp8Pr/RlOlQlBDdxfdhNco4Ihe5MZ4Gf80oTndrby5gVnPBeQdQj
DVnOOLo/MYQRBnw3HLTaACcbCgKA5PEzkqjHm2M9rfsL+10wqtJ9cD+E9ofHl64f
F7uEqQuABy99kVcm2gz1gvMDzVnKnLIdZLHOS8312rB9Zcbag8MvGcsMcCq0T5vy
MByb93XO+UHAzdO1eQUBYx62jEea0q6sQ0XnR7YDsJfIBHLuhcB9sjfngjXea2cz
mtkP1P1ADztpHIQ2XeUL50A4+j0endZbpNr9oNGWLQFj8+dbYkXGN+PNu+h84CL3
QhzeVDS8+dUR94MHjsP0wT4lq+jll2YOF+mU4WZji8dw2I0zuHSQQWtjObiceCiq
1Vi0fq5O7B21w3wnmPARoImrxPvGeoB92SAq5vsDO+CxR/1Iz01QEVmZ8HXZBAkQ
U6AvDKsSgqef2BKY6xgIxhEh2ZCrvkkBp2hKdKgQq4DNkYtxX+bneG/7yDnzYd2Q
ffCNNT7DaKVN7av3pc1Mx0RE5D8x6vRjS4jYijVRv6nXnJM4Gx7Z4mKQZYELfsOA
OEgEZsibmwFV6gISw4PACuu+duhODJXRfMrV9GEC7V95jZg8LVnMAz7NI7i/g4sV
t7fuzDR6q4G4fSwKbi3E+cTfkCGAKkU0x9TsJeCm7Zdi5TKrZujNcbjc59ewzkEF
VvqR1af5KW8E0DmOP58fC9lDS+KTir1NpFKkWIdpjuF1D9kzb6RcvzWSqayQckNF
LzTUCz8eer7AXjtlzBQODBuW9czTIDMRk932MJrfLUQlb2CKT3e4YzFGT7lrAEVE
bRN0kDO+0Vixxa00LNavsbcMCLKqEKbFLTVVZ6SpBnswud35RfTXti5dvfRNaJL0
TL2RX9PMeN4bqi9h3XiYWDd0BpwJKjMAeZdsRFd+mfzFHGBACXQAnJUmOTUZO5wt
SNmCQje3WRxjsahk/lPIUO+Qzek9Oz/d8bHwWv2Fw8yJIRwF4lnm+gvuMEmSAPZ/
NbPiJ0v5n1PI993g9B2yJy5TvK86ZoXn9hwMi0XX0B4tRcBcc7GOrYYyohNShPVG
nw55WhO5dKvlelmXcDqcqKrV6zI3ziIeHLN64earL2yZUqfGCiPWZJW9YWZCFJBN
H8o59QOgfdOD/h1YeJRwSftiNY+7ovXdlbS9dFjqiNT0RIADQ887jPQtTI3BCcAW
KWLIZuocNoW5iMPG94tnnRCK+Y/RJKpC1Ay065mtogLSb10TjvxY7BqKrE7q1LeC
bffXpEFA6KKnb9Kb9FMeiCOW581dwOgZueSw2PKbWpuw8JZj0lsS9cZo538Zrzgo
i4ls/CVQCRuCIaXECkzCnGSuyFzGDQ/BVXgrKNK1PYMbX1aSvVEfE5Zm6/ssDjyG
IKTMpiSR0ZIgNUAPZqUwJl8Ih1eDmju1A+sFBV8htczv5WUdFWMsm7YLWIZGJ8li
V/j/Hvk8PHZr57gn9yMbF/EfOQ1BT9PP4A55qamwyvecfXv2/wzSRIHZGRvD8CKA
oyWRuuQ4EYNsVY/PRPR40eK6GBo38C2CxMZkduqGlaG2jQp/c2oxo5b91McDtWkJ
vhFheWD7N1AU+5Pf064FASJtFRkk2vnf3Y07uNSj0/LsfDCtV/w6NEBsSuyHiiVh
BXW58WZiuVxPVFsX66ogaSlUr0pQE2pI+XrI2NC/S0fv8vVfJ3aRuS0WCU3mKWM3
fMw+NnqM4GPyhZLwwZVX9Q70oqQ9cd4U2UP41oQbFBIOwgv3jbI5enEO1mKB9vq4
7q9uATl4WV/XFdEP7ZjEYIj3BvKZW0q1zFjIfvB4NpbO9MFXnYMgthQIEmVduD7/
JmK9EmWpz/4vf5FpPb6i97AiSvl0Io6AsMohn6soySCVeHfAUHV+4sVE9iwMAl3x
FgiYXQdbafu9s6dfwi1HdAvHUNc5xmPfxD4Ypt8M23eXSApbnjrM0vJLifMV+7ZW
B+KGdMo0ElxoIwy9j5qbXfkrBbQEjk4kdQ34EH3DPNeCyatpJZGaxoW8DW4AcrQn
fpF+nd2xSVZc1cDPKfwrRU8Rur5dDQBW0clXlIMNIZ00dmhvFIkmCgUXItqGmB98
TVgmKmMbyEbvz/X3YAyScYIhjTd94NnvUvVt7va9rLYhUzEfZOc+OzQuwFIBUVUi
96kDLLmGcYRJG6zXeQ2+D3SUkmDHdAlMK3yr8wtPtHBZbDrIaAWjNPOF+EYqEDvC
5O2J1E3MMmFjG7n2MP6jdaQ4hwXzDWUw5Nlj9hEdd4pKNpbMJ5NaSb/gvYtvAHIA
Y9zj9BY79hY4a29MxwYJ8X+aw0Grc0qgaB8gCDkkGy4LMC9fEi2n6kEzhzkHIEPZ
fTrHuLd1ECHsxO0IGAk2h+7amckMajEakEs76J81/87ijJh4VQxA5lgl5kXraTDU
MAELG51Q+9j46xpDVH5s6p0vy1NGvLxgR4oFqCaOX90iyz5Ea4fDUKZze9/THIg5
4oW3XJErdbw3mjOFXZ1Wujb1jXPmtMohhdmIspDV2mf63Fmzi5g5PGlT159oDmx8
7Gv4Dh9091AvoPAC9M4UGCY20G7fK/PgccgdQrRyoeUe3XUHafMdS0Hd0rPP1tFJ
ZBLLDjYWX6LXGKlyF64JHMLvQonj5PdU30P+ngYJWfmy64fHDbKHF0PRDA/niT/8
uA7QC5aMJKCZa1HkHMc1ZVjSWwkLdP6jHbh7f3peV8Cex4tFCP+SlAisdeWJu/XL
i4vv1tJIQFgpk1O7JNqpMYZ125RJv7Ypg9uUu8FAW3q1M0XAU57fKhfyo7Qjv77P
CbpAVVAmDu4SNQLxS5iV73jhu/GDpPJokR2PpiCHT8FODWz+eQ6BYFhYyzLRwdVf
cNYs4XbK/y48A6uHxbvTr4KWFMyUgI82+9ymbTHvXsIWDlKrroodkt+LAOpNvNeU
aGsaD2C8LbcNpjZ5wkhZLjLaBwJlMMEhNUjLWwWzFVscsj6rrsDQdPQAFs7jjRD8
oD3kwBIWKWA4FkrkR8W8zYYb7dLo2JDCwHCvjgNxgXR0KTt9Jph9vTfLdQ3jSxs2
hWQ+Hw5Uh6n/J05YFEIW1axGeuye015CvFz7iPHyOTcISUHnIsc6+clhEg7CELb7
1X5fDYTPw8wA9fKMyA81zlo7TbCrx87+L+p6M/iIcR3swIA/XQn0ohwg92BywVAd
bEpHKYmagw6O2w4Mrjz+4vXoV+UCSulOMegpinF7CIArIPVftQV6+yGXPx+/mEme
L8eZALDI1qLH0Qk2Pt93Cy50xwkOE8rWmmWlQof0QVReqJ57fEMTvwm+VyLHZObI
ckAid7HwBXfhniUMliXTcj37qjjzzwPYqXyRFbj3GWdDqjf+epHBgl7e3k/UCvtr
xA9llQqNWTc822LZeVWf1doGK+FKQpKnH+pe1WU+tMGdyszGKnyUmMVYs2PNQx/G
/gIuY+friswDOK4hJuzh0thHqKMJ2lSPXYRAMDNrsQ09XR1XJTXb3abbGMo3u2qc
932UdhWvjK8b7qUoCuI+0gNuQSCBagCVMSufbK1cWYBlHywnOi7uTcG5wyXrA/kT
5seD8eUAattct4sry7zbVR4CLKq8EdBTn5A0vIKEuW4NVy+cD99/H9N3CqyYRUNA
g1MwHA/O339X+nJcQl6d8k9MsNF/jcTiwrWvf9JBqtAAALEc1Sm3TdPqaN/x6+53
lUucRPVqE4xGNNzhfBQObC4eyZt/W/7RaoWw4nlQ3AyM2rq9myq7R6T6A+LgJo4a
L5yZMLXpK8OoptgXtGRPMkT7RwfC696KcCAv/gewW9k+Mhn3uDaIW184wG6YvmQJ
b+ssmNOntGPN+dmOqxMxm4py/ThFVFQnjp0l/4Bi196kBnuIQG+xPnqPWoGVZnw0
k35Ia3BSiAvqPEU2vr4JcOswWiOIICfVEwD10e2TUnhEsL/9Q3X9ghtBUL9lXNZQ
3FaG+7PCXyZCOEvUQWYhE7JGCQ1jpRAvUq36e23FB/jzAch+tvJrGK1wEOM3ndn5
G+LVkQ+ikvtUgU3cavJOlpbVD3SZg2bWo2tNuqlUMBymCa+2cH2daeiBqaoUs9J8
2JVNRvTpsU126HvAKr5HbCcDR7LBUlu8n5M1V68ry+IsgS0hffSzLk7s5GUhQUJX
Y/luwVpCUsRbH57C7wJ2ncuFNhGbByABAyErno/yZqaGrDp4JIof0chkWmE/E01Z
HsVO0CHtiIm/SdPJHpUsal9Bh8WkgYtwtNUy+P5nJkVjGRiCIiGwFoAMBGaG1t6U
HLAX5UQx/2/l7piniHHbzdM9dUu/wktoxOl69nwVQ16L6krgdZekOrBnn1c9z3oj
KbI/z0B77x6Sk8EsTgO6T5qXmoqwS279gCcOWTAhe+ozQO74AOveTcUN0DUj6Woy
RprCwdU4hdKgQ3h8d6ja0VPr5K7EN2sHsdIeAk6/1l7TAofzbEKf5+XpIOSl87OP
OFv7mh9vAdmXtUZ5gErV5USu+Vkx18B3SMYvRnOZoCWZyDog63PwZ2IKToVWwJ2o
FaTn4k5vGBjhKodhaRb9Kj5GtyqXM/+CbuMYVlaarj++Z8JE0wu5uKRIroV3DtpC
AAbtmfWwQW+v74y+F48p3m+pBuv6iRN8I8G+p+JdPs9XZPappBHMVQJJ8Pqm9frf
iU4vNUyZJtUtgnKzjm0h5bzrYwhpT63K4y7gWAV276zlofcQK0OrCDF3FnLZ880Q
0QAvhKQ0y6Rrxy4YJPru8j2qT1T6vzJZ5fS2TEXuq+5X+HwCk8FeduAQfH7mfNMZ
dOzRf43EIxq6gyhnrBOe24nCf3owD5lLkY0pSqyyC4xJEBjg4uHO3Xo5B0Fd4Rwj
MxYklYjeb3pvihKrfD+JB1P5vzP7kYTpCPMGRL//A7qcRnU6nEg5cxz9NjM/v0oO
94nGbWJ1vY6VGWyUo0O6uaW205nEAuoNo0mWDe4uo63B1P3PWQfw5IJenvvuAFXp
q3F8RYzDRx1BZzLHNRlzcMobBSy1tyahp/81roVuk0SB3qOnU/kBtwS2L3+KnhAe
rqEwWI1wMYmC5S028bPoaG5jyRElYm0U73F3380fzoKnO1G5FJsY+X+IKeifdNrs
G4q5M1wRQgpOw24KTCGXlxWXvW1d8DvNhMyUF1zePqYdYTV3EYw505Mk0ekpUKeR
dSLst+PL8IFeStMy3FDdNWO0phTTmjqjMX8ioChCI/Jdm/KdNON8E+HNWQGXrWlw
kjf5QCES8qev9yPW4nbxVlMf3Zv/AePMqw21/mWXCtgsZrOblGLnHfM61uPo0amO
ilTU8FonpU4XsFWx4tDHFko8aXrv+bKuM5tsBEx8TB5iVf6+rvn95hyYfsLlJNDF
IjSIdlEGZc/0TKUJ3+DELjridQSMnet01t/ZnWe7MZucePCV7ioYuDXmq2H/Yxml
MfqgB/NYDLCUaFjyQ2/B4eSRj0Do9+Mk2GjM/orEEKP8EetVO/i9f2KmKWhez0C2
BNqyMDoVK3FaMFC8MVo8P9S2X/l6afpZ43YFPpzbYa8w0aOsnj++WJt2MCnzon1S
OrCaUfQDHlALjtJdzpaq67VyBI791eV+pnMQnZqRz5Z8a4EBWFR+kh2YMzmMdu4s
HC9r764GhDkq9+ka3hZWsWkNvNOrPUnEX2Axwo4dua8Evit+zpKB9SmtfrYijYiJ
0iLia1JLpLKG4QPIkDEmY36toSsWV8cICQAtCZ974z8rZhtk1+ik3Ba3TPPulIoM
W3em18WIqKaGoOZcyPK996j4VIdvtE/hzGu94DDmjHMnXWu9P4BNDtB6W+L2sXHm
qwbVK1mvL//zCuSX1zZ9lUvaUXSwa1z7Jr3S+PKRC3eWsmKkmDqUZX1DYYTnwI9S
P2FRU+fMpDQglLGm3L/Csz3EgohDHnb+tFeobRerXxdHm/tnjO7fhUw8YOxTT6GC
XcLl16YtFNIaeJrnyhwlzPSJgTd+GLDkYDMLbQZnbwGhzlDjDsxuiZQSWRYJ/S41
vASwL5msSp3tEOrCBQZwIxZQnz6EQZOc8g5zYotw5ryzCnFWeAqAXTWaWnqMdghN
mkPdlyehZb/rFMnA+HP7eIbyYVNff6wDM4yrVXyq5pw99dA8BX8vDoJtFW900IQD
IWaSpmJfPn/Xs7wtan6bT9HrRPh0ZMeJD3H+HcKWpFHOL0EwbQS8nTzCPQ9gAtNG
rYbkYvZUiv7ZHxbJ+/VBfQmxMe/fBXU4dyqllXrR46eQlLFaENtEj9Z+b8eeT9GQ
Uc6emjJkGImPu9GgO5VQ1xiKeyNBc0dDPpz6BDCvUBtGPnb0PJH26tIGcAbPkohY
eDG1+CeNN1czdAvR1MK3uTzgASj7+2YnYlPqZOGuQRtRFe94pmv8gBr1o0fUVYzK
dtE9Fjv6VaVr7zPYzWczqXaa8GGsj8TbL+HqKMqjKSuqfN73v8jeW4B+W+TzGjGj
eFUVfcjIC59aUbLEc+kKMiZEvyPf00qZI1A2wlqXzPzEFa9ozXmraMbsNi3xgsOH
OXC7FNB6nMPHFD+dRh7hjcc5/qdRyxN7qifzNkNErAcFWp3m5jHmS1hI1GW8VZx1
qW/dyiclzVCzLYMsVWG0y4FAwOrC2erwOGeNWchq8OpVeLbEr56s7fLzT9GcMEV6
DckIraNM74xzn7j7450sU+fmzAeVIzofLkB9nWB+UNVKBjcgkFdeHn4DHxuhR5rO
4yMCIF7CwUF0Tx5iKrGmXE8bMjuw5WC8JnA+8BVY+W2DwLr2ttJMXo8324RR8iNm
5T3/2ygmJa3Qiq3Y+kBCkWeT4P1LZVaKP6nc+fJMwxn5F/HDrQz+ProQsrqCeIgP
YLd1bulNd2c4cHeDepyCMVyzr0DvXIG73Zotis0Ys4wxSDF8zyLCIvsioQkqN7GJ
+KXeUCI/f6GCooXjgBEdHp8A62WNYI9U1d/U9A84DMA6W2FKMxLS6B+jK4WtDEFQ
dP9onfQAyGgVuPn/fE+LrJu9a69Ua4xFq+Bo90nWoyXoP8+qSox8XbkjaUoXrN2J
mj4Gnwa4Bwrc/JD+0Pzp2KIO7d3mBdv9aWqIDU70/n3n8C/RcSnyzDu5cVA19rYA
bRq/NUpLvezk8HfFIb5kwVuqdUGZAlmY547LhWWIMG/wnzgGDXSNY3M2csqs+1c+
EZBnzu8CFQgvJrL1dbH/DBjp+eL/ni75bJO9M0cufIjaJP7kVXjH4Pz7LFWFuPCU
5xcC8Pa7JRkNYhenRH3JutOFEu2jcfHAWj/6M2CSUn6620gN1NWLkk8AUfsvoui9
O2jbU9/Go8QUAtalF4V5ech+cfnEPczE/kXUK9TgW6AH/rAQZg441R7Z9FzqkdAp
NedtyXICQNuJKfAp8USDnlkA4kAGFjiE0JtfcJkP1vtnBp5PZKDrBQ0Km+/VAUgf
UFNze22iNAkJULzTZwlWoG8O3QiysF71P733/PyF0IA3JZAbs7uBbFbXk9mMDsAJ
CJFAtGMvorn90cLdhgs0n7oXaxbMeZsZD6UhECq81p6j6BbMlt1QV9PY2hQwtBr5
vf+TzaEI+5RqZx/ZAwN0l/U8eNyO8bIz1/O7kiJb3wozYb4cKcHfkOliRwW1IjC6
4BOIwH+vEC3Cn95s0przqEaNdd3p8X/JCeJgq0UNuFGLVe1dH8qaEvV10TyL4TWu
rkyjjVaLGkvmClJ+gRE24eHDli7ZZrunwnvMGwUb8wlPZsYwqWII4gPkE5afZxxm
SnHiX5HHFyNvNDvq42S0YcRz95qAzXtyff80IDXcjqeJZOrnc8oop24UYsj+hMzJ
PZRBG3Esze95a5lNlJ9sNB/Tpvn6m87iUes+MG0fZyMXeXj/YGzdblV+QKeLEpdj
m7HNQGbOEndOMHGfsfqSMmtv1D8mz0tjhWfF5k9fpR7vy+Ja6Bf1y0iA2s6Cv0vT
4DlHjYzOcYRPz7EU9BhwYl3nrDTg9vuzWPNt0NEp13bavurFM68DbazwhPD9UcKt
+ukiiVcrLclZX/sHdmWEIXxpmMtxtdlmBlvpN1Yuax+SE6SoG/qIdkXyggPpKV/7
5yWBYJ9+6crKusfkdaiw1YPSiO7zLzpTpJ/ruwlhS0wgvzAS0+2f94EHf/6rbLxM
V/PQ32o+sWshpymFPgdpqqWWQZTB27/kDBUjeflNmY6ZKlxGVbHXwrl/wWPX7oTr
kGHtg3JfDKLsQ/acgx+Gz5m6tE7SrySQZfnwLq+1kA7OdVCtTlgUtG+jeLiNHCN2
xPFIUa/T9jGRbz3CTpE4M88GqUtI6YEokmnXJ4mMfYgQ6PaZxEonUDMkE4ZMkxbx
rFtbYYovgp1jGQ4i6F5fibWLY9Ovy165un+/azWeEHffgZbPxr9GNyn+ije+zFG/
vuhlxQCVuBN0+9rD0d6zWgG5+z0Og4ccikSpczbD9kZOfuPKnPNnD8aPwcnavRkP
6hdMk+K2u0uCFV1PF6f1AZwypeJ9JNJq0IrlFLg8VIy3xqBUrREYWEzUxaMke2qC
7iqxRZkHgk/Pag98AVGs5zWYlQc+3OEKiune4iatwCDEbQ1wVC/+/nJH65yiW2Cg
ctyAfCffrCW2T/znetWddiOgyhn74wXj9Ib+3luo0ALk2gJ1IQptYedI9Zy95VDX
Iwtao7hNHYpcFXtKOmddqNh144Ajrv62D/DdoNH3HK7Tr3RZBNUJiWIBIxu0LzK4
UO5IOqdh4jT3BZ3uGK2HB3NyTKDWzDB3nm51UbZFdqGsxt3D894WuxO/v3WDhL5g
RczYFkn5yUapcujY84lElinfX5LJzHYd6/+VM7Qiij0Tswt743suvQ/CIQRKH67R
R+8sf0muaWrAi46xUjrkDVc7k6QBTn6f1LKw/KsNLqR7kjzILDV1SHrTrWKIa1ul
G0hztm8SKzECvuawa0d3OeGCAEaisQVeHbEViE8bLa3AXknVs6f90/VZhcMFIS2v
CBPuSC6Qi65eUz7r6byla+HUx77CLKWeSWJ488u9YiWX7uNPhUm3dMM21hoPGZ/c
/smOw523AOJ/fKAlv48ewUeftXtIM9p6aPDmqaLfMLfz1FUr0NMMfIchsKEcWCpY
heHXf8uzBCi+3LViKHvjWKAiwTq5V8MiLiRioitpAMqnqAbgguMROF6B1C+10VCh
0sshltS1NnTc6NgB3P/kv5xjZoLgEg2g02OSTRIasNqwq+RyktohR7fIi1aS9Uiq
L8pvxXWf+j4SOcfm7S+FRfruw2v7TUyCbYeXcYs3g/12NPeB2rQinKoUlILyh48z
YJajg9PYjChwnJDhUoR043ROEX3ouhgh1l6keIa7UOICXlTE3Xy1Y0iABfNfgQrF
zNswL6/M1MlFqHw2uEcizqgQFlyW4DgWHwf416WuewnhKnbrAF8/l8eg3ZyzwhiJ
EfGBc9zE3C9L/HOL1fHon6/ybAG9PrPKp1lOHw15YAdroWKMpPV9neKZ8flaAy88
c2Dlm6yqLFiLQhQugjAeK2GerGm9cASDXLf83GhFD/UqqWTRoAS/NwzgjiGqfDRz
QhvpADqCp/Tfmb+4bQDj22CGPrgYxNpRj23Axp0kMi7BtyFdPmMs6z3ZQmovnK0J
sDBczaZyRAuisI1ustA1bYW5PywKMQc/UGOAMERum8xllRM3nkPYyML2gTR4iaxa
OB91BPg6urTNFJsOGX1tfuevRKkIyP9/moU1tzTme4vmuVsk0vevX2lSJE8YCIMr
o2njvMwX0wi2+LicZcO4LuOFVYsm3Pq77V1gX0GmjkLOYttWC6MigQWQJ8sKnMWD
C1JKoijjamRGJtN7oU87F1uIj1oytEPNGmLiWE15DwaDwVpT9Elus7/J2D1cZl9q
PVUxHIuuL182IwUk9FyYPfaEhNxwnN9cqebTu4V8V2GG/P7w+jkcUZ2ychB/Ymbu
oQGwliwyRNGTJY9nihr4rxtJu0GiZLwAQHGlqGzKFc9vRTTB1wVJqW8CQAYENJjc
KmC4Z7fir5lr5rQXRiZDvDqtPovAMMs75LZeLmdrPCRavyDgUBhvnFd8GvnChXXc
fDZDOeTQZySCjE9cVzifPG0E9PIPRpaqCDFERwAl9WGUsXqdP6t0jFmdYMQxzSFx
ovfg9yLpDaCOgUERlS/Sg+Wy747IGRqUko6/vriWXg+iqaaeuzg0yUujDR1hD5+q
cb2orMmfZmS1LHt+0eYXXIe2jyiGc9SZFkc9JSBqN3TPzxm5X1QSPE3DLD89EsC1
DihzTkecTudtANgYBFAkRFP7s4j9ckmCiJu2f/J26pMhalyf5XBkbUrS0c7fMx+r
7WlsyPOMgTOc9UJh+Est6FoeoMipsiVaz+88cYlXgp6MA7m72EJ8yxEb2RwKsT2W
zoVce6u5kn6yftfDcMXU4l6+1NCLFyFj/5E96DCUviofwWW6NOK4OmGfhOEHkxsr
9bS+RotTM7bOs3sPqXdNB2kqHpmVu+2pMb2x9c7/5eW8jvX5WPryscjc3Rhi/ONr
axyi4NOBrrFKqo942pWsWA+WuQJe6zQOvp6uyYij7dnXb6ZxYTAUKzkOVOnlN15O
9YziRiQgYLJiqVG9cabcvE2d/hDzFVWihDfgQJrjYIkVDdNvCYE/EOC2M9RITMDm
ZPEnQ/b9gnz2oYQvA4rw5xS7F7yKbd+XTV5Wn+XfzKc154Dr+8yMomXjm57WYOEL
pz7eJ/aOpGNpTe5KjGu13ueuIiNZstCyQpvvQgd9MtacmooJ1eRoebi3aaXy8yjU
ZaXwis8Jl3peO/dNuFdnHKBOSl7JBUJPFSmBk89k3we20ErbpbbsomTrcvMB8Ry1
CbEG2+QSqPASwwLpOS0QoJZhm+6avV+elarwAZEHjg1KosVSzJgnJiUf6gCj3y3P
JkJlJXrVpHWasF7YZIdyX43EJ91FS5IlV/Jm3MCJJrya0DgNU14iO/QMuTZu1JLV
KYdLXhulPLjsHYK/jo2TNWbdNXfcpbfHevZMJERp19cJCdNX2s7KARBVOgIWP3g+
jHfWvzs8G0XliG0Baez7coYzlyYSEUHpS+tCIqLyxpHpu/KwfiwU0UjsPHynD8/9
oG9pETTQlFSHHHsa0b78bNE8MNnayZ6XpPlEjYvthVk5E2A+OL1KdYrlp1oNm2K1
lTY87ORLYOjwqO9yQ/FaqtZZUOv0r2tWcX/K6NfhzPksVsTINxhCTSpgmkHy4U3w
M9etrzrDTNYahQ3WMYJrgJW+VZ0xwA8TTACy9nbqByg/BtaQA2/nCsQa/zAW7sjA
TfmJ0MQAq2Gb6ukst8A/UC/mNpNR4y5XT9CW2dy/tTTDJlik3zqeO2oFEM7MmWXz
4OBFobJiwb7T0/4KPdpOpQwhYU62kpHE02/FKj1T6TVNvzf3GieA5nEVJbgFlrsE
1CvBJegpW6+/fRQoJxgnQFpVEd2tbyxGvbyBGBlDB85Wiuf1yVfIG4icis93PNI7
Vg20XBk4ZK6YCsSPahbl+kFuvuWEWkFPQBqg7qLJqFZp9NIhtlmkDiVPOhal38Vm
8ExoU6pyAJYE54rM+/0XAeVlnfqjpiJGKhEGaV52dYKI+cBmlZEB6Y7jcYytYKPk
XXO5w63QzHNKlw+cdf42YGiuvjdw3GlxACibw2eN9tuzQwG7cT+Mg6PKTRFreLKH
P1+Mvd/Av4JviEx1WudyO43QlblrAFvLTNiLOVeUb1SbOt8OQjMmGTBmeRZIjk9Z
/L/ywxiFGoKZ/Ke1mJOnh9dOmDyQuAyuPSvNzKokoCxjEHr2dYbO1dF7pGFNQUql
PV1nsfuk/8qcrnwN1/EyUOKKrs79JXwg6eu6O33WqziTOpaQSXmkaZT2Dd4qI7Wf
UPmtOACf7a5qM3+/Kdiw8vkotEXpCLv7GM7J1Vxs77ngUmDRQ9ZsVuaetksiHZXM
JpT4g7u9CR+lkGzJt0uTwMWErWqQeMYypLZ0gzFk5XFzFqus5YY/0JUX/5hRGI1Z
mUYAtJaBAX3/t5c/J3xA+t90fpvEKtgSn0UCU43jwuHndX4ZLRNnF3H3KoA2Fzpf
L+g1lyfslrINr6GKuad4pg9SEy07Tgd1tQrwdxIGBfdCck+qZBH9wpO0drHJ9kqT
rO+X00MRUPVp5O/dxGy9QFNT0WBKxNwfWD2Y4c6knLthBFFIDKeEVou5s1uhs5eh
L8BSlKQTzNoNft80FPy0kEllgrlD3F2LL2OUM9qp4ZO9GyU/PcFFRK+M1T3RC8eH
Hyn4LdAKfKjoxGfkjMixfx36qTyoE8qfyPHDC4L3PTC6m1UoV+HSnni4Y+QGIDyH
+CJsFORR6jcc9fD80Gnzkoix+GJ5xcfuiMfMin6QEeg+5jmPjUWvn8ZoD/Ie1AsJ
HnRwfk7SjXOYarhD672vhNtdL2adxB8SczfPIsTAvBSrwnXVfx7Eo3JTXOuOY+a0
0nkaPlcuyDFyDLVlayXPYj0JNZlcl5Oppshz1ReJAjXfXo5LMVKEqzIDuJUKxL9o
5C2cRputX9N7etjS+bJqS3aKlWnY/acwRlJZcexhSu8A8o8Fy8i0pS9xqRyKFNQA
akOwbflDlERNI6XLxKNnQeRhDvgC/WKUP0qRwF4v0tU+aByHSbOTUXEZXwUnBR1F
ezbKtZgAmbO7LR5fCP7DZkJVRU2MaV4OFYKAokmo2dM18Ne3IZGJj2ZLkWUm9doR
XuwnGTMpQMVj7gj+Fdpn2rMifGTVHCwCKv/qFOL/B1siHfwsJy8Uh6hkLtp7U9Q9
9ErkdAz6Mffuk3ghjXijYDp0+UCWKl08A8KtMrviKHVw5ku+tXd6I02u4n4E5u1u
2OCI3zEaZklYhg54rqpu3fZpxoEsGdS556nTm2GtE/O0hkeiSkLPXdZ++IA/5wVV
lJ9JkqWBsKqAP+QA+DyztFPwucGOqArj8JlymnrEutVEb43ysCbUS5o6bQIucY27
qg3CvsjvogxOfrG8TRZTmmK8qgKmclISjpXCD0QzUheGhgFVvPeqAT+jGs/qIuzz
fKxmTyr1f8hXOSO7uiAFDQy7heP5MQOe7SPKxe39dJH1S8fMwDOtqel/ximJVlRl
CUntuhhWMA+m3q72nWxQuZmRr5toS+/TorUrHkmgQCtZyyJoXbasphiu8i7TdqN7
3+o6GCw/GP/jxlVIBV4a5FWVtiyZsk+t+S9ucJpTNlWIEJXfIcODTk47AH52vmO2
KlwmpX1rtr0k2DyCadsXgfvOJ5fvT2NmP6jdfoINQb/QMTIQLsbPLkU2D9pWg3AI
xd3CmJYY1OEc8nT2kcZBd3ZiQnOPv4+L6nwiGmX4uVCh7bRq2cpLWrSUxPJ1u0EQ
hyhGEMfVlyRcRZwQbXKFjyh4hUw3yQB2wE0vON4H+kgM+R8gSUHGfmNZocBczaIY
OQvLebYROqxQtIO/jZyzz8665VClJ/FZ/Ww/7/GlQP89CEGpJ6SMb5qGMze8giNx
iM5yc+pOIwqbZzGa/J/yCAev0CQz9nwnwbq+7brM5xqbba9Iqlooqz49YQWbRB2G
8oExnuWIKtZxKkvx1XCjayY1xJ/Na7VhSfEyCo5NvOVFh2uLiI/YpGS2Qb7yZ0Y4
ZWj6n92AbIMAapzkOuDDN18fTHvWhkluoVsv6pSulF7kcuk3EPz6qi2bB6iitIx4
XCKb9awTwM4vHcqNXK29bAlLqncK0sa1kEBZ89f/kCWCL+OoFWfzHOlJuyQeZrEJ
AmazXooMH091ii0cYvf9IJp82K4SaB/gq3gxPaxqp4s4ClewXuZ1MfVKyCi6idao
uCIQQXKQ0b9FOYnFsQislTAkga4EdfH5F5zsmVX1Aejq8czovLVThK6cLSooYJdB
Csl5pD7IOek5xvVI6tQnWOUpgsyUQxCX9SoRUc3K+1Pje1X7po6DNMViI7fi4CA5
Rn7OUkIhXDativFj7pnP4Uv8bd11MGwN4ZpmUhHEEGad9uGbu47F4kHuv65sVXvT
XvaSZGjosYwRR78I4xhntzJwuzxPI5fsChVAoLhwiTHClrEW0Sjwsvym0vgnczbq
+gcs40NF9LWkoHMicvNE7ar8cAhUHZNsE26JuyJ8g40ljHwmy59N/PegRZFTaeqM
GZOFIN8EMfYNhPZbR/uYNFJOTKTuBe7vYwPOMuICFHceXKzjhSBOaeelclbmMk/3
ueLwl2gd0FpzGCU1pNJtqMs/eIeeBpJCT3+L9yZvgDETh+hDdwhiRU62m+cXxD1R
LBct3L3NNz/gPK/+i8z81ydTXyI9RK35KC6xc1CkPNdqX8a06lS3kTP0/spkLJmp
d49mQiBI3ecmCoxu9JevmrAJXfQniLWzu+RAsI7gbZT/I+whlsbGKUX1TpDBCZe2
jTjS0WXZuAbgMHmwwTCFp4LcdY8IoeRjhOAcIgjfy0lCplhiy9GXwqx9iJ5hnI4x
7e9U/GveoL9Exvoa3dPfuh8DfuI1v7+tZPHVMEcn0rS/Z08Uxgv18w9I3NEM3+/w
I8pLJPDW+6mCvAe5gsHBuR4kCTAQQgye8wt/U8Kn1s/PV+3I0LB/Jwf3kHIq0dvF
G8EnNoRwEq3za+UN+ybpRgtBWF+Vc/OonQFGehAmtvcJXWcd9VxA5q2I/2LZQUKa
NxZYCLuQzSCLpKSOtyCSm0xYM7/ef3jRa1fhiLgrwXFmw6vm0BKCF6/X4gJh5uQA
PdmTTJ4LKdtTHwp+Sjrah7nCGRtRMOaqQqzNwZV4lITCDOE045NtfKf5oCb4Mtlk
P+z4Vu9dMi54yTkJDBpC9/CdXK3lo+nmSNf0MY7253KMN9dt5mthulo+24fK2Dz9
SqJViElQzfbAJhgwvkDv/ENj+gQhh64O8Ck9e5ZJSAj8xd6Kvz950Rcv8RKmCgee
ILfO/CF7MGlF6j6TCwNHhibVSewYsIyUlKlBxD0lA2fn/5TBVxo7oTO/Z9hHGsPq
RMCVqkQzjF+6IYDLs3ZnvMfOY/xfnvzxakuAhWGb1qIpq8YyWINFtHeKhcqv/Vtm
TMbG8sPi581+B5nuMkD8NqCkzPDC6zlKMbD0/WvVqL2s2wdQvjnzdtCX3RlmShQ2
xu9pKZ9csyQXcUTT5LcAJ6anWCGMh+sW++uisgYwPfzBmvXFFYlx4Ux/Ay8Kv8vE
XW8v8EvSFSyPlMfagdu2RBV3LjP/PY7Dg1GNIKTuu8VFH3syh15IIgpducMv4k2R
1S4AHUg3kDoZE9sHlO9/6C49buDSCjtLFFeeDso2Qt/60jAhPGE1SizrKzkkmytJ
9iOJuFqSr4kFWbVzhAHxXn35LMf1pzOIsFJLjYJNhlNGOXg1ioWlf9H9xUGyfN1k
ja4TCunmE5j1qH6pnlfAWmZN/kPnZ7vulEbgC/70ZLpeXV0dd1mUjiamfT/pQwHn
UA/GwZ+0pbsv+SGiwn4Hq7OB3QGR5tVu3N3+ktbHc8QiLtvC6h+YUdolSQLaJIYH
L77MQmvWkuXJLYImzDuasbSUU9dhb/fgW3xQ99IyX6EpxuBy7Wjt/LklbbDwrNJD
N/jnwOhHzy6KvzbLB8HWYA+1cE+Oxt6FdYzLCJgELavSBr3km0Q00gZypfoGtfQi
pyjHfkpGLyBEQlrFb+lIVxV+mJpLmTSK6CEccufG37R56ByRpMAVR+/NXfi82H5c
JNHTXk7gp6osXkdkQHwDNVlW3K9x+ZHldwG//hGJITcgyhncdrls3cO0iHUawAqw
F70yitLT/xa4lesm24QEShceMTqsXVGNfvTMHCpsWyG45dV4J2GULgoepZBogMJA
X7UNKfa+fHzFXJGygITMsh2eCyEBcWelT680CcGm5eLqeQ4V+L/h/5D6m9fYlms2
awy8cI8YU3RN0eGl7j5BWfica+LJYutfmUigjJt9jfD7/XJaie3oc+KpPECBVYxA
fZyAkxQTI3lJ4JvIVYUAcH+XFcqdBdfNt7n75dfACM3trghIg2L4lq83H/WYLMwi
bN4zQqbal9xKePvHyP830gKy7eUXL9jAK22ZY/IBiXzwmjl1U1HKNaIHcDGyMF6h
Mee650F0oUMaEJogMh5HDQOL+PgX0p1ywFQ1V2izSgAT23EKrtE6VJmIa/fWOtf5
KbfLofpSgFwEp0yOKo/4jPqqojPpfDRBUGCTqQ0MHDeoNectexZHQKsAHiXQdPV0
BelDf2i3J/lB1NJVRO+03yYp9YbjRM+9sYprpJU5KJnD72ttJyVcfbkWBDVnbiQH
rrsntjz2MycP1suwAayKhW8PCp0vGAJFjLhHsnxcsVGmC54+yPbbYSRIM8o00pFF
pQ9Zszqwk/7XM2le0TAe2/qQt0tVbABxZWmdfH/D+rokg81mpv9ruHjChFKj8L3U
6ENaWs1RnxRiG0gjrWXmGaaxJPiaVoSIw6ngoQM//hLdJBUkMQKMijF3DKyb2fU2
QS/0aLpOZKgiKQPXL+cO5hK74POp33mAhB9lml4Y1pZm3BB4eCLI/S2HBzE/hwI7
zdzNIlJycvQTXrX8eOR35VZkaeI7ynNJQEq2bvfcl2wy5JOOq3VMW8GaSKYKQTKz
nuATL+KG3Klx46m6c+I3FX8J5uPLYf2nE7BCXnOy2Ca9baxixYxE/YvVQSbjvCQw
CAKgDkpkHapowaSat3fDE019bQwcbmpFUKPzp1x7hPp+kmVXf10t6Cp3fqZgBVWI
1PalH/gOyEFS5YyhGq+xI96p02uumQ5fk821Gq7LfwlQGJqJub/fhrSlDp5R+8Mw
7g4DN0/2qZtnRKLVJG/d0vvEDuPE2VOkjjufa4ftXdtachXTY3uXeI45lFHczE3h
VHbl3snwI7Tau1o74EyfCPsOy7x1RWYx6sqqZzngNkkFTttTR9l6+mIMDsFqEIiJ
DRaD6RqQM7pMfbfB7Yy3wEAPcwChCILDrTkmS5DxnbOrkkQqMwgNqW6ER83yoRyN
6SN0zHelzzJDLWwtD1a4hsdo9nfPElzkRmhsBDMkgh9z47ZrJG4p7APqQnE5oaEi
NqZIgaxb5BIQBf+mAITKrvji/Lu+rc0sLV8FFsTArPH+8Ze8gV9ARKRSZSP+akO8
4TtSWxEAW7HUSwCtnxm4TLCr+/tH/EP5wRezk+ST7HV34LiUk1OaB0dlwh7ghPvl
yUmYJcicqLr0QMkAipITE4hW20Uluyzpz53IbKcEFx1FjvzBuxirA1l7f4x5RD6y
I1XuIttBmrpMSnAgIpXfsAgNLNBZ++se82ID0d3ieumuJKIfclcu+PtPqKxJUtKv
J3mGmRiRdR2ttSPkWVQw7Ox+xDMym6c82xbMPLBNF/2aGa9qJK1AtFBmzo7S4yvH
4sWneSlk0Eq9pxf+wkurTtv5PdKPFOXLHe8mr0yuuVTlNLFkJljgn5svjmLYHi01
et1ek38OVkY8sH3IJ0Qf5GKow0KqySugSwnpxKMpOYOdNIodnKzE7NPvBrWexIFd
RScMui09zT0+wFG6p/z6OHGW3gG4UGl57LnDOpzhnhDDs4w0HMEyxXhvu+FQ9ys8
LNYyiF9Qw/A9a9BCVKQhu9IlYoT5AEoejAUtltjlRdGUcLMQV+TysdJ4OUp9PJTz
Y+wtKOFYqfdPa8KGb9O82PfZ3lI/vB9dbInJKLSkF+CuLSagzeJj2tAm5JYppq3n
0IVn6K5aSsNA4S8KZVmCR01uHTtDfdyjQl5RhUi8awyCYg/sWrCXoBCu0PBcywJF
7rnysb/tYjyKjPYJGcxXaTSVZlH7gFixqU7Xexz1KMxqu2QyYySNpiy65KytPUUO
cHfgcWWNAsh2W8zte/o61palqfFZ+R/IVldquTZcfGQ/tMxrFPEDZpUepnJXS9B9
7fLBGyf5CvaWZa1ihEOsI6i3TRJud50UjVlxUMHLgxP5uPholNAXtvYJeS26dSzE
0EhAsz2X5YiZIx+C/BpycnTd4DKwyulhB2ZNRdkYse8yHR7fCc4v+Zm9cN7vyY/D
R88YUt3TnXxOlgs6kYCWSlwP3v7PM3TfbW3ZdwT3+e+Bh97SfDP300NOjmkOBXkG
5N37wvzMlqVPyTvRAyt+7+tOXC+tllXWC1Q9DU+Gt39kAOZ7uluKhFESXdl4bgN4
J+KjqK+AMiVQ8G4bG01CfEDWaPY/oHjrJaQtNuxABfvSJHIx7xCqv4ZPt1JdJJnr
wfh/FYkswZK8/BdzopxF/73ZQEQ8a/gBKAd/S0vj4xJ+G94aagLMcbT80pNvCqEN
eMfUtfR0fI7zygAItS6SjjdFjKnS3qTIRzSD1UEPSn54EFQVb5Bs7NbdsIjpUZOx
K8apDdcD6PRJ3C6YU/YmeQtwJPlJiD8+y/4sfl1XcAYgPpAKT58VtzJ6bNH1vGYc
rhsagx8N9dfDJEIrL6XzpXvwYWzpozCaPr2kpzBtdP+nRamcj5B+v3S0WAoMhzhh
mXwSiTdexh5n9zx+NBixsPd0DEb2LCYBQD7bvHwa/pVftAVLIhBu9QkJ5i9kUuGI
AElJPsxkk1CdVcZ1gYsWplRKMgtlsLt8eG9QZGy9FLBek5wJa5X6xz7eANBkd2oC
OhENEDg2/WuRFxI63Tjh4F/N7ygKUKx1R8IAs0yXIRAKAyjlAtWkKzn7gXqtE1yV
fdZSqBVRHaZezln3I0XOfR56/70DWfvDQqhe7gAuca6oWvMXpu3N9nGt/X/CCsXe
j7L7xZMcCzwrLX5rlfc3MsKI7qgqSJwJCij5H6mJ8V9W7P5mIZH8fjhPLNjrJgu+
rKBNTF91Zwula6kRGC41iAO2mmlwgQuuIlpW+lxsMpVHOL+uOiVlGX9UzdFvLDtL
5k3ILphZQ2xSlwzLtsbmHK/MUHYnIjETm57m54KG9nuW/kU6FJiP6DczmLwicMQ8
b6uF4s0xyqof+jYMQWkCk52y3Q4w1nVwdGIsNasNvAQN5/B+HXG970QP0a5uIGTg
8JUlYXo49dAoL0ex0rk/9P9j2jR2d4YhAc1AZ64q57FYFj9w6CqKCxYHllcMI9nW
147DWg+vG0M+pP82nWWBHLkSXrlskA/5w/KoaNr5cPPTFEigYqWdPXc+yDySPQcZ
hZvfNuaYu6PCej8z7zTq71qJG4OYGhH4yBmYxTB8pXBZ11Ud4RNjsI36o5ixJIGk
r0DlfyTifyotcGQqG3gNAPKqHbwCgUNbYEXsq5gRKo+BfmNpbFtXbBasxz97q0CL
vyukmxLDEr0c4Z/QcYfQQPFkiPZhWElcDOzIrNBDstkEb4ZrBsTMthTZ9iAFS1ol
dcAVnwm1mZc1rKKkdwldfnBdWKzPzzdkyPSlnJjddMPFFg1fecCck2g1riLl+7ha
yPxTPzi83WGhDDhGMEmmsc8Lq8SjoVkQ/1XnwPFoMJWW3gQNgh1Kec55lylozy7Z
gU69cUuEQRYacsFpDbJ+km2ZRah/1RE9129geRdo6yUMYEphVFtmvvh/ymAJ3seR
AKAgEF06IrULYda3OTus5l2+UB6b8x7toRPjWBabHdnvI5c/CqiDot/nB2pJ7H0D
jU7wbv65yHb/5hvNPObHmI4VZR15e4ATaEmsVVZuuG15Hxw6GGnY0oPN4abw7XGA
/QElndNwY8dU6ingFRGz4pD5q/5Y7nN7kbEo+d0eKJsnD2BkCYn/R1JJ19WOeR4e
if8lo0Y8LA2wXssnPQhGdYipx//1lO4wjZh4aRK6VT3RCpaZfM5cO0h+BxtwRYVK
NMH2zVeLnmVgOmkQmKd0vttaygj2eHca24JQVoBn1AOQvadhz9X4H4H1GQvfcWUN
Qa75aW3zgOq//DJMuxPN2LROq/oCeP0CtqSdkCYUa2FXAWjg9Ls8GtbBi43/PJwq
AKHH9lKeqhbJ7w6Rv0aUR9kzbHGPP0g1qF89y6A4TqZImOIEszrcesXnjFnT+aS6
sRHk/nsWwDRrix4ddAWhxJtpGSEupdLWBx2Gc3mc3t9ZOKQUyZs3suGJ6kj6l4JY
Lh+H1df5SB5PefJBe+66scALzsHwfE4+DyBJbWTYI1f40bnHLSdty+yIrFxSeNul
yAhz52+XHy/htgus/FldyiBnlH71l3yk0EN/E2X2P+sheViZIyXxto7XE0SLOx4Y
rCLkMeTo6or/kiMTdroyvUGUlc9pC763EQvrdzE79y95WDK9uFAlDNasTfLpxdY+
heamAKrssYffebh9AxbrfFKnLoPeoqHREs7wjqFLmnPax81EpXQg1Vgt+OtvhQVN
IQawwau8Ui+HsbBxDYbBxnK0AToansjp9cU0ngeuMXkBp91fuyth7o/fFtoZ2A8L
ufghtcBbzItPFhOgBndV8WDxs8S/eTGgcg+ybc6zd1paZNuxhkjXe3ycs+cR+037
Lb0hS3MNzjB7grjvd9jmw+kdpOEUdoikByxd5/IOP78WauRFh6YMlLR6Yiyx0Zsf
ZpZj4xiQIDJRS7PJX9hRzjX9jcLxYGAu+bhZ+S3EkcCbxjKWY1eGPZV9K5qt3m9X
3ZnspcXQuEnILOfopIzR0xv6IdO9tUClk6ryK3q4LuUGsoyzF/96LR+9nlgQI7uo
E/1GxtFQJ+NhF+/ATntezVz22cUreY+vLvYszjlqP5u6sE/1hxXw+kEU1CLno1dt
WP7Ykw+tbWYeV7lVodpyJXslS46o9chQGBgbuP9sqRY1K6nit+LEeeRryAIppu51
XiW3IoC7w5lcs666XrBh+3rxhd4olrAQFWL2VYnDLJi8kwg55D8yAjfS9kBjO7az
/PBx6hO3C+L7LwP6HzsUK08QWy8ftGc2iGEu0S7e6fI7fCo6pMp8vwF/j5PBhAQ1
k1ujliU9W7IWEwtVgX1D4VKoYFyESgR06MiqZdWFtuHffCxLwLa6K80GamyR6vJz
YZSR9pjw9RsCJt1WSKPXCMUTxKbaPw18kHOnYLEFCc52yW7a38FwpML3XNmbylOy
Ayj33mZsoL2AaVozNKGrDUGLINIw+iUhRQia6uq+MVY3f+SMwdygdWnNoQgALw0S
LXfIsgJc0u1dt1cDedpnjoODm5tzy96xePQRVBWwMN+rFyA+w/OZW3uk2FqF5MaL
kQvjEzZgc8tZAPmjGGaEs5fAwWHUvzkuc1W4DyUQesGSEnfaQJH4dWPHBeBNi0Ut
m+VeYfWbv0FuqcodJ+KlOJ5P15m34Oo3rhDeGE8gdpzoFuYxeN+WSpKO5hGkMaD9
JcLCmGSrStxn/KpKfAICxHRecR5LleahYHVqFON+b7uI0N04WfoDrv6XGtajixTA
QIZGvAQHMOm4mTVpVkhKEdB1SHbsIJJz3xO8YtGuoxRy/3KzEDMUcBTYz3NC7mI+
oPm8DbHQQaj5yKKRdSWqE/T4tMW9D9Z6j98eCz0g+7CoAa8adyBvmXv/J0DB9Tyq
gmUDaizBmMcDipIa22Gvw59GKD4xJkJ5DcDxJA+HcaHakMOU8aa/rkpxIwrJ7WoR
F3KZSg2SwzIzwYTISssSan/1zGPe0fQY2gCcNajSQW7Ik5VEGMB6ylpsfomi4Clk
Ahu1W6lrOXnzhNTylp5aUo19to8fY/sDIgjnmDKYMzlr+wgNnlQ4RFuo/r2lL5bI
UnD+B4eyNF39atnNRKTgF7geY1aOfj1yu2IzXYgvuc5pF4J+WF8Tl2rmXCQn5BBG
MPw3W51JXnYWUK6I+sP/Z1bw2TRnfx47ufbD/MM4ivgjQ56TkK/Q/MlXju0qQgl1
ZagzK4ucqbZGrbZzo305ANukeyajhVfz37/JtoShPC5G2Htea7QH0RRaVtMya8Ix
HxAff/QVHYLfkVTFqO+NwouWNO0NrUpfSKG0/lk6C5B5iir0BzQYa42Fsha5asVI
fsBg46H5DkCiCTtrZ1V8LfPQV/N38S4yXx79Pws+SOrHxrbLWd4friKlA5kPjgVe
eieKO3xrIvxdQ/mCClSedAR5ho7iT7a8nDkf3brn3/Ppk1Go0aYnHBRifVTYsPm/
Zx0p7gXZ1xacnRkeQIgiCWX09tuD1llMjE9HMwYvn/Rc9cNcUXHDFh/3GsOAtOwE
Id8OvSIaOoD0Ju28r5qVgFQCAjUOHYpnape5td6vccmvYyMhxp+00cL+Lx0OsVvs
Z/Jjsb2hN+wedPkUtvb2ingCfORQYqy99YRyK27ZAM7FfzAQRWGMzEJf3MpKMfzX
6OG+hdaTkEUFstHaC2amgy43l66GgsueyF02p9Rh6C6e0U+FLPhXWtYnaRGxT/b/
KwuIwTGuKC/v4Ta+Up22KL+EAI7a9AnLfYO7nb6yxnbhksoDN1UGxjQz1569LqYK
mDvaZ4vj6ySGwm4bjefLZZm7GrY2YNuU+IYm4AstndOApx+rpsYH+awlrqqs0ybe
CRVpg22LLYFrliWiY7AUnScp33MYDsqYsm0psPWr+ztDwRciqpHQ/ZW3z/qots+c
2H5JHC4AVNAGu1vSzExjeRj2LaEpGA8SF0Migp+Ldqz3y//1XOvjAQ7EjHut8W9X
jo0E6PU7/qm0CoVp8/0bEDWw/VpCGpNQ/WnI9ZW7p8VwJSDxlIWt9Gi8YzhQgkUh
IFgKX8SvmtQrRn/MIgU+7wnJ8rzAHw3Dq9kYftAkEOBprPo6zPThEVlF1jLo4c0c
Sd6xno79eWKMeYxuFwDiplxoHuZ8jTKFHI0JLC8IW36u2FTR3YJt6hDu8+qUeNn+
uUxBmLuT2VQuMQ73Ksd58mXfjIN84BH1TQ06af/7gpJK+FPXC4uAMqiuGYKrJj1d
esKXtJiiPA9k/0NK6mAo+CZwo+topaPwt2JUnAq5VblVcUMfOP8ykLWy1xiJvnNz
EsACgv3qFkZxdgtSiPb27CUIiFPCEu5/v75ADl5ifAEh+efNVhObSdk3hbom6tdS
ms/FSZbaMUr2r65JHsMVza5O2jCk6aozNrQP9E/EzEiVfiDKyuqsMLbwu/06D/A3
01GiKNie0D4fONvU5q88APJzlpXbZB/+X/1XLzyr/PfXxG8jeHaKsLj49q5+nKGW
KxWNOLgA9Qx/n4LRsqINAXOHOoQTPG6PqtMxcXeicztFjPZy5U0zskMozG9FM2Da
sKLwA1ATjZ32hS/wTJmw3fhMtkAozvGM6OkiVOWN+cRMM5jD7j7hWKM43U1eLuVu
ZzkaKtfBagWvbvSYlkwTwZD6Ex27bXLqfbENVcox6Xqik2X6lDeCjHVXpI1md3qw
wq3cY2brfFGpSchK3fw1UcSsxvJZORFIATYI4woPr2QuHgu5t4U5vnQ6gJvtQ5L+
T+mzwgdzKRbQAyrDkBWB9FQ4KqjBrCucJIqODGAMl342jkRh+8hYV3ZyWJKzkOXQ
bsO5DkTuIf6oPFf7IBpfU5UiZcJ42Uk5aITRlL4UKxTZPNRq0axZUFV8hYTMMn2R
RZkXf/OweM8w2OFwgto9yuNeIElJTLeze5WCIdvruCINklyApMJ9xF0pjweVnjM8
pTcEpbOORXXsqj3XSBibuYlsdEcOCBg7JavVSql77lGY94hYAy+kzTDwRFhXoOIq
8ZTzFQcMWqWcYr9m6Ub9W35SwPXb9RglqcXv9GaRSPOLounFV7EXGgRW35LO+mAN
uF93/+egC8rBN6xtpCyD7abcksdtUbtwJJwNfYKeHBLKKpmtcY9uuaSxpc9foSaq
U94pLOa04qeBg6YVfxqfkkB1HQTK/D/88y7wNX+Lw1y5R63gQAM8K3JCzGBhay/T
C2ybanUrGL/X2ZOTOVYaX5p/B/tN2gjODEXwp4w8dcwBw4eqGB8byQ0SOBcfpacF
MqalSZML+QPZwj6WjL1ipf2QfFrSFW3tur2wc9wChJ1l2u1wzo+ZAbNzFt2gpOin
5Bzw9ea6Bc1TBI5rnxLgQmMHZL7CElDEjB9cNd49ox+cf+fmFcH2PV+bn0ZSDNMf
KiKZl7fJZum2WZxRdyBIdNHl1594QsWANyRXHxiLo9/NJYL2U37EhChSDDeaiY7G
s7BchohHM3wvW81MzWqbNzawzLouC0UQLEihWu8p3gfgP16jJna6xygtAiz6bPRa
uTQuwHqV+le1URt3EEq/GthNMaypsD4z9UmEHXqyUbdWKWt2lbqRvu2FOQ3jIN7l
mo4zNrlZEZPA8evAAKKudTLEZhz1Q+JqW+qh5tRN9fPdtQUn+a4zbwUvlW1GcAC9
xy6g3HvwbvInCEtQ7YrStkAgSvuCkfK21RnmAIFU+2zlDawVKvCFTiDXfzwckd1S
ci0lXGoITHSL/Nfpc3VR4cdxNoAQ6UZpWM4YkxvPPQYcPN8Z9M6hIVtU5iMfN+tU
wwmTJf0qzpRgRshEsAYznrbM9bDzt3VIP16j97n9z14=
`protect END_PROTECTED