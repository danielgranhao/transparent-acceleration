-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Yu/xym5UAqyhAtGTwWTdDpWgCl5BEVgvUK7rQ0C4cQZ/QYYDHSDJK2nvEwMWcx60zUFS1KOD0xf7
3/hnYlzhBBgdcw5LY86LceUPhULBWfuYIyqLtBzPpbkACy/j/K+x57X1m1bD1rTVq0+e6P3q1sxF
kg0olDewhSsGTZIOoev8M6/eKX8J7Xi8JC/9S4cFazl40B8JFmmKB/o5r+J8YcAR8zjraSi0RzIU
dXq9wcYXH1pIQbp9ZLuP8K/jx/J35bvLrwB1Gt2rYJSUmSq+6xr0XR3eacmbA+1Sy+E72PVuwtpu
s1aNCq7wxZhBCE7vHSM3KZBvmowB+bR0c9sccA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5216)
`protect data_block
vLGpLvF3A5hyh9QzsNtr8WdCGyaFGlhPZZkNuZ64r6zyYfTsc5TLaPkSN0o697oyiIKG4yP3d4PM
txMpsInY+7GiWg1JPCQCHK5R1GW5WGA2NTiJYb4fH1qqPUlWJBNpKwYCfXTZW1kapsRptTkm/SGM
uo0+YYmTSHMcDy8Fn/AIuWuRvlGvek/ScXklSXjf6t8KOLUwxYP3IFYQ5tyr59o4abxTMGMxQVe5
LQKotBajzv2BYt71W9LC1jyVhw1zsI/CdGx1nwOto9zyj8byHATOyHzjILnUgKd1YAKFG7HKtc0Y
O+E/z2QUGjP0fDDk3XL2DXTxbIUKDYXGx1Y5Od7XzU7v1ThBqpHq8Po97lwitTjHK/her9CKgdE3
KzNJEMMfM1cpeLdIDEvBgfvALbsmou8xF2sOm5Yv2jlCUR8f0FSlxUEeQzu9+zXVSRMB8nkLD3eL
TPCq+02nRo2lmGC3XBVoXdxdJM1vZ4n+RS7Yyom68j56AZ5n2m0MtlD4Ex929A3rJVT0eaRaPCR5
noI9yjPKFJe187v2rn7nOl4ai9GqLBKH01wHRi9smdn3+R33rd7zD4F/65XLGYJBuAwWTwF8mziy
qoBuraUxAoUs4S989XJjZopJkOOM7yzeA7Tbx5v8Qy8GZcFG133OiNxtksj4uF51LEhvRLqdcPT5
9zgBXJKEId6K4mP/budQ7BFXPHieTCI2Gb77iJKvnGr4Uxt3itVIjm5HAe/FoQ/mU9GRYwyYyR5M
mqUGhmCtV9Yinvdk/b+I6gvotAZt1QNTEXMXjl6ElRbOqlKuRqeTIbwhg4xKaXsEMKGekmtuAYvX
N/2nHa95/A/LGVNAORwAyCrW4QmoO7qMRnFkN3CZut/pMJ41PFiSzMiuH4ZKJS2/52e/YZG+44Ay
XQDgAZ9Zq931h8APpCPShjiKJ5d9yCNYziyZaKkZkt6Z+5YoBfq6v14gDcm1iQBBlxy7p10yrgsp
okaAmKElMHSpJhAqXKDFEBbgVY3DPq0Ty6/lCsridL/xUbVuIPFhTZCRn79rALsWadOHXnZLTHMM
/2Kj+As9/UiSz3kXSt9N+JoUh0p9q/ml4H2Dcg4OoXOuLXEf0Hq+GwIM0Z6yFA+26ZQBoXuObvJt
E9GUTfuj16FoZPA2RzCtFB++Ye3LrZ29L70Zy5e/ET0hVu4O3NIm5UnNNkh8QIvBU2DQTGO2FO2Y
N1d63kYoE6wuufwPrEkT7VLmCdM4Lart2xVS1Gp6+2El9h6BAIzSFDpcyThnECoKz6qfIHP9dwA2
w6WBPDiTBdxhgnRiRaYGtkdpRGboqaqpbTS+J+bZ9aH46DodkdLmVTgEFtbVvAjMwhcb+oJ1WakA
3s//qmZqGS6bj1u3CsSWa6TG36NOKNVMO/pPiRx9qVC1QKdNDoRTDrl3CPNOeg3SfO2htjzX+ypv
Xj9DmQWEeRgpCi1jd/+Rnf30X2Vk3mdclX3qLyCZ86AhPCiODAcMwDTWU2vAZVV+VWNDI8YGXngz
K4pb4jjG47jBsEpNWaLCmxBTq8z4Rx5R87ZXEmSg7ftsLcDJkW3GrEWuwKFoKokRMrW7frV3g+gO
CgHkmLbBnurA+lQNmnKEK+LI4cwfmMlImbce1DmG3ikyM79sT/zxskK6JeSGwDPKkBmljNTqoC3K
tTJfDTmHWaZGPwMntGZZtEorU8sROtFclxrLsn0+Y7/ypGN1VXdSGQtLQQ28pPepRHOH5xeEzVRU
zkQDZgjACklG60FUf2grf8zYOdArhwmq5nAT6AZil2uFK5ibtVN4RYdsUWGmeLKR8HodDwoAjA86
A5/GJEthaub64XOL4dsERP3JHTfYtLSjuzYOE854YT+IueygFUFJx/fd+5gKIHviILepDk1rQINU
8NEV7JfiMlz9pxEpGLI+b5GoYafruvXOA/4yPFpEjuHixkOd8fPPGyhzIX/fDuUDA1pTGT6Jx6Ym
vB/avZ+Dh+EIYWSSr+blBQHtsn9tdXw+mv/LhlRe+drNpwtr4PmAQHyvjqnVPpkauBLsPbiribFN
qH67llcaTmFQWE1j3NqU7OQU8dDEzo408GLnEE89o70O7XPVbMbb2gAOuWOYOVfW3Yzwz5H9qz5S
U5SOpUtDomxCyPSDFkzQeu0qcZ0mUIS4v5kTiipyf4tW5t3b2rQmTPN5vgKJW26Z3OI/TAUMI/1X
SrPBcqrsLzSLOJ+eJ55Oqz5TEietJm+pAxxwodp/89FfCn/p17+UQhrpunGv//VP4arcrioMzZHv
UCjfhvqzIWnJt1l2D/3+Lvg9z7TdA5Rqa0kXkRM9Tu3LprzovQpJi5O3CC9iwefmT02WXvPoBUbG
w30KfNcx0JcbRO9GjTwswfWeA2dZm11SX99FbLXRz8eEK1JMPEDKG/1CiySh+5W5+DU1tfehkxnE
lrqFaYmDR10cd6ouvcNNyQahEFAAL8WiLmPy/KEtFyTlf991QjRhLbygytE/DbyMhGSYxmhXEkLL
uBq63J0VR0tTUfWtZ5OxrXXE6dM1drkh78vNticdirpYK4Vu1u4X+qjUj/FQWoMKjSo9381WoP6B
+C2Ss6//mZuDkI3Kg9EDL4AHIMyr5i9MtvXZEWFF91eyn6J40HNyx/IYgyRZT5RKN5N/Wj4ULNlT
ye7xoeZR9aO1skv9VufhNXtZIBQ/PclTONzxQ5NiqTOhTNrp2vaRVCBTry1WXWKhmw4wc5ue+59E
fuT+jImYH3Z1kN8YetIVblDithTE7bkgQ4f+Nwts7FH6QJ+BZLwOpyE7zVCGlluK7uKlxQ/5nGgF
XkCjn7I+owzfWo7KXZhcLdkuovxOQLO1bR4TqJxDyMudx+EG4qDVjoSK433ihpuEzUgvJQf5Krp6
196hPLP0cGiYVTzo3ASk8uNhwdO8v25oJkPKsfwfJseecxktWFW/3PlVR9Id2YmKXwd55GkZP76+
XOSB1XtONK5mSkz+MboW+0O1Lm6juFpiscq6dLUsXCokWmng+lOgB8xhf3WrFsLLzO3PNIebwoN/
xHD8eWes0wBDBVaqBSKJ82u+N0UXlNCoIVvPwP1YFB5F4rbU5yLMTYjOrjrVLMhWiE3xWdzO5XQ7
nmxEtfq7BmQbT5G3J0A2Bs/bf+VLVHvJUa++KgUuVs2A9F3q2n0uTveudfW/LxS7XP8yMlHQxiOS
NnrfPEagTbLF5i8zeVvIc3kO9Li7RU4c8QMppbKlZ6lQ8qugg7N8RHyUFf+j94pGu4ggklizxgbR
F+ydUjCLM8UTwxHKD8aVa4S+1/ySEPl201e2bCKuN0BxXVoAVGD0sh0wIG/m7RznkeipZ8MQxr1L
8pkNhb01hZNfhC4ehCfSXX8hanDlMTScUJGsAXPRTgBWAvzbtzdo53nzHU1yhwbGVuIxULBwadaa
d09+YjH2HKOpO+phPpObQ52wwt9SHyzmtkQi5GJjFXv/FaaXK/OKE7CtZYUmjj4e3lVkPcddP99k
RuxLPKH6xIl9rzRdUWiuycQeupQJ8CY+MAf1/kcvqgP5zha2jAWOI7+ExZiH0UOJi3BtwRm9D0ZV
K3bDdHkUh1yclm2geXRGF/1i+q+f8SL95RoL025ag8ifl5nrXyG1+lb4cu9Ru8xBPoL/Hms98yqd
GDtrzDttuZFPqdaJw/y9jgcriUcC+72pohucZkIU9j4H6/RjHPrM5JGt+yY4/Qb8g3zGMQyNimYL
SGu2ID2vPygcGC9eum1qiFKBXPUkx2pGpbQbj9Dm8GWLxFQ7uC/yVsbEzDw/YHibvbPdy8wO8cNI
jTl6Xkuq8vk7tlkhwuZSU1cjuPc4TVHuIB3s4VGVnX3pUSwDqW41OJAXSq/RxAjWZJtx6VhWRqNw
0hAYuVB9/dZsiSqm3zwSmV95SoLo1Lnmp+lXwS2OnNTtI9nBErE28FS9sPgu96TjjnRN8Yw9Tc95
ILr7x5nQJYe3xl+/2QQtdTQr2gxWpfIhGSKWz2lrsAt/23syWu4v1i5Ti45qXbxDObw19glOpneq
zbmJlu+pyysxg9+LFglEaLcxB7zmOH54FZv/eYwntWT7QBS+bCDT3TYgdZlH4ttN1mls+Nij8+8a
VA2mlveaZ3vmup6TE0bDqicX1ntDGq/pkbLbGZIuMbKlW0tDACd5e/nMOLRecIN/mwY6GvO7KKU0
YV7X2GqYcz5SAy/2ecvXvdVlRLlRMZ97agXNtKt6aFUIqlkl2mvVg86mwVsnlrz+wDe2+a9N1513
e+0PkrDsZ/IjvV8uNevgI9lMp9X8adHbmSa9niKPkg/8mP7VlEqnwGzVEbD4cPVdBD/OkpdCfklu
VDx8TPaCdLNCjuhKsJ68Vac5m5EjK1UKUdE/zAAI0bp15uIaAJALzQiddi2JV3b4agX8I1QLu9dY
+9wGzUZmVpKv/6RPe+jHqPG4aDyQza1Fqjwegl2g+GrmFT2hU91jqyNAPfnCZk69Le0MhHIBNFYc
JMrH7NcehX6D3ehRRWhTDkHCnka4zMNB70CCLIJw5jVRvjYGi6XtbqXA9VV6HAtE2wK1k/geRdEs
Bb9d2p+licWuR88sqStkRm1FJXcqVQr6AgCMJ4eD7E52ZsMk2bSqZP/6DCafUjpDakgBWE1pu39w
xTEhZo2Szw6nMPkaJHsw2xLmYH6sbZ0zPZZwuMhQTSa7ZgK27DRisMv6E+U/jojClFBRy/QurLM+
nYyEm7KEf2+dZxMD8PrcQP55Wefd97wuC4bOgnzvXZAOpPqBGGLoAPy9Lx4ZQ3dfl624THOP7m1k
w5u9T2iwio3yrQJxmksAj/Xshy5Fs6LOBcMI9FdP457+PxuZ2hCbHkLlIo0uBMlWRZ/17Ddlfkva
Yy+ZYS4SKtaICOenAmmbGp9rzD1n7el7Kocc7Q9/FsOdyh9TfCOItYF5i8ot79aYUIWCmiyCkFPI
eBoEmcrsEhMGGUR0WRnkiGyKnmmtA4jaFoqwFYRzJaNFlKUK4cIz7M+NLwwJS4040j9RapHSb9fl
WMHYbBre11hQChfIbxDjdQmcm7f61FcOUyR5FEZEe3QqyMqquxqCwdSw1no3/GkxFITQ3SVanXI2
N9EWX7ywltZ1xkLbB/P0iw6KOFuQI8znJJ+2AuGb73627NditlUESbc29DyWb7ASIJ6gpUu+dhan
OrGcceSZ/3VuWpAd/BRPrw1gVgXxBKoAuuJVvTWMixed7ndeOA+UPvQGFQiE/OOW3DqikRkJwkT7
EfzRQyAUTLuTSpBpOdWkWa4C93GmXjuUN1O5d1+bUgJ24zXDs64y5TLGFGl0KtmduphUd61qO4Xo
+Q+j3yWyRFmC0Z6HVe7Ig4b/ICLfeSojJPbWGgj/BsHdZToYZXmU5EMeeb6tP4G2/nq0NvbpIaf+
9WnTytNsjyif85fLSUxdxcDnAwesVrgQgc+LuKQFHYw0YmQpaCxJBlNoMV2Mtp8s7qFhrP8Q8pV1
L2Rf6KPu9BXztNpzSa17KoOIrl05XKQQaDyxa5nCXeHHDgweX467EBfc7hU/jownzce6TzXJl3TE
QmB2Nt7GnutTP3JRIRLmBpJpzlJNZT44GbZudYlxH/9kHm286Pjr/NA9/Rr+TMpNROuf5cCgRmjq
UijM6TdIDFoEjIRxu2P27DZAti8UzEFRSC3DQj//X4NGp1LbbH+QVlDcWuqlI+nPCOfzFoEaiGGE
Z3Tqt+CdxIyn7vVG9uMkNDK7uMjwPQSc0yJIgU+MayE7k8BFFfMULg016Bz7PswI4xViJ5UPfD70
QgJcfDNUASDktGogLNNnRVVSojErsHb9Yt0P4dc6TvA6n6YnrPgh9EnHAkTRwFqnW2ZffviWXdB/
HrQ2QDY0DkRTan/q5iZRVq1+yX45kCS5+Fr78Rsg/HqHugGR5u0AAzkjZKnekuo/cyG7I14kv4GA
qKTDOtnJP+Vq5g8VbT/SDlQ85Pi1MZnV6sikKZIBEJkzpDrm6SMr/QEZ/q8oFihmy8n2SlmdWwBq
hQeqVKgKaNXzDYMCsHDnV9QiVGANRJjVs5gP+TX2io3ugGJnxqKIjfE9StPCNWOFrXU2w9GlHoJp
TrY6cmiU3Uz050fQdsQQoyPHazQb5T7Kf/96NbtoXrEq/8vBKo9T7vmN5SJWH9btKNYVMXiQpJx4
wWtRTVL22a6LscUy+1hTOvcXx/OWnHBz6eIS6V46LU68xvv8pRZwxEYtPtwvk1mOQILLzn8p7KSk
wYrYZlStiKbuXBxUfXo4MIy2PTQFZVXeat2z21zws72W/Jxdp7OfurVsEZ9V0J2hRV3KCwqv8fVE
iRPfv3eIbc4/9Acfa4lHcckmdNLbiB3VKwVwU7NCfRyINiuDjTRG1+UrxjgYgXEow7PtkGVzea2I
yxxWz4NuAc/8rCUAQ73ndFYwMrByXxMIdSzfQVzrYwNrKD1OViLQ5TenIQMk11D5EZJWdDi9IpNd
W7jU7GIOtZ9ksNPTPy5nSj5uh+9Cob7fIkunrM8M36h0mquQRuz52BEfjte5Rx/JUnFExfvQjMDn
Sm1U70YoWeo0v2AcmnnMZEeRdfmanUsoDFvj+YeNGGehqY1ecc9SNl7nBqstwwDN7d/mVftcrt3Z
7WKQnNxho2/OxfsKUw+lo/1Fbnu1jQERFQ9Suvnf/eo+CVo8L9DalT8OPRpORT5crofoW8fWMYMN
DxNfB3pYZBUlqos5+10APThUQ0efDU5IqgUWEHfMaU37+Yi8OLqhlPm9DnE0XD73XXyVuRoPLzrR
PZQcxq1O0qd2ixtShn2xvVEl2FSK6+WB9UaBIWH5SJOT+3J96g4+aQTb4Egf0X3RXkJ5awaBREaw
V+M42Ce6zQtngtt+cqkGzPpTICbeJVUIEYt/TKkKINV4/p/2LPRzPrsp8cAn25tiU6/QOJmnMkwO
gfibx4Sp492HZolgXP0JIpVtiiWMZgPzgXftDqg=
`protect end_protected
