-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fjUAjEfq2GkDtxrfXRRV7uUhhgVzgtv1Frg4jvqxWw+f2T+ClkJgizQ++UMnn8ym
JQXMqgDLA4N07NG2RlZn7bt3UI9xSRWvUNWQIRlZcXRvb0EVCLB2pNg0n/wQZQw8
DlOQLuBHrFVTMbqA2yzQ9pp/ZE07uEU7odiAk3Xc5Ck=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 5975)

`protect DATA_BLOCK
sbGQKXMZ4uo1aJg8n6gIZXN43H8t1H03rYFh1eiEa0c7QRWiZxIulfnwaH0Xo/d2
bM30+abW94Y6YliHDLIqOFYYHtXBS5NaI5yOne88/K8KRhJtib5yxdRGa+E8LV98
iBrkfBFN7CFzabLdF1FzWjY3+rb/D8Mnd9uD98FF3bUPh9SD9cv/tfz/3uVWoXZr
WpWC9vIPiXHP6m7ra6nZpRH2lXymvEDzgwHnx/kSs8e5RZ5eco2bHZL2LZsr4A5T
5UBw0ZBsZOLlOAJgTcHiPUOAyhikHfkmnDKw3xWRdgIhRdg5ZMqjitLMmmI4MPma
yzBwZHA2OBaMw964AthTCm56XNulYvboQ/fYEiYMSB+QhoRFx/mIY/3JAiPLjgJz
0sQNZPyJUy71Yx2W5uxxQMgRgBjvAbLuET+skOoTh8u1jM5GL72954s8W//xtxWG
cKWhcx/nxnPqtUm5jkRk92Yl37a0Sok8YB7QMq2zo3Wiv0VGXOXqIEXkthlLcN3X
tnpKO8hYd4SfrJYasstzSZLd11ffxiNMAIfN14O4a8Ohz+8OAuDd81Cd/9wWPmHp
FOo5qKWAUQ4V5Px9v7A2FtAlK50nag020eNZF5xEe59a71pTz0UU27bwskiBR1L0
QcVDoLiGKJWn+BBJkd69SYvrna7E2wS/1/tE2mFgw89IVuWNrRe3/2AyDOmAg9r/
lmqUcMjHPk7cBoIaDiL1QSZIQ/cfOLwPWJmyJ/UqeT8UjBE8C+JLvI6LZI+Mx5VP
h5NKCG8hJmxIfhhzC7LvYdqq59QrUXPwcXPEbnRxtAfSytVH1s5S9DgolRQ+DH1E
ztQRy4ECwNq4vU9PnGkbHDZJy+eKoWTL32DKCh5pwGVUAYdj3wzIe4/HJ/NCVw8j
ylIEFVH6Dfbuymnc9/Lm7/25DA+k522iToiMKMtNtN4ZwMEm+o6dxa2GTWwZOJ/E
UyXmLXRjkNShB9mBrsJyy9BvmUQ6tig3tfciwopLZcXid9e3KY6JecZExrmV5zIS
QpIsPn9fMBxHq6doq85iGn8t4rwW2ajxDTZIJkvuyBDuMQ787pW1MnF5RiF6ILWl
Oi5tX69WbXd9yedq8IS6WmIH8gxK8Cyn2Wx8bkGff3o1ebTkJPhzMA1LFVG9Tj3c
TQchuykRIjV8Akk+uTNX7Tq1qRp3rwx3pBNn6DLJZLd/vgUv+NIk0IAQrXrggJhl
X+CeZJG8IpQ4+46bL8de+T6LStEY5eT6bTLf8wcinDNOyTcpvQUj/Dq6KIYoNtQp
NRJ6gy7O2/yccrx/k11yTfieq492hQkkS8c9hTEboHfmOFVZgKNPdiwDyLwDbTwV
x3D+BGdfFmkmKmD+nmpGm95H+gel1JwY8yq5uWuu6TkpnOlHbCcL/3HlH/YMvGBM
6bGoS8JRXo6n88fJk8BWY8MSpMhceAgtHwvUhLWWDWSzeOBtZZuAkBBHYrvQagf5
3p74rvbPdmFIn9AorxITBWqsQswZh+/uj0lcb01VyzO69JxqQy3yYRJz2OCDUzkU
ieJ2Fbb9reQ12k8acRKk547khLOjOMhbEPQaoqWy258xSJlu0V088CIQvQTfs8kA
H0yX0RFSvWdM2ba7AAD/DJX8z9SO9NXBpZeOCNQF8bj//uWNwDaHgiQedJcNoYKb
+7QpG6VYeMyG4fVKBs0uQdsN0UogIjHTy9z2zsYOCSErr7R1Q6eDdJyXEqMVTtnE
gwwT+Q3YFbHPw0IhlOx2SWNvrTC4G9IVdLeEja76M4kMsQcG8JdXdHUqqmnMu9OH
abq8seVGOsBkCh0kJbhNMB5+Yicx3FiBywe357eD8BrBzcSmCau0V1VyKIq87Fex
X5vMoNUDYycFFNLuaADx9HBFtEbCo8EP7tDSIzjrm0t9a+kyGQ9LosE0h6HICxhY
oNGKOaG7SRH5aVC6aSaugwzesESnqUhKYKBpCPPc7gi8KqX+zWX8w6XePCY7Im5q
dq8f8IQSHfpu/LM8tSg8j006I4RlQ8w4nruZ1RsCZVd08RNLzdBQf8X8pKjiVVBa
1j2prWbWn1iiUOotmxIjhPY4EjA+Zv+08tfJZUuy5fZoA97vtonfDEodIf7XUM9p
/SDo6jRUWRuLj0LA8Ga1SKvJd9SrogBtktTUHgY7KsJS2vELGZVsKzPQDS8ekcor
ZNbKYRvp9CTN1Wy34F3RlJRzuuJTJVlmjKUWUl8aFA3iWKPb9q6CSyYCq1YcV3YK
Y36YciHLWM+gP86MPxI1JLznddkGao5v0tKZ3GnhvXA57nZxFuzTEprCU8OmAZsK
ULEiSIMEoLdrYG3PutZ4oTymgLAmsoMHUxjfd7/vw97LHYIa+NMHwnTcDjuOcl+k
5k2kul/li56NBeAYEVsEDRcM8RuBCTP28znmBNGezW8lP/MggNROX9ONMOaoLvqs
D988l5r+PyDDv1whEkdkWR/b2A+1ZliwOSXcJ2bBPifwzij+VcLSIUm3ROwA4Aua
J9DUc9Pmi9W/ei7rKO8NN29KZuZF5w4f2kFd3HbV8tB1byS+FgMg/GPxy8VcDrTJ
Vmr6Rjf/6pj/iXhyQQX9DQ1q/ifKy3kWB5b4+4SHtPkvo06mdwT4TN7O2JfN9+JC
F4ju2/R2W5KeHNg74AOysDXMTjf1dNv/n6jMPhBBWyfWPIA/dk6Wh5N1KkmYGG80
J8I23FJ/oYIGmk4oBpVq7fV37GYLPqfsZMqve5Fx9ecJ6HdLWlcOGAq8dAYpItEj
vhqQ7abjqTWP8w1W7Y//4LnQ/CGQTtmjlqjDkInfEEZfoIKlot36q+xki5aoQE2l
jUS9CDsfGOi2qJ3FK2DNnGO7xs8mEdDXTtmeBqUwa/dYeFjd9fEi6O8hwiIaP+0/
MwZjshjug0/2b+dV7vLm2RunvROBTCXliczNBWU+65ICtKV/hbGma3vI7bohVOG8
5OVkEq+OXOyacLm2IsCd5KJgGZ9RgEL8viARUPqDUPlKALSwA+L0XuNbt6Nu0gGq
nSg/NSr8COR8WwGyiDAdd43x/RyivrlxUh4bCtfIr5Rg6Ynme9u44bXPASG9i/17
QHxr978Z7EA5skCxPsICebZvMfBIU1aDAwP05ZWKOriueo6ljjbQGA8Gt5gsypaU
p9kDfkYMJk8HHOAv5uh9C1anrbQ/uWZQNd0g1P0F5Ei0UbjWPeu1ksUZexwvnQlV
pVhyKOzZzg6id5v/AX3+2RIc19MT94vubkYSTZ0SIDqsIQvLaaI0EiNmvkAJDK/i
vSRqqFLd/ntep5OohBAcSdPUrv4FoGeFE9hNIxfu17mBqqN7IcCfeOJ+K8K5QZE4
FDlO/XFAoLio53oONBDnBInl2+dfoxLqaYDRfBA8JzbVZEOnJXxDXUe8VhKXT4au
8xyZSXrt8WVyGPSvlm9OjYEkaqBcA5vZmNgHM1SyObXEiKUQQIOIZhntfCWFHyrZ
7tGrQytHEEc8IcbQblgpbCKgahyqovjLRr7xrkuPIAnODazI0prUAgVlArbLdTkI
hME2LV0cKeIX7Qksl/TNwwV6s3YQ3Y56dhT0Lb6/TQ8JonyFRtnuv/rcM0dq1gu6
RhKEjreO6rFvU4EONB2C2yA8lnPufSazxPEmjUKSw9B/cEAA5xVnbgYzB+YpPhAi
LXvJGa5H8YRC1Xliehz9HajH2ToZ2yYgwy5a26rerhoH/nScxBcOVTMIMOz3l5Jr
1b6z6xgryycyGQHWXivHCfg19wSrvcsczKGBA6pmsANkZDoO0VLX5poT2eysUExY
Z06wPuW3Oni6EnrjulW2UfeBY/8zQtRQ3KVJ5K6CoLZcPnI+mr9qYcNMqSY0yfvK
1aMnKCKS+SeXKkB1Eo1Z594nL7SotM9tizdV3HgGfvWCyCaBp4ONH0Qy8oVRMeIf
Kn2TIX2vHUwEA89v1U/qcWubWjUXM7HBfvq611vxNzwWllEOAvlvANNw4BiaOOTy
+yCi44j1SkkK4P+Z+LoGrZ5sqF2f+h0sRUC/AVP+tl9u8IiRk64Xo5VcWafVQ23X
R44J4CaafLgL9PxaMearCa4pqYsOFUGl6uWzihXReIuNXl2lnDhNJfrzlnd+Fq/e
/e8mj/H+M9t5ndFNA4Mi69tnVBUHARBLXc8aj3oNqp7XrSV/AW0DyehaVX2APd1S
nAcOHbCfjsx3FHoKxMNLtnAhDk/gYO45a+nZbmvENEFxhiQ3ToX081I+lBuXLixg
cPNNrhMx9fda8WfjsnIfg155THm8Ah5cUj1QzohJbvL9yaIqyUlhtHgqHi5j9xO7
9XvePa38ogltt1nhLv9XEUNOrvJP/OnXY6Hwfy71iqaNNvjt8pnlcFklylwU/aKp
JGG09V2WZp3641LCErUwRcJQ3JNBUzymirwLyTW+tGk0XcDxC9Q/cI8VGXq70GDT
VoYtptR7aic3pGPfwqZjHSbezP4llqIxzfqhvxhtMy/twDqaoSPwgOdFz+DZKg52
N/QTL7JBCXddLK8ocilodkVe1wK4uRQVruIjMLTTOerQ909jCMYaVlgicXII00YR
b9rYK3/D3INdWDP3cU8iSzEPCJKBF+vTpdF0urd5K/1RX7U0ZQZEsfEc3nBa6wKY
98snmoXYfo8PoPNnepTSXy33tMZ/noHc6kBOCyK1yaGtoR4SQq9quHiEtzDQ6tuX
wcUW7jeNbBk5CTCEdPIfAH+1xHZwNBIFaSngvgwS5XQGcCQ8gikaN2ZfDbGTNraf
cxBuUCeFIIfaKorExc7sNU957UBDq+UGXS5ail8XKCZb0SuDOlUmmdiHEN0LE1P/
8LriqZv5NvQl9fInFLSgSb4W0flCPn0OObp0c5+97whlTenrFR/fVzv9MyBcxg48
3Wtjt1oAMeWUtHQPpnEzTQU0bkJPSGxIcT0VK3QdwP22pLdWd3uEaUxOmzRgEBdu
IbNjVKyCAwjF2iEAaUMbZrH+1LLZmpWPCJdKU9zbepTj1b7nN9Oh3HSu/dp32mGV
gbyCwk3BC537JxxOwjW1uUBjEdanGZtkWJPgDreuTM69RjlL90Z4sg4B4unpK6tf
g7qox/YmMkAcgryNbxOWiYSmPlrWOvRmJTALWPI3dfADhLTDhVXO3QxBnBrXrA/H
xREo3xr/gVEQOHzbIkuDSL01P/ZFqQFswl26pnK1nMVPkzaj1k8yjkf2/wL14WL+
FIpxqDEGDL9RUbok60lwsvUD85FSpE6b+BdlDUXW7hGmdgfGPEY60o3RJ5nEYtqU
xGEJ46g9kd15snh4fdL1aREZA5/NfjlOlHacL4bmX+jLEoZIxOlinR5M9Z0EpRBk
cXBMVilDguDdWDpiRXkggzgxWXXOSEQRxh+Hr/19ZtqVap2iy0i63V1AoCyEOl+7
ky6OuQvnQQAOiSgpV3q+96x64BWXYMJOKPfUz5YHyqtQCuj16/HBkcBjp8z/h18o
7ukUtaue28hlUFYKClq6P0e0/cFH+/xlUxIP5GQ2u7IM2ab0B+TDNzrT2SPVF0nI
Q9aoZzs8pb5lMh8wK3QLH2ofAShBwQh+/mLmdY8+7J79o1hgDNP1PsslRlNMKCmn
h3OKKqE/AtLHJJTZT3gS409SqGPb6hzp2EMZV+bNDe2jzsf3L8FyjugPows1loy1
VO3yGzoQdQX9/QrNIeVhQw2iwxX1rainhJatuTc49PdIIhtnGO/p1Br7O3PVcYNK
9AKSbYuclw3m1uHI4UnWdgNaFPhkulv6VetXM3hrFn72YUM8giH2FcuyO0Ew57ED
7+Y7PmzkxAyNXLB6kQran2VPJrlXoBSapNT2IHWRWLsyAGf65Vrg/A3tzOTjeJPh
OVo8y65xdzMM6M4Y2SW0Iw+pgMUsFm41KRHL1N6jqn9LATUiRIzTC4/bEFC01DSh
BzYlEpjqH4+eHL0RGGtfRpeQw/qveqIZPX5oePgw8M6PVVlMLRm234JNY2ggH6LQ
6NwX7YS/cNU+4jK/SJa2E6v5wl54oWLPOL/I99nxmOHL7VqKh7nArpoJXoDpjHKe
MdhX6ZXkLXCUMZyILdS9TcjOZycaX1BQVNrChpab+E7Egbxf3wWc3Wvl6wNxeogf
HwzCuR7E2p7rzuyApBdIHu2mhSNZVgUFNM2Cv2C+PA8VgG8bP4BRUILXWL+MVu3X
f9G/S2e7zXeLxXcR9aji6Xl8qlnmqJRlC0Q4klpA+HCwFq3wFmPvBIIJVpjRhLlY
danzDqYSxLyf6P7aoBLMJIOUTlU7ShoZX16pip5HQ1NMKaqvbVvPdP7rUsye7QoJ
vxck2vGkWM8573b2nIvm8pFv/S7erkneEzRPgM7MOJDii/lz6/d0gR7cIJf6/wHg
CRODd2U4WuXusOBkFUQJHXslCH7k3eInxrOZ/ThFdIvNHlLdHysj4T6eRJQ08zXh
0jDe4r+CiOzsY96HuuEIxj8CorYk+3KvLUw7zab89EfAKrs4s4A5GU5MBEx6sO11
pLle03Ews6LLic09KbnKret0YkJZKkwQNC/SXFANiMYCZeHkGD9pn9jsh9hdeAMU
YhwmlrSAHHSRmLRE8PZGmqGEFqkjorOIfrAbmWle/PZbvyfaMuDKExb116GCCXDe
4LQk8Errshe9Q6I/QRPuhrn+eWk/2KJA7WBtobufoXv0ndGogrDaPhszUSkjpvd7
9/64MF1zc7W6x7TsHZXTBdUIOtHuiV5oeMEM3lme8p4JYQxWLkLCVaoNa1aft3uu
pC4sfGsUaj0WeMGJLj1q0PkUwGxe+Qit/DvhkpNAzjKtVI7ZwTBgwvYlLFDqNNsE
YMjaflNb1tGonYV8b6jhx7H7GDy7cB64OowSLmr6QpLyJWxB118N6VT4wWhPKsVI
sqvIptCdkcJrnYHep1xUBDeatEshTQG6YLRqjxSZdbXmnihKRb0MukNvRPhFBH36
6LD44rZ3slILRkRkg4UcNr5zPoojIVADwaQHs79sA7lRo5ljqUazVWdQcwphcvHT
WWZOmtz22pevTzOpjKMAuBZPOoM3gSWFONHADaT0aXEIA6NwcYsNQgAGG/ieBi+6
zWNTcsCKu1haC8uvJHf9jTFo88hEeLo3GYG1p3BcjJBuOZiHz10NaKpdo+S8Uz7M
f5V56Zuftn8Rex8IYwoNAP1iOCGd3y71xESjCAA32ifYRUi/7lp4bkz/4jH0TlRf
pJRkcOiYLoHWzbT8EQsxJG4rS1X8ikFvbYUFxwqdFau+RAzlsDFVeOFxbwXsjgka
0fbhZGv00ASR/kWGuhi2byCAyZrzzdBdgwTpEsHux5qQRIomqXyXbVt6EzpqLSl4
KP640M1tbNQNbM5gcICBJ8HpJU2YeJ/FkGZHvoETx+b3kNzU0+QYOwQr7C9GDjn1
ZCzKDvFvH7BWZz4FZG/kvr98d1grdAT5NT4LYHf9zaq36ZPNIYI9E9XQX16IS4RK
i45h2dLYPyOozzAPavhlHau8ptdZAa+mdBrfABq1GBRiUf9TJSVrzkM13RKHZR6o
4i7eJ2eKTEVjq30UDldU6lbK5/jALSkIkpkFDCQxN80MbudciWpJ+71P/GAF31la
ZA46OV6avORRYdkDr6Rh2fVejtYilNlJdDV+D2ULvDcE6aFRgGHD697UMuQK918x
8Khf0+vL+m/PTfIprNI0Kdxk0+xuF7fH1tIkBRWLnJXEw4248TA1rcQ8t+xd1x5P
9TNuakhhVVggV2iEDfh5GmZhP51aRxy3+0GsQG3iZyWhRDBO4ZN57Lhr4PsSwMI4
Lb9s07Ija+XkGGxZcoucFiXrRQIq0oEMFZ/0zeXQEjyJb3bAi+sUupVcYtlZF6hm
QXsONzj0UMFzxkFijFDdwOkjnY3fm2V7wq8+ft4kyYfktz7dBVoGeVTkSFbn1fHF
BWP/WRx35/UkeX0yl/ZhqIFmzMDQboMgKT3eaEchNtGxGBcQPA+jCfmUTh15DhHj
jOOBaqKHBW7QCfYXxeVYM7b8uTgXznmugGlD+4LaFUHJeNO5RKj8h+1uqIZt/GN1
`protect END_PROTECTED