-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
eHILAe+wFmrEflXm2YfGJ0ytYVLgabOsxjXWBnEyhhNmeU2LLZlV0jef4Z9Rr46Z
DCJDK+FAa1cySaUMuSudf+bQ6vh6XdPRwee9QPiWuAK0s5h/+ZG9SiQZrJS8kPRT
2G9+MzIklE1avjJqcTTPK9cZD14u4T5bCyUwo04O4Og=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 5184)
`protect data_block
0O0aHQH5ItPI/x1v5XETji5aVAxR+Hjz7sA62MpOIDIgEZAgwOTXvVbIuKm5BlpW
9MdBhovnvwsYuWL5ZuoLeRuQuqHjUUxspRZnye/K5s8/YX/3gPGerXDfun+tG87Z
QUF2DELjNDJbKiuotPFWxEEyFyLnkmpd2DFGAjocuphk1oYQAjtZ1geoUamn147T
YSU3zZ/GngkVUiPOaVyr5Zu1rGFPUQVKxVs5e+iOK3hETQE6UQtOV/Q+KvF1J+1b
OaO6MRiic4dsAdFGBy0e//V7W7z88NLIjUHOpnxockrfwBmhdb+zKBVsSIeRVN6C
20Nq/8GFFOvrrITk5unPdpUhmNCRLCay9AY51fLwOxbzy40q2v+4hi8uIpnQMLwW
PPEeDHdUOmeOfhzflMJ6BH5USc/rIMm4iVT0+fzwZDzGp0c0gO4EZlZ2nJpcQzFI
05JEJDCz27/3VuRQ9K3Uqhijm+2bJnMaOZVD7UTdNA+NXBRiut6z5wefyyN/u/aV
d1bYgmPxT1hiobRkENbrIDkGodZ8PciL1tncOv+8YIsPKxDcVpUt6tUfpmGGnN1u
zFwsesHaePOl1gD2vzDO7t63xQRyZpCgY3EYWfEcXO5HteHgL7YZHkJGbBf3JMGs
44ozkE95rizrVhLDTwFB82p53JifslkQfHA2HoRAp7/SbrycaQ9Qypgo2avzYw9y
T0lt4MXe2hHfUFkzPOT6EsM9iUJjpCzMTY7oT0Pfhnqsed2CXo4Tj5DPyRrwdwNE
UCpHAGKJYL7lLvhE7NTEzmac02pRhaIKVfnSzyRUtPbNOOjN/riEe0oPzzsvkISA
2f+2QkLscYtYEBmsb/9M0gOp/d7dtuMCkiNYfSNALGHFK9kcVmtg5l+cIBvThDqk
X1UehB5wwtaM2B23+X2SbfASU2PmksemuGwLrEdIcRjIcX7YojmGfCKu+6ByjOxQ
EzDEljQoy+6A/HVGAeifAKchsGB9kFxuU1ae9fmrlH8sq1JZ5pDEpfs2/U4logIs
ZLWxNvFqTwZFSmQ39axG9Ohw55YAfwnH139N6c+hKulkPAJRWoy1bYjoKmoF6YYN
Dce3ujfyL66fQFvcXnkLae0K1tW3fD03Glni2BRT7WIwD8DuFa1p02K6DIDvfpB6
tTLXrPhGHE7Bm75DDx+lftyXyc5MhSuTKWT1iUwHxZ+eubVPNXYYVR4y6bBefh2P
SpIozo01k+hkbM5v6ZHNkApkqyIHqxIiP+YYVIMi+CU3Ze3FdzvZbIBHCDWooYfy
E6WsHGTRFXw67XWhAF18d8qtBLnsswQ2Fvs1XRT/d1E2Dn+aKLCuLKwvT8YnY3i7
E8L5NY2zVjhzsIvMEtQTLYHxHGeCnlQ4rGUlAxzYaj+Fv4V0+04epFfFDD8CFSQn
hTXpQ249gVy66sg1GzY7xR3MYvE0zo/UtTzWQr1OpgFWyASBWYKNmpDQ8UipSISG
l9Bq8YnGhhBG4E8YyTo9OWLBVge7waUEqOjUn/qhQ0qLGga/a7E2YYMe+a9isbAn
onifODTwCxbbyRS1b6LDBHQlVxy6sAY2IsyA+h7VxB1hMaYi5yKM1EYHdDUOPTZZ
COD27Kkq3yUyUG+4HUFJPa7i/y9eV5JoSLiy0IUULLlNfWKfe3A9CFNQHG4XECD7
w0Ki632sAk2sSeCSqx0MIwBn1uf1zP8cOwiNBL8vtwiHBgmtmf5zvcTAkcLwOvus
VLJGByfwBQnol3CBaxTiA6xJFbqcupiihNm3zskdCDnP45kubOsvBdSvlYvRmc3J
N+lwhHx/fLxod0e5oDIh70v/VI/lIQh7gpApHubE+KK4zceMFGwscMQ/I9+AIr/s
qaeWc1UxZ4m44q6EwBQQNyrll7IpGu8rGJHagY/vUNOVWXoOgdJgm3QsAvWk6HQ7
TV1YfnVpwQkw3pnnfsUV4t/Ufepl/QV9lJRjRVCt9csbfopVOAh8hKgMChPytQqC
ajbGR4Sml2RYWVrXhwJaCidLDHzY0CXvpppypFp/EQ1+GuQ3s19lZ+H9piB03yLZ
EmG5rSD2rAgUQwMoDFUI2mMfP3JfGkRPkUKg+rpO5jrGHQ53tvajN/9JQGzW65cR
7sTRVxeTGhl5chwrykRw+tbmE5R93PpH1cTfk+cRdgFjKPNqFcJkTZ39a7iF9nHH
lj9a2lYXaVMzWdw26LM1/7vYpFZoxpdh7keniU6YXGI6CjY6Xv/uTWATHDwZGNNC
Un5vxkMBwOATrKeapqXqSIBDjV7g0T9UjtDthWLKCZO6DdRxFw4N/CE40k8jeeru
KCUNFpK0dt2eysFYQxRnFXwY+eHRT0X4M6PPw9C9HnXtg6oIK0Fo9uFH9zDrgfHV
r/xp6hPPLrR7QKVGXdu/Dtlx4K/PMBWm3LWS4KZLbnOia5opG6hJQU+V2icwM69w
C2u6dOtL9WooGAgCVuPoBOhSYDtcUk38WcByIJwDVlo7DgSL0CrlI5gsnqa1m6Qp
X0baqRCuFjMl6P3B4VtduUouxHEPS0ZRjcK1Ic+nM2tJbyINksfdd7c15bgbogRx
VYEhOD5LE9Czfb2fFoNu8irpKA7uNNjGle2Nykf/xpeSoK5yzcb2ORaFOwgMxrWF
cac29ZyOLhxmbF0nguHAo82nVoYW6LbQa4Jf3ogPqUdzU8xvNdNSacnkUlL42YeG
tIM2ui8tWgXa/Evp40slDAnkUQNaeZudiQPcfS+CeyEyNK8mrb7uCk6RiLuFZIIX
r6YKaoJAHOo5VtVJ0bqEIJfkU6x6UaDuE4xzzixuivJwn8ybtrmKxgR5Bt26JDiB
M2/6fx/PXuE6gmH5ytT690/m87hKOJObzD2oW64seeur/JrvgCiwzr+H/+C6pE5J
XrSYjJauVqXdnfi64ChHeYYSCb1Lb4J2HWUN94U7OtxpgZeEpOFk3MKl0WJf/j0E
uqUTFZWeP+r6pkoZNvYyXRf4xlwxUj6YHM/tdSmNtWTFx0+XYZ6xwVacv6lnPMjS
VYUIjnepEYENpXzu9+Ed+68nJeh93gp1YuCySbtY22kyvWqJYtDtqSykAjCMOydU
Qk7LN0EORjyvq+sB28BKORAj5E9I77CzRXKkDFVSgx534Lg7mMWebqjdqrnDTeQH
iTJtymMgTG9csxpGLSS6ff8465CswUulRAg25FgP5A7x8NfNmzcScm+ix7rkI2bo
Fiqvm1VKHSvFrEq71OMZ0p6mxT0G6tBUcdBT0ZMN1XjucZDSPncDdcCW8wxyCUES
C/AYwsXPeTibYQoYMzJ0MF94apo8S3xJ4sQJwJSZTV5Qb6RNylV7r0mFvR9BB3qY
GJq1HWfqPM61BVWOfYi9Vk8ZbOpwYBBR5BnZl2McgW6nKW5U2GFD5ewp+MMA4Z4B
ZwhGuLkKnb4frX6VHXe6VPfe5UsQN5flEQA1VkAqqzRsWf0+RVaedCh1rlA7t2HK
L1oe8nT6S0rv7osMPjvXnrZfTsyof9sfrKTdROEQpCrntPQhdnnKK7NLnkGlMD6K
xRHym48yWhe9jT0TrvjWO97RzhhGV85QKjhRACQv+Jwro6BmHO53Xi9sbU7qQB0k
S77SIJasOKeP3382bfYy7umFT2kRhSs4Wu6pJ0FafMgNs4Z+jcD71BimlyOAnU9V
QX5T8vz79GkmJTsSv5qpPY4h/zd/C13XiEgyOkm8hGucX9gN7GQuwEqFWojpwSBb
XqJVQqQDFquy8a6f5LSSTPzh0w+e8gbVIjFmElnoec4NChU3ubvTrAftfurVqqLE
tYs7KVnt6wVEQ0pylC0BP7wPJlS8Xzc/B76i1OvCgmsJ5+rRHivuLzyBMtVd+EDQ
BEqonK7C1q2hNna4/+3I9QIIEYta3+lg0Y7MIgWmcNsaZAl+ycaQ5/QBoffJ20eR
aDqUx0M1DvVelOh9eLhiR0HLVmoY5MKAEGUrH08FSdA1UE2roLAYvJ1+L/9/AZgC
pRYCnD12ryjr7ZqEJ6ZPH2e/tKbzV2AcugITR92LiEAVRJ8ePDxEyl2gH9Z6dnBf
4Eh/zRRdk227q+g/srpFkB9wkMlGAvVJ4D4CfnDbeUVM1v25Fgrv8E3e40RWfjX0
BteoM6tRzSklwupoJ9zAM4Moe3sjI59zesDqC5JuxxsIPcMQMSDp/fRCjc4jvz5D
9H7QySETXg4KjaJNYiOhgSZ8YTl3tfGabKGk5V8yuhPEp0QHM9DtmCyqp3iW8tgF
nrssLBDjn+0p3Q3NdlKbEOHc7tqpT6xrguavy18qbtrMheCoP1HdauvVmQkzTnQR
k9NYm8H4MPHRwSM0N85GSY7udPie4SrXQkUA1Kpx13C+rwgnOeD4JIzgB2IA9Jus
kJzMc7iejhDaKqzK/Bn85rwk13sNtki59G9OZl3XpfikRItlC/uGV4zsHyAyXB72
WgLlw1IyaDw0jXRZmmlToCrgXkKFXDXJDhUTPRgB8JI0mr1IPBEZDJnB0pG2nLC3
7uGFr17a0hVzXNJ/XMNBWddZ+TmvBssIOEDiLppWkJUC8lxsoFGZuCo4eeR+m9bb
0FIEZwi5LFicSVDdAM1a/95LMPIzb71N6bpuvM1wlTKFWAclN+/+HOTXtdInJE0C
stIHx0CxZCWm/WLh302xFjkXiPbz9zDeBhbJAlaZ0oi+O+SnxPh2A5drVEqEWT5y
cFGi1OoJbIQuza0LPR0N9odCjY+Fzgwtb9galYPWRdUcAKt1gL88Q4Z4onZMrcA0
zeoNqpvstr9zyoob+585nwQZjDTuyDzBFMfAAz4vZhrbN51Al2G+AbYHvKArM12r
dyOdYwL4mz3OdnYcUuFR8k8V41W+10+k/NzYvcR+QWMf3042XIJmYb6aUIJ1U3d1
w6STpO94asRIFh0zEEogf/c0tRfJpAZYek74WGBc52/jJy3D+F+QzUVlFLVfmmHW
lX9SJQ7FP+ueaDnPBcJMsw4D0YVYFtx9B30ED+tOhUxuXZIdV47zHfHUyoz/oYV9
jf0A28yNBm4OvvxNIs1Dd4ym5yiIptcdd/PBqioLhZCUuGoDZ0OY4Ay1HVIz+nsd
Qc2lw+mC2rSz+de6CKLrzZstplRm1QFMSYJOEoKkMbyRN0+6rcRcjeFLsMbhGVN1
vdRv5Mjx5AnKd12/OnmEFdEjViPW7clnQx1/VKHaCmiH940Gms2FRHL7OkMA3ElY
m2U/BZ8Pcs3LaKcy1bHQKGunbeuDfCbv4CBciDCsxc3wwOeXWNevodezofyBoL+1
VTXdm/O4tHt4zWnfjYNtGSjv8tdBt/Fi9w9mtRF+b6Q3r3JOVyfWUWfc1+zxEYQX
f7zXT8OqhbJ0TUHnaGhP/qP5qHftdR04I9MINb+jDnqvS41QrpMRBo+XaH+rGgRm
tHqh0vC4mYiiIjWE2Hq+XP70YqqJDP5i+H/1ZF9WQE1hgDlY4WOx1g8IV4y+tBnO
cGiKy4O5qEWDvPndFq+cYc3SqEKwioguH0HyP0q38g3ITcYK2+fsALL1qqrCuGlx
JrqxPheVgMi2NFf17Vb84KPUG+nJOLbvuDD1nhamBQc8WEKp0GJEX5/NBYhS+tt/
PIHpIWqCbrB0MAydeh/o+JvtNP8CQsRCYGQXDlsjrMgUfAL300f/G8Ker1tFF83u
vDsiIw0ITmVZJOC3RvwDEHK/+YMqxJMHGgq6HfoucSK851Ce1ERIaxBxOQCbGAFH
Zs8QsyoohHC5SIqqE/hS0GoId59uGPFuhkZCTt0Kkwhny/F+pdN/FT0EkZWCfyb4
S47I+tyDCxVP9n9WTW0Nrg86CtOWo/rpVnpox8WMdVLUmfz6usJ1KBdqS+jMwEZO
QrXmDTix5oticQE78uEU4aAiKLKpUWhAqHcY6MlWwBC6Z6nhESLgynD/J0/Xt6kJ
SeJtbHtas8pfZYY8yHklbvR3Bc047jT6BP2lOGj8aWOslf9ZpcTSYdIpTnhXHaIH
5Gudr/LIrhlX1s11Xr3n0GlURH1ghTuubs6Q6kKlD7GH9ge9Xmu/3lkztk6vbXuu
sW/AGhlZqs6HrlZqOensMLgdG0fJJtBSMd3o4QcXfyrSko8wqsh72XGdVMqUdk+9
iJX3/Sx/Pyogf1lgZnMwf84MhsElxF36dPptbxYMX33h1ml2gEUostULMX5p/YcY
hGJq3yr7tbpGGvqAzUDgQ+zUH3pnOe/C5/a4G5Gunxopk7L9xmtIc8HClJzcvbc+
5nxhC0E/YP1iRqFvERAyzwNd9/VPLtL8imEs2BiUx7tmU+X3TiHNfwaaOB+VvDZm
jbWlVVhfRoHmqpKmbN2D6Pfeim2jSGIOaXUFhSs+pY/KU4eikd6mijCMpkixUMNo
LBbFmwhjwXfouZW8bndLkK8Uls2xdjNiBF22PAV3c98S9OsrCPbPCSlKMsYPX9xv
Fb/7cjV4TWvwKNm7TArfBtSV3K7m3GSEA/Ma09LaWgNJ7+6hwaZKX43AXm0zWWEZ
5urIg/d1UFE7MI8e44iXMyPhuR2y5W+aU33GG8NNzL9tZVYJkSQRNWbAz/0Orxip
oQss70YOqw29Q2ExQVE5eArymKsFg5oqXhUFpN3UM3MlHQDQ9nGKuxYpRDAN76BR
PxxOCZ6qU5iehV0QuCnF/JJ6uD3qwAAbbDSe57WVD77vgYU7EQnWFLFXwTgrN2p5
mfAnlEsXfX4/7hFRFQKpYAKb0NrCqtO27TieOVWE/g899la4aTacARqc+bUNov4U
E7piCSjqzzR5Ezenn9OQ79/BoflRHNBQhRUr2llngoV7TlJevPcJAgUgzwZ3BPl9
Q/hn3a0rAzU14NVv9NJLw2Y+3DR+cJnCmVaZp4OZ6sKUm4NK/CtOUyPt/OS/wNex
4qYmN0spXVXjoO9N7rDMKXoymPL3w2WANdV8tkG/L0UoMqfUW+rcSPqkQeP99pBi
`protect end_protected
