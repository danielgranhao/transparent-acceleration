-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
Pp0OMP8i/7n3H3li5YeK1h9ceNUQn+p39EZBzkOJQoM1JVyXlxDNwqNvULpyh56k
YIMg+zNTJwDBQmCwB7s3JTuZ+6PzZgQo4cTTg0+o/DJp9MbPaIA0lfUcMl8+o9V/
aux1jxrRY1YcxWnR4zNg/gNHKNC2+jyRHywnfZHfjGbXo0o84ypLLg==
--pragma protect end_key_block
--pragma protect digest_block
s2mzap287nZh4t787eH6f8LtM3c=
--pragma protect end_digest_block
--pragma protect data_block
EYnhADumDrT6zQpZj1/XDO3D1KORwSfFA9ePF4kYIKw8vqFY4g8bH+dLn22dwRrg
IoNU3nr2X3cj2N2gCYM4WgA0mx61/qsOFt6E+0Q6w8SBQ0r14BqVmiV2FcNIouQ4
icoyLCNbEZ9DcQQAJr/jDBfCu9TQrrSdRgEInqSblRzm9UNcW4LdV5QT6kmSlYgh
8xAtSPvOQLKPuY2o/G3mRkAdV6rB2PA19oRbXBq0v83GQ9TB3kcyCEgnEu3419gR
0IME7r1apeombioWQDHVA8f8+rNl073PHBrtJvGqCv2/PSoGanDdIL3XtpgHyxUN
YVy8jpR7LlsQsM6gVTA7O8wAICdo1n5X///MQoXj06tEoduMxoaX1xfdHDTqgT0R
hanc0JF3I6p3LvzVoxUARE15rgSTy0ozlRXiw36xmFoD4lYtPv/UW9cFoaOysqIO
wwhCFH0Otqt6876ANpTNvqdKlxzZc8p1t3P+WXAN+xLiuexx2wAGRPOTx32BZ6AH
0vQPJdzHc/FFsJ4yWqfqzmORbt38axu6NBrEDSeyeEB78X/bsFXgWFzM7sMvUNKg
OhnPYqR/jcgxrSX62f3a4YuCAUCz666QPcRAjPE0Udi9+MIsHIwDV+jW3mX/gX3i
4MIIzexeBn0UPObeDmpaKCwv0zYybBcWWoX9Jw3uYrup6HAA8pbYZX2QiMM9fnZl
Gma+vhO8+aljfoc9Sa0iko7AlZjK5v7urpZwyZHbJiqfljhqMlKjm6weCIoOm2Pn
Vu640kft6jD8ckV3+STUoSxfsA8b0FvWgqewNpNnEMB4EqEqGnQyFkpNxzIzady5
GwH/QJAyP3Br3PGr+HMbCPKNcPuXD4AhGuMqxc8k5DepVEPSVmBktLpeNhtNOHyI
YIq13J5CVmBWjwyNZjC1x6tF+zrTwK1C3zWOvvRyQBHOuOfVmgr+8kWIGmp1TG1f
7bl6pulycto6H8YZSclL4sBTLBGthxoQyNRwVUDsnLUmxiPpqHzpVDllz5gppVTi
6oelGZvBE4XQ46St/zANPCJ4d7bSpy4p3vk6KPPsj5GcOHTQ4HPyJvQB9uVNdH5S
LBiV+PW1b/H1uNjQEw61TH9EWV/QBpu6U2ue29gfiDnXett5YosucFnfE5FNu+8X
PH6YiXd4+WnzxVhFo86W50MmNDoGn9bmkp/b2b7hlwygnA5AuBIV2BgB1g94Gq2S
uY7zWI2rx+vxV1KMGjBi4bVe4CpECRFArn2bpHfGma+WWTWjQumGXWfNIifM1e77
EVpThJWyPiCyFrVQtiw/2DaaYmY3DotUOk6IHm1YrjHmZcaRJD8w05lSVgVe40iL
H7e6FtB6+vc4fz/hhgp4czcS4S/38KvBDrX0z44G3oINw17PDlIWK/nP0u6InrKi
kFyIUiEgN+bUSUCy5sPKmBR+/CWmFwPAwUB2D44HHlrhJlvRva9iZarVS9QlUql3
fkn6c0IBjwtTYxn5y35aCyKJQ3kDyXs25qli9yxoj3rFC06Mq1GclZIY8oUQ+2AT
mIaqfE8Bg6S/s+BFijJN0Pok20pxHJQGifCFel/DH1Z+kuXLqIRIBtfYaIly7bf5
XJXsJmLvKZWtL9RzJ5YgPJlEu5n2V7gJGaJ6X+k5KWVtlXYnhRncNu0dbNkUx2Yb
wE/3rMOHhvCBbPEm5fEMBeI8SGcvsLVBl2OQV6cH15M6MLWwJkqF0G70h3r21j3s
wtCrfNmVke7gwvrsqkhGCoewediv4DznZf+sT7uvuYNtKjy2Ycw3lU9tWxv7HsKj
4Ov8PfVMMmcgQF1/lEWrs293ngb3L3kwhwIdKn/nEZxX0XL/Mz5zl8Mk9F7hz27d
e0pB43yX/b4aSl6Hqdh+v6vFr/DiF025qBCcMkEd+Y2VhCniK4ikMaANTZDhVqQW
sUB5obzGNjaht2zZSHu/j/ZnR9mrMn/Uu5wCUvXwp4AN6GnkncxO/Nt84MwZpc0B
m61ohPzl0crB9jSQ2mqAjk+A9qLn0H9YM/ZOEvEcRpdr7jGsPv9X4F2cB90y2Cca
wyhLShqBhrnEh5Jagqgt57GGT5CfC6WKdqBA71zkORa6AzVzAXYspeQzBM3zKqJC
Sh5EB1yjeuw8T4bxxMvGeWb9hDK+JlHviObmQNr7yj4w0Ix3NAE8paLVQtddYNl/
3b6XrRGjL0os6wYMMPc8PDP7CzCOPtIOAtNMfUGFhR6QbHOELyYlkz+XIkCR2w0q
QOiuYvwH/Dfioye+uwBNQEkyCNTxltGPSGc8X+1tYDbOorUTxfPzcFIUyl9Gl0fk
sFf621Y730vp65+AsuEmMafXjG9edSk3bU5EEzeZzBHAXvj6Fvvfo91O8E6DIO5u
yt0gZu1WN+1Bunw64/d47lC1UX+x32bvytlLmc3Pd5mlQ5WSQExVk+TfSWNeU0iX
F2Wttr8Asqoo8sRDYIDOrSA3Zl7gudpIX40NRzvXAnn37h1m3EA1ioJLE0uhJi0K
bt1i6Hd9jMH9h1N9g9rKVcxyGCehOSIwaMMvSx2QH7s0xmEF7Z212wrkq/MNGC/C
eLQ3wYayxUkZQyGZ4jzAAfLiBhF4+UUCSUmM7P88LOwOUlQSrvIjMD0xutCob2R9
Aat/4kGL6FfViuDXlTr4PYORx3dOXHTc3Q4Womn7WnVODr8AAfi1onJktmdl8p4c
fnxoWKC3yeSyWJ6GmwibjXw1TTqsv1S+Kw3gSOQXA6gNPVhI/y+cP3c/pS4ycILl
/wNqeASufYCgHNsGLaHht8nQpezg8fEPV+7R2QNcHf+YxGs41jfqa+D/xnSI/ycs
13RvnVHBnynuFtz7PgCnfAhCvYRTtHUk5M7EKmVZWfwv4PNSb0hGXzqPnpeMsALi
dM5m9hPN4aIlQWl9631RoQhFT3X4MFV4jipgYen6zyR3FNGBTDwdpzsThHvEeh21
k0bGiXSKlWvYjaE/jVjomNJ9IpdKZH23BUWN40pTiM72tEdKD/34M4qsNlU8WbJx
BvdWvT0VFFjwaWhWQqLXZPJeRB8+rmwiA6PPRZ9+vwaljGX5yO/h+d7dCKE3gbj1
XXueOD3rcb5BnJXoIDhAYDsycKowk6VRY7XY2QqZi33jNSsAuHlkIkcXicHfv3nt
6k3n7FgGCCBCc6yrrHC8+vxIE8GAOfoWnlnPt4Jell8mkSDZ19dtWv3DtsiJ0C/e
aizawD/POBB+GYpwTj0zrPSreF02CXGx2qZdwxIeSnHjCM2Y8RhrAtbi94sICMcD
siGQjYCbi+XqlYJsP1Rjj/ZO0YQUe95Bo4udvPmwjfjzDPdeuQNeU9fQ35tG7KzU
EMTv9vhpKNPcPPpXSJFSLdbb57jHK0IDiSjY9IeAm6IxMbqzgUMO7gryW4u/mzzx
esV89abnNwvNqMyTPtHsglCI/Vh7tLh/8hFhbDoeGv+wJ3vsd9kQoXi5XDNSyyvV
7EtaAopNRIvs9/brmLXbhhuYqgzEg/EpDY9LOxijoGXnBifDgyqIERmCsmM92u2L
7dL6CGfIj08ZSflT4DhtQgsw/HdLaKm9fe0jRkS5uvins/156iyPITXaFcfTs+t1
fJW/p+WWkaj9hz6AiB2+wDyd+4mr4E3vyHle3lC7GSBqUrPP/h22+CsdVsDrgvIP
LtOfer2WKm0wk10OkFxWFoLk6YvaVdFnlKQQ2SVhcF4RK7OF3ufpFtJP7Ni+ASEA
MCuubXDD9EgxzsmRyr0A39FwigkZYsXaxUPlXMq2PjPbwh+H2Bge0yOm7i4Zb1Gu
N+Ft45m+bsxH9UXjcaQQH7zNv9L0HqmHGXUV7DgY07+DEuXDewud2+EspMK0LCTa
xl893Gn3pIeDOXEvOuM89aZ6dwUKzlGkVjhPjr4xRITlkjO3pxxLXPhAxtrWlhpy
LWg3Lwz2PkKhKarLagueq3tn/9sSQQkuoBPJzL52LFii5PG1vB+az6HSkBBtiqKk
zcI8EYf8vWwYb89+w3ZJmS9QuLRuU7ePdw6T8oJzFHnTAco3DAxPtgGg0E7D8dlT
4dd4g1oZZeW+F4Al8TCKzTja3fUxCbCnnPjFmldc3wPkrsjUjo6NsZ8PcVZlktPI
ik3j5+U/MmE5V/JGgU/8ssOVRHg5bTHctucjQgxYVWMIjyMh1+N+5h3kkOUHvHlB
8yHgvB+DnNk++qo2J1p+ZVNiGRvFMNETZRipXWSnOYfT0cD0+0RHuUq511oAHOTF
NcF5DPxltyeql+2/2K77yB+X2jImEiArObz3Ug8ZyvM/zxlbO5A4LRSCr1kHf3km
A7SCQp0FV/0jYuGU11XRfKe23tR1fqvFA95eYX6eWGU47VZKrz2ZhjMNUB21o8/E
f3UwMA3kVi0s1qxcOI+wtaLpatzH4JozhSBLfe7AQ0BxNpWH8dnUB2eKJNu4+3HR
cOGWtrr+nT8cGelndXvaJ3oe5021eRXziAT3KuE7MBo9cGO1O6M2a4EBDgscAi4O
JhDM6mxiithlzpSbtgp17Yj3k/DwVh/0ZzZ7rsRv+ibGyXXb3f9aUTHLTHHe4TdL
/ekZdL6y20ESwrnTWfYTLjQ6F1JNLWTiFjCtyx8AzWlKuZ9WExGlsWUltKuS8e+I
hXgeIvCJH9mB5ZfbpZDwsyW1/tDEF0cRONVGDXXjQUn1Q6BTMzDlvaG9ygKjJj7Z
h4HmBHdYP5Ghsg0WxfYTihoXTULpdLGbIsN5AalV26Im1lpN4wd1Rwkqhn/skfSN
5Lg6FmV8htq3AgVslUkRq2Y7ye22uHOjuSaJE+LzQZ5VX6AyBujeLigBea/52iXH
vtvhwrDjhrcbI3KbB0A38djD2lZ7VbOHC2FSMq6Q9Bfkc0PUw2vD36lijdQCdOiI
HC+iyX1rcMeaSS737AG4c+Z/ujDtAtl4ZAbwtSbPOpuDXsyiaVfAsWhDQyOASsmr
MQlwpP+zDAsXPc8/3SrQgqYjMFOqGkoM/KN9JA4EuHTEctCC0nl4CwtOOEJMQhUC
eGubPGMjS8p+a84Yo/BpJaE8twmQQf0/8Ftj4niai3DPt0RP0EXCLVlonviPd7K2
D/Y35UrjDnDUdk78JfTDYlMUhB9k26adR4LGA0UK6+Zj2KcrlsgAt+vF0vwI7ggM
UJilJP4v4xhXhYXiawzr/cQklpNaVJD7J4CNvWFf2TG33i83rzcJQvbo8G3wUTJ7
3cwqeO/71xVDI1Zj6s0eJr8jsqTnhaM0d6TIUwjsgFPUVQiTTlw7H8Yoc/i0jpDt
5UQekMv+HCQ7CteQhPmcroFRyCjN3MTUk7FZHud8Q/A775cUAgUwPV3z2NKtPNN2
ve9+fvj8z6/HxNof0KpBsKyPBGppBhbHrO2d5Ek+dOA7Q++TPSlD4lTbKxMj4rTx
VqCb/2GAZj90TmtUvk8QngpJiSEC1FLe9fvt1KXgMf8HEGTzTMsLMV6pj8i2AeF6
fhPyr3FY5tylzd8v2+w5g2sBVctWLhXKv0ers4nmXbFAiWvZ6Ftx7xL/ADSls1vy
Tb0HFpQudylqIiT7wJGOLqJj0+aJ+LRa6anLKWt9o1x8HksS94UIXE8+jFFLIPO7
5BKByT19X+ORu+JyKnKTHCM4UhDbMvcH27ZeYJQhOKDuD7Biz+5Mshic3P8f2lr1
k/TAXQMzYbQokuQTTe3djyXz9N2NVHxjD55FEoFrvBIAlshn0WrG870LiDiKH3Pj
Re3u/tC8dXo6pL+3OG92K4eyVH2/FwmJNbWzERF8MPXslJSI6ij5UfIk0JBm7ecf
tfPYQgtMNImF9JxbWuu5NYiqEUl8yzBE0W+t8o1A4hM14Mg+4A2SRu0Oao4skETb
smKEjVUM/5kGjVTJetTuI9tYaAH+rxvLLV50ouT19JYXDQBHh9xk8bKalfDSGMf6
yexXcPSNKOudxnGcPjKvnoUdO/9WbOsgDUIWqPPFEk5Y7aVLNRCSIGY4V4EhUT9t
J4vbYeJiJgwy2NF/fQMP1WvWZQVPR8zodixH0YRV+j4d2Lzt9OtqReLOheBjTrdA
xu+pp5vP3bKo2i79HjXCPRC3wwS32DswfZG8JcjXap9VnMkhAHzNE+eY4PiW3u2t
QOVZvB/fSJX5GKOJZ9ztBOzFQdHURGOtwo6XQcMYiwSejSFHzag8m+ytEQbTDMYj
yFOOlzWega2bV+tUAFiAqivHRJUp4Zp2gcjfoPx5pmt1xqvlFyH6Q35BDLt43ZK+
suL6fBFcs6+w2WFj17YafDNSmbAozWb+XQSmowYxmZXZIqU0TQUk53QQyAr9Dwxv
dlD13ZbfgEJzpG/IONfpHayOhtcxH0IE2zPu4McqtSX4di/VKO8M4IKVdLnS1PMJ
Y3cGOZGFJZtJ3kut+RszFK/ZFN/PIbp9FOBKF0P/LHCLVMyh0Ro6Jrr6BvqtcExy
oGYtJMuqwKEjJ6mYo2nzkiO49uSp18vmBziZYob5GXgdH8VDQxSYN3fZKYUSKT04
FyPrYaItIFS/Uh6m9dCM+15dM/20LDPh4eaZAuMQZzngq2vMurdlms0kjYjoTkYL
i2VTllQI9VN1zNG5Of6tzNsJTgLTI4d9buo96bDTtn+IKwdCqLUXChHZxkSzXQvr
k6nHAiP3ts+rKMeBQV9UfOtsMI3r4MiKcB40XZaQfui0dtL2JkDGZYYRIETJGCeS
9lGs+ypZQ4X4MCkMWtqk8zr54p7+K8O1GSgYeOV5XTvKf/xxEPa1FgLaYSonPtld
LsJOZZ+We3RPzp0EOsXpzWa3AnPjreJ9u75af9bhFotw7rMP1R7RScorxJsfwDjU
sCb494FRa4SB6+neKbdgJfLaFnnVbvaeGrEG6lrXrZJW+myXKPPNq+UWUuNkGZKR
KMak94JbHy7JikA9Gr+XKR9PGQSc2tiuCa19ZasINWUpa95CNB3pPy2x0n/SXZL6
8fUZlCduMsSLwa1PMAQi61BzTSHyuIrUwrQontI/bVmbWWptjwLsRrtKzJNCUzqr
OEsszjQLklQj8a8kVe7mOZ5ha8JpaHDnSyBUcagM16ZjvnGCiYuAHa5AyFguQakH
y5uclH4PXq4MyO8ENWIACImoyR6oJpcnReaUHJja9zcIVGdLaxpsSqHUtbO3uuli
2o5Z2SICsCHPgMtcBCPekOEzipnndZxHBvOH1wKy9+vTA9Xb+esVZNIE4BGPyv6R
NhaPcBwUvxCqTMlV8j5TqEr8wLJFmDjvFyTsE/c4kOPIkFjqc8QCFUleESRLT48G
8NCLV+CQIaqans+XefOSFdHIb4Ifk9ygS7msUXJ1K9ORgwqmXsrPCUgj43qp+6wr
yGlW2SV/G+ZuXIFt58GqU8DOPf1bkTY5S42e0IreN8Aoe7ukQt7RSakrMz6VNj5d
Eam1IvCvbWd06qBjB+P1HbF0yEJtXO9Si8d7C+gameRCg5tE9xGQUssC7EGLoOUw
jZXZ7eW6hZ+PbeXoSKa6gFi+Ey2ZGaYduRCUh6r9Aa6qDr2M/D0ChDy0ie6frMLI
8mii58sXdmfCF0+fkXhlxTYnD4gU2Mb8U2QJXM5uJZQ1EYxm0xl8zRU66o8PW7nE
lZZ7pFaZqsoPZevBH5a3Aa2xdtnJ/yBryDXl87k2+17RQo4dajXhU3XkxXJSrpUe
21TRKS102UQs5kuF09eeDf2NV8JOD7t6Knao72nf3SDITfMmAJt9Mr2z/DYAasvT
fCoUExcD6gjMgMaR3QojImgj2BqYR9sQFlwbT2Yk9aObmzaqBf2c+i+uwGdu8g4f
UIXgzUbDhG2zndmoCaWfB+ccsxcCjcgxcTw4D7qn6GF+567wlNa3Ia5uxwN6MvEK
YmCRb3t1fqOYQHbNEkSNj7he7xty0TKp9BTJUYsfyDjbONu0BFidyk3aQibR5qem
CNWQSqPdupvTfewNTZRuSSWIfcy4ADdpbbHMt62CxAA6GKeLBQwHnN+/lwd7NBwo
J2Uxiu6ViIrAcQXXAAOhqGWI0DlbkDGy89OLNF4+vIVWcBQm6s9j6B5RvOwNV6oQ
GgxWKaurcTboOzbQ5vOS5bpgGLW2xbik8Qo6KAM/bQ+QXPXXEYUXsEmxGVDpEmvb
Kl77YBeDwDJm1P34MhBQp8JrLcdZvGSuRIVS9q3i7f4FgM/JI/jgowZ38kO1IXp7
ffs/MH6bKogwDPS5NEg/UxNHFMK8H7WUAwRZnMPQf+83yiOveL7QACLsrcFeXW9I
0cX+VFEL3AL4UNszrE8VT9Kj4tz7bSeX26NYe4AT15F3CspL1nKG2H8gQFyel4fr
sYzDZn77MHczagiztq3PIPjybhDF1GZLIflk6c/iqqVXIcfLmqGu8K45j+vY3OxN
Dt92A2siyXCbiTiFmZs71frFAkPbbpTMt7bJwnlQ4VrP8H9P6u/zI4UsHpEjjMew
ohfBf6w6eFnfnLUoz2CxmLaQzQpB6Od7rNTaqQLiwIQWk6yTdU8oUGUMZ7/pBHYM
o8PcWapcG4i8twfPFbdSL0NAslrv+RNWMb5uCuEzxfpVNpz8XBxBajo040PFhW63
k8bZBmE1VgER3jdjJnHR6eXckZtOKoLFUu2o1oC4D/Ky3OM1mF7g0I9BGasr/VnI
CVY7woJh/lodjVGuN22rQ5wZLAt0vcsYONxfhgH2D5N1LJ2odewHm0wShSf+SSNe
iaNnN733mly4RsbadwkUmWRWSoP0AqSjhF8+9YEcS4oC8auw6+aPN+hMCKxNyFTw
zFpIuP0FuUViGsavSbUmxZhtEiW5YrVkB1sHwjckc9cR9v1XAwjKP9kWcpnevTfQ
tTpRtxOUVr+2rOE4uy9+dr2yvKIzAjI0OM10wZ3c2fuO+HpYQ9XftyD8wRZaUD0G
q2RwmVkKgEsIdbcgD2NPgz4aZu6OW4o6tlyjQ0TmtFtPVORVWc3cAJIMtweUSFiW
vJSkvY5cnP1TVeAPRpOixviAQsl1b2Dr5CXuBJ7jE0fZNR2x/7KIkBEQfmTPHTh+
gDZWDP9mUX2LmdKJKS0g4Q4oTgq6o0HJvhtKSBLuutKuPirYkYJqt/A7fxE+Gk0p
sQAo512XEw7aR+MDPNLYrt+jLQMgmQ2+vQ3CMSPvwxi3LX7Q2AXuNTs8YRoiE66h
F9qW8gbhiGFm7yMV2SXqkI6fqDNw3WTUdtgbtGLIV6IzzWtgeGfH24c1Vs9ayVm4
YPpBxwUalfV69M5atfPdY7i6neUn5WnRfceDLgdNztP+HPFk9agoHOgtW4/GOHFO
JFTzg37eihH++EeL8yVyPaZSUbZ3onPXpIFduN1A0qlTJpgs0zOmp/2rJEWVuG29
6wQtd/ScPQPAG5Kjyc8L7CvIlCfmob/CZAc6CU8Zq/j6WrMxYD0xv2UdCf7+cLHd
mL/69AxCXXEtnaxRowB9qjPweWhuEAZL+9hHtq5OxaBvQqneOKlfI9dpicmatj5g
mcGQvUXwzQd3eRCwje1btfZZImNpUPpnMHh5+5NqULqVLSP3zDl2BH1qWgpR9jZq
f0IIACus8JKXXNcmfbD6IL4JL7hvsmCoFdcv3vtjtTIdY0Z2ggn1twmQOfQAOvaQ
+b97Ywir0BTQGoSJaTpxMH+Qiz2DgmGmqUtnrCO59hug0ZnPtQFIJbaLmYqpRs5X
n4V7FeoBR5eyTdqj2Ikeu47BVnu585/g0tnWWrufM0jy6+fO1ocrFJlndy5twYpr
pnpVP4Ga2WiaxyculbK886JweosrREEEAazNCJKOwiQztMe27bJCdHf4krzqX/+p
MHOc2MvQKlkx6AJEg4WuUqN7GUyUVZ4FxgXAqohT4iQjlTxuomx2sF+pX7Fuodtr
QMnd0F7G65fZGkoRw+ZklLSATtGchDdgake/pYsUNU7wyxMmvGPj+mDZaF2J7fxR
bzRstY0r1yrMcbvvkSdAciES8jonXWKlnaxJFrGywubdkq5kYzGOZKZ77e+Az1eF
9SWCygpsjQ/pLc2OaNLQH9bLJOjoqlAxwCri2H76II/0cEGt4JCukpyugnCUlagu
GRuyHklVXH0YphEFfB3CV7+Xbfnh5ydiBFWnHaVTcjWLM4+1U2bPKLxpYjZklZ2/
iCS828cjHLxZLJfKqUUd5teybfkd3eIzQYw+xIx9/fzTwH1l0WQNt6e4B1QJA2Ad
JCasA57mXYP9sNp9f+D9FfBTx+VjkBTUmLWeDZ/bpoW8XIJ0dQNiGmcSCC7AEvl7
b9DuNTkgAQMVlBQaU9b4tYY9S38lCyjR+CUNv+jU/JQ/r8rwx9z7FSYW1Qgmys9d
i23AlkIzSqq23WxPyatFNquXeR3edpqK0zk0Gb0vGweALYSKZCql0yg4otpATPkO
wMZRhlAnD17HP6xImFMRoYlaR4dco6F4mFP2bJ/gTGwjv4bHp3W71m9t+4FbHYyA
L9Adxyp+/NYBn6MIs9I+NHSddno8wR5tE5uqtMPBMN/0lJH2Blc65jU4DvRfhRGC
nRV6psK1Cm5yM4pN+3N8dzWsZ7kgaulLtB6SYwgHh07lj+McgQzO220+00AWB4BV
YErHRxDinBBJKiydUioRQTZd8XOU5+AtY17f9dkh7atGdXpF3yXGi5GYgQV6QmaK
V9MzDL9jxVAcsl20ZRs6kp79rn1BNvSuAFR8ueyIC+oZgNYWoLC8YodlGmL+oJ4p
e/Xjnf2DWnkBr0CW8TqXvNvVkSu17tKnI+NVH6TO9gBB7Ha8xAPhCb+1ktz6KqTI
7swtyeDKkqFeTwjhtzOLCpyfkgVMVh5Vo22aczQ+nIkl7OMISojiL05BfHD56cY7
7zWwCydaAuKsnx+w+UBoyoa2OvuNd0//kUbH32zDjce4DX29siQvFMDjASRfhuLA
JRoeB62iQwX/GOHbzQNjdajcDeArpPTMr74W5IZNEm5VDh+eOkGy0fIVlKNC6Cot
sAeVMDNreZIknUVKj+5pFbLKbSZ8oc5v2lhPB61b18RP+sfsVD13alJl+nuTMW06
+K5kM7yZGPAe1498hcZzVouyCdBtpZoTmRnCqVWP6GKKErJw76gZLd4tCNnseA42
WkNZ62yR8NJof3AqqwXEX8hGNcbAgEmIaJTblvBzYi+h7u80xFaj0CoA7TRPPkVV
u3LJTC7KVw3jG6N8EdjfONBT6MPbgOjq1tL1ObWTrfxcTKtPdXDCqsVA0d12yGAI
YdrWKuJ20Km11FSbB6HNmM31+R9lF5ivXYVy8KZCHC9a2woGCKigzFhMuejnK6Pv
BgNTL0YAozxU/95R5ESQx/qFfiTcfrd8Vabh5m/fISmXWT/5ER7BhSJ8KusjW7Wk
kfyIYK3S9K122NudlePyHilwQ0LsHY0fD5XaHosaShAyng6NsU7YDUWGIa6PAGoQ
I+LPynD2JbIdUmLmSrGFEck7HOXTGdd9pisWnIcWfaw7FhUXPywJaShnrMeLCnQv
4+AO0xiuywzaj4O9+ApV2gRym9IdYRtGG3AAWpUwvVYyDZlQ1c2eY2YTq/8yq5Hm
AUYG9vhPKSeuwelJp/zwqXzppVwz1AjS01DlCNcpBEs6vdfunhEyfHiZnE2VyQh3
erArcTOR/O9F3kBCeKaI27zM3Ut2GR0PPMhhZjP8TU5UNwBIAynTK5vnax/JzGS3
EkCXoKaysh9iXSMwqheFZmiq0dWfOBuIpJrIi/vCldtZSYJOPGB0bst/5mN1MAT0
tGF8wrbKrMcMqxp+ugipGyvGDZlyJY5+BGd+TffpfZbgOaOIjAkFRXhyITh/Sps9
GOFsC1P1MNPEu0w4wYdGD7SSkWgqBin1ekYh8bkW85BkukedGmxXynMi74IoaAzO
gKYphY9Zn88ocf6np50dx9yj32PiIQtgLmgy8dVWv+j/tufM9NiIX6oEG/hgON6r
H35elPUnI96RrdjSe6XHXmC2gFE4O+lXAw+BJqUhPOQ6ZbRB/JJH3saVXbnjXKwB
p6bX6O5h3XPvc7BE49M1Afe5UrcOLpfQKNBvAkZksy5IXtKp60tg67Ko63/bDt8W
l1+ZlSyj4FudyR7/B9v0Q7MKeNKdgpe1uqM6gZd2ZHJLo9O2XvxXSo0FNrB46a3S
J8L2EEJqCXVRoucfylTs5Xai/On96Q0udkhYIPW6w040aErsRHN0X/u7GaoOTOj3
mvuGboVLI9pT6dq1gow4KA+ahNQ8uh15cQHdgSuz8glMAbCOAchS/IFMekPtnTzy
haYgf8hU+EhNByWHQ6kzx5WL/0YZknOWRu7+SjBeCcTm/fjmzd/7klYskdhmms5Z
6fFDOdjztLZv38P6fOQ28oO0VgZXDokIXvoRSTfdkSsmMYBbcCFVx+jF9sGtb5nC
4CyvHRAIfOYF5beJRJpP/RAznVX3mOJPS9A1SN41r1Y4FbWOJqKTqQQhBmz5+wvB
hII5AX5++65ZASF3vIjk3ZmpQR5aOLzmSPzgDmQ54y0PF7uJJUNMhfgkTqtgjlb9
lPD3ygvGamWwrGIoAM8ABlFMfJuJP5488qdXT/WUO5VNjabyelL4VvlTbjA2f6KN
EOkAijs8FRDjYi6PQtlMyQkbhHbDwHm65XQZ4oFLN3frlrbD4dNkzNHpFwBlD6sK
UMzMixNa4L1l7ceeGDuUS5VUR1+D4m7ffL6atOmeNHIaGjEY7GU32VvrVfbVINP3
TMp41wOYv+fhI9P6wwV+azpaDQwDyoo1C2XsA97LMLpw+e/gwPhk3+Z7/2J71Fbg
XVst+ty2nPNjFlAh7r9UPsyQ/fImvxxjIMjrDMBfPtBGN26epuVky2Ist4K0sldn
2sVN6PtEDK3SJyosmS50mv426NYEolQyOQtxVDy4BVIMBEc2XZxBG0TnQyPGFcd1
rLunMWvbNj+DVl8ZbQUfwGDSd78EYXgfm2hMS5pf/mwr9sfU5pp3uNZ5UuGpYkp9
7sGWG4ZaR9vdtp5kQ/IMK74DFTWxgsY3TCD576tKbzT3FgGJeGZSdL4f6VLWWBeq
OI/FgSu/E8UBm1jIwgT/GjLVqK74KSQP4ZJPEfb/WKzD7gs0gYIulAuYvvNZKpHq
AvVx+1RzflltJJRvYIEqMk8qV6EA4AjmtV0JYgBe9XgDatN5+JN39wkddH0hmR2Q
T1q7Vp07oLBKYYFSZyQwe9hSIANgha0TXm6mu0V4ciCSdrz+fzOO3ARYYYwaqk/w
DN5ZROCd5ptI57aqWwtHxrHWnq0mQrpqwviHPDO6t+lGDDs1uc9bFLTFA1GGWU5x
ksNGx4cCF7H5/7HaTfKCaGNd4S+2xIRqaCRRijMom8GHz0cxnpJdvGNwcFWLQhuK
k/jpxxGImEg+PRVyvRs9n7RzQDGzFXyYGeL+J9+0bvtPsuk4u4OmDunVvpqMrkDO
ohpqdTc1jJ2ReZIk/J7JZPS6ep6wRT7j3trAZFvaTX23QEqBrXMZW7sUqIG0X2ot
i/vuOkT8gpxbd+CwLdeT7ZFjA8FVY+J7ajcwmBqNcNUYones0aXFjeuJC/BsFjC1
oNipNdfXDhYBNJegkvf3mFIPErHCYhl4JgwRQnW9fpmI+7CerL0b3G+UFwc5m0PP
iErs5n7wiiz+gsBfXzuscosPyI96WE1ZpDladbxu9Ql/kQ/CZwH+qeQOAWTsxwXO
qS5Q16b6bzROVMEHHGrm4wzHw7xpiDylWfZevzhjM0r07ubNCdW40KKaZpVTvGYm
8N96QJ1f852xOv7QyPal3rFjiHTaz1lUmLS4Wvx9G1RV2UHQB9siKS6SG8Am+dIV
BSI/NIwHdcU35/teSB5GkJ2zjQTFyJs7f3GUKGjWq++XjmYHumbdDzm2FS9rliv4
q5/1dk8U1yt1CpTRZ8Il9/uHVt1FBSB3Sw6bnM0sWdMYuRbW7BZ70/RvKKRU0pTo
TVNv9gmID1+vRSG9/Q0Uw+4ifBpbfaTIryOFbUpQwzUTmz/XQtJicIBhGBA600GJ
uY9TJ0+QmQQ3YWxBj3cq1MGQyy8NSiQkQf4APDtRMrd8TTCeXTxP3nHuwdvsQs/F
g8RfytxvrLqOgoptvLrmrHLrS2SRcx9TxMjgyoMvaXA8vujWQep1NX5Jdg4A7eoN
DwkUdDTHgw6j93XBBXVSCv4QPzVExNwMmAhKF+8GDBqV7+9t1sebWtJitv7Yh/Ss
Q8C7xokn9DW3oE6NK8TQlk14/9GJWqotw2dChJfFV5uXrFZC6Vqj2+yfNDUmzGTQ
R5oMfkTaHxiGuk46p8Hy1E3WXR2tsnG5qtrP1JUlulx4tKCFjUFwtN5Gb7T5DCGc
puTWM/TtBy8PNUqYNXCS4rV6ZDFR2WrmPTp9a4uM3MGJr3eeR7Xw37GB6BVZ4ndF
Zf36QUOcsni2USilDOySqnekmPuV3RGQcUYVAOXeI8jCE7gEfGE1qmzYHSgz1JwS
yYbFM6AOF90Y5/Qzkzp+A4zbtkgN3KOihYD0d3HtLD89sMoMRJBSjFkDz4DE9vrD
ttSXtaVnTg58w//pJLnNbNJSeDPxG5UxAvG7pZvWFWUPWHTD/6O3baVzVb/aTpWX
giomhfuz7SmNkk2nK9ua3T+P/GK+ebCtjlLsRNi71+OhqqMtgTwQyjVFdqbGyJKD
hSgwW8n8NGXyigl194J5HpB68ITsAVwTPbsVkUwSh6KIL26gRKak+V1ntD3RBYGg
CygfcvSvJo7jioEirWWjuUrWclHv63boVTMUKYfvVcMofxfGeu8iDv4sueuJNKCM
YjXnyJf3HKxyXQFP4mZYNVPOXQTXI121yQbYIUFj5t4A/cG9ilA4hLj8pr68WuYF
2268lDub4rYTYExeU+5tXg3KIaCCWZSFZnshgaAJmcq9aDuvvfj3lAZRKYMvQFcr
D8S6ORH78Vgoho2MZLDc09gk6ce7ckCwh2eNdYbokqk4pdktRBEWJgDQLsJsc01r
X39BOi1dCI7BDMWKNFN2gM51eOjy2B40bJVeeBLeB9blysFeU4jOFQ23mo6ldhRn
OaDtEnjZ84/ONGA8lwCXwDseC/FoneaJk4MWsPIWnq4LUqmz2C+5IRG7xFViCOIk
j+Wx3+SvZDTF6Ay6kZ8CwnyB7h1DKBNMIGVxlF+v1hAI0dCRdlAu9RY6dDJz1Ovv
7wwU8VEh1+jZzOZkI6senY0ySVufNxSXQpzzyWH2CvcCS6WpzhvKwy1aTyo0JdXd
eZb++6N26e0aQ+Fu/bKfPS//CGHmpA8L1C37SGIMJMVFrDUG5gBLlPmYastwQphc
omBUNO4H74A9l2Vwx/Vh7G+dJiQTS1XJ8BkByDPGppen0rbJa2Ec4vvD8l7vy0KA
CI8KFuqJqbe/Qk5VjYkWjmJo12LeJGfEzSN6nAi2PlnIXG4mWoHTv0XajzQhyjEp
yO6xz4PrCtS4ffG/cKxEi7mTdWxj6K29ouLdLju6te5D74XGfSnu4t9yrXsjh/Gp
uHDzBhQctIlz4VVIIlciuohEkWRsd4ow8xA4d5eT/9cs3TZEXJAxR9flFPdhtjD8
fHTIcxWclAfGZQ4p6S85uhyUq87H4VWp1uJbkOANQg6F7jFeYQfUW+LPwsfdTZz2
Yk2IovyP7XZzu8uRLQ46ay8SbEkc0HqOOXF9GRS+t6uVSO7jbixZ2D5aVuzprHBz
RLvCq9BNiA1+sqhkUhqkbtMAOzAcjA3OmgaAkgZmn9rrWgzjDr+bZnzUeH+TQvhT
SKDxg4H5n1Coc+F7clKsyMFjGyx+VCssC0hE5INHoDot6JQi/azhD9UxGs24ExcR
yGTXOg+CtTRY9H16hqjMoHsnwY2Ac++GQmEyF3t82y0HPmNgKBXSuFd/Hj7UCA5h
YGipAvP+8ECcG14mEZR6hMLQhbwU0cNgAWpuyQ3K36DZLxc7UnXw51UIRohjcEyH
lkO+UwIb44Kq1si4ObfHhGgJmbjWtVv7lKnULskvEXYD3qv4uKHack/Ey6c8vQkT
82x4Y40qULKVRg3gihGM62jH4Fidx3MUlIvQsHSvKVEET1N3IgGRptVUqsbUKln8
GSXE3YknrofYktccgrA8bX1YbWV8mbtgcnaeTZxrWJmIiJVZ0x4PGmPoLp1/nVga
YxkHMse3NQvDeFLrmVfz+UJ8kg+TnOXy8wgGqeMWlT8V4rPHvUg2mFBTbp2D0Rqg
KUZ8RBqWOK0oraqlCIbaV33qh2WG+qJPyfD6CJ0nhwE8VwVjsVpbBbZJyZk/OF2U
hCH4HilRMiZW0/zT4WTfN/OuD34n70mw3nZ/EhvxZKeY6LiQlrFo7Iy3/5fY7a0e
ho29EDPWxZVhqBSU64LHBX+65fCZ+SosHyCb6GinnuaPR2HcWdnS37LjW6pc6QGX
RABwhctiqb/DMR1UkZrKk3/EUWKVE6jbZC+eISvznmf0oxQahOTfmKudIlrA/z4S
sgvJ5yzhMAEdYOBmybry/NYoSWFIU3WHf6Nvd+X+l8zdPt53wDAC4uAJQYbawnUk
JxI5zlXevATG+EK1azN7d+Fx7/4kF5dpDQREF/y8wQ2PJTugwsbDgTSuT2QPklcf
i31KRNfDR8EwSsfYcOOIcjeyese8nLnsXhOG1Fe6JLj7xKP6QrUv16kEGqXKnwJh
weHnH4uIUPAkjmkb3jjdlesR+9P6xvkUREYBblwBRNsYKo3Yw2q9m/dVVQFEV7qp
Ddw9WYBUd1/XC0iA1XvgZVjuXTidma1uJWeQ6ngvntZ62LEqBOI4dM4idnH/N/ow
H4xzq/psrII9wOazI+lGdK/e53VTUMxA07VG54wJcH2kaF2+D5lB3NqllnDe22gO
UKN2ymqO39LdqOO1sk60Yf60Bio/LjEmQV60iR8u5L+XRe2sTKo3hwG+mlNAo/CY
rsQJVYxPDrvSx4gJk9TMROyIbNmf9lqQeTH58GKHmyVnoFSrETk2rJupQYIfY8GT
5fkZoiqEnBGGurl+d5w6LTobvQfE8wbRbNfziF7fKn3RYwDw6Mc8qWGkgUaLAjRa
EUiT4WSnhdoz/2inMfoerhqiAdX9tN88Stercb3/gIE9ORqZC/+psO400dxQlkeG
ujjw+MeHuY0AtxSX8rMjlpPqs08oVbvVlw3CewkpSaBggOaduF+JmIWGa0ErMxeC
pXWHTJexc3E5SF+xaRP6+PZj45aWfACpHo4Jcgzi+wJis3H3yRHuZVL510UVzPGG
DpqwJGlFqq7m8R5PDZD61hqyYj5wIAlfN3nLYDaQ5h+nJVBmMFqovHsdZXPFcecW
Ka/zcBL9XVpAiuJXi33llzqn6mrkgd9/QL6OBo+uCnIh7VGukHoRkgPuZxHmP/ym
ME5SNMfvuGP2PvrQE8fo+AxTE/nYDyJBJEBvebJRSvdKwfEqIaO9G2c85rewmqod
QxBPWvzpesAiI3TehQyOGpzr2V01SRNUYHJ/JjjjH8WXIuvmY3LeQYNfURlbJzJ8
SeErWEuv9iGhMs4SXFkktOOBI03cExrfEKPLebFK5lNpswlUDT2rue3gCdyVfoCc
b7o72PZVQPh9GDFkhJmQ93sikDcFX4dwkq9a4W1dR+r8YZg/KCBciWabP2VVw3t4
1mQm6c9p0LBBFvYc5oY4PvqKrQDDAcqBbNjQ0Ma3Y+f95/1Cg0X/RbEQ1mEupQS/
2qMZVTPVr+OiaYzVPi8H4F4qjx79iNFAu+IZGtgZ/JB199S736A+dKBxEecJpaF5
qIDP6ribEEK7b71OsTwCZRdUHr9WkF+gvQU2iTNCIAa9BqN8WtC8uaPp+0ljIAKk
U8Frlf6WBuP9fT9ZIXu962qRcbU1PXO8RotH8vctN7XkE7Fn2hN4mjYrqIZFwCtX
vQWGVimH4JIYUNkBFpxDnC2ObA3Ogn3ngvlKjv72dgvo5vvnwX9vfvqqhVvnKBti
okaL+4V+wCOzAVk5B4hOiGPD12Pjn0uf9g3JFOAG4th+zS/+/bCWA/KgOBzDGgt3
t9WlL9iUj0VMBseLEkkWSELH5v8ONdAsV/wLczGNz9fen1hc0WRb53NbUqVSUI02
AX4P2EGxPHAtZpB2WXWNvlMebVDVS34ZBdwkwi01UB6GxldPe8/4ogEZNoSaDRdw
ur4I1tg1efxY0zIIahSBHl732S8IYzt41cch6kZ6WAGl3x0b2ivejPJ5wvLItHgR
xkVFA3ZsAlebmz07n/TiEDv0XDGA8BAMt3N8A5l8joTRGkEqbtlizijHoa8lYorK
pLnf/ZnUZQFKkxaSwmdEa/I6xWaUzcggisx+c5U310WOHUZEIRmwTCTppA6wQtBa
XuZjEAvqmRwvmY+SJEIFU07AT3BOJLiw1jKt57bJSTHueulPh65PP+3s2cpsdRdB
cj9FmcX7YkYE60Qzti2msqzNxZtjJaX4RRC7Ufddb57qfqKL+L6PIOlKztrhTPqi
1ZGnSMyT7VGsuXtf8q4B6UD352x5AvCtg71ABV6N7nnzImQ9GhpFn3OO/wGJ0T56
cEomLXVlj8fcO4znoo2JYq0UjwPe9/UxfLElLxQUb2vdkTVwhTqq6zoal/5POU4r
UWdp0aWsRirfmPfXKC+cF2mQSaW/h0K2UpikYHY5PSWFdvf7tuhlQ9wYr9bOPxY3
shmjH2BRExPHfR7ZHVSp2RYw83rajO606IyPIcxFn8kqVvCyz5f9pxkTGODMYZ9/
JIRNhoJIkzfbBXoyAqcf6lSYmB5tZJA/JeUyb3az4N3aPdAtxufA47aYIibcj02/
WVwRwvnsIDwbQElMpEBj32ra6IYdj0IHlAozVIZQ3eUeG3lx84HonB6CL+jTbZK7
ap1pVj+bS7vwWuaaVStrCzGbtqxim/jvsXV+T+aWE77TYo1YkviVLmEn+vGEo6/f
lNG4ypMaJh7LYSuGid/pAb6QvqzPPpOhYCtGl49pXXtyUBJHbCEOGs0sl044qHVN
aZUZVAUbAxqwPjJIai35k3Ecz2GGNlxZgJExuhMNC7AqJWU4i693vXMYAkpY5edU
hmrIuE0qmnj6pJ8K2xJGx3dEntBn34rYHQBcG9koKJKSA+k6Ww72y3c++7Vw74t8
uGFiKqFBrsUunfQezJ5POxZvlwadV8KLS46MPYNhyzaNk0Xzjcb7zBW0sms5eV90
BLWT+SXtqORC8t1BUXi7Tayl9imozdMK2OibZqpAejVCk/zxpZ2/U+W/G7lL277V
9BB6KCx3KVic4Jns7Q/ZsLRBxor78R1E7vbeoF7IIadS74Dms8sYNICnsaKqaJy6
nLQWT9TO5SwXLZ2caG4DcGIe82wG/RtO9AQBdjGj78trm3bVA9mQcNRfn3HLhNUX
tEY+pUNQWXEpUCV2M790nw/sv+v53aMmzomxzgVcE1XUR/OtDQwejUKFIC9jq9nE
OV8f5BE4kujWXYxRteWW3+/b1fgYniOihcFErujuqcu2fu+J4xE6n0qqSNf3tMQQ
D3KXtrqP0Qc9DaZBBHPBHfQ1t4AVg0xPpN75/QLnoMUHMf6gt9IEBh8ZFDCv2GOO
k/xwK3PUbOOOEag/AaQ3HPFgcJ6eLvtmhM7bzaQTTGzscKXOTnDZsyLaAN+nLBMn
Bwmue9y5k2tQWDvenn8KEsJt24ghTgAl5K53XcY+uHVh9hg3BvASrNKkiFPP2b/9
aBim12SAXSimpr0NsJRVnT97jASMv3Sue/ZoqaTmv/OgMJg0XCgk2NfwxtON1IGN
zWbWzf1dRvmNGiW7l1XjlJQ/lI8taojCFkuNcYpatWMaRQZAnQGqqHcPG8De5S3R
sUSoD6IdxoxCIzuqzxF4i8ClyhIODllCLEhd6wHv1h1qnHzAlQHDeR6B7Dw5OhLg
Fvigju/ytij/TfnZ0PZTDgPKBNmX+FFLNbs4aOHWFo/PSayNKDffsoHNpZlC5ZOs
uzKAsvwKR/dCRMGhBHWd8OZoj64aaFGAiulPwnpLWvLkhrQIv9cGUGNIVac6lj2Q
ofanHbNcXml9DXyCNmYaSYNZZwsdQMpgfz8eRslsJ+H8UoZXI1k6Y/awg+hNxByh
piFb+o/SgCotirrWuoJY9HPQsFeHU+ADTZXDv4xAvUHCTuebQIDQpjUx9Ut3mqHb
jv2kM2Imx7Mwhs9eF8FeuRS9yYUPQvLhF0qvEyY8G2W292Im1RLyHFlGk1Bq2vJc
DXClTU2Tm84u9Zb5mPs/BaIoiMnwRdzTB+ZhY23cLApeA56uVFNk60aTMYvdMyIG
i+VaCm8Lzlu7rYRIfxHLrgazYnzRR7QuUZFWx4XLQqw5nLSfnbp15UooDDu0GxWo
A5LQ8lzIlGLKd1DQ3PNu3Sbc5amx6J0vN+8VdCPGoJrlo1nmoAA9ZPmH6CVGIJj8
U4CX2x5dRLDDEx9M+gV0GyIXftbD/09B5wteR3EZ1JxwE+NK8xncuqTiZvIPhvWl
pbO26Vut5e7stg6TWRwFjZzz/2qPuyI1LAzU975HgltVm230lT29WCOQomOjrJsp
0jcNngYb9Yt9wQmOrkVJVzOzytK04d4RCTzvnlY122qQGF7/eD+Xwce9hoxmS9px
3O6xJLSW0bdX3Nno8JGmr/2vw8NrXNwXoAlV7g962fLLzZ9wQGRYSj1O9n3t7OWj
anTit1lbq4pV1rXa7SMR99d5iahxn708OKxTkR5v18ltP6lMFdr0YMsAslkEIUmA
IHGnBnbNlt4Lt/T84miP7F5WRnSdRr66ZsCZ3oIDOEumQGvodrnskRdJirCJczB6
C68s62wipP0SIzESfpNqPmgoehC25Xcb7dc57BtSbjrxWbDsmihzWfNpCqkHt+2P
Us6tNJpYolO2zWlugfD+zXhALZI3u6hyrE0by6x4OO83CIwsgquLc5waqusSv0QD
Isg4f5wAqL+laUt73P4IliOzvuCAEKtBCofalMCcSvY76catqJCGtzoII/8cH2b1
v3J4qU7bbNgWQuG/Fp3TEw3VXwEd5l9UudoGXlcYjKY4dVPu40BLpnnTIog5RKUw
q8wifwRwLDYNzKD44iYOdA5WvOMF4zBkOV+EC+FmE3u5ShSeYCXzBHE4at7rQQZS
PDCdMDKtahMeu9OUhg72nt1S4D3NPSvuVPNjVHrwnyE10xxuGBRQBRsbccmWWApe
H0XjAUI6McKIOAxMDjr2HkpbIx5IAvDjd18BKMwtDwaE7T+ky37gkwqqdjildQpG
Gw7jfhTuM8ixZepKimYKwjZTLC8xf9i6TGhgLnWGb+EN4Xzi0WO7qDbiNGH3rreH
Y0tT859YhW4gde/YWRiDEbfgDhowdLzunMgGh9HbOtmRTTmGpGYc5zCNtGPaDt4X
qGwTpzMu1UL3jSMxMvINW/iFGEuSx07ctVqywZ6TfiTolYCKynwmEYqeRzCOBaAP
AeYVmzAErR4IGAa/1d2msvWu3ngbspEMuVbv7nabgMq5I0iKBplrb0ZccVM6D4+i
EaxIPunShGJCUHLEwxsuAfseSLeV6BJsC16VuUAngfHcVfnwBWtAfP12yxL2Wjx3
7hrLwsZfFU5OcIyFZ8vE0mLfx/vJGaAignXE7c0GntgoLSv540emamv2hG4uGqot
ILKPsPFCywOZWhMOzwIf2VKr4KdbdVjPMadJsdjiERmsy/UeC5cRZ6rHTRGRPdte
KjMMKiT9KT16fne/iR9YgS/w/zbb/ehxv8B0xvNZ+CLBtB+qWb/RgYwK29AzrvCU
Ey9UXinuI8orz4Hl8ZGZCtHpho442LePMXF8V6kavYFZ519vo8fMDtU9bEP9ccYF
qOF8bGgSWhnHqjPFIGlRTKLma2IMplDBg4T+tmftvrheyDVpIuHEy6r0gkwCHhAi
DhrpPunpzwYoOcuYvnZRqThe0E7/hBNH7viRwjyENgq+oD00kpHaxkqXW/03qWyx
OFWBseCNOGr1GmWBCile1H7Z8/iG62mUV5yDU4x76/qbv22NiLGH8UvxyI9dg9Po
QNvSC8eaRGztuxxTt5w33dWUj337w2UlmRgbcat0T30fHQfU4cSKBUOecupjnh+n
PbQnJK9XlKg4w5txdw6xkR/zaVFMYQ/Og/G0DNbdct7gvsxWIDQAbQtwddTFTCzm
Gri1PDMOgL6Eau2L6G/4Hguj/tONzHLnr8I9KNLwMZZ9DP2Nepi8RsK/ANdu9iB4
3WsMhl2By+/9icWP5qvxZqjfchA5EpIeNX2b9CHumFAvtsJe2JK1K32ILU9Haa0S
FFxFZATlNTUAV2F9vQbEriUrvJnGrUCqSzAuNgTM9uSu/ybGJb8nRAzDC9XGTykV
IFEexRx6kuRHRPv08JAO8GpdieXW+FgDasVxwmItVRoFLxROcjRalkBXIDzOCW7G
KVezF/ZikF8q6hm/HUL7JFdfmLudPmrYIo0COTZWuBc7s23vIif8TwyP0khqMhXT
2Zd1ZqAsB7TIL8XS4sf/a4brIG9txX0gjnusmdTbDvUV3ezX4mJH1K3UbruzC28a
R6lAWObvfyeqVXUoqEertiAFgywvCO8/SstqC5gMc70u7knKsmrrV3FAMDBexQ/2
m7F5a7t6ThO+bTIoqMcYrRflyMnT9U6mEZZP+1/XLRzCs7mbLP7AZbVsdRBzUQ2h
sdbvflmFiPTAczdEVr8GNNRLl88/rFr6CAXOLJLtTwkvCUXLYKKqlbnSoTfPNnxZ
WkyhaDcvZUnvWel5xPhuhDsFUlaWHOAv2AyhnE6hzl1J9JK89jWVemHR1clTwveZ
6SeBm5CW1elPish9UzsbkbVJ2zLyAZf+qLeZB5BGrQzCHOiSRyGi/z950CvTaf4N
Kv8RpIO9Kr7bsF4/sS0LOLSMnLZe8ru6b9DDpEnR80dnXI1iysAsocNNTGOwjyV1
xMlFs0DlNJxcPUP7QrwOBusIBziwdPvzAVCWiANfpUdXgg6MSrUmWI/USM3VhfrM
VRxPQu6wGQa+QVnzlRYV+J+uZCz9hpRuoDQyxyPIslWMlkpLtiOocv8TvMbYnB5B
IE8L7B982qApaT1u2sIUMyr6Cz9H++DY87LsAedghFtbuxDdNrmuhIZXPDi3xqcx
gZ/3ATQydALaOnqpO320D39uIgLKbjzKKVGTf3pW6En6JsTQUpukmHYqpiAQ8fpQ
2Zsf8/kTBy7quDKYFnou3ebEcpJYeLkxNi6Er40o0ZjocAGADEv/XDaxSnbFzYpi
//eiZyVTxbOUV+DXUYZUric/Ok6/BSDM5WfBdns/5YJKb7cGo74qzREO/8bTLNrV
f13ZLPwsK9dBetXiSiCveypRjt16SIcDd3mbDNTDvDjAV6VloZz0Nv2HcU0jFS/I
mkOyYRQiU86wZzFBsa8bp/qtSAfKL8xFffJwEROUBgfohPKWwKrm9AbQKBZWn9PD
O+6Af9WCv44tTDh9W0UttCPaSZid4l22iGyaS7diq2Mf3SKHWKbsF4cQGpYPgIck
1gycS4fq8uZjHd/IqiO+HG0VlM8NDi4Fa7FjGuTy1SzWfzaHT1vHk6cEgk6HAXVl
XR76Qs3+PLN9conkmtDl3ymJViVhmWJKVBmRXPROYR1hBXlDn8f23h+XqQtgPYAb
iJgCLk3YgUALyv/chww1uQCT2929FQxsZV3HmLPdhYqojN7EyRKT4WL3p4aZwTmT
FH0IHvQfkwqtQiUoWASHRmjAR//GGcf3S53+/eVJ8WaXlOG4Bli2a05gVWHNRErJ
t2SPrAr/MhiOYQQ+MqrQrDxFS9GPheFtJd0xMA6lUY8e/MyzikBlOIRIYGFpDlt/
j4voOgG3Q1/g9UzkxW42y2aN5jVFInWB97DLDBHCI9tmGgKZ6h2mPT3fwxUs6tv0
MvFae88HwSbeBiyBGgMWE5QBTZEIdtwmuJ7rhYE2rbVVvTiSCt7kr10Tt9R/1oAI
NoxYnq1LvtAlvV/GC0Vn8pUpQoFQJn3zSqkC65S4zGeTapEMplbMLAbIGyuZDPED
Y0mjvyXdo6jducenXdyWuY3ZV9DsXL+2k6d8rQob8KvJt21QD6shjEtGDGtlEzxR
xeZtKciMvmj/XkwvDz20x0QKS1h9rnbavGj0miyiSxhDpKWm5aMYBOIST5c0Js3q
KEmutQnzqrKTbmArgj66cckj6SoAnFUA8UkEaFE/l+gAeeIumK8poyF0Fo7GN2CH
z9GAmNhpP2YA/lrdP+lHl/fm5C9vSZ9MLNNnuqkI0ENiouGLNdb5Sl40SRa3lDEj
MCgDCauS7vQKj1pm5IYFLsrBOt7Lpp55XKWHwzpLG2v2s4CTZNTT6Fo4oNxj8BX+
Xcz0l7YfOp6Vu0fdFBJWJx+wU1zs+OwR5hkBEQvkA8Y2CwteuZ4c08QNW+YmFO7g
6SSLxsGcdWsrrCI5tJY1CONLxIRwzsjqlq1T/B/dvO3bC9/K+z74AAf3Hkn1K3hV
Pa/NsIfQVHsBZlpDY6z/cNh7BYXKzvniVnjyp6gJe3Jr3uLsWGPXZfSznCDwtcHA
AAXN655IqrJ7TkgkTIYO3nL5fr4sGlLd1HjEdH1Se3q9VsggSRV8A634xP61rmla
5OIaCWForLNF5cLLQAiS1iebkuapkz7fYPd3mWzTXOEsiA6vsM8bZMs4H7X6YkaX
I7ryoYb3qtxuIb1q4jueY9JKsltPYyKEnTAMpUczHFmZngO4COpmnm43daZn9u07
+43MbgEHOdEyBWkONO2abUHhcD2n9LBoYWA5MacLUDsTMO/dP7LUosFiVemfyF/v
t+2tUNl1z6jZwuXS+F/yprbYA5ahLxLeKGaeGZrVQkEZbxM8lfJxsRFE3paCl5A4
LpUNRMeMLygs+eG7WHAjEe4YalrcKdT4QCe5B9ojPKvG3GnHIyEqfJAHLfGdF2Ol
AsRi+idn6p9wl+Wn5pFs2XlQdO+xPjUviuNFy7ZD6GzisponVuZH88LL8fLG12Z9
A8j+uW6X2wc86SpiKn/vxR64Z7pKzyOP/EFhgc35zoH5w9mZvkW10o6XOtREO+4s
/9e2jzVdi8HikZZARk+kquQ3PNRbEUzqhoPS2jdlky5bF3B7wRg/rEXhpXcI9F8h
98lDz5OEUvuwmg6Vn/cGWToT21EYMLfqeRBjl4MOvA7GRAfsgo+xIYjocCVTGoUd
imJpqHD8TCRhg8BCdh2mmRRBaLVf9lq+J+Xlc3D4QpAusyoaZlz/9Ae6GAtZN5uB
Q2QqKWJjNbe4E4LgDL8K5JdI919akDx0rS1DXsJ2i7tNcP1RdJZCt+SiekrTnNIt
g0eB2tBHaz4j3Pxyr7nwOeA5ydcHDsxVi5H0/CU9fSf9oC31AgbuiFuWX4tP2vNl
+MWrr6gW5XATiwglOC1wWUOupMHzTk9Tkb+4nwt0pR+/p6LqXEM/lvvVNMVCym6Q
FXKuWsASBWF4nngZ1JbKqlpeQ4UlPm3lnDGCBuQVOhsVGEkuUcQSqPEe8Y9B/rWd
4WTqfTTRfPXmhkJYPsZtTQJkY+1Iz7viMkGyZKluo90yjOPbwnMh8vDPCeR8XRG/
mjSDjNhDNgwP2r8cf7m8nlRdWirgju20eYTn5TJaHuD65ybJvKPwrfpi4z2ulZon
1ldR0psp7jTiUFbpQAyeZ566I9Q1HLHSXMwxDsfbQlY/6I6gleoooPjGOV/LlsUc
INcW1I+q8sQZq6GmOzHQXMRsvHW5tovBAw+1B7OMZ1nuRFuOfC2zLLmu06m1pO+1
pfpGriqLJj/bMm/XAb98WTQqVK+IEdCbxDxXfUxtqx+OhWPBIuUx9ce1k0CRmZtb
uqvaqo2pExX85RNMMfAyIy/p1T47BUN5JHQoCVt+JHnRIBPW4H8pwpZl53rvhXIA
th6YJK5jC8yTSU+dyO9mw96A0J9ERqJyFZQcEq+N/u3zfue8XBguhKKn/6TEwvzO
aRCW6243EkHp20IfwSGBKJxjS32gp/+jkYdXTWu5uKEV4dEkcmpAHg6W8PoiLFLP
j7OxauESrC4r2K/zaiafr1SY9Ud94YuDowFuW1yAzY4Dn1pcgMmk0k6j3ZIqxQnA
CGr/WGs8nCWM/iOwhTzty/ll1BQxpWwhfRj+xRqAT0+MaXIApsv16atmYBKxeGQ3
x/4uLhMbJ9J5nwncZ8BRO782v2J5atuDFqLnxMx9gomFoUVhilQ394U+ZcDKxTTV
ct1f4M9cpPDiHeVgFTM3gogcml0HOYmupwFA66YrLipgNPuICRjaJIKYsKXc0eaQ
54ehuJOHNcB6WE9DYk/OzGruOzsFYv+OdXkjxt7070972q/NKHXK5Kb6CKU38kKM
XL9Tmpd8DOOHGdOiS8WsEcqb8D+rjGpCXezfCkmbfYyD5mzwK8t/kyRAbBpQuS4i
cNpKIvRoZGIWbmrvWju2HQDoCY7sRcw0t0hvTDMqGxaIcXQNtFXehp4z3hYFgirm
ccsKsBpXznP0QpMpNG0kxegqF3wqkEJB2EaRTd0AoR/KqdCA1x6udcwW0j//KFUV
wSFfMwuyzOxUurLDZv+C2sDGQX6CFk6TnCzEnw2laD3QkcmGz8tHz7yLHmLcN72K
jH/7JLG1+pLDlacYkKM6jjam1ZlvGtdbIcMcYAg2mpex8kwu84cODjQHSgptgap5
Req0tZHryOL6HK94w+c2Uxrsg8jtoqdjWEzz6rG5+3+iM1S3NnWdZTtifhz2Zmhg
NRwnIRw5ZoGkoDuzERgl6PvT/Gs+hddvgaeA0JMFD+VXzB649SfwKf4zMZ3JkNNM
qtJJkO9Eji9gv21pOHf1u/cyaANWzAr8jdgq1lDc/dCe2IOA3nmVVr/xl5pUf3TP
NeT+SQXb+J1z7E46Bv32caGwEnX5809F1JbwQmTXia12203PGYSJoAZSIzTzg9dM
oyYpNlwk1Yd7WlMX8YSBllbvNpfsW2VkS/JgzYnbRx9+u6BLiL3tAjOE4EaTC5FZ
EFowQ4kA5jJCm06bWddJcAQgkamfC9/7cu+Paq/k6fFFf4DaIJmPsnC0PGvo7ixc
iwAvF6rQKQwVUlSe5OipwzOF1cu7BA0L+O7m+I+N2XiglGhBTdPS3WERRhY+AXza
lPN81wj9bTOCDzPvdH4OvS4rZdHNW0fzhfyg6dVdDQfIKI56KLkyfp+tcPaz2NHj
fOsWjhKmjfzsSk+cENkoo76elDCYL4UuaoZGMgUdIuwksvKO1pIHeby6qXvyC+fi
Mi71xrgVii0VcdkLZNAQoe5ENWd0M0jslDDBFx7UURwGg0/5n9XIpoPM39oQlenq
lyFq5LlQ/RS8oK/zSiojsDE/tC54r2IGUoQgNBFD7aTcJQW9nFfaEcmwTEecN/1h
OZIS4nOSm4PPIsi5mdpxzudL2Cc3ta7RjQ3HPTR75/Vnpxd0Z6X3fBtT0zbsrICm
M+e8isLITPibwZY8h59WG649Pp3KwpiIs+EHQXo/6Dhey3576ZEhBa8Dabex6GiK
SE3rVhF+UgyyeeuJOYk+aZDfw0f9VSVBm21ieX1cHKq6LV9vkj7SICbkhqLNVYVY
r8967xxEBaWVkrjRv6jP5dETX8OVLJFROAsEV19hfA0hi0IUkJizoxzfGCTdMHLD
9oxCNtC5/EwaCXrbPDO0vaT6t7Nhtz28Zp75elzL6wUSeLm3iaCnk9SsBHghRlbv
hwF7Aw6qcaIxzkoQwAnlykrzt8USrPGLAmXsUjaZATHVFoFZw2sVgOakGHpI9EwW
XGtLRPxeDcCGCtB4k5k25u1skUxSKDaVtTQU1WCpNHNfQSRCJAHB/pgtqA1ijdfz
oOx0sW46v2G2k5QGqHu3pxZufmoKqg9kGLi7lAu/kVlSShXJjcjTxhozT/5nDQnY
ks866lmPJf5DQuafMjZv/+jwxM8bNPVe253iSx0/jtTV1JdTU3pxZ+R6RnSizu7q
SPiDdSEMsIlYFLK43PasiEzXNI5KzFUrwd2HRH8SW2/wnLwmF0i8/FTyfSScbgVv
h4x0e/DhaWe8LhLibKaB2lGROj0y3s2f59BX/ef8bNURDTSSqY5islZeggndrGF0
0s0rPyKltf72mhEN/JPR97H037B85Nr2t9qxNELdLIS0NtZPXvXnL8V0QogzmQgn
iWsM/oObfQO80JN2N53oNxFbY4pZqGXqExFwTzUz5b/BDgpZrHX2XtgVqeOkvrrl
pULtG5HfNeDlOTaZwBv4EFJ+s3X39nTaxNmnAh0hKT2vJLN3hzsh8nrnj0cXHumh
Gbut7OVEmIF9HwI2gaCrzry6ZCrzZ5MPHUMjDD9bIb/Wf6eWJBYC5NFCo7EHPgD2
b8CvddVBPxiZJOMU1ry1yOLANU3Lua9j+3VdmnvbcegkPB0JjAGuaPKiJ5oRLwl5
u/DCA4ep0lJXXXTS1llg+Hk/NDu18heWe6Xs5SS3acTBmtomyX1+sXEO6t/I8kya
7rd/kek0Dv13PuCBqbOY6Ff/6bYLQp3mTtRxDZLP9rLQFnPBa7nldpqnjbxbEidW
oRaAUGOS0k1LTg8NgtjMvyYkwPHjdl3oG0NI5zgZ0C+DhKZnwIFJGGt2tQ5SLgL4
ogjSvvQXxOVSBBmN/YklpJCJBqhYcMEZX8mQeMNNfbiDDge9Qw9pIu4RSXP03XD7
fDppLPLC1n93lzjlekveYVxbBKY61eI6Pe245t5Q2X2xaARY3AiXOxcOPwxrWMz8
061V14B2L+D41i2E3F87OiSdm4k2ldbazlv7YKPcgMFewBBb/8RnQWsYPdE7PpLJ
0qydZNlr4Zjh/04+BzJ6az3TXxyVa2HH1g4NrhBftElfqdJI5zF+RYfPkodMIyBU
bzsV4lBs3GzcB7fM6pFzvq9F9kmoR9/u6IUiNU71GEWXTIlbGKu01Za2uN2Qhz6X
NP4MHPs58a5iy9grgkg4HyVRWmwGeDgQS6mbjoWna4Pq/r+xDHrEbvMn7QQ1nhZp
cZ13UmkN20kuMKkzbKaWBEznwZJQTcQA4L/Lzo2QcD+Gs06ZLxFMnbLj0R+6s5u0
dpgXhLtKAsEMjJG2pj8qFn1I8hY6SGgAQwx1MDqjC6f0xqmty42jCMg5DDeJGNVk
R9JN6NFyAOSu1x4a3cE+mNu9pPrj4WOZtwFsjhaPgmwVscXpfpXPrgEGtPJBfxL5
dzXGJRbj45223cbMKRNA5JRHmkuCItgVg9neZOLzv7dVZ3VtH825pSXZDBIQWTYR
7DdFAGtfTXemoOADz2+rQmwwJYMTXCxcBIe3MlybsMG7T1oTi2wLzoPepl+PYPfX
ydFVXELnAYv5sRMN6aSqMBuymNFf4N7ZiiuBkXRlZBp/BuK5WFVNN/ONdODDE0Rk
Dv2hpda+T63Ir/JHeDTQY0m8iMBouePiU5hP39QYnPMR2fECbMCEnbXVyFLuotgM
yVSdLgl4RH1HbiNm0hbVQSd/CzYU3luiF7bcuWUaEuOfAq3GI2FhX4PmFyjRdaFJ
P8w3EgnwfyNiJp6KkmeW4o3Cqc6Dd8TXqfSNXoYFnmUBvAyXUCe44NPFlKgHinrW
JFI+ukGc8+nzbMdPQkzIh2Mg8s43wz5dObtNp5RJlkZoqyOqjtcbMREV/sIHSvQd
WKJV/fXeVxqmD4OoIbGYGB5FomtvGBBD3u1kk9LWxKGqxud/UN6dWduJ2lqsxs7r
Z1+Z2McAmJXpk9u0q1svbhFhDL19G6kpWgnKFjT47tcpye3McC+Is7TH6IXFQFUs
liNopVGMH+mZ9lK1GP7wWEt614eu+vkCm87CpcMI8idebeV+ghvR4Us8Lg2qwQ2R
udkvGm64oRi6ocra0qmK56+Vblxo3DUmRbh481+gAV0ltdw4CxREuoZ8elWBJghn
E8swITfm0JmLzw+r/GzCIcWxjFbQyBAH59RwMVi3ldMCoU6zeMGe58keKEKtj2do
y7B+o8trCIP2vOGakKInZF7fbLjJqHUYCqQGkLgqVZ0Uap5wHRRlWUMPJujeSPgM
85E3NB+Ch3zRJzoGRA2xeN3df+ppYfk7SXfMlCLTEIZ+cz/fOPeiBj7T6lQ39uUK
d2/9Qg9kMgFwe9hjSmkCimSLhEXUeKC6z74WJHy2mJVYpSUmZr1va2Ae5twked3L
hTCfAJzuai3Kqd/iop2N3ILfZXkHjPlw9aPYN6TlBbbcVJoOB7769mpM3lEQYItQ
kH1sUUfcUqWpm2GnSKXGTOrIYq/QcPDiy+fMQT4eJKxPIzpMB4Z92Km26QCHIdEt
dsG1Zs0C60PwOC1QIciKUxLbfGRpkAFzeU+ZZ8oVRgXvWsZ9lTn3AFKyZhMDx9it
EGVusn4l+XLp8WcVXGnCk/J7XYlsTu8KyvGaJ6mbj+cDlJwFIp5Bn+4eokR/sJdC
1OuN2qyCBri4VtBfdpe5kObxOCdMmEHZ8QWNGZkgwha95iJvAS7IX3p26O7wBiXX
pyKu3Q19GZl4lMhjtrLXrT/Tl2mmgIwDy2WSzL3cLOukD3QPNXK14ktBc0chaINl
OsayjQZRkfTCiR1YWY0rtT4KFCOR2Xallp0nAiGzDqG847OKWXiFDqzWkwByGWXo
OPiYmojd4OF4NELah3w0OFhlpZYgGNVHSFPC5fN5qIUdqq4uO/WC67Xr7lKEg+YF
FdvmRffBrXDQQraqMU+xbaGe93iCdLDKpCcjqFg6KYnpv94d208Z5xCreoDtCzue
4MVCiXz6dqzD68QLMuTT9oagQX9MJV0Rod8q5URZVc4dnKmpN9+nQHInbuN+Eco7
TZsqdX7cxx6Ocmis02nJgNTwjkbKpTqNdUraoWafjCsUe0sT9ypl6cSjsDwCPP0E
nRUGYmHb2/OkvdGJPwf0DrAziqlnr3vEgg9AMDOgMnvAuY3befwSabbMcdlI2mjB
tmPzGpgCAXop12r9aDfWBWQcx//7HaZgWD4vqpj1C99xagSh2wfXriAJHY2EWsbA
9mqtPu69/cMoyPISRIu2Pt7hR8J1ZfpnbwyZ683nYSFoUUAm2v94xiQfkckHueiF
6lAt4JwScJFYY17hNJwYM2p/+0kFGGO3kDeZW6MjzaXlhga2ku7FHfkP6kKGFAbO
Y3MjUzPQ+6b7FIA4udP5o2OhTAGheRhNYtHwf4ul/GBLaYcMJyzDnjDSgl2CcH6M
8u3cWmEykTar4n/Ic5+0ODyiumu+afg70Ll/qV6qHogeWW7TjUykpwY8kj8ft0ML
lndYcxYcT1faUBq95LmXEgUlwzVuaWTbowMEqTkDdi9P7tLHgcyTRvCm/IjXL5Un
wkGPrw1U0qtXkNoM4ADG19Stgo9C4W61NwmCiyIYGJ8o9ywpnLKiH0KpCLuZFIz7
BFqEkEZ/3VKjgmgfPPA3BtBb74Vtr9fmeUy52bPa9Oi+PLdRTDuuIJXN8J9uPshn
JkfCBzYyslgxF/7LFSw9gXQH56zl6y80sr1CaCbR6QHhjugDYudaCYmx78cxAl3N
5j0G1DYCrEu+N1u+6txph5fGOUYTkLM6yvtwW8n4yuWScZ64vHJSRsUEwP4oyOHq
g5Xzb3SPnit51SSmav7FBqaLi9ZiieWQGI43CN79K8DhkWw/0LFm0w8u2Xz6MFae
Vh8oGsA2MZmv6Vu5U7U8kq4CW6yFA3G9vihQcztLyjQ=
--pragma protect end_data_block
--pragma protect digest_block
tRnJzH8+9oV/qVtkt18Nz1oXATo=
--pragma protect end_digest_block
--pragma protect end_protected
