-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
htRaVnZWS8hPJm3uU9YSU9ZPo4hy983UlR8TeW2z84Ox7vV7mzD2+6YXZ9lauAkolYyRvP62nZbo
HMIrhkua7sCOBd3VzaRqZBND0nqDSQ6M+Wu1qWNqt+wSLBt95hQO95cBdcUJl+5H9F7JlML3+rH6
0RmyhAtWmLO+RzsA1zybZTlFSP2EDUYlAl1B92YvWTEjklsE8ysY4UvN1DPBpsutnS7KI1RbRnBv
31UGqllhXXsMYFYZzMp2G8FKpwMAot61STfW2j0diBcxxq/kHTNGOtx/0KIGHcx6u4GEQxfp1unU
6JN2gq1FKWIFKv6otb7vjrb+g3991NNTpbMLlQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9504)
`protect data_block
QQG8hQKErnbmGrFHATgrqnD3yyniOZJgDl4gkKEmr1NeWHF5eA6AmuYnxijcSOIvOvEwm6ZXDzBJ
8z0OCtcdbU4a3cH9O7cVo9dE1aFgrCExvVSjf4FJIZeg3ctiQBOuniHzunOxtad23fZw2hMJAzC0
kpyliZlzlRE3ByE1+xSgvPHqLmScbtOxolyoRDHbkzAA18Tij0R4ggycmdD/Nrcoem1UjIeWRTK9
m+l0Wrzi7YCADzzlVr28cUqyUheAAdc2GaH4Xz9gQuS8b/1WSVsFGn5DYFN7oO6q8+fElOeJ4T+m
/ApYe35OMOiVuuz1Wvx952VxoypCZsIbcMKZ0RCY7v/oEBe/3tV3+a5sAC4dm9Gi+VvOe0kpbRmx
nRCfpIV70EkuBs3SJxyu4jfpuMHrmZgpFGRpwky0PtbsznnpIWyLxj5nYZkJPrWILzpDL7wWcxNP
/0i8LeYLxmfzQfCDxZf86gjFYCMbtTgsYBcvDwWxMDslfhbsZILAghX0c3E/pNbYz0b501zbSXeB
tmDe+TRQBkfkd7QOFu+lHzxpNsMvGxw46MSrdCXuIVP73OYaQDl/4NblxvDlyqtrR9XwMERg4kxm
gmsfO3SMfZmV3o+Q5IRT0hWhE8WALzxY92tNQmlI96FB14VMR6FnwYuvY7K8flVl0VMZ1YLVvmLV
fjgwWpAmKeNLP3hJWqliNXxzT1uRZI/RclSqjFhNvWTWw2COKI2Qff2zAnb9WgV+BugXStxbx20B
ByuuQdjXKb9TxZC9YoEsfEZaJZEBLoJF4janRIy1RYbNmNTBkQl0qqDsAIf7QuQydwyN/nTED9YP
tReTw0IfosskN26uePuEXZ8Zyr3D009b4m389gzZ47VfrUu0u86fHbR/8htp5i2dZJXR5c/XRLMJ
tg80cV8uc/70Zt34jT9RaaCmIyLCUyQW76UDcXJW3MvutGeOvbba359Sxlm5vmkukNHmY9EsUnMJ
EHyFykX7mh7obe+KFQd2v0qUHW5FjhiIP3lWWRojNWurrzK5gc/zf4t2KDbBJesQGb4nc5n/0Pz3
wClUZi73WjCAKIye27fw1gwNGmVEubYlqZuPR+b628XBD3NfVRjbY3vw5vhdl4EDOMx+AZBpSjZD
EHcLYBkieuEO4bwIW5+ofv/h77Km8jxrM3dl7BdgWxGuCH51lelj1Uh4kJPCUMk93+vgkdyw2g/k
YFUFp6Nxhnydrs1raEI7ZpkZxWLeSPJWYqRMQY9Lu6qKmEt3Ahf9WDI/Qg8UBERUK83bMIoq5wKL
W8kADKSgI+Bu2yRpAFogjEWB3FDeJiqQW9yO16aAu/nznorfwGTMlWbXi1ANih7cleTe88HQIpi7
a5Q5v9IibxeA3MPcOySwiadhjJPBkWGoDnJ5nQtI8dFtJPe+u7leEeAStdoHqXPuwCxgrxzlNg7q
VUBvcuocP00iPE+lS2B2QIs/qioMR0ZwLMTcJciHNlJ43tGI5TL0J4rGp6bwdgIqowCPL95W3Ds1
lktVrG1ei9NzKWWmOJO97fH85cJ1oomyUzUVUxBtXvoyWbh4KaODmrA83cCfmaDGtszdviz3aEOs
oiJzI/lvcxWR6JrmbSSXjk9tcHzHTa6AnjW8Tj/xCS6AUHhJulnir4GkIT/MClMRrveZrBe6jkaS
bTJs8DkY4OFhZEyrKor+u10FWkSXXi337fQEn8w42OE401ZLdP6CAe+mdpED4CnK42JS7nfRUFbC
bEBjwHGh9coxMG8LZJ4ibJ+02bo8rHMOI/XAmDMfVWI3ISmBd+oTrHow108tVzoqOfIs1PgYwn4j
9cvCTzOAvhCgsUuBg4HbhucVxWdAyXPN78jFqz511fB5NgecTQ8nQqKAZi4b3go2qRzU9EZ9PGS1
guZ9Cj28zqd900p5jMFkZqDKwyBaSf212ilIhWlCA4MjSgQ2GDHxY7WSWNZhH10Ob10PgQBpAlW2
V4uwJ+oRyF/CSsZSFsWWAuuDGZSa736FOWx9XGZlX3w2agrwDP3Q1N/hii/wpTGhRhmNBW2BwmrA
kdecdJgliCU+Xg+MsM1Op7SmLf0Xg8aZECEaZLHvTmDrIc2Oo2s4i1hNJaR9BO7yhX2LKNAUzb+n
BOpbYPA5wLhQzy9/COwPF8lEKZF1DyO5Thqr1gmVsNIRHog0By7bqA04m2S676m4OTu+5VHgi2NN
l9ZLVwSu+v+udXQLU3WLG0iAIiXgk+Hkyk6aSzJzxZeo6xQL1MjB/jDhiD14gsxe3uRFPS/50zNP
qnlksgZa6c2qtIwKUrH8J9nAQ3bOJN/BfFrdCn43DDrCnvLQ25qCzDsSxtmutrMm2GMz293exYxU
gzNaKo9E0ybeogaOJe7H+sDbSsb0NTvNRp9iF6vh1z9X3BwUikCsHLkqmT9xbr6latYG+N3IELRm
Q1EHP9eu7NNlcDLd1oR1adqiaRY5SJY4lnThWqNGlm9hEQTsgjbTfSrGNgcJ34Cqt6g4djY3E7vy
ZbhOo+zyNlpKKjO52egx2C+35cT2SmQ8+45kozXITm/R8oImVn9hpV82kPNjvSshLesBmg84KdSZ
mJ3mjpOiF/PYNGdU4Hts3Gv4v+8XvBDmxdvbWll+TcOHZ1fY3u6S81B/Y+JHVn4X9CV7y564bQcR
sefdIhg8i4m5wVfIpFjXZ3lBGSilPqmnLWddMZzkXh7Td0v1WIOuqiFpiekqiRu98mN9rpZmh4Hb
VlEnDXIGSYtqO8xUbPJRVOggxsbuXhZb+MK/f9ECB7ucP00owpFXckPwquvgWrDaFE+SSnwjzE4s
ASGenhPI6BLBAnX5CMaeaSi2RY2mseSY/43zxBCWULxDChGxWqAiTPC+lO6YLi23Xp6PgKNDZcvs
5gdr8jADMUXTxMte5ogDMdCdCGUcqjgd7yeuqlto9d/NuZozV2btcU8TLHKnMrYf6e6352LTeFvx
hVbiDWgPpF+kv6+R7nFGx4JQbgITRZvFkVJfKT0wVaf61G1WvazLk7mqVPimfHoF+R6sjgN2Hk/M
EAY87omslguIaSeSUtb5qNiMLc/BzdBULpnSysj8ncqVKq2kZQ0h1TDEQYEHD640ojl7UtxL0Ot7
Gzt8PbBMfudwzpSqc49nbZIsVIb13zIailXXLjf369QvVp0cGnw0hIIwiLuJSZ2S8EtsuRzUN41X
eiUHi4fOiwarCsvhxMnOl77cnO/j2GR9IeHjGjQapMi/dO/zYmc9lZ21HAJTKNxcTk+9VVCZILMX
lLlSkeUsOAHFkRwsjY/8PKg6gAES9o9GTn/Z6bhu8wbshBsXkY5i57U6xcoMG0RTVvPwoEUtr48w
eIGUg6BKIzN3L6bQDxaEErFmKA+wZs1seOnqpPloTDZsXWkmtHtogSIesBgLkqEkw+lPsCKWAfDe
yJJcloHfQ02aDhfot6wQBco26eSwWYaYzrGhTxip6zbbiVl87BzeRrDfFbsEnAYogt7tnzLf2nLd
wfRXRtoRtxEKcyG0UgisuttHYEgy1p2aelM6WwjWQ8YbouM+pIUdjkzdQl1QUVWSQDNpA1i8Utay
r1yOhShVDh81nqdRBNYtY79mfD7+Ps+ljZ0CAPYbYirDh/VqKEk1spI++ubVVkO65NqRhIwK8oIn
gLAxRdQNwlVTqiHbVasysKGGiXKPddpilaDPJW5iMffXsgiyTsmsoLeaQYfglhH0g44KTbPIxbLp
mVw/GLU/Y8XDafHXyX/SSIa+cT9HwCYJ2TdMDJX/7/Xj5TsUC9eKszM4T66Ar/4tJmgMocJ24tYy
KQNM5IlSeW8dtWrpLCxoWrNmX4QKTSlY1/ejA2A/vcqTsrv3GjPgTWabj2Ipz4nSwifjeECEOHjZ
UApjoisbU3b9pyuOcv+QfnBWnPEmybIDe8AqDQnK8Rixa7e3sJdGYx9/qRYjdnKErkYZVAarM3UE
rXmbUDom+rKsyur8x04NOiWcSpEYt9Fp4uSkPKx64q4QxvZdAsEGTjZ1OH2o7QKmicQXWtBZVze4
yuaBgeX4Kesws188Yk6m0+LiRKfJOCpSNdaVHfN/Ug5q97ZHy3oNmID3j4rxJkGwiUWO7ClKfadj
YfUrHEKHa6DTzAV/FwANELZ7OicoJFtwkq9rK97RAzwv8W9uVywt1CEW0cRbfQrfa/2XkaVci7/r
U0rw7TNuik8oSkNMwYReAqihF/VR9tYJQDPnj+9BfBDQHwdDZzTF0DuiT85kymWdFwaoB8R2+sNm
vcOCg4yb7TggQDjt9Kdu8m4lE4re69shbefuSUzDJBnqNRzh86hXS1tbbw0tzNKTtkM+m9xvz/nD
OQgRSrtybFKMDlLXGiXkFTjaqqfR8drpSwO5ZWXzvOacp+I5LMMLVxYYoph3W9BlopDAfwZgqJRi
Tw9fOs8sn5hnH1mkyKeIuv5fDZRvJlHbhnbouwSMyMmKlAP+Ld9wpTUQjuocSHYtwzBOglFB7/kR
3TcCeR4BzHOK8t50v95qT91FNccN+ga6T5NpwoiuoGGrrZf52zrDZPZSySUzpdDQ3WPZ14GdVr+M
G0VZyUn1LB2DucnZrxG33FwxUrsBeCdKcAp5dGl7e4o3aC5ypaRRoQkohA8e3NxLc7WHHe/SSWHl
PKw03jljfrpAoeYbQxgYj5i3xEH9nLliCgdOt3OGxBF7sGKKsOfiREL2wh5oKUBtrVqdmDWERkPn
F2T+1sRoZTboWy0qlyo2JmKyBfYeb8ekRUsiPJUHg2UK1KoBOpHzHEmv3DJ4G1g7JnVQMSXtry6+
4iIcbjkS556Nq24acp0lqWvSqUO7JaIg+k58IXYPZHNonaGgMcxu822rnaOfB4kiygv1Jmph/RMK
uQUFHFn2FDmAvIVI5w/cNX40hzvioOzwme+8yWURhmdfDizElonthNuGwrispCQc/X8ujbazPgPy
DuQfgdm3nVnOsdIXpxrAseVdBTI5vgErCf+gD4y9RaOzTs/CycfHPKWHWjcRiqtX4vQ2fMOxwnxK
uwo0YrBfKPPvXXSMZRJdQVnqK6LotPf9++4FVAjc/cOimffyXZ7jJGhKMKwy6DFh5Og+AWzkZZLX
B/trbDEmy+QkhdqUMXOwYbbtRiScRI4uvVULORtzAOsGs5xIiTk6hr7loik/H90Id09RDY4aG5Es
Y4And+IwuvUfAypXCdJWq1GSFr1/mbeJEP1tZzuxPSlnXG3TGvuIc+LlWSQ5UFb9kxAyC230dAL7
0w8wToOZrPAomDUcGb/3G+ceDqT7fQDz736oRW2hBBIVNyGDSmEZSEKtUrJdFr2yJJPwkX/62Aj4
zE/94pmPVGcypgBQmKpEioe9wvsedkLSDSbQQtbRaU+8MVf2ZKKTa4n0n+ArocqiOQxPAvYcptVM
dQFI1XBK/M+cjbLreX+X1/WguwL+yJgCBrzkCvcleI9+PQEjwWl7Hzx7EtwTVrKL0Yy/SukaecNS
5P9Q/9Lpm4X/GBXtiMZRw3xsBUDcC6i8oBZlAuIHzKwz2+lpGL2OMWSqISVvleGwYXp34dfdrt34
i6fjzYiWc6LyalvbsB6H50ppcwFBX9XQ+Bvx8dDGtTYxziZ2R/xpO2EVeWEvMDgUjqk49kMg7MFq
O/BJOpFN68LC4G9GyWFDvDlbdI78CnhsOIWrXUbqi5t03AqGmAudW7sZvnjIdPznIS+RwSYA7AEU
+HxPAQp0H7kDdhV1uHXFSIWkhJbm0zIMxOAdi8Y4DDrJ7vtfb1r4//RzB/ec8OU50bMsAKHG8U0X
dlA5zyZ33WWt7TzoYvrrqnVnGdlwR2/NuFJpHRtkIThakX8na/PERvZlVDKJMMdvX5zUu+eVHJaQ
EgSFZcZ5rjk/eU1AjW1fyK1BxF4bSlDPcNKrLGF5ji9zIe87MEyWNRvk+NsT1p8NICfCafv/lBHe
zvLVaeEzG9zLiX6WG0exQjkfEItunaKX6mod+QiBaUnvcWnnGA2epQ+v4Y/AwzLkrjtFOFkKYeZo
qEhfHCI8zE1NE6GZlggi1u4efuR18pi805NKjAQ7/6fvRUSIMVDttGcuG659B7NmvOAyHZiKbSJ9
AsF2iiTBtJK7LiCUpCV7U2EounAdyRgjwZi+YAMPwTmTmxowLUt/BY/gBeE7JepHw2M+7sysfR9A
GHf7BI/JmuOrPyCacX2jscwkXdNr5dxjMlDGggeU+MCTmJaf82BnTInaxjuF1JRjOn+ap2Lj6jM3
nODMQPjv3pTLNgnsj/kQOC/Ns9aIBFEMsqa/RaqeAwxDNIbODPWHaXf7YhClr5IOcih3iv1sbbVt
oVMzIyPrU/ribkQ82b/Q66sg5h64YpyObkchi5vQAo7DgfB2QDJIJvzSGurRZBYK5pF0YJheEOS9
6lLuVwbKZsQK2n5v2DelA0hcMckph5BXIeZLDa9P4JmyhlMsnnDBrJBWZWlMmAXrjSaAykVaBEJn
vvQ26Oqw+cTbAxrVdB273pTn12F75L68IX9ZRLZ8g/JjfQbvG/2MSZsxjY4bjwn6NSbDOW5s/sRz
6O8Sh8UJGfyYvQ940a6RFwoPwafewXlzYPFE32uUoQrPz9AD/SJyxUycopPudqDBUHHdiCNXGWf/
XAaGGCcVPeQzPi0V3yza775wtI00LmaH3KlRTowpPOsU3TdbY/yNb3cSL80CwspyHWQJ+OGpeZII
HLPGswa0eRBosOD0RD/hY4o4LnGGnlpTHiRwBCCghf4GfUuGI6V+LkU0nawCNeuExGBUrcaIQlC/
TZw6AB/dxV8aKn/hiS755/Q+ZKrchZG+D9SYPw2eN4V7jb8ex7tbR6YoNYBQyqwqRReZHBDdCTc5
SCVC9ew28OJtY/AQqzP0tn2OFwvxVz2Y0aZpvoJdcR9R0yo8G7Bk6au+E6l6ZszhOuHvHK69TWj9
j0hCZBSOi/Qzpce3Sg3XRbW/hT3aYP17n1/6EkPZwrnH7NZfZBjxVaYB/zoysKFcIKMtHTsXdF6k
2NY2vIikU0PisN0tPvmCbKKUzbl55vg6HbPoBE0r4j3L8X9vn/xSa7ByoOIkIHnDv8HTAM2TNpZA
ceC+zdeHuuIRIinLcRvptaCyd/mRSTrV1ZPoNCdt4itEluSWOQCZQInEROYMUXiNBO5kOvatak9q
9D6yKg9p5ZEjM0AMJg1CWe0dUGhqiT7W/ZdTn2jsleJIv114fvpVUXXNZLP2bvNM7lSWYPlPVs7L
JJQvVFu+gAprv5HlXQ8Km6zyPwZabZV6Yqm7wqJJ6qXpLEMldq6Kw+b4X6erPqLeeBl4taoBpAMK
Z6t0/PQ/BeQz5M1x2gMVjGflJj3L57ckASKYQd0tKm7MH4OAG8UBTnlPoy1rxCoN0OzMWvtSoFfB
HGOvDwQXmUQh1xeFkVGFICdQRoyFvOn8Tnn+XXXD845MGVkQiSADghE4l8Yvres+iLZjN2uq5p6O
ewlO5MBxX1bjSNC4XGeu5PTL48/Vro9tUg+n8NCVTmJfPmztB7rsztnFalPMQgMJFz784730uF/Z
BSYhxst0pl+8cDy/wkUMOI3+AWhstSBMPKdFkomB8biDgPo7oOoPCEDkHY7SsTz8embeV4uoebJB
IQ5kHRe5N5MzOQ1PbhTXNJAimwQgNiTKletkMmKhO2HVpGlb0H/VB2cAWmBuBWBP15fDjHzp98jH
YHNApaPuvkcZPPFjugYisxiPFsTlFA4eXmT4yeanAnv90DFmeQwUG6WpW4vLLEnF0XQCCZ6r06pe
1aTl6Rzy9sdwSQ9HI4fdIjlSqxGe+l3tqy4OosprCQir1YRhPAZtqyiKIAhrYA7aXO2KUUX886XW
MdmwC5Y/+P3UO4eDdafK9TLc8s68h/V7cT8q2x6uxacA5gQofksJzDM7gUDajETGOUUsN+YcQH4g
vGSSGZMJFG1b6bCxRzehzZ2puPH83j3PRfpLExwIwhK6+52ORhZmG8+JYzRgbmytCrXyu6cWGbLo
n40U2wtbjxLenoYgnaFfzsdhLbzJkcSqKWVOETJrcrp7WifxBQ87ONcz9rl5OB6x9tznS9YYSLIm
pSgCgT5kqLcURVlFJLs9v8pLpWtUzx4Oj07oxJZtPQEUVkYK9wlvlneVdfRLpcGroVV0WQoJ1VBz
UWF1VAwgaJJaXgJnyW4nOMzg39d3moN/X5wQ7dIperwhkW1wtoUCyeOwQvpC0hgIRhnfu464xHqE
2ftcDXiwqKuF/qLzDSBOVG2qoYECEcMzNl6k1BGDMHSnfwjMx9Z8o+ShBA2V1+Cr2AkMv3APp/kM
Sgrjb283u4gR+fKnMZvdSoHKMfFXqwJMzyIjmBXl1IgLOg5FfLL3bDip3Q4ActrGBnEwnCoSBy2V
5jJz36PkuTelcFpAPHJoI4QO08fPYhSpzWyB0R+A7eCeQhiZlM3No/MXANaRD0MhLNVJ91LokPIc
C1CKIDi+cn48g9IJ6UuS62ir+nDUv7wEgPyQ7W/ZR9HAKBO7oghdGoQX7RNdRBvo/1+Hu+Dibvv7
J/SXAj/SC2iVWQY0s7eaiPn70uOt/z7w9XYtbxRKssWQ0viN/rMj6USXdhsFgqF+R+gQA87S0/dc
u4rZfLyZayuJpUVtXwG7uJHVxn8ILE+d0cbmc/u4CW+Dft3bU57fEcDDnQHKtTWN5Xn0JDFEAS20
uTaauUh641ngBvUeo/Uy/v1qAAgcdXIorbouAPgD+IzL4/oLE8+CeqI03qCQAIt/kC5xWhdrURU7
NIgSKH2NpJeMDktF1fE58+sAJV0XDZau89eo3aIyXRtoOXZfw45DkREU6ZHHJfYCvcbk4RI8kDhQ
/Xz65ZpZOHFlLzKdSF9zNntSoPTQ6NN3F4TS2ffR2lNpEYX+gtjgGYvJ1J9yTt36Nu55pIO1z/9K
fviwStV7tPssKOwtxl4HdH0rbF+9qcsBn4wRxOklvZm1kCd9SD8AKdBlaix3ACKWENcHWJ4sGY7V
88Wdo3+57uDawv7cT7aPbwg0KLyb8wIFrV1IGMRJEWf9IOxB/BXnNOz0Kwq3lFqo84NZ1xXua6sY
IRzDwxmna86OVWW/UKkJ0pkUKeOU8LIOVihQ2O33CawnMoiG3WmKQgVHS9N7+kTms31ixUjRJpru
F8OvBrmv3Ae3b+kdswFUpAgwjzHxo5wB6shxmxI3WPPAzz4IAqLHAp4vOXwa7xAKWtUlOmYsa4Ta
Sy+STsAUWXlXG9fiCslfE/MXXcLEg12ta6EzU0O6P7cirMUgC/ZtXG4e2aBj1ssoKMbSfNXn+q46
9oT5qT0qGU+yiSX1LipolNLo+3/7+lwATdpkz/7uwqqSFEU0qvhZYJiIzzopGhcnFudhlX6ygW9R
axQgVDY/uVR8gwXHsEQNa8M5r/Rn2HueIH+MxuJddEoC5pmlff27BlqN0anCEdM4qELcicExRewK
2o4Z9XqP9aiqp6Cl9ll1Rhm9xTm9hDBe1ZLZifSCcHQtgwoeZC48j4+2x6qKLeCVIbaD8JVrvd1L
pv0R9UPmKFFHZD/SL4aHp+5o315he39D4bm9Eg+ww8loGVxnaAPxbM3WNb0odtbTadAmDvw05iUJ
pPGTTSi2x5jNM7hxylfV2/igcDRu70WKXWFfRvX63P4JLS83SunMGGKrLvyONw52F2y3Y593U4ZY
86ubqYimUqyL3v2UxrOms6juXumKhNjmIekR6kya5a9P6BZVCNMHU26/bRXb/0M2ZZYzj68oF1VL
vY2mgAvx/I6h7nYo33mhfdGSoVmhD0iuJkOQ5D2pbRCJ4L7hYMWvHltRNULWoBkWNrcP0I3AkvV8
2YrguqY8gzz4ajncP2gZklFhJBF9eL1Xue+TWTtdmSNogYICIvgCt7zheIBUkY0OEsUtNvBzeUHK
7RZWasHKc/WGAyznIWmERkSU84CPk3334d5XWZRWt6Bi7AJn0R3yqoO3g4AUh5p379PYGqE/l0D2
AOO8m/arBcXVeIx+3OtitMjCGAi70pz0lrBi3QcFLi07lEJkPVA2VzRetGeDXBlKasGgZ1gKJm7H
h3xgXq6ROJMBTjCl+xKlCRdzlS/GWPxoigIrjt+zE03t+bBzx8nuiBRGXkcDUZdGGDwaSwqMsMO/
u2Vf3OVixRj2BIQYZaiCN+0+POODbobVZToSNM5o/aUE3LjF6MLxMRDPds8dRa1nULlmpxVeO6A8
8hDK6RWXImLdos7zSLhDmft2EWPhANJ2iMHSPKSdO8m1s1JiY2ccNTGmm/XcEgbkZcd5un4SOCvA
l/Gtsiz/FGon4yWilofpE2ES1TvpPLcSD9KrcAiKNC6PnucgpqsEQgwzULUC5BllmS7uJ/58ckvs
aenZLvqImAN/cIC/5HH0YlUEB8HEJcgsBR5eTPLNMPYzhQWaMfySGkSEfp2EXTEYrNTBOENqZcQz
fIjA6+2FOAyvwpz/1PEilDMHxBxBhlbeE93Jsm5efWNyR3UWkNSbrRw0KvSulioCFcc4yjElaTuz
Is/xEh+TpuD78D7IZtfwMy3t10+2XjJOIUPBGhr4UtLyovtQOGpxZRY+WLhvxSiQtHSZXdV1Vxns
OdlWYFZdom4n3i+q6yVbDxONH3PmTYcX1muNQxSlvRlYoyUW8/vhyhScN3KSDt5U/aJ+ICBmxV55
gNKMomR3pKE6tSTlsK8gSXk+TQMWoGCFX8mq/6wOWighspqb01xhJT2JNkubT53OkQMfQxfC8rBN
NBxggb1RwkEKolA5wQYsUiuTR9OiXdb4qWaJruEZvL7GsoBATRe6l5jI+Cqs4CYPU3Qe7hhYGyur
cP6RdfD+D+FJikVZ01JgaHPq04IJ3b2CrkkMNJH0bwE2WLb8pa4H5chH319PfdsdILp/mdNVB74n
lrWFkX3o6vh7ThfdSJgvBDD3Rx9Vz19nUKh7bdCDjdv1rkro+8p7V52ZfCWx+Q2P41B1OWAkk6OK
soQ/4haCVclUXDPOyGmw2NCXElLcHe0OVz3FmxyQ1arhlPYYkvzG5WnLEWSx3deDEVKaGFF7ovvj
fF+WJQnYhtxu1mXTQGbPh5mbuyp/Ucq6RCFnnksiq3ErxOqWKNpmB3QhwDWS5RkHe32RmJ7hI6fX
a4APV3oww2hm2hJl3zGE/7YNsm2O/OitPIn/8a46dz/MnleOfPrxkl6ynRZlh+0z1rGtS3Qv23Xw
f2bmkc5Z6ZZgizxGhePUrllWbUwarT+1EqpJ7fie8hTNMPH6jfplFUz6+/PdrPb/FCb6PerL+ETP
Xdg+Ptcr2xF5U8bAZeU/6rK+aHtZf4uv915tr77xKVt0KbNc6UaIa4Z6Y/loQz0hagYM8pwTMmis
urN8QubbQ8dx0pT7ApW0DLQw0H3eGrPoUj0I2U2JN4J7hoPJR7YvvDnyWay8+MAoLVQ3k/vmpuf3
Y+T2cHPukjZuUgWgDXGhfqm35FVtPWgDmPFFYDzuqfPB519Rye/c03tOcBvbhsPNc7JMxyoco1kT
IF2wTOxC1zU+Md9e4rDNkcwbhZfS/dvku3VQLYGlUFrD9LLFwqgOL6nWARJxwdoFe78939G/OQns
5+gp8m6NXhEk/h98DH56beOnAEPklGgoaChL8pudUNSY6oVm2X/2xkZfUBUnD7+jpFKY7JC/ETc/
YztMxrC549QAPMCPlhT+kINC6oHQU2WFkZofXNcnDXXnBEvhz+7ZOy6hTcyzBWT211T9lLT/a38A
sXGTMRZULLhMJrvuvPoDllQxPAWZokNf+9nTJie00cd/72qSqMGnmRJwebBQS50asb/NpvsrYnJH
ZdqDP4NLhtFgFuzTaaK22Mo3E4RjCHwKRqrMq3KFNiTzfhG+60Y2TFcgvOacnM+86NiwIYmF1o6a
ewEQyEtLuETtcKLtQabNsG/0AgR6kqgqIV/uEfQmh5RXdAhIOK5gEGlZeMPePPKWm6bWBx6NRFlt
4QFGw5B6oObbOFxdo9mavfUiYGltR/WEhVjovmInYQ4VUR9I6fSWTSLpVaNZAoBxmP3HnYl93JhX
r5YqmCD7El0gow4itcd0yS4lEBCXLhlth5F4Rvj9HpjJKw6gX0Yurj0pcqhxwg+DCElxQ3yjT6E+
W11lVCP6CD7BuCNDdpeF0gbY9isw6dbcNb33wz/sfp1GICOszv49pj3l8M97Vek0y7tgCXse03T+
LvcRqLaVHyCMoZT+RzfBCbOiE+QMrh2FtXvVJpy6fJot/ZQC+u+wTiCy2BbYnnsB8zV42DVHhTPP
1+gaW3zJMX+cO2jiDgoXbJkDZiNOzbGDJgIUOcyosRyCtepgAv+jOQeLMwUMjSM7xsZ32EQe9nEV
8Ja3pANriBemvfgvUDJ7yEbWI8L2ecWEshnBKRgrVmhAPUe2J0fnHhxYvXQUlXlehhb0ewr6tUlA
txEQO1MstcDSXVOmoKAOFVetmF/jyAbZFR9D0b1z4SwrOB895WOfjLQ2GiTNnYOScRSsVhFHBFH5
Ufkv+OaMmyW6vkDWXSyPxd5by0ChcJgT2O9mDsNOgjupXOrtme9MfNiGS5ZuGEV/LjcV1zhXO1hE
JlgsfcmAlRU6QGYY7DQEZCsGvK7026dFXRALkwKrwXwzanOnuQgObjr6Iv4/wkWdItFJ6SCPUNUh
SXi8KaN6DuWAMljKUjX3exY0GxFYcL8rrPjB4+PEyNnA7r4+/bW4iIQI
`protect end_protected
