-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
tQxJvU/ijelUN27a898LHjpDiGOaIMqmFjuWCmrF0E+ZgCsk5HH549UeS03eCEw7
NYBCcnDvdtJAhSUXz908rFsKMs+cy0VgEg31O65/EYLPZobZ+Sl8F7Of70O5XEZS
xFeq2rXBc81mAP2AaJx4sip5TyIjo/d0n4qc8DjqTpA=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 17152)
`protect data_block
9mRv+WqgZF0QitFh2wPYTybjaPh8Nk2zyM6jLXmrcHY6IRTwV+0NI1Jkc78o28Qt
kWDKvHXObGpOne4JwlzpaoYqFjNJWnghyF/kpZWCKPwMuPsnylwo/64IxLDiD7HM
RoTpeoPn+Qt0R+5u6L36UkT+7ANVHBVHQtrwcRXsKnaIg5Swu+kaQXkhiR4CDEdi
It9g0y0ZEl8E8wlIzJ3ElLdnqQMuFpQBYd6jyHLik7ZHFc/aWydhAH0ivrAWuXdX
yAT9X9eEPVARgSuxWSakkhdLk6wfE8xb6lp1vTGpMXa4W+ScH6cTZ1uy7Mt/hvBd
IXJdg8Jfg9Hktjv0xCo7tg361tFlU+KqXUqPZrnAx+XC5oh+pjwc4+QQB9OXcPt/
vGmaoW20vt0u7dtYNaByadZxRCJ8/v4uMZ2H444/KGjI+UdZYl5SkXfAX9mOWseY
QQtunBM3yMOzC4oeJp+EG2mJvExygofwWFCz+Oc9KZAJ+J6BZYb46hSIMLn87ZoC
/6cvgCeLslQfGcV0sHYve151NtSxEt/YN+LWLr3BXFsq6YK8AA1AuOfAFb+czGJ3
jj9bpBBpmJM1CuzTVuNfDJLm7eSK8DtICMIdEanV6kWv2WPqXz52UiMgCgDNlLAE
zFmv+tbna7YpVDD2qGYeROL7XHib1qMtEQtdd9RAk+NCpIXmQAcst7ztsy9TFkRW
YG7qVb14gTjYA18aPCX4Cf9F0qr5VNs73rBFTUDF/X5wCUPYDn9Lq9i2yoHGoYuW
5c5mZSjqIpgmNvwClbwzh5ju4ftjWdAFBRDZXGBfUqYK8RynP5NHyDBjqeci3Aim
fyeuLhxK9Cq29rLclazYx8jQkOEWulZqR4ijAbWWkCcDURyd0DTaPGo94v6KtBDJ
LYcKLvxVgWfk1sI1MUQdyxBgOEueERv/0+resqDBFr96yxA76dLDm+TiEbINucK0
UjATLaEIydThoM5eFV/X5mCJWctC0ecRGkvC+HoYkpu1YtBVRqAuHT2OpyWtqAZe
rcmkfH+loSBlk2fyKkdGD17+vN6kc3uniCNkkYn4VqCgJm3LQcMDFfs1XiLJzLaU
7hR8ATkczNDExkEozGWJlAoUzaQt58FKmkVE//nMcbiz7fiOLDy0zRKRJygFANK+
pLkjBBgfwyRfjM4h/Aa4kBg+BC8ITGLovVBOaYsDQhe9euS6EL+iac4wylpNCGsv
iXtE+dGClCicROmwOUp/ZEv+Y535/VRyTFYyrmaVzT+p1KHNgZ4Zrb2JY3Shho8s
L5zZOY5dgNc0sAUqJ5zdeGZBZCouCg1EIjU1SJwhT5eAiB5GMHN6NnWgTd3TaYAD
yyoYMGSBAcleRuXO9dk4BPJ11G5zKxUSi7l1QuQdaoT9ku26/2q6AfZZloJgcilM
3ja9UzzDQUbZe7VptfLKAqC57+62A6C/D9e5zOVqT5rxv/sgIIR+J3U3lPXczutQ
Jg+llWQBBs9wp0l8+fZfHAPkJQIQ56/e8VhwJE0EyTce6kSB2o/Ud91VQbjVP1Fe
XPHB12kS58OlkgE22fQcB0lLWk8RRsmjrndnmUDY1Fv8IGjcJiEoz9lURR22yawC
YRGyl2qbLwad/Z2oEjuUzzEstC/VH1GgTTlPl2KR0mm53JYCWC/zE2TpGeHMf1DH
HICNqYYo5SLc8fEmnR+TJd+knGGQbOvLGwPJeHvoM7aoycnFzdkN47vbmp9UDGWC
Jh6v4lx5rB6+pGxCrqNICQ9y6Z+LGr9dD3aVQ854Vf4+NgTYrURH6+MPjWsvPpN7
CTijbIc0yzELlTGccQvRuZaYxDhGqrjaPkUrS08cTxk8ZIeYLo4eGkhze5FqQqwh
U/QWynhl3AU6rmBVabH/0Ka+iWhLiXPNaEqU/8Yn+i//llfMVToIDTCBsaT/OIlE
rbBqJBVfaEDAM93bu8Q5Z4GIBEw2oPJFZG4T92hDxOTPP7xyMTij1Da3G82GHmB0
9J+DgOpE91xLm7WB6yTAo4+KLZ14GG9myxsPnAvjkJL/egC8uaDwdun5lwSwV2Ev
PjPqYJ+pSZvORHE+DLk21S5oNxaFDv+5PCDEgCYgxiJbZDYDv76mtKbqavHjw4A2
ibQIuIxwp0Uto9BTrZdBoTCf3wOS9MLqhREoARun/SNSnwOevSi+zfIyxzpl+pY5
zHxXb6DM8V1nHqMAJNzKaIQqe5YsctX2WgLKVYaCn7vwp4zdfweB41cimYNBB4eI
9JQ2JW6HmRLyC+CGkmcRfnIbOSSzLvbvHIqe1V9v8AXDV40AVln9WDXwCczFaiEn
TgG1/NGqz1VAtQwJFnQmwa7OMxgdA/JJE8og9m9+A+EpnMQ4gMJ8ZIZKKuhRxzED
3exOOne7WK0TdKpV3XF2FrkVcBNuGCOCAjxLPA4JYW0yuLk0uMsCJwyoH/OVWF5j
OUybxE7/RIvFHWE++DnXdRiAlHnmGBxxoHDFz/8Jm3kx63r2tOQMSihVoWAn9nNt
DfxXuJ8we1Qdl25wMhVDw42pHcjNdOXu4/YcMk1NQ6rjjhmF6dltrbvWAmDGuZE7
Ywyjjz8jrGvR1LZ5XBn6PSGBYfTEDFyoqrLc5GMD4PIkbne5iBdXHInDCaU+xDAQ
XYa5iDlepyyiWPEqUMpGiq9PWGBeFvb5dyXAvkp7ClE78ROBPazwQpDgzcLHSzxP
mTvyvElIQNH9eYyAeSk46rA/hRkcv0Je4ektnQ0fofclASo3agW7JiZeDBDY1EjP
wNScl1VfMGTapCDNBX3wPP7utFWqio1b2vLsVjc5hCE+Kgkr1yMOxTEGHVPfIMBp
VkpZ35JJkZWZCmKAtcAkX2aTnAAGT4z6nsNBBw83dx7CQ61FRzF1BaPCBdkNCrQV
hBORiWnMVFS2yxO3k3kA3/lSdWrxezYDcsVfh+gOfxA/brZyCnyhT50LdEBqocF6
aYmZMDEGvo4ypv9ezAJ4gEatCNaZQAvLsUrzwH+DS/5JNishw5KhdqgygZ7xA179
0aMNsmuJwYxqchun5u6IQths/xqf72lKloPwipq9r4+4tK5ry9VD1mgwQYQjATy2
6e/N2uit7S1ji473Si7qdEFZXPLkdU+Q92VBXpde0Wwcqhr/uWmdTMzjaL6mGuUI
NfkgPbPZlx9qph16SPDwP/j+RwaYE1tnbU/Z2C26flPaRnqXF+VQOCXvTogPWrxU
dpxADDMCm8D3kw1i91oyRbnBfXM4FKfy6ABNr7B241qMs8u6sDJpa491Scous35T
r4txUZSWil5EnPQSq5i55jedzifWZwtPqkVpEeomlX3PW6ZjVpQj8oejfavBrZhh
3CILke40PXa4f3oqOoKcjndUloclxk9xr986nCLhRWA4VSTPlqBpRaBiIMd+b6rI
R59Mt3N0712B3f8Wx0cr7NeV+rNtpVUo+fMDXF2Ave4PIId2jqVWazGmt6eOqd7I
BZlZlFQhEpaicBUi9T8Wh4qMzNyLJmH3ZzqTyq/vXnz7wOsFRTL5PvUZkFCrm1AE
CL/rgG9z4sLXpuyFis/H1Qai+Dvwwtr3c24o9O5FWVok6yMiuX4dDqNcFYf8trDH
mmZVtHpl69ypPrvFebrhMyHsQlhCxlABYEdsmK3DeVTcKIBBwnallnof3TjsOEZA
imJ7ZnZ1kCoVeY34bL8Q0c4fsmyOr3QJCN6+sRjf/uOSqzSgXCF1v1qFTKVZMjL5
pG6FxLmW/fe8KwuM5MybJn0AZSAczbj/EUcAHCLFA1RJIiAIkSAJewQ3hi7MjKAr
fczUpXwzY0jyxhXN9/A+/b2BEmdB7UkhdhscTUV+eIMDHVxeYud8Go44++nHGF90
3zobLVoGEaA7syzs8AXSLX45xLlB2Q77PyvvnoKaqFhgj5/R8ubsSlYGEj9b/ixl
JFNLKeVVtLzxELsWClcsBzL+6aEL9ijqTe2ohtBdr4pU4DG7RqppbaDVzsAZZg48
+R0SdF0WqhFx4mbazCjrn7OKTIi5sx9ycujNJpxzwxhBmSJnnm7wl+Egdh9QkVrs
Vgi1JW17v+bgxFgdoZ27gKcU5dkJxhKonwut18IApaNHVWL7wB5HSLadSKoz+h9/
SaLOF1SBT1nBrpaUUT7QlBOldl15Z5gWNNrnIkmnbq9KUtoJ3MGmLEx1Gpbwy7hj
ZgqqCNmcM49rP5gQmI7FksIF11Amk7QFaYXwYx3E+7xI3W5R4tBsAzzPynzWvlBB
KZWqG3M3siR5gNseLphmOftuDecgob1U4Sti9hqKQbapPcHI1SzBU4vIC4SBNCG4
6QMjr+Dkmh1mEB0nf1ycvolGd8WQegUe0iP1TP1ISGDhrXD3qb38kn/h8rKZi87m
ayKFtvQL1ry6DKSHMjothgxGzdV2gAHoUpnnICCGRJl92Bl9DyQxJbdFWr7n1rRf
yrSch6KlMB7j6xwiNzphxZrcZBUP4v3WMBpOW4eDGcZVyeiyQndyMXDESnAe4eRy
ITYQKP/xsAkiu5qy7gxSrP8yoLsmbH6cUHe64Rxg2p702iNEIGFvrCDnWur2cG3x
nsAGB6eqCTzVwkKaqsGoHSuS4jjhZbj5gWO4pjC+PKPkvjcr+dt/hKUQRGB654vX
G3DYtCUUQB/lG60/IPIM1IZvUPB0aSMVz6aptAvABS8ZppWuKgJvJVZj5xP3/VNM
C863EhphWI6hm6slRNurfyvbMAnwgfkE7yv9tNOZY7WsULea/u9KFQ+Y3OGt0wHV
sFkQ0s2YBwZykb8zFw6hfZ5WRnYnywqLp/49AOA74HSAdTVbZ/vrInFkwFHoRYlb
56pVRlUHLBoWbstJKFagf7nM93IEDbYI2BWuQNLIuozXIYj+SuLyZKN4SBjjvnvk
rBhfoNM1ydQhc2OANk8LUjI7OWNn2TvX1mcnSY5G0vN4oWGyjpiAsZFrEU291XMY
J3NAaymoV45uVoAkSkqiuuq3A50IV4ZGwVvEX+ZgOk6xzWiEyGKya1zcUana3bHL
/oSvzxorMWnof5NKJDPW9m1qfANKgFo0GbUFCDvAMqY9r/iRXtAbYG55F1980+2p
//2KZye1uWq2xVzP8XIsms/kDlwBWvPzy7hOQE6WNP+trpWEXf/6P3oE01TMBb8E
lbpigPDEg3VK0j2mHs4O14oByaQE3OqqGDhWOAJO2RBdBmNIVbaPUaYI06aJFnGD
W4RkE5TNranJbEycCwJDdn1N8aOmAaJmMcbta6Wl9kKQSDKJMPINQWleu21REAUx
E4bdqFeCGeyeFmGhQ9NN3CiCVpNTa+f+K4GHaAzI+dqxcTpQP3TfHukqknRjyabz
m2D6YFNZs4HFtDQAzA3SfQDxlejkaHJuDoIFDS6XQMbQ296Ka1U2v/1yvRQSDWZZ
XYCIhZXo7euZu1Y3DoH19fhteip02VdlxKItkAXZ8mD6ExstVIBBszKkXb+UOvGa
/LX+xrNDwC+nlZ8kRDmEJARImjaFLRyRlipF+8goxHBQVA3ToEbxaShZw3yyFvrk
RxCRKB2Dokm/YvfmLG7/WLH33gKDecBvbH89hmRbvuPnIuIQTi153UWBkwqB1RS4
8LHHz3m+RNmfhfnOzXqqqbneK5KCAEPg8YawDK/5XB1dej5lNKaYhA+jpWfv4yqx
NJJspgJ9P60/GnwR5oC6AvpxQdSluv0dXgH+ERyNjY1QB9D2MPvC8t3pu6dWEMdt
2EuQ1SAV6Zqh/A5kcXa/Hs0dwiZoyk/FdpNGVEpnxRM+H/jfbNcUFddjy7kzEhYu
tWUdDraGiXPFlG0oPKLohqcaFDo/4MidOrg+maQf5uRzBANT9qhNCjKVStwHMYD2
/BCxwKtKVQAFWDc1c0Y/fnRSVJ+EfsdvIGhGXbJg75S1/xeHeLW5QjtJKP3JJr5b
SaZZiPui1DFs5DkelQqX2KAqmImpVvVfWo7aDs0/69prE2GToWCWxYFiM+7K3XPe
NDNtU+TkNp4camfMR/sif6WDl/iYMf/PzdbvcM38z7kKuuIp0lW3UksXNd4gy9BG
cGAye/u9R9kQHqIIb2wNWxy66OANsKcZsG3OxytnQKzXHx1+Do6uigFJPHrK/Q0t
pVlpJhXvUAHhfZ2+b1qtKeQ/GVDhecwCBVZav8+hPBU1pw5BKmVMtHgxV4TTyKes
iRPnvMdLQ+sczjfKXFzaUTS8FZbcWVLWjmIkWFOcTFLu2aJJYr58bpa4ksGQ7Trl
aIASThMoxojijPJnsB3UDxZ+ai7VJjQaNWLHJeKZkKANo/VzAU0yvhObr6zXGVyy
+rXzpltZh6kVvAeX5TwlTtypqKRgvcjErPe91oqSBTgiTbwxnvBFcYngrkukIGDi
c+qdJTZa1TcnbhTatDEki1qSGlhpbgGOMZDrmTlIbxfD/TbR7+nRPD7fRf2xl1ao
PD+vL7ze8yDAEzeVMkuhYL2ABKLZin9XUB4C8WUKCQZD3f0opSU5wpshj8Ws8erk
tRTeLO45qVsp+6G/1thmC3dFNBf3ICxMJhXH+Qp5E/SHIM8+vl2HCfuRJmRBoyTg
b2pRtUZrG0AmQKZxee482Rj8YcK3Xw0sAvolSgVTrzGQXObNkOWYxubW8hlhmSPt
thPjusK3fTiImYiBD1uzwRt1KqXrt6j1hB5+MVp1mbQWmo3W7PmxyII4lNDpfNXm
AEK3w/WeKfE9fGfNVuAVu7u5YpKI2LeuBFw5eqY2q9rH7gMWvU5uCjq+MjaKNiTC
ZVjQKdjW+//T1OQKVI+8NF20glGaEOhYumpwU9QVVVsIB4xDn6p47DQjd5a5IAvx
cxGca2e1rffqKyZZVpLb5GSIclAz8nBa46osP9ibFq/1MNWhAFEgI/MKts7BXpR2
RjxLi3YlRCfUsnYRTmkNKkIjVsVlHW/P8p4xFg1V2VErcKTuILaAtPRdsAAQVGpz
P+rM/K1c8V+nPBouWtQzhD+LopuWAlTPWihBCUids/uZN4LRBTgzWYnmv4VYZPK7
4BpewB3P45R++b6+yx3eHAC+gwPCV0ci+pkOgTlmEMC1dvRmWcV+zG0/b/aSVStk
5nK5nYrdCDu+8JbF888C4ox42J0s/dKNRtEXiMbO01sOz8uVUyGvD8Tlbcw1WSQs
gSBIpmyDo9iR6YYW7AnsYR7LZ08SKjUaVosp/gKUxlVqtirMbdWDSAqMF2/3iEmp
fRbjZTTIeCGJSjha8ktzplCnYV8MSBnBiPEYCN/PHHOvSv4yV1aBxHxceNcBUmy1
aQuo79YzljS15bdxv9R+uBY4RJE1K7wHKXJ9F6YFdOmRZiHfLmRgob9iksX3kdd6
AzttwInYNubZgnsIUSuLFYmZh7/BwmLRfk49ZDnCob+mCf1fsGM1PnQ+CG5W3dEV
HiObpSS4T+AEtkspFK7Z8eeBx801qztYrsw/2dCxO7fiJs9HC3+466VnE2jduJ5A
P0MNHby2zDv+1Iv/+YrPV3GUKyun0STZxU5UyNlm1GOmii8krg81Dz17aaV3KiSF
vxtGGVFpFMJlEYTylKhI2L/z1XuGJWRqrHZ0X4KbG/gKmxsjKVKV3Pds6lh+kxbb
SJFyy++ATCINk0vEEXqij8w1PuJxb8+SNTQ8RwsQ3AIYftwzO+xcyycUWy6G24FR
Jt5KbLTxrakbwyrr0qKgcIRpqjxVhgoDga2a/0l+2wqNNpAMIrTIvvYZl6p3Yz4h
7Wx/jpq5I+KMfQ1yNVbFbGdrKUIfbcC9if5u38bc/gpCSmilfJabPaEzglXtkrNl
iG788C8ux+vW6VZOi0Evi/vZeorDQ5Z1yp3UsIh/iKFIsPfShIUVUIbbdD7q26pU
MzFn2emVvxeQqjBiKAYvuT7c5sdNwTyF2Cxv3zvZXXxzCC9kkHlufN3eX7eEbMku
f37gMMVA6rKzHZo0BKbF/lhKwr3sYivB/9UyARDgbI2Gb9P2cOWgxqh1hAP8Spxt
M3irZLvHKm18hTHJ/ASypB8YcVEiCoUuFsj7opVLe7n3G5Dh8SR+tNsil7Xt3HhZ
DLqR7zkW0aGSorpJ5XLultQvJStdG2iKviuXsu4NoHc0o9bGGddEKaZM1H43qmQq
IMoT6rQbPnbZe7TrX7kCa1C/xZ+vvp3gqTKVQEJ1vpAG1VPSs+2hldqk1JhDRqR/
2rF8NnWONBakw6Qz7SeolqOb1jhXYiqx9mGkeXS/adDkex7u6q17DvsQQ88d2+Y4
lwUp7nuweFVA0iEFtFLmypHEWfdJRF56K5izW+qDEMpYDjZOM56glhFYGQ21pJw/
z74EiSYfwjuX8dwdWcOKsTP/LX+2NTw5kPGaznGDVqMKcGa9P6cpCCj/bFDohLGW
YPJnfDErEMPTvOlX+eqDKlq3woSRjg7qoJfLs0HxBgsnkz/kXrdxUOhJyJ1cWqIH
/LVezowuQVW3YyxUb86xkxa69VNu0FuDpHHAosgyLQUkOMZ3mMHXzC8bl8FJNPaU
HzqVeCzZKgKgELporKmMdHfO0dviAaY914eTEcv1Vie8Tsj/kJ4EpUR6HWFXVrwZ
hvtB0BXjNuCKe14PWd9aGHqnnMkQ/1kC2bLvKPSgQXBsZtFlXNILxleBESvTiZdT
6nxIMQ2GHoq5eg3JE7Ds8w1ZOjBq0WFPDdQaUU/WpPKbn8FP54IIklEXS52UgfuD
UMR+0HCG98hJSBzppyws0Ix7mw84T2elaXdq0N36bHhK0bfSqrciJcKYrI5yQfxq
OZ1Rwt0RkUqqhc9NvUnqJvjnSTDGBU38TBvi5gq50pZJFn8ZU02394qnWFzqgFTL
b++FTBzVAn+l+5qN235O2Ny9/LD2S1YhistfKAchK8SRFahhGw47D7ZkaGRpz91I
rYMPDVcHENsDOdYtJApeOocptye+m7QzQYYfctfBynnA3AMiFgvNIqpQcoDf+drk
TcqatIY+7/3EqY4GquFhVKlIPmdY4A+xq0x1gQvjaNbWtdt4D+IHvOh33uReiwSn
VmMDZRA9XIV8V1nUYNO8nmgcgWLnY2DiACMUp4U3updiYVphWrOaiKQVq1Rv8BQT
os6Sd/dKZodfMYNsxJp835yLbHrwosHzuA+n/RmDnlPAO+OZt+sW+ZfAhzbtEpoX
Glq343NrYjvgMjXr68AZGkLqPoeTmyIt6rywMbyMFcfVPDrUUU6ZAacxRyKdAYFW
ylVMn0tUQHmxU855hbCf/nlKogtEoGn+GkdhVGL5sz1+AI7b9ZS5MAzlBffhqf4x
GuEidZ3x+qN147KMXJb/TzDN7mUtpy4V9WF0mZxlPN1ow6frocG3AYPEDe4NT+jR
Q5UHx/94B1G95500XqqYNuPwWXXTx8BTZxiRM8AeSrPzdsLTN4VzKUtV4gswMbtf
SmHe1cz9kl3HfGEsxuUuiwxYQXTV5hZ76Vm87b8luSznO2vNT0VJcgxmwWu2f3SW
Df0R0TwNODrSJbJanfLT4ZljQgCR7SlKJ6KBLgycUCfFGMPNHZMCYZcfRh9G0Tcn
yvN5kVZcCdUG1fxyefxF4grqr8HvGmiWF+GoUwr9/OypvPr1ssZXkxDC8zJsMvnH
ffzPrhEXkdTBjU/QqW7uS32ilwi+9d4GT8PGkqv8lOZUQJVnkg1wiYLy9KYUIToT
Rq5Z3Ifnu5XwiiHCfC37nbhTUL+ZX3/REN3wRQtw2Z4ABEQiYVeXhZtAVRz/iFJ1
JyOH7h5Nos1nPFM09f6rw7UvNKocTHaMJfw2pLA5Ajx+UAMOjf0cAjZk72aH0tF1
7SxMwohTJ5VFrQhcQJseGyrBUzeaJNLOfjgFOC5jwUkRlFBwGKNy2Sk3tPsw36xn
mKPzly35GBcjTJqrvZGq+xpSCrOiT+81Cp+/VDlis3wmkVuyabHKjuqOzwmwX18W
lWceo6cbxw0h7/l6VH53IwaMXGE6D//CUc0E4V9aeSg8P7bJwQKpzbn4FEIyOwBv
YNUFsNWfQer5+NsBHlfmG8u/PyPa9ny/nkQ/VBGpCnMHtR2f0J2RZke2rga+Ed/z
7O1mUSXiufT0X52E9UqeimEN+9iGNn7nmIboHrRcjAnGyngBmQKjj3do4+qQ4CK8
SWP50MxC4O04QKeBLc86lMwxw12nkGsmt8hpjebNAgpNFnisWSIpM1XaqD+A1gTW
sxEqbdVwGL8MT/ePbG/YOPB56oSjIZPHgAobW37J/yAfcRxJr2Lj5XboaaO0Y/VE
7I26Hsboy3LtKIXGJGW/ewFatRn0ovq2/MtHLI/90kvUKXIH+rE/zfht0al+s08C
MYAzT7MBb8ZQsyYHRwhDx696rXjIa1AKD8LFpZhiqAZkM7jyuGDYq4e8c2NWI3/V
6EAuZ1jhyEbTZgWdnSb0X7r1iVR8hPXAhWMlp1jPQ1zaY9n8tXYtRxL25yMXnu1C
KfqHO7JP0JdC3Ndv7Bx4G0wQ5iHkQOW+AhCqTdtGbwtLeM8w9ySn0M5upR+P/hpg
99qlHfCQPrL2qOfXFKUvUGeMXSXQTH6IqEJJ5NyMnBOPOXK/3/Nlv+14jhxM9o0M
YjY88+3EytqYSnBfXHy+wYocj39jixSt9VQdJdkncBtVmTy40FoLAuL18hD9UDkx
nZZRSd0NI+HJ1mgLP2cADl9EIGbWjPqh73CizeHQDbLiK9LoDDm7Tt2D87l+bmts
UE1sCQZhIMaVgPeEToTepq6HQGzCLbDpV/tQDEL5MEbNUJTHsm9Ab6x9bfTzzJaH
gkgLD9a2wIAl55U6Q58NhWhJya9eO3XxPz2M63l/MuU/1aIAiDFJsetIYr4K971r
u0MBuIvj6dyLtV9Pmjfy7AvyKg4tNSPvDteqjS8XgBYpe/Dd6PbeM+g0fK/U10sA
oXwler88Tj4u8Hi+izCASyM0hJ96VIEH6/xg7a9OcEwkpXwOTlg3rL5VYA6lB2Nj
mn8EgGtemOiIhKT1Z60zYTHA9e1x2Zlkwc+7ZovlLyFw6bXfqh5knSTtok0uCohQ
m439i1Z0RIxsOAiNebLbYFo+aPVGCMDukpHq1f3FYZZs/ItLESJMN+Wzw2PO7ZWc
rdyuULeT8KTBSVabZBpw2W9TAnqBVB5a3ZeThAI0lrrr5C7eW9L58uwYJesLB/Hg
Bq8HVxC/+eYKA5H841Ucq/91sVegiUnsZAIOtspWABwmC5wD7dGa0zBhQS15yzaS
BvPPc8P1f0AGxpuqJW0Eh4qQCirKyDIHX585rdhk0tE/S9hhEEW22DcsEPphlMtf
BbOfyV9oh68Vv6CIaNpzWntiN67zu685Kaik1sK8oX8oHvDpi9KdnrbvwjObJnCb
EZ6n3+WYM51BqjmkchBEw1ASqdJGEFebISkYIGjKP7wcIXmbfX5WGZ3+GK6Q5Ih7
LxBdnOocYMqgWgop+cjGTpF0W+dez1eXOiLjiNJTDPIySWODpFgb5qVToMUNo4Os
4WqSsPyZlNhB62yuFRMdV8tmYQWL1P+k/jrvEPEjMUitEef2Hfdyah0LgcOmZyKW
p4NDumwHfpUd/UFgUnWns3iTl8Jbn6hZzXRFQHTgaL/uVd7D4QMXQlB0FnPpuySL
rPZSbZo+6d1eFs9k1tuwCscTAgC+QlQEFcnDmE3Zty4OL0i6r/ujXz04YGHUbrIr
7aJf34a7lTzX9lgDpx2GklsFbeVK4RL2AU2UdjBWWiFFmzmOaoahBaL5HSjeegVk
HaMeeuIlsUiaAiZsRFzKqKerRbIcWanfL1hYPLgTziJwjRDcnrbzk5Smxtx8BMzg
NWqvYkxtbHYNIMJ9j2W++urbfyUuvfHFpSOAM/fQyP2TQ9IqaFpk57aaf13OeVCw
yEnYYn6zHs+Z+iE00Wv1ix2DAV23zDiGL44tC40C1huIihFBEV89ZaPwIxiGscWg
+psnyn+s06kRmPDr5rxAnvLlXMNSN5mNAt5PlVhLX2VnoU7ISTelKjTclGL7O/mO
18NLCPZYnT4tzgKS5/NdQsDza53vyIAd/E4wEluRMWitXI6o4gifBgR5+tl+EGEq
4Oef+q0d+70m/s5H7Z+733T/JBja48oiLx5yf4ecDwBpDzYxxNUMdt/Qe4KaRl/k
WAWoRIg72jTG16wH6VArLpz4i26uP+JJF326kJoKoQ9Fukcb64qbrtegi9wVpYNw
PLN6ykJqL6a0mpXEbR515muc7V0tIjE8j2K2CbQvMrBSK9w0Ty/THs8gnu9cCMHi
/Y/yvf0P1dRCCGP6ITdn5QaBpOhviAOXp6d7ouLmXRi+/aTpXf7CMQ/T/Dq5p6CB
2INaOvCQA06zlQfUI6FDE8oQXmw+qfPjL22A8PwjDRqjmY0FLNEjbAok3/5UERGq
AXK+bI2dXnwwHE3NUtJrpfekVIj1EBu9aTHpjksL43pKz67mWYAKyBi/zrEelOTh
jc8rQ0aMO+ecXY/4qY/WdJef69pfvzQ8nxZCj+zG+2hdq3ApKwAubxt7zKDmvKp+
g98p2VznknlWPA9OpyBlXp3RWLtmHHW5ptL6UaWKlu54DTjab/QdRLAYkBwdHOm2
9eSvqfzbrK7jn0+8gXe0uRjQwSDzDpfxMTWrPNoxWEv9ocPoaEeylEw3ihLSs8D9
bZZ1WsJqv2n8c7b5Mxoo+dYC6Gy8Ygg/qHHPxLOtpw+3DxnOaQXX5CIxRaB51u6d
/lTI8pVJdN0CaTV+sGBlvpcL3UQXSi/dy/p/Z8N12FCj1Bfo2TvKkZs05dlri7Qz
c/gLvpd9oPo95t3VRZA3pTakgPUkuYQXbYS7wz9YOjm1bRnwyAZmENWRTovx9zkC
fp11H1EFqDUs4m46x/xo+7ewUa6PWinE8p90p54ypECaHz5DlkSBeGTeM+r3LoRG
Bo/RgZ5JF58PO1rApo77G2vwymvFg30qR4fY3leJCs0DvX1NmU+5vvfwqSOzXp4c
lJhHIKluo9WogqmZesOhLxsga1qHpOO1ozXnhuz1odNdShMY8zmO7Y83LE4KcHuK
PSp46MrEwjWpR0jy6STtaz6kqR4t6QpI4epiPIyKwUQbsVLNTuDQEscUECE9sFQp
LuQSuydc2zuvzJ6xvvMITYRxM6EnrvrNRTssMoZOgjhKS0l4o4GHLBb95LYwAcM4
cFrWqVfpx3YpuiYU+bsR4UgHC9gTvQ+1M4CGO9XNc70nC8B5uEhm5q6sEgps/a40
xo8at4MK5U0dH5XyidcRdbyoLwRhmZYasf+nzk2LEZ3qLuAufmZJyLF5rL/n3pzC
PlPCiOa3R5hmy5kshr8RIzuk0UbXmSYwUNspVOz/cT5XNdWEY/ElCHb9jw8eddgW
3HAg66VBJ2qrcw/ZiOrkh5OrtftcoHGIO8jNKIapfl8AencWUgAM34LUvV2KVN0K
/7t/XK3FwjeUANdc5Mq0vGLUm9bbt7ZIWWij63gR3YMA+6SwDjfTeqREJY3TUDkP
Zq+iRAA9AUo84D6nQ2rjdo1N7SAxUvHK4Bi2kgAk5Yu+mHafznJhTr2VpTqEqpUi
BTl+4WyQ7QD4D5eEHp/2HZPpYHARXrmGrGBeyVGdR4Ri7UcVyc3lQa9UupglRyhL
TpAHA73f0PxL2/tF2cDcOUTHt+5lXrSf+GpLovjBLeCnXQilpOwRjPLL/sTYTaF3
QQQJY/JlFqz2QuC0bxSTdB4UFH6af2UuHOb+CCBQ4pHPFtjLRwo3N2xJ8azzuFc/
fLd3apHnRhGagiJGcap0fXkb9YkDDL0dcgSHo9HLOE1zZGS+uXybLHdSkVi3iuT8
oXjmops15f+UjlejIurG+ORlkFuwAtk260f6UzmOPnAfL56ThT9PLTvIxQUX98x4
FWFmaVMln15AMJonjrlHj33h7jd+Hk+UKMkUQw5qinA+MaGwzaXeeGqan/JtPh3F
Vssqp8PmR6nyC3qrjInlMXVOWoyydIQFetTSRKsIAi59nPksxAsFfh8wmm7YGBEb
7HRilirfS/+k8Vjjc6UZPYDCV4bu/n4a4qmhN34HiErzfkh/NxrfvC6dVCQaWjbH
NuxLnGXdvvwpTeylFL1zk/KdqcdvMC3Kr3NjNCM0gQKRPpYBzLzKUXYlB4h4ytrC
IFO6pT3+qTLqvFVpF46lLB9IZyH3YLpzhPdAuiosc+jW5XpgxE1Pk0edtL/c8NJT
NXby7T7ZJCKaeRcGsHP+VDtp0SBXwnN8Ueu2E3ddj0ki+7x9iP1b96x1c4JKqIDz
904Tykz3AZsvTdK+UYTN+SyyU2vywviIwX2GQsDU+mxKcc4QrLd3+JY7+8QyLn7e
400kNH9UEV+U3Q/Tvg4zwVB16dkOS3xG00pzQz5P63fUbPprG++31uth29lTbjRg
YzMwUBmK3OKe1C3pFjysBHbTTJ5xsmelVSnWrYKy5HeLDcKmZixntLIDUl4DI9Ss
8CC8SyAHEGUCgdMOQEhjefMZXQssYaeaxIOLdgjRzn1mgVraJPf5rxjtB1HP5cM9
yeqrit6obPIA7u0sgnlld/UhFCLXHVhXCgMT8DvzWrZ6aSqhMtgh8P3oGArDlKng
cR23ifTKSGppB94SO3yWChhz7UPz09e400Ao/TQi0LGsuqLU4PMgqB6BMLGe39D4
Ke/SXf4VYZ2xG0yjsS18A8CVTs1CCzuR9N26vNxcZOSguMeOLB2e6OBHYEXlHN7h
uMHsjDos+afviBhUn8DTfU63tzcehBVMqUUvNm9lmGzvOKM82vjGO00PpG6zzWZB
7byzquZz+corOx1PJINtMhNPWPHEpTzr5AdZmrzMVi/OJS7Fi+LNwgTSO9/V/js3
miPv2uduES+7mxQcgNC6chv1MmUKUnT+T58fIawCXCgIzeclc5F6aHu55pu3oGlW
U91thx7+RtvDnOQXa867HP7X6NoOwngAW5Xb8+RZw+ZIFFVZ7chryndaAna9/sSG
KeBHcbb0BmbzMok2lT9C117yH533qolDcIXZy1gFx7UgcghHfN+Xnu+fyCR1o/Ry
vUCU1S5OcbEJo6CCaojmMoLCjLOmSuIClPezLzyZxJJBx917OIaCyor0SlkHKhwC
B/fJjrZsSwVIfY1cftw8WZ/S5LZE/iNHwiT/LxiPT+spYHb5nb5eZrg7smzGPdr8
NdJ43gRNMqKkyCAHXy8c28do//u4oSeA32VGDoPavcOo/X/Ds8NBNYPBExK5THvj
lcZ774AOtS0jPICsGgJ8NzW91rOxRSNRynralFuhVdn5ipaChsHBrETjLJZ7jhNf
TEpVrk5mOMTj0mHEKrVRW8EwXqsfinmPBXJnH0N4Frx2jSu/hqiW2zF18luH+IhW
FGjWGzAgnKGsBpECsoiu1/CX6YmMacpiBBYKOJDFbk45M5qQM6MexFgsfH878mdL
AtHwycBr8tWUOpnOAgkypxHsZRknOyNsoTGND3D1fhUMKzEaJ3Rk1VsxUOtGHK/z
7oz/o7wfO4SULk0jzAQyZTNcrIJreE9cP0BvgTyMN2Abw4ZHxC5fWbV75+mxT1R1
+TRTn7S3RYE432cwuHYgTAPVKWep2Ax6DfQOI4iFIsOEFVIXmEyeEWx9Jl9a+a4c
9rxj/A0jj+HFmwjq57lXFlMQ01H60XE92B6QiR1xwlp2Ed+IYGilfzAArUGBYvih
iLO8QqU5BW8N6Kw5UNk/ka8JLIoDmkc8XPOxJ6cR2KofBSYUQAoWCI81aN/G26jP
i7wazKuIDiJAgN+WsvVx3f34/73nPZVsN1HYNwDUEvwlgj1xZdJueCjcIVijC1/W
W+bnqg8CzQ+Q3lLrIeLj5/E7Ie9/QIKqDozXNYjX0trrX9VwgyRhmyJOBRMONfu2
bD24za8/MKx2k6l+CL3oj7yX8r/Wy+rREvBAzq5cUdPTdYBAcclVDBEjGa1rLqxf
SC6SBnYBDJOzkp+2JdV1Taj1UmeYD/5e/4nN1+vP14udBaaTYqHgZNKVk0UoY2IO
Fz78H7fASugeFBlQndRErAyfpUwILPmNsNqou1D7hLKnEECd2IG3+Z8+VDOsE21n
vkx/bYXTg4EZ2WJjqWJjpV27O/JisFnAd7W7j+Nq8lFnb4jfR3sUOka08b0WFGDF
wYgtpzvsbKHVZHippReoZo5HquAwYd9QUMb2DTBwnt4KRTxZ3nvaT7PaCzYLcs4G
ObUcLVKw6moP37eM3Di0qQYTk8Ar4IBiNbv6FH0L964lZcFcW1RR15h675VqmXRd
WVgrk0EWJ7mqTT3Ax2xyYUjnbsStKtNBVuSXdbkdmyXM8VoCHmn5DuU49CUboN2W
m8wxiFnHAdK6AFCKpgH2wrXPXormGvJx+w9OpbfKfKl+xUom1KiItZj8dpVljXNf
qbOwTbZusSpwbgoN1eJmcAPJbpYzTvJqLAU+mBYj6txQOvVIdUVCIbBKIgUSvFGR
W8HhRjBg1910EYrewVPK8thZEFT53s6ISwdZkWNYICRk+/EITw6/MnhkzyDbLxHd
tjwexgwza38sR+eImOqqk3E8lBHy/FYd2PNlTbrP2H2PiGb9mpe4PHZ2tTG76I77
JD+4oE6qiqmHYLW7PSZWnoZwHrowkCCIE5jrkoIys18WavBOoJGmWFWAigmvthn+
2QX6oya64tnO4fu+70fWSzEOavlkGAnJke2ZdOMxMcIl4kMa+oji6uPIQojS7BId
PLSYdiMYZcSod+JdlJwuD4hQJStsf0X1nxoOhjKmGNYT5gntaqDBk0YgRlvTBOYQ
Nfyc1JCDUfDwZgMcDe6uQXJy1Qi/1br8rMO6MXf4Ptly+zUvN7rSt9YkotG42Wap
+P0+QrYopHSyq+BrMIYb+JHCfoRq3VQRMPKuL+Zpb2ZQjEJQaT/+qGuH07M5oNNs
VGMx9NX/nTCM2BBAsK4wAhviAwzbdRwToEN6FhDAUVjpqPrYRqewz30FLC4ldcD9
ijpwioW07ZLarpmuRTFJJ5tR8lQ8eO0ewtJ9kxffBA+4AD30kvaJDyo4ADan14d2
F/5Mt3VtcoOhUa4PVNi9XwGbDdijFAbb0vey4CYW1am2iarWtuOkSmuFVhcG/yi2
QiZxGtwd7/0W5MLjMy+yCARWkHlMTPGYfbYtezh7KHKUobNCe6TRUsN0G/mFFw+o
8RPTKZJKIjbWorP8F0S0B227y4XMAffq2uOvJK4uYCjBHucyKJXlt5+KvZov3m2M
qAdvBHvHvShhtXAueGGIoEdvoHrFUQ4lgv1vUueM4b+TpCagUchJFcn3ldJbmmQC
OU2Wy46GyyBrbPyGtNfHQS230nuNRfhTz02eTJiwsCEyj5MBPLp1vngYmvLKF0YZ
6j/ooAEbb3TXgjT6xpZsCVNGK7fEXuHuRRxn7LAtr7gPauBrKbGaWx8aDByi1RAO
RJbUKzzWlHHOxcXFK0uJNTjMJM5unlvI1meDrPz+eCITUKMzlnJOPEfstUvFUzEr
gZc7m4Q0IA92IC2Rs7NEs0NyCjf0sCAc0tsLfebPhLl7NDnaIy0kAnmBZl1FGsfw
I1XVZHbht5ihuD0tOngR/Cj2uJ9PwEcfKLFgSLy0I4fi8YcLMicZFkzKzE+RCVJ8
Ax5P4PPPFkKU0r2yOtkjUoVxQ0iLcT4oAfhNaOgmhgPZIwCWBp6dJFWVB6GCIxbt
z5hvavRBGwtQZ5o2TtsuxxvYMvdxOx+zDRf6VOLHcvQDZgw8D2veTlifyB01nhlZ
WQFjbi2uR1BEDsl7R5AVkJpwjcmQUwuj2qj2T/OuGXtcUi4iYiLeNOc8tqOhQYq9
fw9qBjmxA7uyDlydS23FYjQh8EA8rLReUFDmJ7hJtNbKMi8JHKOSt0ghF8U0EZKK
U1x04XK3gpaFUXaNU7WyekFa2Y56Ioni6Rw5UFkt95Is5efvW3BwmLagl/EQgIXC
5x0ZMaxvUR/s9z4udmsmXlqtjBXQegT3zxvPgcAZzpmjICOXXhgr43EnDdhX+LxF
Hm1nEZasFM5zq1CPTTh75liXwoD6QXKDK9FkYqLyVQOM6rifJVjhKgKJlc0D5apf
0Hao3cg4UQWVo0l1hB3Be+A3hhVwY1nY+wVgxWX7a10bpu+n+pYMOkvuQsPgQE4S
h6fBWX5yDvZsBiCaAoOjrYZmEl4cIHl0DJ3fbEYoQymzvRXxTcBSpDZ4eNmojHUT
TT0/oNT3C05AkO/o5BOGMgTNzbVNCwh6HOhOwjYVyFE37FqlqhNv62D496v+0peM
AW1lFwQRXTJ6ijeLOlUV3c6tytTi+UhSwFxxRoE5y6addLfKqCNBWSlNmsBnEGsF
9VnYgwVzd+R6DIf0PpOuInS4Kvq1v2l+GdiIjkr9J+vDZ4jrPepCWDKE4+asRy2d
gJ0y4InTfKOktF5d40XgUKJQaZWCkh6/8KqdgfEL8sQI90XSTH49lqxrknlp+2DT
JXopYFvX7kQUrLMae1BnMbSNU7MpkHMfKZiQsbotzLlq3xQYU6tAGc4ZQubR2EQc
V+lpJvSQ/8r+aEmoou/BFVm14jYwS7pFMgDi4vF9DcwOFCGaUYALoI/jtpkNHwcI
OO2WvDabNtPjh77AwfkFDpSij+7c72DCsknpS4dZzsETOpTiH2KZFby5rCcg+fM8
LBHW3NH07c9dIifXTiN3aknERl4T/0HTWg+LGPK2OrGct+A7VarQ2K8nDHOto9Lm
mlW+cRWRzEdN/P0M+FQKJ7rsF6jQVrguMKxENdjtVymZ4lLNcWR4z1SKUkv7G3tv
vle7tvAfjKaI5EYAgG68O/hxKN5gNNjsDawdctSEzqHeK2Wjge6WpSDOut/ngoat
xE6sgAFzluQDu+kshkaCblmBIJVXRoWt3g1VsffLm0UdFqDT8o35eWmgXacOOPWz
07Guz3eN/I7NqHXQQ/Kpf0xG2mHZlehO+rcGqSUQUICHkuRTxIZAI8aYTLrZ+YJv
QUmNSHQWET3q1OaWNAX9mzeZGYGuzd1mYJynZ21/UB0y5Qj1ZI3KsMudKNOlDWD3
TjawhD56rTG0VulPXk9SfQSppiJtORA4FVnCNwjffYdEbM3TD1Pwf1TTYgiikdun
huV5aq0zGQqviCuXAgLqyMoSkcJd+lzzqUKRrLFBalJE6o+ysOZRqa6s4tPhtSSW
Dkwcfu/jwDT13HRYdVWIEVBIQzCSbIRuEm4+IEbZ+werVliNZQJD060I0q4sMoGT
tSQquLPdF2UgRfnJvqK5Zti7aicGd69U8XDuOb1veCUi8AxN9Yc1hly2YkW4uGwO
rKU/MeSppTmpgLRCcU4Og7LQDUHlXot3XlshlT4VPJkx7ML+OUx5G1yGWsEp8JyK
YN/C11mg9MVjnJjk4YwuUsQFntDr/ZLFBoJys+m6dv31nGtSp0lbXljPpsjMuatj
JhyEvgGcwlW4OT1K9al0jFxegquuH3nUy7bBk0W4Yecgmxe23qzggzBHkfoHsTdS
UBKFxr/rjZ1KDpKzXNwwNU/v2dYFKkee1MeOC0pBaH+jFgVoLurWeUBkympcRusV
QggWmfQSx1naZr4UKoUL/7TTL5sZYrSDKnwmZmMvSrwnwEZRk39elEyFnQIwai5S
PKYww0V9j7qdCZ/vCUMAxkc8c5p0yjcrx/O6Xeo4UoEBm/ieFkWIckrhLVJgV6iP
3tjzs5+4ORBZQiZa2gbzBlAC9ZxqYFMC0YDbaQ4nESSm+o1DqXpVOr5h20j1AwOq
WhE4Ze0uI3kgzwsOHtoaMAPkUGgfR00LGairmlomxOSOTVl10Yw6a0RLObUfNwCO
EaJyNr/kpnacXGwUpDnJFo5eWdFCTSHPyiYxLQQcYTIaAyoUl5evVT1nxepKk1V9
Uy6it2qk4ogYrgkEKxs6Zr1VeEEJcpKsMRdgdYo/pceHVKQX4EcvO3onSoFh8ymo
dMk4enik1q7xB5cxbaIrrLRkGOMqTVszPozIvetKqKiAj9ZIlfLRoRebYZPCzLqS
00ZccV1GbYUc/rIpjjF90n80VNtFCIqFsvX+n9MsNzVFhDMbq4xGFMP85vIYQLXL
pfTfCPSUUshfFSt2oOwLKOQO+o6f+y9FnDKb+EFdQW6lh10MpaSs1hIiX6AbCzTx
VpJ/PwzzV2UUIs0mKT5M0652wkTfuWIUuHC091lpPeCfphG6v4Rf7xu7kYfjEAtV
m9u4LdJn2TZGKMsUgYhD3MMkOwIRFU1fmARND54bULlIDwRXtTPAXu5VjqIVful6
i6AOW76FWU3YlAUfcOS7UQam4SquC7gJ07yi2ybGU5C+UNFe7crzdAMAGrkrl1U0
hkx7kdJnZVqt07K8eev1LYZ+F2/EbfVVr5ssOpQZ9aSdfdh3OtkZmkT4IPl2CfWM
maApjsAo2KmVNDXQ+FzQhPqGFuwUBStbhFQLB3OGgE+Wu3s+pjKL7350ea3YWBgx
8zMzn5o422rA1sLCXlOeF/dFW5IuI44eEttby8WxL+4/xvurZcsU8X6Up2l7St1c
0g0PS/n79MybhatWzL7JBny6+9U1edl8Cm5hkL+iKt9wP7qo8DkEd+wPMusnIRTX
tJWNRauWwwDGxtHZOQpLdQoH+hPPefxgERu9uvGqyRgl3lVWR1vlwLjqvH2WBedA
IYzUJM6UNk+1y1ZBGXH36XMMAn7B+D6fLIBRXgEMJ4/7Q3NEnToYOMm8RRaRu4f9
I8i+UNCD+Gug8bwOb5O43OlN+V8IWRdQfayJgLZwU2wres3TGBYLlcdvy8eq9Q/C
DAVFce6eZcY5j+WTOqC2Y6/xKlcOu7EYXiNmDsG1tACspaOwprYfGpnwgkdZrAKp
hBW8ecTJrtDJJ+DHvXWho6+WqXj1WreS61oZXm4xLM8z46dIh/DDkxu1hVnoahVg
xkO9sJlQa/F1z+/D/TXTIHJYYyYLJODrWpEZXStUWj3B/FWuuOW4kRoIrqoNrJH1
Zan9seThCya7xxwYbnaQGOyHx8fAybhOgei2mzR4r/YH+9SQB3E6frHIfhwaiSCQ
XjXQLXUSdwOR6wspykWRTIfeLBTXgexjyESjNUgcuajjYsFtXv1ymtI5bEf0o5GB
JMdYH2KQkpxIJYyz864uug8jsPV2DGv4Oz16Hwldh0rn9bpHoQ2VZVl/jwstKfS2
JbY6AM34AAWpqtjhVHPy4pJcuCd9a5DAhN/dWeX+QYNXpxdrnun5ONj8QrHbyFLe
XcjsmYBVp5NLWMNB2rbkj+S6v1miSjyVsCZXO21vy8jkmjo7xUvfJb0f5Zlf5RwF
QiiReYYUpzmyTHGS9djuwVzeXHik6XGkioGpc3/s2Z7eE3a4nQrMZjCBXKzNCofs
dEGrNY1J00YqN1hMWyqkdPN2kYyPx/qLuMy/fQuiwkJDQ/dytgdE8XcRnqfzdfP1
oNqhzqVI/7rPFwkZ2vmtJGkuulAvABz6PjWAFlMgv2hWR2LFpOBDgvLue2KT7T6U
dWnzZdIZu9VRCORAcl1VVHwHm008pAcQDBmYqmWH2sdAFrRwhplzsUkuMf/zSuKM
Ebab7i5ey8XhZBr70y4prMNbytqlPT6Emk/8SivPOrxLs3NeCE2fqdTUddQMMkky
by9W5oGcVfbqBf9MEk1cMKuftx34cUUxyByBssMKhUarI+7suEw/WT8y8KS4Jaqk
mrn/RDSzkOs9X7jqnZ/vWfuMfCYY8S+ei/NL9E58Al/3Askvq6D4u5NsRdM/w0qp
lPv+Cakq0qtBQTnrKH4vCTprvZFF+5I2/LqI4xuMxNewTkoTRDpZicv0fLMtgXKv
lxcXuUxFEUQhnPY9kL61cn5fznq04Kq90wA9mY5xw1Cg56Mn/dwVR/9/i+gt9Tn2
9kdPDNc/0rtv26WwsZAwIWE9n4WsjWLrBRBtHL/hKt0t4lBlj9X+ybJ3gIKadZXo
Mz4Ge0/3qb92LSsg/DC29TrwOm/opwAP0ztQ+WjVAZ+WeKikMZfYdHclNkyq3SUL
4QmUGwmCZvqTUEPfw0N7QTORV+GKAHpDzoSE6bYy4gdrjhqzDbZLAitGCuMG8/Xk
AJHE175UfLwpMS1bJQ3b3w/loCbiK/sN7QApO6zo0gvzG1VX7sEo96FPJcJoQ5RG
jCLdCVCGnOeyUeSW5MIuECaIX8Dq7nhKmvbyhx7zI763t5C46PBr1PxB/NmNnhgX
AF3wf86zJnOjElfAxPlvXw+HOvYuHBSh8JeTo7nsLO/MEYeLn+1p5T4ODtB/rFuL
8P4WRDVrFTd9vMIJIcHLAE42hjXt+lSAvD0WfxUMJ0Wm7pIbrKxe4qOSkbRu+SZa
hpJgztNRsdo+hKiu3zM/LWivBKlvzaGOW7sF+rxsvFGKqZPYdrDxxiZgk+copO9V
pDLQ6USvU8+yfE8ykPrfxoGSxBKeKX9Gu35LdRufDjnDzgxw6ICpUwUbXhDKFony
4/TRMlbfjbXnel2hZ4hZDoF2ecxIqXyIyYHMVROSor1RP3PvEsp4p0u/msVn6Anv
tPh5UJ0yTgelB/MxFWkL7wzO/YZyTPn8YcN/QSybBtvrdIys5R4WqUbb6wCUN/C7
qAzmcMj0JRcfSeodH3PguAj62+84PRvXhkwsfjW0/6dh7if6eVerZqvctR9PUo9U
3s/oj2YY/mfIXZGDyG2OEGLkNtmVJn4flEmlQQGj9h2KUkTgiNoua4O+Akc2MBKx
XMQwz2FeJz1uFt50FohowtSYlk4YOnaxo7bSoWm+gef61Pn6WB/tHabHWt7ERKN7
zTDJLJmKIvz43uEWjSZP25R6EtsLON8wvWcqDeSDEYxbTAdn/c16zjtXEzXLI4z6
R8mfVGq6m1/OBtoyxQoKferCnM7fbChNVHBaqgW1x2gTTgS54viT2KPk+Jqian9U
Aa5w5+pyw2U4T/mkKU/S5c0oCoK2TdHyKmkyBlCbwOyU7FAvXrMRwKgWL6+3k7Mq
5mdjISI2a2WwvclROcu/rxmjzs9P+8w77gRd5465KLZ7oIqUf6mHHYuJccE6nifr
sjNn6iB9sPDNf0t1EUMCMA==
`protect end_protected
