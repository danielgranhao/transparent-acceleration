-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
2uZ7XPcO3XCBVyk2lAJSByGFhE5zUDcM0iYsTWG+8grOpmPy9ofznTqmkcu/97qX
m98HpgilQAvPdS+ZZKsConuTZXzouQWzvIHzMTdv7jPyfJ2p4DKfsJ55U6LjStAM
AWQtngXeHDMYSY/i/2/kcwtvD1UJhm7UUra7WJyWjNfELbPcvk5/tw==
--pragma protect end_key_block
--pragma protect digest_block
ibJSbFdOPP8WY20do6LHEQf144g=
--pragma protect end_digest_block
--pragma protect data_block
Df+i1vTo6Lr6aECv0DuU0olcF4mfDc8rixAXh+JVU9viYf5NsIwoSBcRfXsRZUIN
XCKRKwurLUHz7qIbPsj5UxG67GmcvariUbeJffQ5wM2EoDcgDEHjrutYvx5YOV5A
Tg1krSSPVVAglagM23HzieBllRaaJ2Y6Gq93qSva2uHiZdhtkOKG9i91aGveSs/c
sukTciuDdWd4i+9Nse3z2m4s8eCl3MyVI1N5t0H5bxhmiQutINtAn5RsBo3KH4I6
Y4uXMXk1jFnG23XgxOjQOpWu0x8VzitTYR2o6t2Ud3wWw3sc1DF9Od0gSE49Ue5Q
UETE/fUOEBgWNd0mAQbJKfqIcrzfBqbTqQWRtRpOMVtb85j4WpfUxhfymk0fuMho
s7zHgWB2IMFscuYQor1yVmrAmz67/xL9g18i51kk3qBePIncqkpdZKpUHZTlXFoX
BEc3liCHd3qbXK9E3x2qxkagehgdQkDj3BSoDBa4Jfy3NfL/jX4lUn6+M7j+rU4m
pdbwDkJycTszJ5yJvJ5QeUccEmXXYefLxxSLRvTTxSRSZvFDLoq97QikVm4ULHLb
XfMdLxKhJHrqwbptdTakn9VQpAQEuCIYVv30ZHAkzsDXadoa3SA4ZkM1VHk40H5W
alvuMIf2nz3TafRc+u+lRtlaS6qjUOGKG64izG6RR2Nuw1i3fdQPaCgu/tT92gQ6
EewtjHefr219VFfNFyWvU7lTWpJKwyesTfh9hVS6ZJcKMANdLS7LZY6FKnCDImxJ
aSBimLJjhMegvCuzpsV/SoLgIj0nASQbvsxhftDjx/Lp+Iwm8S9SJz2MbWbo6VV5
7kFex2HT9bkW4D9UAwtBpmI6UEfnQruawmGrJIL4azkvx72vyCGHfZeUDZlnGiSB
t6WhF6uhtx2QSeuvCpINxN0TAzZ8I1M1bmzXt6FeJ3dw6pna0EjdJnzp5fgdDJug
N0unxv0l+W/ZbZlXwmu8K7XcQRmeZHLsJ+ARmeDviYCvrgb1BQrz2EgnNgr1ctCl
HgMwqypT9P0sPLViarAeoANqry44E0Pz3alEKekNNaGzMtG6Gkm4Ltg8O4QJkB6S
fIyIW0JBKkCbd/Iw3Tfk4MM13ppEem6i1u7LgS8J0uF4V0HByiM/WgayPVijoJQO
q5gi24X2aHi92Th4ThbroCBdlV1A+kgvaBAstmyQ2hS1Y1lUtPlUsa/ALoB4tVIZ
qnNpzMbnSnaZFVfZgOTrO7d6+3CfaCR5FJYqG82hkdSzipLY/48wOTa1zRyvUJrP
UOOQRN2+Mk79jwsecEi24dgeEOsgWmYm06vN8DTBNAwqrSd+K8Kr+5bpNbPB0cp6
IiBFG4nMkJ3QYwbMjnArBj6DaO5w8mSsIl8EvlwMz3EoGvo4A0Q8EFE8tJELmw5L
lo7kGjTj0whwjsBq7qjPQuHxTv2N8F/iYbCU0nQ7+AP0q5Rg6IgdtpAMAKjtcACj
OfPHv7ebKBLtE0eonQoV8PSqw9xLqOY1Z+Xi831+gp2TQnLevRGFYX6yAk75IWUh
kGA0t6NnHkq+mU7ESHY6csqpqYKP8M/qlVsALIMnmOKjR23IusP0dv3ZgH/JsNED
v+lgnHgEnGix5dZGYYnPk9Hm1TiiZYNQvPVL6aDunfammCQwxB+m//NYSKp6r2i2
Np0Mee/VPfDYEi4QiY8INTigSDFv0NUF3KIBEIE2IGZpe3Oxmgkn4SzrsSLZ99St
+pJjEyC/r3QzpQqg94SNL1LTHqoQo78bBtKA9huvx0N2atmf5RyMDzjhh0eUIRW9
J8D//U+lMUB24QwdsWCTySm4RXFDJpwi/2Y+cSaiauDKmcRWkNPe5D4WMK4s/avO
3kJIoLQZtvR22eO0HmffMAiwfg0pXro22VspTt1jdML5FyJGQ/APC68RsGV+frUC
4Y80lEtAvVrwYbqNahFH+uK6YEzIcryJTVRT/zaBBNTmEDXfn+2P27hrm5K9NJJG
7knvURQB512Qw0Y0vxLPqV0EQ0qydY7Z1Wf1IGFgqfK/xrNi/pKzI4DIUKzdtjpr
UHg3pQds3TjZni/fcGaV2th2nysHMq0wftnKpIWDvZB+LQGnPiG5GXvt/JHRl8rU
oRsZFTVnltrLbjlCBLx/kwphIunXU5E0zaikoetUCzZwUypo2MRbFtrhIFIfycsE
xGbkOb/rnN01hwD6KlZaujcrpjusUpDfaDE5yj9X0vbONjR3oY3y8i58EqrU1KXm
FtP8Gh50TKOym71wnDLO051+YsJMmDktgCv6TQjZFlKjLg+t43pBkvXHk9IenuTG
kGE0VDvxq4y27Xc+ifkJ49VtDE7xqvnm2PRRWWDDnVi8iE9mGE/Mkcc1Tw1ybODC
WwmtIIhMumP6oXRjaARm9W/4QAjRj0Sjz4H9UUYam/5+Nq0SKFMoyBWodwOi1HgC
mIyu/6xGo3RU4xzf5NRpFyXr94CE0bYeP9tVosBbWZg8oyvMjMN9qUly3TaCZGfE
8aoi9/C+qP7mAzddnAjGfhYcYuGauyf0I1hrgDL5vzA9lf+UBdBeQYm7CLFLCU0v
UWQOEeQmmUHDw7NmRikL7y+WjRe30VefeSWvE7L/9qiiNBY54YA4F3JFXkGFmRJH
DtyghfVt6BfyYWd3W8AlJNaMAzi0CNIALffdQDjOC9mb+DvjrlTBXlcq1+p9vLN3
s9iMHyhXyvkVEXO10Mwv+UKsknyk/bv8JtCK6fyNZ0P22vGuNqr5l6cZ2/6lc8nJ
g9IuGfMSWcDRETVTqnQVG+Ns4zL+0mySjf7CMog/B1m95hWLg1omuQuwFtDedNzN
g/OVBqE01t07sIA+1ZAL4ebkbcDysi6ifeGAjsdz3uVOxp3FdOJ9PA2llf5g0LGv
Ssl9C4oLAdlsB0N7xL0AxCzjmr75Iy8QJCJ/pURZWn28OiU2gJGSGlBtpFcfg3Jb
QOrWt5eKxQzHN6leGk7IriIEwGN0rdtNG9UMRw4KLsiaUS73LI2nbexiCDD5sKzT
kXP1cJSKdYIH+QQZfS/YYMFMJqLtuFZRY1coJmJiGaSgBbGK/09qGyCsFK15ZxC7
eWDEfsmwvkP3+YEYBS0lnCkzL1X4qAC9z1NvS4ssBNJXVZYvrl3Ef9+51VZwJi5k
nGhb+8QsGTY5Po2/OI9CuP2APeJoxW01PE9JoKoBMPKt8L31Z7gH33QVrZteR+3c
rgJR/TQfFkT/xkk9t48rOMOGuBxDXfX4B0OZ4oWBXqvRP8xfAbw8vDctqmsHQF57
+Tln4JEpxsV4PuitV6Y7GoPx/aXDXTq+EzyLu8VU2tBI/ENa+LKdDsclRC/3FT4H
UWHz4NltDOK52Aw835M7N6SDUKtW2ShDbxh3M2T3MBI1sei1DC7FJmquAoAjvPcH
W9eguI/0WeBEZ7MS0L/WmKj46yjGLCh33OUrV0fmzwmqbOgca1LRAI5hXgtsGn3+
V+dykf7pICQcMCl6pEvNYkqnZZyOu/iH+BvPJM2qtQLrJZAuqjsgeUcAWkgF4eX/
puAbRnjs2K4vyjAw6GTHsqapzbtcJmB4CkuELem2j29inJJZaYX5CrBG5vRqe9vC
pFOuFGgLKXjv7+ZZaFwFDXdpTBr4xkTeVRfepq6TPb1FToxFNbW4w/OtDKHR1C8x
Mu2LgEvhivurksz10ZSTOkDVaoI+B8Alc0MzPSXNNGvwCppl0Vi7lOrCz5wpcvgA
wEQVvPRu+N8beSCQptOQS4m5J8up+fGCCTUqWSPPrj0+33f4/W38Cfe+VQ2b5zVB
UMJ0euu3qy85iFxca877iqkaca6UXmJZmO8Ln5imoCjEp1SQgTMnk6MvpiKQEkMa
DI0I+Vdo7md4lXZRPYm13VxY8XpuMYQtHnCSAjm646EDZgekjuJWtsSA6RbuxiOW
+oWgl7yirv/KZBbUuyZL9zFwxCpGckY5+4CAvodfojBhvj3WNseEG1CS2IQovfnk
zfaENf9RWvBrksz5lBGPftqzmabKw9RtGzQvB3K6SLPhJoMhUoXai5D4j4KwHveT
+hPpgJ8tcXRDzSQBMl8RW4wA7GR/9hvmiPU1DYpmv3Z3zN+pTFkP35IuEJNj9h4Y
nmul7gdYEwLp8is9R3Dbe4jTWlC4qfDXgbI8Z3KcG6h+NRxkmqmWlaGY/xFPkeyS
dFvVEKv67JjnifadBYioZVvIYUA6ExFio1JyBDLitrtwiPWdB0nOjrb05apBmjFS
/biveRw54H+a0eQQy0u4OJlUKKLjuilQLAMmViUPatznCnZ7olGwiEwc7Ob4I8Yw
2QRIxU0/aIwOM22gck6k30p3EHlsfUIel/Tb56JXuRYyjaXRp2499Wx3f8WbVfyt
NKXlTM6rE0hVgT/o56YZ2IWWqR8XvkwAnkVNn/N+tL42NkXjfwCJaqRcUvuBEUpX
3AzufY3uUgqJuIKq7oQ9jlDyhQMBgVlOpU0OrkNyEvL2LFa0zna3DEuv3jLF3hgh
sRrj5DMU/M1wuthcwdRtrvEfqUwmCGblIE3CAV6TPEfMvfoLFtmY3xrK2IYEeTUx
Q7cVoyGR9I1+8zAeRR3uTyFMBRl7QhOScjDZ3v1/3Z6hi+KFPxGkvazsW0Ra1MuI
wpC/lcRM3iYHPE8pyrwJBoBS8cg9mw8Q6AlXshO0srYsDo/k0vI5UBWbdUVjTbxz
VRas+ErVz1VFmRCTJ6PWO9DU2QgqoggjHo4kZMJ42ytuno4JX7mQrxkiHf8rKs+L
6YjQP0WlOK5dwBuMhJl1OR/LSx9FNwO7+jmN64Bgojf86BLt100GwrAx+t9P6roS
3IzrSlqAwtxOU+90VC1oofs2/34OIB/5DDI5py6kHmXdbpcjEcC5nhAg8AG8xKyU
tmdSV88hWEkT7cSq52wE+Ob/Ob8on2I/jDsJ3ukFuwiFzFLJeV6pYiIUiGO/dOKM
/zVe8ghaCT2R83DA6oIMxdbUxIfDfXfryuvO8AQaIzGtbBrMkxa7OV9wCvLcS73c
5B5hrrX1t+Uks9bBtTHPKT0KP3ZToKm1AWDAlHxXqutBbyJ2idPL1I0ocwzN4mpa
JO4NR8deRBUGbKwxy9gssLiQmVGMmyqq21rBF5tnex0XWRzENm4Rw7/A62QzKDEl
50uH98VYvOOQ9fwOXMEt84saTer14m7kriyXQUc2KIBOgg4pXjUQfCqganVpV9LL
3gttxZM73BRfE1R0pkhKYFKL2JWoOpAW0ckHLJnf4XJ/96WJ6OI7/ZhaOqxQaNLh
pT8Z7HPolMObsTs18ijltPwVY8Ybkr3wRr999ls1Wh3u5FWZSv3Do6tOPN/JSCd5
ig8sVsPOt5rXrtsmn0eR1Os9uBD+hu1nh4IqjwWFblHt/csuoY2BSDaJIs85J6ZH
SHYuODKs1qwQtr84Kw5J4V07b4B1XWpVn81DBd49loHmxfJmtJa2agA5kKNW1ujN
aMH+UMhm6WA56PZ2tT43hPP0+fiLNAuHjyTfpjCl3EGAlq1Uz4rXuxNcVlVR3lpd
sW9ob7huLtgoBfEV8pgFwUO7vcNEJuxBIsQdHzmj5KZuazcaWoN6q7jfoef8XAu3
RvacchXkrmLvC3fu2TeFVx47p1DKbJFYicE+qruyXHd7WxZ15YWGsfYjPRTOmqYc
Fy7UGLUPs8RPggaskAkRiJWZ3N+rwoNd9dmXFeRf+LRgcwN50U4GOwa+6Zxcljxy
p1fwyz1MdUw31ltk2J9cT7M2OBRbxWSmDNPS41APhz4isvgTt4nDGshEEus85MVH
jFEk+/NRhmeCupwUsx7/66IfZMbxLory0KVvlIZYZ+/BGfiSMhb/X4bX0LTG7q6j
GhbwTM4KpgFSfFw20bgDRKIbxPQovhPN9lfyRZXIRT3KbUXVVMlO1F/112CMsVvE
f5ddFoD8E1xNcfaoC1CeGEcAfA4kHGj3e10E5lYHyn+d9Gf9pAFbckZfbiQPgysf
7adWVMQlvJIIE8X5czdYpzVP9bqFNQ6+U8U+Zk2zsq0duFnygmPmNF3wRzwaQb5B
bMEVn8cmqVygecufNXJ5bwaUgpi6jgqvduQo3aUlA4N0DZzk0/bTLb29gWbIiyrh
Isoo1/rWqODwla64FE4FCgthrq8KA9P6a259OxdKycD7K7bTBbXZ6/ApKMZT2QW/
HGuPBKUfSDsfUymLmitM4cuTgILYmdMmGvnGz5WWFWr+PHecvlrY7jytt7AMwOi7
jp3sQFF+NyyFYmOhlFVtPVP+bXpu7MF/+X53Lg7/uLrf/CkKRCjvTJKOt/tSYihf
JnE68Q+KNzaQVbZouJnw+GFirEWl4cDed83UmBkiknVCfsuxZz8zTvTqPtni3eOQ
kE7nqbPgWndOEQJ7lJhkGbyiM/3kfZpw6+tV8lG2ybVpUGpVgRAZbnvyTUMXQmZI
nQiKnk6uHFFEB0cYieO5Dw3zwnr2+qaTUjv9cSciCBXi31mk/AL0vZQZHWLXxcpX
Jy0tVP4ufaiqrTQlsIuBpSSIS8xGVpZ0jTU/4k1mEEjh55jvQp5isRH+yS8nT/+3
7m67GaumzERdFekhJUyIwRcI7RZ4ifgcgTGmMQXKh0tsEJWjzS1YaXWJNGp9Hukp
YhE5EVfYuCiKYFWhnBitr5AySZ8otiWS2/1EX2EsoIQc/1QNE/Bn2TJjtGS5T9r+
8dAWXYnB9VMGJVXjSB2nsjAX/QWemsqygRfTeTJAOj1YCBDvfEg/I7sy+D8ZNVJt
qXjDFAzTHfWD4K14jQBT/c+jtsksZIlp0zgA2++k3JcuR5SjrTM9DAMAW9mGtg/Z
EMHLfGHbxtmkGgewKiMMHazLofUuWBO+S36HI5D6nCGknodfl5OQsZ+IS8/2bnDT
Ls2LzXABQJ8UjiLX02Ai4sBxc2M/8bm7Vbr6mVqszBN0eDogKRRJGxOkSacr15by
D9eF1dXLizZ3GMSkI9IJRi01wZjRDvL7YGmupaYQqr05n4J9F5jvgohJuLFWghvY
K1R18ldEw2Zx5zwtRn/3EVboGKpaL7/dQYy1TdMewWstspUN06OX9sTr5/K5sKBq
a98t9HEotPRINOw3EbzmJMXSQrWbpXOqT6yvfyVUlMLK89VX7Q2UdAQKaaZYibpp
csSgYzt9du0MqZmEWiQGqBGPSA009zhViJn/vlpCMlFaOuulON2fcYCNfftK54qw
nF9gu+93ildn49S74tedIQfhjGk4XyIeAFPaOJ1nzRu9SSaRLOy4eePuTjn/QWcb
5AXm+Tz8MfYcKW92skto/Ohjk9LC+nXi2q3zvHALPDYN8zm8b3fGA76NJr+62wuI
MPaL0Ix56A4eMwmUELd2yBPEpqnhsHouokxW+dm2AGuaDvlY9G3vrtlTYN7jnuCV
L4oi7mcIbPNFZmseRJiOIfBJnO+KkKQ3fV+MTBxJOlzBcC4FntIb0Cy8LrlOXH+d
yPmYkrvq7sjBlaon7kPCORb46fH7fl6ConslDoIJlRmL8hjMQ7g/xobVAt6HdgBi
3MalChbhqKbqjEEgvXiAnOF7uP1ye3GUq7P87277fDwSz0V5K+GM39fTi1F/v111
BlMH3THoPPw9rbpzh88XT2i+62hnKPCdXeubV1puyrWqtshMPmSrQIGm3nForwiM
yDuBHgVVpM6IPys6fQtrmMOQcebDWzESuI536CoFDBHvI7kfp6wsZTqqLp7Soab1
mgM3iGQ1z8wOmefFtT0hDOynI7nqeooXi6afp0ZSkUA+tjFjK1ag9JriT1/2Hhl6
OImIniZrHo4mUo51w2eJxdrxTxU7+fAPOYpUT2Aw5rtG6Z9OOT/i/aRsceppKBI2
br6+PPfnNNvXW6xoXvzT0MVNFFscnlMR2mU4nlo9UN4dgDWGkZgXbsfbRXnTrW4T
7BrzagOohXXRmpIN5fTOzGOK2mgaUWmGSXKrCXv1aiDmzJFl5A+4nEh0ZmFrhsSt
LXCth2qhIfZPs8wUxDPy63h8QhiiCsQTM1AL3wxWXVaLXRESGs/+SJh00i90s4SZ
uKwDDvNffZ1WHhR/eGOAeselTr6zL6MFODxBSUNoluSOLmQOt4Xfkq7mRbDVLkIe
8STL/y9CfUrAXFqbsrsd+vlodn6samOqppGTWT98HBivYn9wHv7MS9+pXZX8jXiI
D2SAeMHt+FP0g0YoO3wqUSDNMBJCnPa73ejZrJscZ+7F+fKMJkECci2fMpV33Yf9
d2wniWwIliA6tb7EaKg13i9IC886njvXggdNoGYfIyXLJIxMfAzGrC/fdok+4Je7
F81MfNcPoHNg5at5CoFpEjPUCEQTUzaTI4FkkLXEfAWgHQP6Ka6IQfSCC5MsqpEs
RlyNIUbnn0I3d1pYrNB4UU63jQDhyyKKkUrVAXPtvY6zJEQ/U0GuLUMyTpRSpOpw
rJIglYckpReI/xzM+VAVd7byCt8qOVGhwa2BFuFKnyStXxi/81n6VyK/30BTRr30
kvCwZTW4s8eGs5mjnuG25+K6O0wCSGplY+dCrPzMY0JgYN2KYYKqaocuMdztr4ah
xB+TloGkWGx/lWgra+zEenI/DzoSYIDDJ6/h7wwaXRWGyvsTpRS7B4I/fz4yRxla
BF1JbHVUXmD+rMXN+U6DRi5HQySNVB2cfhFfyN/7nTk0SIL5cTs+1gIn/4BgCpFY
dZlLyfLgHB48SHOvBWVtbnw3u4ToOya92FbLS2Q5tCYD+2dU7aidQBHqqCXlmFZo
tgXYI4fvhCisZ0zBOOvmFT1fKe7bXdZBzJwTzLaQLqzgsIUVz+YDuWbBK10wKkVn
f2cBT9DR2cvN8PMkQlqBINeadwIjM0Sn+GwXh+o10hm61UnfWEIyVVP6B8RhH7+Q
bgq6bXtsAeP8w8a6zhORNmAHzq5ny1D4zqzP6xL0qgLY+60jtG3eigLTPMBH5frd
qfXLWKaw38GFaQQ2r8MCjaiZwvxOuUd9poe8Vf3r/8PuE87XLuUo2kIlehAh0bSQ
HH9eiDrapX/t223TU7KBID1D5cRu0NlOxUv+pNMqGQf5OQhNUo1glK9ORYxsTqOZ
M9gSIfQnz1JH4xgHkJoB07JK7mMlZ4P0ar2wfWKc9qKtdec7+sCBls7pxb4f1Mbt
VeIyz5PcfBZRs47QK6S2VPknmRSPZUg75l5a4E5vGY9o+Sv8jB59KiJ4HTNr8u/M
BWmJo0nMmGJtvWk8Tn3Q6STFUvtRkS+2yAgNho04DS71ZJAiWWNnOnYE8H61vTIo
C3O2SapyjKAAGKuk03c4yIen42rcDpZH0iOUkKmedATwiF4ppRiiX/mwX09SSz2i
9y7Sv7WvcdWjFWkW4zni6aABZaOmKkpfDQ5eNswpvk3OY6zUAGFwpaCkyfNzsY/v
89hBmlyLKkNBSoxynoWNslnfiIa7AJ8JCNaEqwdB2pqD9vvIF68/Zj90vNG29IZF
wCg1uvZkgzs3b22LrXZfgw7YzYAshfA/8l1jde3Fv1AoaGdYi9nNN02T3d1FtT7A
q58SG6bUvtFEtPTNFojPhyBNA/lfBHceW91VF8TjlfhxYHDxZnsGZjmvFGgiLGpe
8j+XgL2MHRVnYlsMdPWkYPeYJlVqw9K+B8yAcdfU0WouI4r37unOSkQaxKB96B5X
VpRBdXh2IuO7pNMnkzzWDmy9l6tyr1wKLfU0oC2D5Ar7wZCWMIvYAX84mjER8+QX
+NDrE7Yoqk+VxvDNLe0qqcgdns41+/eJcj5+GxPL7CDFyYerGW3EGKjvhgk8hHXm
x+KKSiRvB3/A4wpvovkUWmVLdRB7GF5Hz69hOXxfBFYbFl+kJ9d+rArop406ZBnP
WYqXcTqfJczsrn0jKE8ljZ2i5/zF0Yot5N/KOOmVWkhOL+d0bnqq5dpqqZAqG0UV
8xc8VNwGbzZu/gz8/pRyHbtCeBjPCY0VBSsDqlIC6q2JIdsPbjqTHTSGkMbiqRxM
P0qtLJ1p2412ZmJ0atYCIpULSo7rS0sOun70/Y0LYy5doVRzJOTsP2hNDyQXu8b5
RZLWiowL7U2Mjl6ds7lGL61P6UkVBiF9k0zdfcJD5e67HyVEYpbC7vFWFpB9L+yV
DHu4Sp9BP4WoBONdeTKmAugIVgEwtuoOu3JYu8gOUz15spBru16P7AbmGTrJdSWZ
XW4YabcYRYN/K8YdCURrGHgCrRw2ZWZF+5YveKy6G3jzVJ59ztBfg6zH/rzSI+2H
gh99F5Ipxu8P5OIDQOSSXFgPp4p8ySHVSWZwOdVrWmw0vr+gJxNgzxzyi/VpkzOE
ASQFVtoVq5XAzQ3RW/ELLgQhV+dyN1JcDeCheuUBKHMQaYvZ6hPYRcMRN7QWTy+v
sIym6wTMfauBezQlIMjLPtlN7g9/8WQBmz4iO2GTfJzOnRMTXx8H3zfMleHqQAQD
z0pt7x7DU1GIw9Dkh19ASL7pVGaMAmrH6Z1IWw66cd11YiegOnKgJm5h7hNGGBV5
4OvbWqaSWlNK+Fw0/Lp2KXLHmU9XEjjYuQzDow3IjpHs4GdPIefnbGAM3EzdbLSx
XoY1mmNg6Zc/y26XXmVa4Xqd3abelHbs2WodhVWNtRK8Y9hHcwQOReA6lFJutQvj
YKgnr8mpbKyyKII+wNkLWMRoHywFo+3ne5sXdDigI4YnsS+pUnpP6IWz2tcx5FxC
BNOyAzxaksuyOvtP2mjhVsrgAlDZrAtWDmDSBvezTntSjtaTUY6XPZVkjtvDLITs
MqMBJf6xVU4/Zpj2mxOHUbpv+TC8cUdB2T5zRY3eLDGJ/rpX3xbjmWaUun5QInOh
zPsUwBgfOhB7pI1Q+or6hroOcCV+7WVQvANpGYErRZhSlVrrB8xgf6u9Lw2EoutF
k3VjeHKAdlMGuiy1dv9NhHKRp/2P8EDct4X3TQ9JJ8mcDGTZS9yvVzexjtsZpBb0
MmpImNU7VrwZUnsyM/QZ+m11Y/qr/wn7/N9XaGBrtoyR2MD0IbOK+TYL5atv4Mpb
8tS+tB875+uXkF/zfsvqSi092OfIWOaaQFg2pjLx/EEuuTgUIAIxMCqF788HclGy
PXWJvQus9GG8aSO02kgf/uHHbd2KayGUKIHsawTunZ0lLIpEtSkj2CIByuOAKlZc
J+i3FyXvxCxW3EIar8Nqt01CvTEoGl8vmW31bBVEq8zvH/bx4uxzsPOCRFg90c8U
AUXnndpbhd9sxOsc/MH/NzP6r3wJuOkmzhQ6C3+BjQiIuXIqquzY475IZ3oOtAKv
/Ro5qrBxH57c5HjvbyG2wVnbgiwMy5Zch2pRmYjGWOAmidq2MCkHO1Z6OLkGtN5m
T3IDkhFKKMlbRjblLl+Z7dfGLl4oblcXRRa8EwdnXBFk8fND9U/8qwmLLBJYVL3+
rkDaG/5e3AyWgeIF8bCv7aHEbGjKlmbMm2FCd9QMK7dFwqIcKpt6pFpeNVF7kSNX
SazjbUYwoh7D7qlhwRMJDkO4oJD7ZGpCqX2l1J7/pzKxuFAJTrDwp4AdM8VeWgUe
Hr9LOYvWY/hxZM/5c39FogaH0HvQvuMgguUrnZog+HUwgXOTbHuRt9vO5t/d6I4R
dnM5V/5HzgKQS5HLbKjGWoCGWMQj+X+ZL7HxSixaS5iSJMgBeHlqUjBi62s+Sa1N
R8p3VuDL54/oxGcfmux2+CpVzvgB4Icfd3cdJHyyhXnxN8STHBVxIgdyEV6+kdFv
ryjT7icIhklTKRfkXRH+LVuEm2snStSziw4qzmW5g0uGarpXxM9zMAaownIVq9m/
xF7L6AqpvYuMhUFbgoMEuPY+mSTObkuynhHysH0MQhDzQHKPl7ibH6fbnNtUdM3H
sWYiXrEm5MGq0YTx9wUwI9xvtJ+4Zff7ea9CszBvmMlGKu2IexHyuBehpLH/HPJN
ZAk3zRmzcEONgt+VNlGpUvoSsHM61km/uUtGT/dYZJaUFl4Za+A8AdVUhhelMCm9
LX1f3qASBXo8Hn/w9UD9cJzWbEzKKpiTj7PTZBnG8CwU/ylwF6nu1ATvfgOlJhVh
L1a/CY0Qw7Wi5KVYspfP6wYa3kdZXmmrhpQXgz1DQPn/qz+OzJXw0FgSMONCU4V0
2CJE3bEzljRfUaIHvnpddY8MlHRjxVHbqSskzGNLi55xI4jJE+qMECiZk/Q7SLqm
3dC05dshtCAMVg/t6MrpXdxsjST8z1uINdSecVP/ZFzDQ8YGLCwn3SNri/miDFXO
7RP6q1Nb56+hiEUOpmTgqFWTdLqv8U8yksM9H2du8h99jc5W3wBDY4m1yaUfZJPN
310EXXxgsuQgQPeucQXyP0XRBWF47MHS2VxhG/jZCOFB7AunMEH4hLzNr4FU5k3L
wmEtOOcgPg6kNWFOww6ILJzbN8hUsfom8P0PJPdMmZ4gjxDXhv70GYyT3jDPtxxV
m/ebpi9Wst8XskpYgWmLWuY5UoYFzpPJCKmgi3K5MBiecfxf7GbYooPWs3X9ucwE
DQB+KXbdcQjVYxz3PfEKu0ZdMoy1zfHzO2Fp28UNzi4Nb+pU4KN/N7Zzi1auTIen
q7Us+d5+AMPOonLU1XuYj6htFejAy64/LN5PJypFHAC3cqaowsR02o2Ty5Gzsf8l
KA6WFrJBj8zHmJmvWcZ1utwKSIG3M3YYaspWD4IkJMtDBjWydEF/RqBIB99WPAYA
tEI+cf7qq3e2nYS0mlsDh6xID0v+UNzTwnep0dIfS0inVg0KAwqFujji3GeTIUPd
udZIBh6aP+KLORhfaiYu7TZsIhwro+x1qwVbyn/GUM5lDHCllEHumOfXYgK8vLUA
JpqvPt7sMgN7JUfgQc5CfHXt7DiiDYUYpeVw8P1RbURgI74YiShmlffpXL9h4WdO
Z5kZgYIeKPKrm+JT4CGS7anIi/761XECjoO2aM7mb1hgyzNq9dyPtHsHMUPUFfRs
bP9v7N3xUut+21bOt+9TTXBe1uzismWOxzVFPBnGhV22VVyEUdTgt+xP09V3OFGY
79yfoxv0frbOMyeGm7tRttZ/7558nhhZwjOBG/eCJsiQrGdAPvGzVkwmt3fRzbae
Uw8JneLCK+IzRVANCyak2ur/XRQhdNNrwVMHEskP9a/ZxAm1Hdtv7hCr8jWMY5I2
VCk3DIgmqG3Wvaq4xe3IZTS23+YZZ1gdbUFUDOwiUOunFtFHaBJI/UW5YU4J80DD
+dYnOYcDQwWc5qkF3iztCW+78+3yJbKfse7quGStn2b6BALhkbuRmeBpbpmPxpmo
uB+ORwjRKApbpoegtsdUYV1WrS6Kxg2WN7GJRE/e+ahy2G5ybiovn8LbBOZMy5nU
1PjwWwSkk96TmhdXBX8138ASLUr2dCzOXgPHQvK/7WkNujUYA0I5EsVLkZ3MaWwH
zAkZOE7nLXnS3kEzcQXurRwP2PN1scDTH5HW2CkdrvSuOC1R7oquUxNrj7uCGZjY
rtsTZjwfsUIz33zVzKvZFJrRvREqIz4tJLxPae9APnmkw6ptdSJNfW2LjfHuKPy3
0JanTlcirsZqDDOpJHIBmuitYWiGAIJHxCntcBduDVfOdK+cV4fDWyUKyHHduw5m
7IdSWN3hrrULjjj/uZm8GVpV1KlTsxQq0nUizjVHXRK0nTuRxlkb8AKD+iAhiNiV
sdalJKitlIX3N9c78vpQCi0FMwon4BhilrCQRDwkeAREZYKTOIPyz7CCTp5PThia
/ecU+Pfi3NalhjTV0OSSzTe1PnfSAPDEpGpN5cjDjCfOPKuxBiSE1J7YxdNJ5srr
3G5bxjEX7SZFjs6teyCV+/Wig6nHYBtrC2GbxzsJWRz/IW1UmcsvZ3h6t6GZtfyD
dC58t6H0J0B90VNoOG1aAsZSKIvVLHHIXCEgaxdIP5ug3ktqIHvYYWTgvhrlhwAu
gbhlM+4OQAstx8yBBSzJ9WoSxq1Vz4IcbVe+HX+mZeDMVsxNjAqn1E5Lnshh8el/
0RNFvm7DItWdstkIq9+VzfdDwSHWkCKznQSPVkWrpYVPjlQYgmsfZtBEg7TLHCF7
zft9usR5MqcS3xVFVtZkbEcnkdykpPSewaIqSIOtWwOsLpJSBxWm/6Pz8bYFwDU7
7JM65Y5EO5lqAVZ7A8/J/6l0vNfQHczwAvMOAi7XpIYPWktIiqYLe4ve8D7NswIf
I4NsnHfq6415EesrcY2wckUccImhK0VgLQqKjrcRuoYH1oc7o3h7fZMpS6kL/ClF
4viqlQzGyUB1TaZspnwA1abTTratUKszOAfQvLlUnYHz04XigGpeSMSC3TfzsQLJ
AbA4ToLD4/fKW3KmqyqiEJHOVzWVh+R1zKJpZ63F025wXzVdlSCO2de45F6pBu8N
Z9AzAKCd9OH0lnwxJd878IapetH3Lnva88Y5Ep5ZNECp0y/0qgEzWZdt9oK2XoeF
wY760K1b2BtZe2hYRz7NQ80sLDwnIXXG+UnPKftSE44H3r+iDh4N7wrdSt7mZUto
eqGsU0xtNpsQzNomckN+KWR3Ms93hRpPCtHyJBHvM6llyw6kWf/nPxszfVj63MPh
oiGTCofyXkRXk2QNrlUdBNW5q6z7ROm2eGYojsqZgS2CCZqlgUoWTLMG7W84oyt1
XwV7mc+8xu9+G3eLkZUhqIXx4kKtQm5FDmI6+tzzJybrVsmn8Fjrvb5ONUy9+40Y
AY5GlvbxLzpLXPLa3Ep2JdplYTN+N1QSqyhNVoNVmhPJ/Vz58KFXOwZ7THVtwOXa
csIYOfeTvmt4li1qJSHWbnNDQK5gteuLDUH4Edm/YXd9rEOgkW9K1FHIupMDfuaS
Bs0vKhd3o9HM/znqlZT8uJan3n4k6Zqc2lE4+rZjuT5JWLFYK/62gSXDautnv9Ep
D56zZYS8LyS/6DHDLG9T1ON8ntJ0A6ToyTeo6LrQflsQGziNi0B4coi5YND+38ay
VBuj8T6OTu8s4Bo/8Tq20FPH97glfh8Yzce+n/5XWDfo3dpwAyyrH9gBM0g9OYlM
tvBm23aYS52nCQAp4nQaU7IxYOC9ACoN9fsSX1NX8F/lAQ9VIYJYcWXz2zLu1j+o
P1q47xEQULDEeIBb4GiRjiRDe4X2mQu9S6D11wPOGxub9v2TFGlJYlI1MrVQcqsd
TiaeFSM7fYTiYT2RVdpac5JFAY3Vpi8P0n/Bd9YWzb0Uutn0Wd7SvIq9Ct5SLkLG
IKfs6ZGnrv3FcCVY7I+oSvIDhL+MBFV9SiUxHjYdu/IEv1XNOmxUKepqzq93ONut
wnPgdRsI2lEeoz4iDFmNVYjpBA1D6DtG4WFFZHsaVyWmXzSjLHyB7eg8kW4WWA1z
arJJ9r/TGyeAQREHHVq91uLBgkQPI3nzLfnCeF48aZymqHUsBADPIRouYurptStl
Edjv447QQHRZD/598tBKoAjt68M4aN1XTyl1j86fxJOXTZR4yJ1mscU7gqoRDEvm
YhOp/z4I7JU5imJfZ7HBmJUH5FEyEdpTeXZ+efXXigxc3YwK+fAsI91wMg6g/vyV
T7ksh7ShpjmkJPvRgO3sNuKxiDNnjOLV59RbkhQy8EeKjZN5AH61D5LHrb/D/VbU
Wu5kEVMcLJgjwWggNY9/546I9HNyEFrKJ0aew5O5wqkZ3oh+Y5vpKyCDWeHdeHAo
Id67QgSTFGN3n6ZdCbxonjTOnXAyFG1EfMVB8qsiPBh9djYnmXtXOWIfc8Vk1bsB
iMMSK3YK+nY71JBg6AFSohm0a4fikVl6PWvqL288LOeA4oXQq0JfwXbZMrniAGPE
PQGltILfuKs7PUCkJIs2TbEKjBNegqVt7OVhscH6gaSjTMA3Ci3rM+BocCLwHicf
KWg7raAytPhnSk2KUJD2Sk/reZnFaOa2QtV9DZ68gLBD51nQ3Q+Bmfq7G51mFtah
Nrw+ZkOCItekHLJPe+QdH4xnd7hRLO7ZF/SdIwj8L4Ri8Hh5mUJohEMzB4rdJUTn
Laql/ZWV2rZCvD5/eqhV2ahlQEun1KA448TfcVAsYolEZZi1Gh2P4eGszmx+Hw3l
Az4qmk16ne1PXKW/PbWMSiMhBrtRlCr2BrLLY/KTUf2OKaEVUcQO82c1Zen6/4Ky
iOSthJUiOlHDxG+YqQcXDf1YoiCBYDrNnV76ywMBFet7vYknm2aK4+piHulF2D2J
8X6ImyPa90ipboIjd8uNyeLT2z1qKZILBabdvoM5M6j/L5hpjfkv0Z9H2PvFPWLz
mDBX+t6/yGduq767ak1xLrRv6gWUxHntaXUAcV7fSaKEpcCEiDicQaCVlk4zV29i
nQ5MVqvL18fObzczFSTSCOJ4v7rXQ3hJBmOfPFaeAOvndkXZjKAYtfC1amUXry9f
GCHsNbH4LPY7TU9OaYUD04lU7TcODTYoHR9G+RlXICITA4leNV3+m12tSoYtAEWK
4mce90fS2IODfZOeWvhllmhAqhbqd6PGbUjnHqzLknBcd0eRTwwmUH/EiyO8xYTv
iq7S6dlxAyGbLwclKkC3UAWNqd1CCGScB2ipcMXTf75ItCaNJRH5pY9PFE9HWUaY
4XqFtRiS/kaRxkTLzTlmAFQyOhdm/H6ei/TIMQQ/DFuL0rAOX0EBtQP0d4IfCC3d
Srh48eI48HH5M6H2O/2ByCpDaBh2Y07GIDgXeCoXYyfQHOxrTiP6lXU2QC/xgKu9
Mbuq3WWu+yeNtWe7GHKniZbUvHo7A4ub0zK0yusgvSANfugxM4pWrxTi/bqMLjQd
jm1FHmcXH9pfhl1KX1uzW87uEG+Ae9h5RSfBrV6/wd027e5rhn+gpDpZ46IMsH85
mOTX5tQTf+XQKVTllmkbWX3lr3uvuiZ+hpFBRonxLbXsfls2VhRAyVIf+5OgnkJI
PJxO6bRMScgfU1tEyOeI7Yuey7c7gLrQCx6M+Z/yFAiooIdnqTcM3ATc8Lr7X7Kx
45Xn0VVsDlxDdKm6Se5EqNcXzebz3JBK7yfxFhI2DmAroaeucK8MNz+Fai9VuO7V
cnOec6lj6EgA4nUtNr9bw/CahVejAru/I9UqBkWcnm8bvVSB0S0T7y0RHrfY7QgP
sAqkO3q7huJ3T+fcvBvMoMvrhhjhBFQY1I6hAXKf+ZqftQAhanu6b3QAQFZzJBlE
nc2qQbPHz5qAJbELhod8Ke7XItzH8T+NjrIQUwJjfbcPjtOu79uPQhwCdQOVRjUm
OZzdyBM5HAWbs4nj98Fp99ZGBCPcPv4gC4H6Y/uRKCC/jZAlJlK5pFi2m3izbXns
tDo2SsldPGbiew6a9Inf4Ttdc1vl8uuzmwZDVzCIOjxWHLdlsFrHUHpPLRwtrAqW
/nP3B5jxCeudnVRiZyAKI4amGafjJyX4I0SDICupO2WqJ5kP0GyF6cTUHkCepveU
uZnp6gmCKr4DDU0pd6U76RdMA14GY1A3RqLCSwVEPKXrf747xDOv2/YUsPsyniNy
26Ie2yuD2MeUxypIsyWT1bGypi9XpGd8YcxMgaVQBePNMUiTGRp36oQGd++gY3YF
4KmGyGX0TZ8TVoY7/+q4cksEB97IxNIZWz+5o0QTqhnlOdtdSuOXZF6ph8nXC97V
UE/dOB5RPqa8onjM8vprBu2qYYEK8vwWOAcxt/z0I2Iv9wElXTl8gyOD7TD6RKOT
A+HOeEa/4gYb/o1ryG4M4MAm/YpNmTQIw8wVkDc18651Skv3fidot/MQzB9LwPaA
OQZNaxXuXMVB0Qy5lXRBKeinDt9JkrphrQtgAK2GNaqN7vk2NPyAIepqvZI6iqoK
w/BbIvLf1X/JLehJSUoS+e4zrpm0GenJSsDxmxvVOIL/En+ngOmr/BTU0y0x2bSn
TPT20MLu8kyVS5pEiJku0IczcQsov/w3GEWaKBHIV2y1UwQymHA4nTZ5rRbTUYix
VowIPow5BKA+eZ7o9kSnca8FJZoCOBYI2w9OEraT9Fz43tjivqwm1qgHuTT3EGQr
l6ZH7p2evXYj/pZ3G0uRBuhPDezfg10Z4RbaXS5JXTP/a/G0iWG+0vDdw5yOfoZ3
9RgzpGaIitIP3WnQA93sYfek/nLxqPH8L06nyYOZ+65gUJOCHGTXrruTVG1gqRK9
ttChn3+5FokbQfcYFVZDn2qURACFwe+PLCeyJc1d1Ku7iAtdWzJXDqj464dEx8hS
v+wm5DO3hYROQH1nESrCWGejTsmCUYO2iMio4EOZRJmQGXsH0fo3Y9T8GOGhvDT6
38fmWB6VfHy7K70voJidm1txavwH/YXskRu+BNo0E9cJ7KRkg+7kNUe/RlXR/OWx
1iwOssEbD42t9YjKUSRCFPdXoI/ggh7vs6gWTRf3XMLeZB2CYlalQRDwszC/cmA4
0C/f2swCU5nzOK4ta/uQKDABJBWiep45O1yYV6m65wFkFGpMdd+ez8d7cf0GPq9i
/IUpNBYk4w7YgUoXGH/CEPLr+bgS2LssxeO8sShsU9/+UZ08aP+dYbaCIxePgXOB
1j+LtUlzYEtC5kjpLP0IoZTk49lfOSgmgecdU1xDkMO6g4CiAraG485paPconDtf
5csJR0ciQ/FW2m0gtu5BOevXkiWVot+OnHfHDgC6Ng4Uok7QeNSfGgtphqcwhaty
TPztqHUqn3HyMowJZ+6Ude8QF+e8HMDdpppowyRpu4VUEpjRvgo5wRNgCEB3Pyt2
MegXh02GY3amqkKAyaAdnRLbXTWsCi/LKLdMcrBn8pgxR2jiTPMAThoJPKribvO0
npyVVAayzhBZQp7h4dmjfSemH29kxvAfo3ki6f7HMWHJuYjOMnAKhVVJkFAEXEc3
s+ff5uBdj/69xcZNvC99WMXkWZnYINyzq6zee2ZHZM0B9yfWxscQT9CKVM75/XNG
e0g+KezbDA1vQ/gH0Rv2BMA0gm5dOXKf8ug6W3vhECPAEkpzXCHxdDS8+n+PMQHb
ecaVucEC/UHnkSd++i9wUY3SamEsf8YfySbsuPu86Wym95pqt/+f6QZAHLpwTNvG
UXW/1cBFrDvSSTpxbARl+ZHPF2ZWJlaVapC2qHYoTUjRMloUTn23OYerTb4FaWXv
Jes6hV2a9ZXn8G72JtV20jM8JUiFmu0IJGf/XrGmmlcAcucynx8Gono4Lr5Wz6xN
IpG3hfC3eo+/ecWAdgBkS29GSO2TwgBQfYYHrju5uZX3/XIO4C47wdQGIBP5JzvQ
z1J3PgTa7MISr3yH4wiOcnzZfotkUHAZ+rjDSMg7x2bAcNtL1+paUewYvN5+oVC+
jQoy3QmkmRNm9ZFiB5s26l1urHxwm0Vx/BYMVEZGEEj+jrdqS6U40Mhi3GpMHAcI
wq5xkRP7dhE3Jhx6nNq6h/njqkXrBvgc9qub/XwiGp4zFEpcIq+m6sXJAB7lg3fZ
EDqu+YFUm+RabyeTdRe4xAOfeJpJ3dOxVpXj3q3b2Emrl+p0mgz1jYB/HeqULLA0
jUa6zn6lRu9aVlj46zQQV06o6LXGf2FqXgmtDLIWGKHVRALHxVOSryXaIIl0rS+i
MpfJYq553DELqMvtV5qieZZ7p1M8wknwRBRcsiPsDxgAnH6TDl4tnvlNK5L9TMAf
SAELaZ6/TNEHSc0V+JKwEIW76qZqiYGzgDFQlpZN3UGOkyIvkGlDVdvuIt9pmlka
IuFkTVzYuH2qoSAEuGDvasB0O3ETalj7dlXZ/2+ONf2S+wLA2hIWrgRpFdtmppmY
GnO9sBgLjeTjCoke+y3P2Un+VxNiwYwHH7Pv6KokWtSh1ZRydQTwEKuIxHKRqzvZ
/5q/Ey6Yx52GGZChn89FTh27OXSqlNiYo5SNLys4VNIPNSnA341hdIr8CsISIh7C
VeKRAbKQVI2/1QrgG8Ku611BoW7p7dLbo4aK6dakyy+oWdy8KdBz37MNPttZs7hU
XSm/iJWE86FBMiwAXFqYRANIFrDrvsraal7B4vK4ZOkw1Pzb3xCd8g3B3MoxpgNw
TIOI+eIwnLVC0UxnrmpDqx7MKY7sS4c6aTsSCehbGRBJFpiA8oltezbui9VW0UuR
vWIDQczjg83ZNDMENDKXCE0O9u7uWr6koN8p9nUHRwPhJ4GSklEqIU4ELYgz0rZB
zn39RMgEIeOhBQHimZfh9QXZdE7WU2A555q36SogwUidp+8KNDfkSLRskgwRpWoh
yPGIlhIxG3NwhBnyfZLWNZHyhbdu5D4J7rJoMeRZph8mBinbSSa8T3ypgACM3W+x
uBQt6s/4OOj1BtKqAG4kw9qkA7dn7m3Zfh+hFknCgp7aHeE0VL2bzdic5OelPgSA
3lsuxcEvZF8eyohkAUKXN597t94NmgJahNlqZ+A564zsNHQPAponIduP3U/riYkA
NP5lC1qqJ7Iz+kEwuj8ZeiZDmGy8QxW0Il1c547UCMToJAk//E+1+CxnwPydinip
O/cSbgJYmq/bmcklJt32n7F5CJI7SSWYxlF9bYHqTzqFBtghq17Mn1D5wpsGJuQX
8XgpfRK93pi2ynOyFHC4Z3ZpbtaXQCnWqypc7EYk0Wjm8hbQ3k6yh1XAP56ZeUUS
WJIBohyJIub3W4higlpIcP05FuIITacE8tOCHojWejHA0OKoUUEAcUerRnzpctVY
PErFXZKxqmcu1uq6egfjgUTiPKxssF3FxQnXPB9ymPUMikwOvzdY86CxTIAZpLzO
xOQk/RLyoHoDgVDpCE8+/jA3ivERGflKppS5dr0jcD4Ho5db9aboXXFUlCeg2xFW
mixL3qNLFKLXrjjbfsI4A1KtOGHaJ7dP82P4w+bmKvJhaN5pLAtibcrH0oZzAVmJ
q/ITeaLEX153hjER+dNIAWbuON5xLYIOjWvkbi3RqG+rYSzGsnuP+0F7hIdChxo/
I+ut31eEBXERpkl1Oj5rDE6RXWzsDyqhGPFQr/+95UK+bXa1biGcHE2dDyqDFaB6
HZw+D/wIAwaZPO/+KhJtKVLUhwxSkNdUk/IQqxDD279JjnZTFRWP3RfPEikbhHtY
Edx1oHhcaqj3BYFgpPeDfFrzMdyW6BCNU3YxioxS7mFMSbdHsBnagqatAnx4qq/4
rIj3Qv6llRj+43ox1uXVuXTNeKhrCt26ABqS094BFgENgyiGduuYspQo8SjkPRWz
15qWEGWF0aGVJu4ZPU62PKm7yPqumLuPXk3dLlX/VUU3HUHA716hro2vy2jz6nyX
c2oJAEncUZSWH2fwFy3h91KhyYRtJsSlhY0trUQP7IRCenXpCm1S8KXw5lCz7X7f
twOGy/OM3MyfeHOnDs4LAblFq+GmLSudzwXxeZ76jjh5nrCXtY0zm2xc9mLGRO6m
Anox8X0BvtLm8wUiXZ0pkBUTU2ChVhEO7RKcc0PV3jihGIuZ+7Mej6a0o7q49WGD
RR+pLWgW2uU3SdWfu/yl9Pb1m4cfb8LebIEOy01+LxItpjP/lb9fEo3heqdC9aJi
tfGrpsvnkkO1mTNucpUVhHoCcp/tvdpuPUbftR0Y15ZZyvHeWjGhvKrxt+DlKV6n
DtlZyKMflSKaCdikaXdXZLnUBQqSy6ari4yXVLdndIH5tjLKi7ogfIRfCP+5hQzl
RBt7RUDBolvHVwtiPpGbvCI0egXJE5HZrmv/Ydecp3HCAHmqbQzzfO9RxedcHlWA
y0Or4ASms2dj0RXrYwonzVeeKVoQDf3SxFEzQF625g4HzS9UrBsuJksrkq7d6XtG
R7a9oZ1tSV0lafyw97U3uDA3OdVypG9z2D21tF0Vn9KoF46hCYJp/qzqwuyLLmFg
AxaMsfSSuILVgMoSwN+OpKdXxdpikdBExb+ybw58FdlEk8SDWjAfscLynBPmpf16
YbjdBtT2V9EqWPZ+pL8bVNVYQfrvCfAn8OyBL6j4SPHYsBjARO1eeE+NSvIzdBbh
FN5efCDKmdAymhl1SlX1oZkuMRnzA0/1j5HImj415EYFtA5N3+3v9dmjvXjOBveK
Fz7duA8HGCwqsKshvvBCoYNgmOSPhEWDLKCQiZfm6ec5CuLUSpzqfMhjpoHAJJyH
0U1MmvIFcYmLy5PTCqPm29l1zdVQyYWwSU10hfAhJZq/84Iec9yHA9cz3asgyYFd
dHVg4f8Jt8trLu9gP91m0oP2jBdtOqRLWjmEVgC3N9ajJr64XzKgiAwhY6dNi0ys
knldPUjcDchdJpWEbYERu3DMEn5iN+ul7TRW0Txp5HXOT5Ob6ebBl2ml+ax1eJor
pSVC7Ir5fpBzXaxk6OwY7wBbeH7G6RIe/YRj8y/SSkWphWv7ukgLatPMPaEVBovz
u2uGfbYUH9xrfDrbdHSbESt7KTxWoKonypPKLCk+t4WwKHjVUJ/FxU475g7V6+b+
KYBb6h2PbgGep7SqhsG+DoxZmvQ3jDRsE65GOFclTYJFEb2qgv8839F+lNNrgenH
orzjQaAO+PWcxoz+w2OWlyYmCLwIdacODKBoMaMvUi0tYdc7YzsuVAOsSJjRqxF2
kiKbmHZdn8trOM9XPB7yeDu6tErJ3wJm41eEO1u97uIuxrxbPBBB9qwALllOXifK
EuiziD+ZEdHXGaPeN9nK9eqjltM6QYz/SJhrLVLL9NL1wcqGpKgIZwKLP2JHKeJI
nxJVq6ZYnsmgVpc9HgW81QVb3V9BDOiHQ2dLmd22gUNJDFKj3mWPreGXed/zTQye
SA8FCxYwPXHRU/WK3leaRszu7eXcw3JVB/d9H3OU2KAy0iAWBkfzuy5UAEdT0gTu
fXsy6qvttrUb44Zjuraiupg0bIZhydst+X63fBLNkSeoVAmgDblRiUay71L5pECh
cso5vpQw2YbMPSsCm27DbEtSN7wBXuyEIkEfZ5jQMG030kFnkXKfGo2iKYhTtxfh
LPoewUNdC4mKnqLgk/me5mW3PkLrkrNNT3SY9u/voInIQIM6PLqgFY031LuOWKCF
X/FsbLP20FULdXZv8G7qdhxkjqo8+oJWSN4kFsIjLDInTPZwxGx42Zk61laCM0zG
bnGf4E+CNHk6e/fH3MOQmIBPDp/WLZTWlllIrqPRnwrlyBi/4gP4DU9gpfc6Kobp
VU+9gL+fke2XQX0lJW2g0xlefYLWKNK2PuDUMeDKzO0tsq+tAGxEKCaAZNu1ddJl
ByITQXNVW7VtWrEGXp7DynhUHDfhMRTnJJ8GWX6V9dnsiGLk9z2gCY8OdcNRXiNc
frZihyJJMyqRRVphaKokGl0X8fCPra5TTTF4DmrAhMLBvPK39GHwfx5EZvEdT7i/
JNIv+4koHjCHsDh7rlzQB9YWAqmGQmzYBn93zsn3H4xhQGT5F+xkzNSVcwvLeRlv
4cpeilbk+hrzmMr7tALXcH82j7FQf7lrk4njbligpQCf9ogY9/xWMfKoLv7KkQUf
dmNUWbetgWnpWwU2YWvpt82MV8MbKbPFT6hIQ9yQ12jH+I6RuRwb4b+mIX+JFROT
lIpCaFlvBNvUwdxVyO/jA/rO0uVkAvTdPBm0vP4AV6g8nc3UD+cD38FJRD+mSbtu
IaU0hSBNUCHHBwQM9KvTFrxxlXbgFUneWDAdmXcC0pjIPSowUzacyx990BDIciPO
nAUv4y/ewBJZ/MogOl4kFd6jv7oclDVZUzd8sROtGhNgKsZpCYEgAaQ6vxB7/wP4
qBlOgjaKoDpCnrE4yB8Jor7dsgZKvWakayX+WfJaLcABV7m2M6c1qFRR/nnF5UOO
2dZVBPNR8zVMwrqinssRP0SV2+UDsZUHc56Jir4JiRK91EOCsGFzzMae9S9pAseT
HVTjKVWsE8TU4CGTAxVCBx89LMPlgfRovOgXCtwJcM2GDftCKPDgkfDkZ6qgLLtf
FTqJunTziUmUFKwPK9m2D1qGK+U30hlXsSS8OjqPsV1CLakp4gG0odCq3UVXr9MX
8Ylp+Xo9p0Qb7quVsarLKfxIoFfNUkvIQsXoGok2P+GJOZBb1GRiEfjPSXmb+tS+
fDDViZa7oVS6+jsUCpGXZJAJ1GN/5vUqFuQ9JrVpQ3JcHTaV8bl9x/FWreNeMerQ
GcvyZIJd4kZ4vyoyx0OYS1SZv0ydJsgh1bWzqnJsE4xInq6+lNXl4n3uUm6L5fhW
wbkHTzkidNOob32UygYx680y1E46szAMXKV/lTJXuNGmmSFGxrmyMMzaIGFI4tUY
orzfR+JNkLtDS8VGgbiRnshj/kAoIvI+WbFdABBqpaHQjOL216ilnKtcvX0Myp7A
8GRjVd1XP5PY++sddDziaF2Wv0aoz2+JPV3YYKu6hho7Xpe/tnLyF3vC0gx+mbBa
DBwcPCSTjPWw1VYAr51YMdlztfBDuuFO5/BegW82LwiS9UOrz+bJTpDqaTevxqg5
EMQKmWwH04EdQoC6zaBVpIQn8MP1UtzaOvfNVpHTXZ7ICqpls0FNPRLHiAa1lRR/
yL5zPhWam4vOwM3iYPLygc8TOXsii9VD+Ob90RqMVZyxvaz4D6eL2gN2SQdQj7Dd
iUqlawxoQDAdZjeF1P+dIkzm/FVRf7BcteMUNXU9JvwXdLRgc64psWCX0IJO/Rt6
fK7SYCRkDOnIoLoqeBFcks92K/H1E1CHiNKcpCvNDdyXfQKlAXxFKSkqFwSKnzGF
GN/oP9NJsr9dP0JyMkShT5EF14EELVE/qSIFpzpwmmVz5CPlBen0gTsCYbEqIfqE
EGQPLmMkaxvV1JKC/2G8fbr1lccHNeL9zKi1SZkIBbrVPSdj6drh1DkiOD+rZZkM
68LdahyZNwWyG78rhQPJyNMD1hXmL3Lb8jlMPk169xVY+ddIdywMYJfqSDYOMh3h
LJmh/s7cRaR7EnePiEq5Vjdnw2A5I0g7G9ZKOM29H1ngsZDEPrr/mIcgTrHjqqpN
PsCYfGnGsNW2IpDGPQsopqtWIZcAbcLv2Tg0NXBi2axFooHQRsx1EvzXPY5oWFZj
AffYvP8uN1SBhJv7o20I+wnEAk3NM2syAw34U8w/C9eu6j9qZMf7+WV5zbLj+QiH
6WCH4y2zWhx2oGLpVg0abPhlCKxri/a5kDivkTUkVR79V5ZkFYhbmvLe/ev3bK3J
BWGxyRg5TOja681BqHChHZSl1AJyzJGwLHFNhP44S8nR9eOxJHnLOi3LSjEeWaw5
9ZrL2N3zZmkBx0Wy/gIUEktmjz4kYcQeiAjeTwyiHwtPG23yzxfugXRbeTOrx20q
5c4us1zUMmRDLxukg7zKBtRYLSZPFXek2r/7OopxWR3OkHWLtI6AhpKCog13hAOE
8jNjrO1gUlxdH+ViMiT8jWuUEu0zXzKMKFdaWw5kpw0u0n5LKEqOgYA5RZTYlcFi
gHOGtXoIAOXlxa7slLL5gkDckM310C67pE36yzdPzE1rRQBzz2EeIcnhHRhF15CC
vun7msY+X1w0vpVpLz9vNUklHCBc7G0r8FbalKAguz09RC4+K6owmNABrJ5Kitgs
VLDDRlNSTcEmpLIkp4WaIYCuUXt8dmQX2M+HgJZUmkF1lRM5PwlRMP+56FbON56q
6ChA4dLdkVTLKWio3JGBKkjLMFEY6FWy8uM1Oi7hsvo2qC3+bg5idAxzdPX2sK1X
5/ZW+y0PPTHGYdn7XyciX1UPHqCYy091Ut6z2RUk3PiHU4hLS37cuttcOY0icYjK
hF5W715mEei+GbGmbKp9Yw8FBhJROX0eN7FLFj63ubzS9f/g72r1GG1yyO/0SMb8
3YPbcQN6hvNTKrdPyUEdXeLEkwDA55C5BEkvPs9deEgHHmHhMGZZZKejX/Zinz52
uvcyRKsY0+zyLjj9iwGGXOeMuPJRIfekPGBflL9HOMclek4uRlDSa6HGsF5DQn/B
wflHfPFe23cfKHhb1iKHWdQHe22j4cqWqhgRouOt+nxrizzr4qzZDu2vWcNslDEm
QL52Djkp2edi+8OO0hBJsloO8jZJ6+qLMYMAEqPLhGXBMS2z+19nc4HI8HwZ4DPS
Oa2WaMDtFomXaXo8hom/csvlWBJlrbCk/EteB/qO/WFMjKLLyIcw7y7YNCvZziE2
WSk7crCr1SXy9zEhLAS6VkKpcToNc572rnpwtlm53fR6P57jm664+/hKyFQADlAQ
k09zgaOVWgfp3+Cjj3oyCTR/ae09SuOWs8nVZUIKMTZWtSYLaKLMBlO9Euzakjmz
ZyDZdcFAkhPAFDwHApbhcMQlL2AIJGHJIuCjD02l6+tn0RGB3HLN36YKjYEdTZ5n
kEYwVJ9CjQJtrSpefZedy7d44P70nNpSeSLS8sM3GMLcAqoJbCkAlrabIzoHKxuD
2E0/451j3/QjpnoOlwRiwx/e/P38K8E+S7xC9+XzgUhR2Qjsa7VvoMjoD19O42Or
Rkrde8iLJkAr7LnXuEypqKx+CApFPdGfUOgqajcW59SZ/CGw/TMD6NfTq3uZDu0K
hBnOhrch6X23afbFopCD5v/taYIuUFYM5Rqjml4t5Ieo+9uO8x2RJF5JNLAfx5MV
wKAXLxlTS1Cmxajjd8rq28wU/cGTqMHhPBqgD1pKZaRLnGHi9oxOdMgcF/4sALXL
YPhwMhCn8qNUfEQTcnxhv+GTa/0ONKl6klMrbbYdXjhO3ZhtV/aoeQE89lqNZGiH
sEg0yd8pmJbFAzNj/9kInT+QyW0T+gl+818QUtkpb13l/2npc83G0CTZqtzoKemF
RPCA4ufkg9EY0qwfxzKXTZkpYipl2ljp+a9Rrvs+poTBs8gmFA5j2OcpCor9b3+w
DgW/Zpu2hZLbNMYKWrAaaSjCuipu7CgV/mGqCtFQLk4f4GIlmpx76qfX7ctr10Iq
jI49KzLt+DYEcBwyM1CxqBiB1G6TLThqqiWh9uDIN5RYQGuUuqBAheKOBLiakz4w
fSVm9PNFLdxPVFV9oKBSmYjmTrp3zngGdLY2Bb+T50PmK0QgVdt2BF2jZSdJJi3W
SAJn81bRoYzKRNmpux2qoiGhVjETBBDCBkH5NpBWdLaTlq+JEKF2VHxdvHZKx7df
kww/bb7VwdHVK0vX5YWFa7ZCxQFNxOvrcEjg19nx/euoFywOPyLZ0lPzVZLWECnH
kIpEVZKxaZsJsLvJnbFlfKTH+2k6vmNHhuxBqA1oJ03PdxBzKWcEoIY00scS6Enb
eXIrpbXrubzu5t1WoJhLHP+xiiPRZD2TQDgA6BqaUR9zM08rztkBZXTa0CbNjyta
FO8sloOsHyDA4JQ87uAF2fBDN6Bk1Hp2sxh5ERQOMthJlqoo66nsNPKkQFnSZnc/
VXXIxcIB1ZCkllndxDv9xjWKOvAXWUrbamwVhb9dLmhTf3i36EgogKp0a/jb6ixe
XybsPFJ9nSsqTweBPLmteZNooIfF5MEX9K6mV2oyowD1aWXDCpd2Arvx3yW3uN4i
PAtQltchfCqoTK8ilb3ai3L0dPBHpeb7c9JXXhvizfLyn5IvsmBmdarAgLYCQp3L
74E2vdPr0vbULxOYHYcacFAmNfNnyk1Snioq09SccVA2/60g/2ktVa0G6kzZ1qym
T3GcCu34tunIlJt6YxA1vGIp8ERnwgMOJE6KxNU+E4oM6JKb+WaykP5oHvNEN5QM
LmJnrRhv5R76pVQat2gVKns7jgHGIDL+GkZnYG4n6GVxAVKld3oRRKIdM4j4Bxpt
F6SyH8rcpBuT/QCLEVU4ZgORBAomePF8DQTZYLhHV/c+DhOAf0Y9aiiCvNK73mbT
QmkwfwiZ5AiHAOqUDnKc9BdrJkaGi/mKHhOqRYoVDFczt8BTJyvWdBEnImayQqQX
s9rwRSmWpuiCtg3PcNpPdmmDt/MMFsXj4yabApD9Ume5tRH1z1wTaOxlogBK5AFQ
/Qxw7Fgr5BHhxUH/StiHk4y8UhRa2uew1WUKsx9Z5c4mBWUD0H7T3DhLestVa3ct
yGvrewamGk0jbIBBklgLU1hqoEWcHdwvlAQkB8yTR7DTUBtcDPnAVdTBVdSAJXJj
L/deHJXXKovzkmV0aaFiIMVVV4ltUYbKfjWU/S3O+28PG4U13yQqG81x+EGROr7q
JDLMmI0AMDpPIKzS7MHjLb50MLFQnOrKpujBIHGAerSMNH9VSw7xlouX89ExLqbO
6rxISEiNQukIZ/6wg2pKP8rvkf3+ChIicNIyYZe/p5QMttcq60uGGonA15FICNv1
3NepybH9INqzduls9arFMglxjBappjh2a7E8W/SUTrumre03Hb4qRve5y4gsQMCf
kucGn90cTo465Yvwg+j+qeGE3yJPOpTE7rPRY0rMdPfKMfFg6+b6Ur+4a/3z2s5i
Y5LH4+0Oe3qzYWT0K+XeJh6Npi4NMN8VyN8uP9m5vjRdjeG5xVglb0d5PHrh1rXz
a9d4iUvyeKZzcHcxmaJQX6cc2Y777rWKOGLpBTiWnFsZFhHnen4Zb708aD24cptb
J9pC/AfMqxXiNI12Fnt+fG6ZnabU/Y7KdKEcQujz9UOpGURclsyP6ItYwJC5vPJq
RZOuTzxJ73KCSiSrnihvAu1tzgQ3+7SHAX2RiF4m8YkVg6dKUkL5p04ZO636UF2Y
x6r2GyDUDj58JbKoFfS23GnCsyozM1QvzYTLIfpf44tVuqH4OUnx9EYsa/uHaRtW
OBYaNN5cgiZ5FZd6VSupUyKLgh1dHH8nmOK8TTnYhMpYbIROQJwfl3xnt+jqwJRc
BRBh16OEpiFCaTr0Ym23PvVjnJX6Tof31u5Z9T+I1LbJgGo+1HMGj62GyyAk2lFt
bmj3kNyBeLFnHCJzpN/XCPULkXjxr6kcJ5Rc35gKGJXaPizv3Pk00pqhtq4twigO
uD1aP2n0zJX1gFpyZ+1Z3y9RmPPtWCoEpIVBH1S6Ui22kAz6P7kmEMdXNSyI5iUY
1pvZ1iunSBFspz5k5GfRJBztY7eQp6I42+61NcDIOVTP5wIlOhPzrc69HHteYx6P
+hpX2XkbcLugfAkU0QmHO5kNcdyAmieMYr+vgD1mmu9GvpQkh/Zzf3OT6TIMgTAJ
J2Xi4Nau6vVB6yuoz6XzSu+Q2S7sVDL39z+/TpsIdGQ2Zp1s+FhV0n7V+yfoKO2U
/uQ7inBsKHftZkwfllCanawXJ10Oz4sf3waZwPCWaER2JcJXgp9c/F67V9GvZEAP
YpytiAD0iC5jTCZ6h6jGFOFvNZG+rwm/XdKfyU4NvCvAgFCVA+SDyPxlrKBeSTtb
QIcTrDAG7anZOSO+mgvwvBLBzg3hIxO5hdvLU+h0/wmF3OZyarjEDSSDM1oqTsDl
C4MwuxuHiBsKjO7oahVed61HoWQbA9eOs00yafb4XAn2oL25s2Ja+HPGdBfXpjTW
zx9lifnBxz83OY+wC38TFNI1mtb2X9uQwIBkB2x9XogQWpA22hlBTXX+AzWQLSQM
Ji/z1tIyf/QwgAiBB7Z/zu3Sz26zQf+QXXRjsywi4+1GHNRsj9Fo0yjEIYtlxzmV
fdsVhfaQB6cQSISpIFVzyy8K+rl1CBJmp/1SHryUc4RD5XiIGv/LeCHiiZzlHBUp
eWjY6adweniVqw9hBN7vgGzawlN9CqbMhS0lQ39o4zJzEXsan/guytc/UUWzNY4w
ZA3f8+8Ufb8ORBJE1hTNE3JUGkCPe5/OTXTitFoSpzlgcddqE8p91UJg54dQm1LP
qCJgOmishgSFmOPld76wBVOUoxHJOcuA3pFJhDcqkjvag8yk9m7k0kIl3bFHnrbf
SfbnvDtS3WfXtu7ZDlBkVO1VwJsw3H26/NFiiW3YZw8NlYjjBee1JGPogkIEyhB6
16mTuD3KGIk5NREW2nVQil6vu5GNXEoa43jTsQXu5GBJewwGqEeoIcxrATMXIDpf
2uqauCLGpNPlDK3PdD/2m9MpyDrQxvi24lQ04FO3nZqCsSpiw2ZEJtiGuT+Lvzlh
pE3mOGfyYaxXnuPrcCDV+ZD/NzOMWtQWt3uqnNn+4hkvBfxh2PcxosfpATkvjASd
Di2DILu9Y3fsOgPu9jVfiIw/+41SR1k7ETOe2hW3VKvDiAaAuZULVvXt1f8as67j
P8eQ4PkC0GKj0yNFL5VALimtsdtYOz8q5vPHblabMS/b7+fH0n9ZdISpNTgaAjsB
iQIWwfeaj6B1eYXpO7FcUDY4VadnitBs+QETXzmnlGPWxUz438ZeHz8UPJhANy1J
zJawPKEXim+mVSMa3fnV6mfaOh0tbRBJtEUs+Xgar+frdEdvBJJnA/Iu1uZtllk/
cnDxcS2Fz9zQiG+d3mWjbnLkW9Q6jVf4YAa75zlfKBg4vnOOmxYQu0A8oSu5Y8W0
bE8janf5ROc25rm+gpPHOoZroNijHvTsxskBRAdj0VvmhXU5AMWFcMI5H2vUPMa2
s354OyMmsnaSk50Jg4DZWnz9jvw2PmVp1TuwaA+3UeX6BHFfEhi/THZUKEITou69
8VTj0+onlcgFJygCo5Om48QqwPOncm3W8yFGcvoUwx0VdJp8LkJwnwPxmgmDFYhD
4UC+dlEUKq2JUBC4lbonRciSlwPj5sz3OzLFVwhVW7dafGSNTNUEWYN1j+X5/48y
d4Dt126Fv2DlkHmquk3RHMDJPdSJWZ7wzhLsnW5DbFTvbISU1sKGm/PmRWXfazVD
NWQKSVUVtVJk53sHY/1WTNXx6ebNhkWNmjFEDto5fkgShprYGOMfz6BPPida0i2D
Wqh3ZW+PQ7/B0nKR5WZ5Psg4SUq+FyuQSCcNOFXnLcktWD9iSQuUmoCi8HfdrWcn
2RaeZudYqQq4id0MyEfUsQCHtw2/YKpacWHBuiInFybOWsgCYGmetOrwoodFFRcZ
Lhuaw5Wyrk4lEjFFMx6qKDBUDbsvtvPQPhxoHZ395GrhHA2l1GHG9DNLzNaAW6tJ
L0CwaxcZOeoKzvvsod4QpiETyOFDJNqi1n8wssFHs9kXBruoNv3Sn6fBqUMi5DXa
UExyhuwN3TqURrvwndP5/6+DPj/ALD5Uc7qe8cZ09i6e18axtXkj350HEAD9bBd5
zItwqFc0wr8WpTMehZBhbRdvUCXX3KMoyX6+pLoGoMomHAXW7gljfvPbbD51mRh9
ehxYAu49n7O80Cts2KDGnCDzXt00VL3m9CSRgDIScAGTEJjqffumBjliT7dIsVko
8XaePxgN7qx3h495BIbNMm4LM2BCaTYOqfe0tsqNXdfUpXMXxta0dBuvVyK7kQKf
N1YU0D0Ple77YZsOLVPvspNvzrSaBrFwD3DWkjdiZTzEhp99IC2RGZvsrTqAGfGc
mi7BX/bzgWwjXgHr5s5A8dJtKgJHN5OccKoJJjU6U+OY1gNYZ5rYegrVL3ISVL17
eYDBwLn55dP/Cyc7ERnb+NGejTReqFbiL57OClvhP4yANexMtwVuxJdKVVnSSQch
YbnAQxkNsxvbmxULOqYEMX4orvl/DUx6RvDGx6mqmKErt9WMKzQxdWrnGf/hRAwp
y8HjqOZk2ISscymYlc36UU3lW/j3au1ryeC7ruKh5B/EpxGbfeMuZVTI4HbyHS5o
m6t4Km52vVCtZsvWogkwvc1WEl75g4fUfRke/kvv0+DQJTYdRitkiI2J2vj6e1Fb
ZwgHR2DgWIC9RAf4pYuzhv85gUytgUvxkkqGbFCgUDw/lAdsdawAp6YShF1aWd1M
nTJfO0QIPHzMEU3SsRmPEnG36BrrXndWR/q8pHPpe7h4r/Gznf+jXp65TtYVpJxb
o0jvwiHFTCqSk4OSUiJqs7SkqXhh3gpwReNGrVh1Klb/WidIc5vpYMAmUZgtF2yU
JDhCZUqjufVs0D2K3e+lDtpDo2kOpryoquXcez5peIucFPHkBquhFTFJSvfYfc8V
LXJPsxNFYYpEI6ku7bh8SHWGOz5lhIOSMbICBhLgeKS2gdzq7Ejn3Y0KhRPW5rsC
SQrAYv+ekgXfHOoxYhOesamZ2mTn++0B858SnPu0sgUb0a2tRppa1BcZkXYtGh0M
KLXuAIvPeFOrgO8u2fZDCLq6hHGq6iDX4LoeSUJyrJ24j/Z7XdFKXOPeABkhOMPj
VrNCf6+dlPN01Zu2yUM8WggMFypMrdVtr9bV9jybCegJ588evdx30smbXHzQQF83
EJDCs+JbYJ+/CtOtrXqRQCPE1kHtSfUeuLmC6YqkZXpUB6GLswZ2a+l4yr4fAZ2h
8L4k/EBK/I9e0IPzPabZScNfwJwCvxODwsPPsJvLA5e6a6+9f7cDPxzAE3eH30lN
9u3JgJOIKIWzEY61NzvVophzu3vvKMuIxH1MhtwHs/aDx0PyJLPsQ2+KscYnW07E
erwx+5K1cQR9TL50BoZt2qr3fCkKl4NbkpK++i0Re2pfUvwDPmpWq4P5VE5ncUrO
62H0VW/vBYpguGDCLAiYTPpDW45mMjwnaX9Vhfn595ousPBcWbUosSrWv3Moi5GQ
gsziuCW3hr6VeW7Vl7iAEJJsiH9SpFXdd2fGJg13a698Bkfef8OHMF520igjZ3UM
FTMMWY8gNux0xYNLMOXoXjbFWx6rV6RwufFO1luLvQMnz9m14hx5zMhw0e8fwDMA
jKqaml7nXnRwuFO/JxRVrXt+z47GggEDCul2CjmPePPVonDLOFdihW62mePwwMHw
dU9TwMdy7obGus4Y4dymAu7GvjCIHGvfY94P6RfptzkjBmGTiBwO0VVmJTrUMv31
PCfjZHyde33xbF0pZgNsTa6JorgwaoG2tqgYW0h/pzKmPR0v0xM3nyWBzWOk/NmB
2ZBXPJ/+TEiETnEu8zv5FjLaQItAsSBOQ2a2yFnyRHqwX1ZKzNZDCpJA9v9On9NN
x3jHtYxyOC9SAtyelAwHdH+jS05MOVQ9pWpEWfIrJRsaYjNuiRqvUgI2MdTw1sRR
DhYonbtNPwNbdGh0pIdg4FLPmVaaV63/+pmA0tN4y5zF0NQH6N9BSDFwrrJ4Es3a
IT0rVqI2LYnXoiPzZIfxDsZ5Njft0oXyAKSZbL408Rn9wPGRK3RcsgtD+eZbD8XO
E0b1QuDN1Xhza2TDMNWuSw8VUdPpHw4zF4vCyBvI0HloWPN/hFH2s/+purIZOgTQ
i3UtA+3SXTm9xfjIEl7k76Gmj5bNif5JJWhNb2+35K76ic1f8Il9N9ytCRYGUfGL
w6GJSdm3cyZu1pGNb0zeJmZ0aTnc1fgM2EZowTtUhDk7Rd4zvPg5dphzh1WGdrTQ
l+w0MnMVKmMjNFJPlxKt3EDn8rd4+y+m4GD3+KX6HITzXUp1u3vytj1vbJYriwyj
/eY+KEMVE4PaY2EJk49psuO/hQZugsAXBv2V8qnNIlqdEx7ffRJYr7h/+r8SUqbk
5f4eYrVV/NunL/4uI9nMK3FJodqucEOlxoPgrDHzcGALFALDnDvvSkdF+B6ivXOM
J39rkhnwPajOI67bonD6umoxAZBcEeiwkWbpLR21lDISVYbX+y/ssRWaIdRw41aE
fVuCLyzNY1KCr735ggkjxpG0m28n1RMjUEA2KZ1a4tbks6Kc+SP9+gfiSLiB6miN
3Nm0wj3xo8AEWHOt5SgZ6sp4tnGTtVd7qrN8lGv8tC2MrfeIUtsp5FAydpJBs/CP
E87bqZ7hxrspkcqlmO1/Dv2KntrwRm5u+c2SMW84e0+WmnPb+tNP297bDq9zVm4p
TDojVFEFt+6u7IXK5QtX1Pg43Wvl9QtbYCO2RipxtYxeWe12NZdoP/8BeJuAN0Ta
FA8Rpyg3XtN92eAYlP793lc/7TxgaHhbxr+4Y9ZSahXYeGGYXHAyJmucpy8hzxB+
iCr1Qq77muW83Zj7xhPB/e9Xcw3x0A71F9OIuYij1Max4oZEwBtAdeAaP8kx3CZI
ZV9+UXXEqFl/0vKig1/03zpxyDzTJDmRuFwy8SACXpDYQaG+9EGPU1+9oQa5GRDV
SNY25I91wUSgOPkvGZld2h8MC3hzdfivYGVoEr3qdlvNiXoBQQ71jxAK8l/i0vtt
jEqb/n7qVIwTvxnfzqUBw7gp6NeYRzuWl3WZ3sl4vZ8f2+aacH0qhFsOZkpqDk9d
D48EBSYuYZW2IiAVOUrlZtDadwWQOJ/fV5m87uV9hE5vMY9YBS+sc2hKBmcab4YG
CYu+8XjAzPeCMlFRAd1By6xkK3W+Iu9Aue5XNc02Vq7H6hnGDVhK+hmv0loWc3ID
aPCeVnRT5JJJSEs+2FlotzRZ4r6uTCp4pcuVbySekvF+uaNfDPBnEwK4N2sDYFYv
HkIegd9F7ywY/pzjcugZ8KrgGmV+nGewXKWx9ySycNG1V29yHIrMc0+aTG/K5sJN
a4NK2pFQHpdgeeZ+shBrfFmzfWqndPEKAagGQq0hUjIHhXmL45UBJf0iYtf9jJzY
T5RL4m0st2Z7hv8D3JwX16e5FqHeUVp2vNZAmaBX5leiaO4olS4/sFxoEThitm4X
S/zL/fvEbUECFG0gkgXCbUUkwkaH6um8Qzlt5og0h6BapjzlaZORCVfOVB36FXlD
PYtEVc1+JdLRqUqiLjosR/f6MlXKH77CNQnYSeE87L4HAjogK/RE6xk8zMO1QIHB
d/SJBSNFwT2O8TPfVigk1lFKIQ3rAZkRxqMNmMbjZlXgzYbYvMQdKP/qjX7QpDwc
H58fqDhIJsPO3mO7zMfkXVL7LPbu3Kb9SwUZrj8vKYSXgUskV1q782LSOjtGn58Y
dxpSZhUeprPsRNgvpcldMqRAXIbZbht7TbofXIlctfbQoSK95B2z+QU3unuTib7n
nXBKeHox1HFZZkwRkniI4DQVFMsdfD13sa2PqbmqHiseFkVRWJVPxx1MpwsohSyr
jYqrfDtIR/rmgFM+BJRP7d8kuD9lEQ02Itix4o+c/+FQhUEM7skOCjemS2lk/11Q
IDEbc8x5HQb3D3dVY9krIZKlmQ/XuiwXwmv4AHbeYEeBn41i150q6R7QmO15vVHU
b0kZV+unIlkMi20m2tFN5g4aeLPmsbl6x3AtzfcdPdPuZM1uErSgQdHgUs3HD9+C
Fm1679SxfExJc6TxQsMBGgNwko2VULKoxcYRj3NpLZolG8+r1+h+9R2iAna/Bs6R
klpgObdFW8qV42d2VtpHoCRdgdOi/qXAwqUcUNuqSWHdqkJmu99DWcW23fIQ2itQ
aQTF/o4TnQSysW2iMwxnFWSaIDNJ4kwXJ5IPQP54CPNm6co6/Pc8oG8xL4MGpS9b
Px7kstjtN9lIwaoflaEGv1/tv0Ks/feIiqdZszA/6Omej+0HUt22kTheSDtdeZB9
u05m8O1xujd0aBVEnMFabBxl8H8GPKlqU1Hanft50mm3jW8+23eD7vBK34tx5FL/
K/kKulYwzDgjskjRnaYoGJvMMhP4aYg3FVwuGc5fjcCC7gqBZrH+/aGNdu5cLyE8
AnjgunPpEcQOeVROWYGSKhJK5zNgwdBMocR0d0wR8otK1HxaQh/1GAcoqPExg5C/
ESDcpiJ96mb7HPDKeomni4z+IfzYUDy7G/LNaXri2DQx9+S83m+sZ3TVTWMJnLLh
l/cDq8Hib4YO2FEv/X/x3c48tJ0bRZOiHmE7+yWZax/LyOUvDwJQ/3b5zkEJnKEW
Ow3xtR2pRik5JovdAFUJZxPfJhbewgCI3a+WJXjvfaGz7ov6n6Wy19Hw1x2a4CTi
FVYyaiyBNjxZ2/kKHAz0f9xcYCeTOBjqRvEW7gR7g9A/PyL659W95EUJH4NtF8UL
EjyMtLJmZjLuN9H6o6UFSmLwxdxgzs5SR7GrASSSBg9oyaBpZ74gpXV7GOtP1Hou
9+Wz7+iRU9LVq7NQxYvjcEwWgK2rc17QItsZCSWtlu2p3242G9D63EgxmC7vCdS5
0xHdzfFdRxOpVTlVgOXdwSQHz+MOCDF8XkYKmv3V3CyQS9q0eEDQ41A67mW732UL
Maa3lcrf930YFqNluFNGct7QMfFNugEt7vpLf+sFrNuOVIFDNlFBfCOdyBqGUBYH
U2PSRhkI8rdvSLgKRYCLOPAA2vif1eSOrM8bVVW3TmHciF07dvTffnSS6YqyDA6x
PdeqdEfTQsVwRIqS0tgp/98f1zWDRS3aF0qaNl8fdu/F33eknxKtjZIqdgLok/a/
gPnDfczs948/C7z388zdSKIaV6/VWlCbfiyo0uv3esnLTsOfHBPlBbSDyKXFywZC
C+ciqV4iIDVMV2XN2PflpSfU0jiWjtcBaAJatCy9GNOWEL4LNnw+NdqjUMUWJMeS
lKvVeis4sShr+8CHZjMrjTk8gc2WHHdyyKReajjCwS0uVEnlCeUWNpSv9NgmrIcE
Ub8Z3nqbGfTaWJ/rpR/I+jgqZRO/GKUUSxbVzNS3B4JTUmCi/zAIY8dwygyMrS3k
bIvZS7imh2bsaJ5dRkGzoLnYNASlB2Y316zWxfiYwhn+lpCSNkp3K3O+39sKYJU0
fkakPO0eS6J/pRsfkzy667kxRd4LqXzjYhaUbt4cdLXU3JDWQdSzWjvMG53MvpPy
e1OuuQkHGRTQHkABnOrEroUVSmrEq30hHykW9zUnAq+zY8g8iIrs6KnY7jeOujoH
yMqgHMLOBrpc1gimuWTxss3+cfczeUMFlxDng4H67ckhCDUbIysswmzqD16i1jDX
PwIbWGdxJeeyK5TWM24nVQ1LkNXozbmCNoanUwNhpXa9B6KhurWYDdLUK/5gN1gL
wuSA3DhEv+d3vJNqSdpQ1M6Rsgt3UGRt8SI8GnJ/nhbLvxmIrwjMeaogF+r3PQCJ
9Gtiy7ZYfTixzmWHZKaaiGW+ghXMD+/bJ42eGCQKvPhBnZSNNU3fogaxQOyfar4f
F0J8Hd0Ur7XiJkohcFgQqNGIwQKKqLZgYFqA6BZXDDvgM/7LnPlKrs4uMUDJfzK9
0L7MEhjKANBAytYZSNPCLeFQRfo7DUkxuyJn1WBAcO7L3WoVudlcnpPIPQxuGD81
EtR6vAzeThZ+4kNb9FBAF/BzGFCKfrNPlRSqi1hP4KmNafmTEaiOj1nQPpCsrQ/U
Z4vAu9zZfMXbrRu6Zb0jauzaDqa8lNY+Zfvdxgi2UYeirYQh7qTp2+HobnP3M/9S
VQv+GbMYjK4O0i5tUBlGOkHNJIUqp5GBtgVoOC33rn2EcRaegZVvZO5ftK4e4/AM
mcxzia7iZCSwkRo93yeGOg+jv5ioRYP1YaQQK24LI2+0kz6cv9conbddAVASSP+g
q1A5H+qFz2hMZGqWKvowNxdqL+T7RMyL5qRNCtPzy/Ul1spTUuBVeZCi+f237Pbc
4iJg0Kt0u4sTKSC88TGgvXqInSX/ECR/I7Bp9cpazohF7Mb/REjD8evY18RM712B
64pqEonRoz9dZW1+/QGxd6DimpMcNpXmleMbTESX13/g293ei1twnDjjdDcrA+L7
WDUA1M4Z/6M3tOZZ+LiTrGDzex5MsYpQ6gQfbKm+oSNHeWslUONB/P+ilZlnqYTw
aaKcsERgBxOKX7FAIgyGFhFZXR/LerT0COvqsDVEIQIZOT/wxY5hPADzYBQho5NV
wELgb2tISQyiUV8MPtH19e/vf4bu0NeqTjGREOPDvz6B7nReSVs4Pe82dUZGdMep
fGL72oz11uiUuvWMmXZtX5XffZ5NB/fpCt78PZ6fJZjtn6Ddpko5Hzbqqn1GzjHa
8IR/WcUfsE6rS17lQTiTvunjcBCF49x6mmmfOviX0NKopkdC2RhulnLkqLH2gpN9
XqQZmksACW0/91ILeD4Ho0v+wnNobIdYX7uTa2+sKXWpYmMVYef/ava+EvAN+urZ
8YHMlQoFI5nwjwBh8OZvKU0low04iO2AskfAJkfoXn3xaISMG+M3p9VbAxoA6/iu
9CYeRrikEXCDvGxHhPL+6EMxralc5AV5X1KXzzQcIdS5HVT4rvSAKwoe9G44/tmA
Q3C0TyvmDSWN6UgC3fW14RKH7H8X0M91t+eIo+LNc4m4RusEy5EP3Zse56sK6cyK
XQBMj/jfcQvz3BaHNQA45YD7WEGSIYqxHvX20b7l4sSdvQ1JfX5E6zJlGvcastGQ
LdNcVJHwuC1M0+ehpnB3vK2biQGXaH4R063cD/7jOkzOURMuSUYtGzdifRuNiOra
4wkb+2OQn5YqB6qSv6hgFVveYnPSA979ld1LydZcOw2WNUTR97nhqlGn3kxvpaDh
iNmQsFe0vNjejT7BwJ2dLYtktuM/UVfvnH3cdaELX2KsQuMdEqCCzDWttTyZO4DM
xLqmB2XUKKlxOmvmmtbF3gNhRpFtW5jZAZR1HtKJ51RFYalmWoYdJnB82/rbWl/x
WiIrLDt8KQk59UHG2x38fhsv9ycRjDI61KbG0eaF7/LBCu951lAiWDE9kk89Gghy
RI5wksTcyc1DRzDkewFDD8aGA2wiZIZbzi1/aI8s4nJqV3Tww/YL9ahW5hY8Eyla
xIPZF9J8g5OgaaqWeytoMhNPJ1SoFRkPlRkB/OBACP/h6aUgKX6PPjiQu+DT3gH1
eCpGDdRjzYXaGl2wzeL6B4vjDWdgshLM/8fpUSJr5OB5q9VVPWjWPLmWhB+DuDZb
PUx8SDmmTJr2Bk3wGmRIau5XgnL7lgcxf16PqYUXIQ9fmgQz/TgVMD3jF16OPRg8
3WqVz1obo7kYQm/p3IGLlGFzjOTSjlk19TPtwURknaKrb9qJLXxc7+GGyhRNRjcX
DSX5jSFsOM6tQmJpz8cbyuxylOGX1OPzViOKE7NCjEurQ0EbzeizGii4NbeTMu9G
MBX8sYk+MSnElZSJOEKmBB6yNM2KeSDfojBYtYoHE8hnag2BgC/T1Rkq4yxxyCPQ
QobHFZGupLbJA1Fc4uSa9VmRbUkwAdGfdCX16VeJPEiflGGAVYzmd2JNVjrDJOTq
omZJFLzclOrxuu/cujyvTo0D2N+sYex0bJBrvO6CatYnmuKeD0B6bQ02HUHm8hik
SyapSC4zTp3wJa3aSsEGD8aCQzJaFDskw96LeTmSPb8PAWel/m7Pq4j/RTcd1v8G
g44NUdpal3As79h3P2zwqw5SyDcFk9EPPUdXVn4DAsiLZoyp1mSDHEjhSHd7WBZN
pn+hjO2kGMfy4v/WbWCpEkkEL6XyEKxhMiikUWc+uKILAfrojDzls5tE4DIyr9aU
UjdEE3Atnn3QijXnBFCK0lt8d0sRK9sgxflEX8ooobOt1WbYMt4ddlO9wJeycekK
SG1oKX4mBWTzeJheRz/e/5sXFgHg74pOKqWxXIIkM8fwH3ND8WNgsEGEpeJLGOqD
2w9FIOvjUkl4QtVCoNMOIapvEffvov2PjPbVYEY/uPVrGJ4NFhvyEYHhspWQj0XS
1eiP5p23TH2AaXuJ0Nob/XqReYp7Ybs1de+yEL5ySGom22ucbdG1bi8nl30BhEe+
HwGluOYa+mOrl08+28Do6v3aPHNQiPWe0gJmUDGlBcsuGmvPe+BGl7HPy7ywkiSy
GBqL2gQGehEB/P/hPvjJXzDZ009JVlNOSs5+/EtGNQgDSbWEWEKxjGU69gLSJko4
s79J9XEuAPfrXYt+xhatvp9Ifqi/Hlq5srto2EQODxpZ5TM0SoONnS3PX0bpHtm5
fBOyfxZ/JYIOagcyzUfjrHZW63o9+5yGA0ih1DNcxwMDp74DMCbHH9Jtg2aZLEZQ
2hV23bXKNH7ZHVfsOiOs83yr4m2291xODR2RrlEi2ae726Q97A//jQRoYVnJHc/O
sNhwm2qBlHBck2eUhSNLhQx15W2MAsjGV02exxvsmfgS0rhoUHoUt0wXjfSMWzu8
84osqyonrns152Aj9YH088ZHvEGtTop0EXkNrG76gWaS7nUwGazKVcOpu0UWOXkG
KF5jjWkPm9Ft2G0tV3YFmYQx0BvoQKFukn0QVSKmh7FmOQO6Xk7o1doy8Qo382tc
UBRAK/v9m2yw3hFAoDqDT7cSXbYkez4FW8qWdzEHYJ20FZf2eCUI18scbr9ahQrI
2DOtygt1Jz1CEYIbIxO4Zfza4p4qNh8OUxsDoCDnpnFdeKR91KigwWikqWicEZp+
i9E0ENGOvX+IStfjp5DBbJNRrncPWqrwNnSJLDaX4tx4l/HdB83it6nS8Djhv8ND
CEhM7ZL1nnmcrRzDZXe3UyMc6Uh+teWW5KWOFWsZt5mxIfinp1hPY5mET9Fml3Js
sZWbNyZPFtPkcxyMoTmx5dOW2/M4tTVlScibRMpUt+9hFDBPDNEGK95d0uj7XfdU
3VK9jYgEYEKihGtOAUeXT0RG7VLnXFF2Xz37p1GhePcyTYZX8BJWRkzaVo258yiZ
gm/FdBoaDFjmkYjR9z6YKD58DwJ6nD53ErbIJ1ejcNr5jZJ5XTytSCASSrWnOAyF
bLxANLSqhwVcIvgr8roFX/F9J00ScKf8OxJRLxNJnHbuJCVsN60OiGkd4dcIqD3c
90HA8W7/MpvSd21F7e4N+Nzbaqx13QmM3bLu3ZEpKVoOBF2p2YhqpLiAplRFNq4A
sM2CTFt0JnYK0w3YR8ShN0uWVjsXuh9gTJelSsFW6/xZlhayxTWzhEnZuKIUPlTr
JxPFxIbGo6xuKGsSUvCS6/zBRH7GxSlOIgc1HXasfa5hbkxQ2ryceUGXG0OywOyK
vJ4cD3vu5E1Iczn8Yqa2e7oZfcHc7BkEhNWN372w7Udn23ruRWA83yNmogp4pOpC
k4w6BQplXt5b8YSf48L8gybZC07+aEr1xpH1pdLBGjXOn+wNW/BxuankuYfe+t41
5CfeRWv9o16HHMfp3mhmHf8tOCGUVW+Ju6U2119rKRSwMrusAFeeR3RxjpUrXfw6
tXtMW+iLiztRLbAnt8fYgXHhpziJfeUDmw/BtRVL2SBab2jiyqDxIzifOBgPWLjD
KGBQU2SmFAWqwz8gz9k+OonNdVR8B3mj9ZR4GuMAfjlxhqxp+iJ6WRjiik4u5cYR
ZR4Xp+ev5mFpW6GiF1eE3VTiB0EkDtg5btza31VhB9kmimS2MpuQJxbwv3DI36vz
LYkqW0lTcKn+nGyaawvWKL9jf8XeNuU3crf7dTmOX9ZETFW/glebPKsKkhf7MyCc
9aTWVB+jIT9+bbD3mEPn/0PKba8DXPFUlOnx6t5oBYLKp8kYyU/awQpKtcbB8l4B
My7PmBR3zO29De25ikU5978ALX/rETIXPrvwDbf/kDEpY48611FqEkmC07uYGKLR
hmXnsWiqE6Bm5Mr9CRA8DakWrkY/6VOMGSFaNyPfhJveMqDDAlVbANQ6FoKL9nYo
Svvm05hZa6OPmujcARnl7aYAX00zx643jFXvmInYVL5ElYtsg15xARI5zSChtm8j
fnmYhOlLsRSxz1Z2Tt1FiUcE23KI2pVibVdUWCaaGkAM50azBnnDW2B2YMMIqsg6
da95JFGNFOZOZQo/PKEFQiTA2Y6XRf5YKEBBVZZCohTAzROEq1m8BkcejJNzZdYn
uhpCY1iyDnY+YnHHrjyXu6eodx2OWBhc+SvFpu6hn1bYbXqJuXgNswKJ42qYJfRL
L0KBzC/QqWXH5y+CVSOSXLjuu38sZL24Kdmz/gAf3Iwj+kNvLziyEyLKM+9F5JXR
2Qb1slloz7TBv4gS+uz0mbkcr59dJqp2oMlM94dirZmpvTyt5bGB8+AeLaFO4pBT
ouM7zbXYRivADZgD3xyf1cK1GRMXzK3PEL9/OAAzZaEiG3P1lRu/rftGYIDZFeKH
1wYRjgThJFRhofLtApP5k7z0IQej2mocD/Wrj/HyzX72gid/BP0Odo1//vEziSxl
haYB5gnFeNFzNM4Roo8z3CiTt1vG6MStlw9F6JWlvrStGnw82c4x3oKZZEW1n4nq
zAe+GZyYVknjng+OvallYop+/ZmEdv1l5J+o+7SNQRLEHC1aZO3TTQ/j/vxIRrtm
e1QQqTDnS6NTwfwc9tdK8+/E0gciuO6AKF/TWSFDso/UYHKlsBY/AP2cJNNBCmbe
w20p9zQwQtynxOHjrm3xT0/dQN5Cm4H5CTO4yDHwC2s0ebGhacpt+2M+CwbApxH6
fpnq7HtS2kP+rAN+zQ3AfC//rS0Nzx2yBK4ZV1CpOIm7TuBz6dOxZIxReo7MKc5h
dQaeQ7kYh/717SKUb6z/4O01Tj68IPf6gwLJfEGR+siOtTlz162urcT/nUcGKWs9
Uk6aIhtpP3DbT1fKUuTwNIRsqAqyJlhWOqKsZnvfnKspRglt5J/xo2BbS45wcz3k
BI6hb2yTezcZyHMU/Od/5MKUujZv78dcPw5mEQh/oMQQHEsPtZFckASFYBhfu7J7
Z2AAJXif9VWhzv0LgdxzF0iMg50IveN6OeL2SOqhzJwLst02IUnZYgu44TojooSP
ofDqqnjROsXOdz4JyG5tIEE8dBLsEEFRb09TcakLx/IWypl+j9b6evZm/GVHViru
hOTCouzyMX1YxZ5x0Ueqb/cL/GSoNk3WcTqMCjg/dmSJ2krjyLIw8P59Koa81Ktn
XdHnX00Z0gYqLmNMqYpMdxWNGFZVbM95xEslBZXyk2rIxD1FLLLM/uZ4om7cxVbL
4Boqc0m9tM4sLATzLaJ/IkOTDCG5METg7qJSlyLQ6iZA68Y2F4vZ/d58AZy6Err9
quVwNIwYqNqvjwAqhEMsdrfv8xrnH4ekKbT9o0vAjyiJcOdiJbhLNKIdNu4gOrgK
qQ41665EbdiBqJC9dYFkUHe1Ygux9XDoK9y2ES1eIsSoT5bNjXpWAwyCSr4tk0pd
wI+Yiw74buR4RmrMS0Z2LL5K5O82ufMJ4EHi8J5Z4cEfF/soymgLWhHRczK9h9IH
Dw9/BSACkprD7JN3Ps2cLQ0CqWIeGYmu7KD+++PA07zH3hIWnod+NmW6o7kG+V5K
j6xt5PJR2ZBkUk6/CP0IaCysr81S3orIHTcxfcMKpbFebcWQol4BfECYtR4knnpa
qXYuISWLiEvK4pvupjtw4XTbfQsaunWFpoxcQbddIBUJ2WziHwjCyBCl5glpx1VZ
d4oJ0mjT4IZkbH5MXKRz8dn8SajGXwMszQvYN5QeLpQ95Vp59BPGRBEP+kevQnSz
V/OU+uqS65BE+KCRJrXQ/4YOXOyDudG+ZGc49krhQQFQ6A5SWQ+RTtrdRTa4mgLO
dfhyyUvcVY8HKK1xIKoiDXXu8tprIehv56cxv8Rw/D+KcO73/RjQ4TeEzQkrx9Z7
NLg6+QreXHzDlrcJlI2zqF/1G0inyxk/FPhOZt8Okhk6rl5SojB5QuJuFqZjtk+8
NmEH4dduVIngDTlvluZ/uedfxhFGQjh/6mUUh3mEZ+dPuSoE7r1Ac4YuMHMksw6Z
h1axcKABC1xO7Kb3gKXBWX8uoG32vfWrusLCXKA9Ocehm88MzllDKhLssfE53EEZ
6IZlCaJu3XjSihV9qrrL5txgiy/xLOkGRc4W9OZBBpiRrDuQqbMMAh5osTTZi2kk
Hji4fNpgj4E/fdXcH1sEKX9kFd9E22V40KPtMG0oksFiuMChv+p6OuIzPxB8iLFR
IezA38vIE4to234bo5apkDB1LQ1oJ4zRtANAsSCyOIR+ZxQ4b0Gg3AWQdUJp+G8L
RivNslzn2Ka3CbaXMZpAenlza5mrGHoykFw0bMkgpMG1NUPSMZLoh6QsId8rhxQo
xkU8VJCqB1Zrk7xyfWuf/A61GRav3pbe2zX/dc3sm2lLKWI82DEU5DL+AlH7b+My
KX32gyTevd/HW7hNgo0zPRxquMr26JWWKu+F+XEW53HsJ626MTrcL+iCd/isk2JY
OkLIYduST4HjhH/tefjSIZZJS3oLjOjg8bRtVISfCbkJSqSKMBC7dNU9VSxwSQgU
uQNYYJkKMnJRku3r5RWo5b2Te7USgGR6o83pwZ6rJ9kJd0luhGqBalYVcuH8NvrK
uF2nytkyHMhB9kVNtzKZaCszqJo715RN0jlFly7QFH5ioF0p62Mj8tZqX8qAic1D
zPHQVh7PJM2eMigB2KQa64sYg4/w4nLgnEO5cel2p7jbgpKKBA4K85FNIYKDVdbO
mgdbat7q97azPN+pcMLT/4R8Cs/0yZcR1+9PBN2L2r4xWGsoC1jn6gcKoLYePGzT
A69tY5RBH0pNtbW21+Ute8P/j9EBHZVHmFvAZ/eXaay2S0dTGhKQuzbqbjgw+xBK
brvBDRNmN1DLWZH8LgLRgRMFwz6y9DXfbOfhPibQQ+9HPBlqIGacKv4maBW9wx1d
uR/QycEdgN2YORoSumwcpN/xdBrZ4cAxNjRU/MY3oB4I2efMOY+sW6vStKXO1xL+
gxdYPEkron82RQB1fJ4+Zk88dWHWtXsTdwICGWne27FVZNGnhz5p1qEG0YXXbvII
0WnJJJz6HugVN/aIhHHpdDnaQA7AhcJlWPS9tKznFLmK1SGd8kNRnWet4X6IXycL
TTyKFbPwdnYeGzvLdgTxpv6/HxQHNYBVWgIPhACFtd+VA5tB5T1ESBTEXX+r7b5I
AgT/H+MN4yuIwokw47QKmgT+HxwNhC5hE57Ef2wmhisNP+l8DYAN7grK/GnJg5UV
a0x1I+vvl3NIVybUBRplj6Vurokv/jHsGSxapEmWFaaNmI8cPi4T4bqqJ8uF+ucU
oUYvmYNdzaDrrwxHwmqgyDB767N9WTh/Po7ogsaDykazHfGkABIso+WX63F8gnBR
fKMPQCua2vzbbtDjGIr+6IJRthH6cy6ptDubR5gXxhT9f6XONRXEusmne9lvAxx/
UpNXct6wT7Bv5c2Ttf+qiSgWbEPkK7AQr9izXj4uUIvHICGpTVDZGDdntgegTYoF
N8LCAkbyeRx1YU6jG8Edi0HIdoVvA6WQqzsqWCbjWzAL5mmaN1iFQWO4Or/wG66A
M0OQzhHCVZdPWxiWDGQXqyjE3Zi2liZU3bt4cCMeztZGYhLXKTwA0bQk94GjPob6
PcGMDGajiOVE4uGqfiPaGUDVaRdiTHxJW65DJkIKV92xsxW3fSMmAEfV4FYykO7/
jmru/u7tp8yVWJfM4IKLcdOkLF+dKRlnmBFQpVaUImrZgSCpXQ3L/W7ZiKCWRc+x
k+jTVAqnTxtXv6Oj9dLrhQIGwitulXDFmWXKjqZIsSdwIfrYdDMbAUl+FqwrPA8G
0x1MBNuaJmizrDfCEkqF466kCXojturbZjLJg/Z1bNEOyNiK1WyEj8zCEUWO+G8U
pDx/z1cZJS9S7Zl6IyJqxhcEGhlfsZwOvVPwHesBaAhMDaS9qYaNfItE8yTiy63y
zDCP57vkYMq9WnULK31R/DkNFxQRuSviWTTTWzO8wmzoLWO5hIS3Tu2PelQ3KDu+
GL1vqXyYlsTuDk1RM92B93ard1FmtTRc83fZ4HXXmECMEsqVb+rHeIgbKeMXq7+8
42dDhE5O0jAt5Z+EqBAoHWGEMgq7C+w6YCdRpfn/Q54S1KuTpZcKi8xvwvZp0Tkq
Bfo4XN6H9pq8u7vq2ZJXeLDwKbWFk7ZS1sq8MCw9T37rElHLez3SkWuiAueESvlD
wI8BUtAoXnnu0Z2tW7RC1Tb33Lba9vBTEXSJq86PayaetPNF+lPjYDeolgJDHRj9
3OpgkzgNBKv2BwqpnN/6lLqlfEX4/t5Zoml8UK9MIVYkAdd0inlCiBJH/w9UnnJn
1YWFrU69/iiYACN5BUrMnNcaG4BxbZdcF7zP9UXijFZ8EdKd6LWfiFIdKLjwvDkW
vKjVN4EKz/dQaoqia4wBxDjPXnOxFYGHhQUHbM4BcjIGPvJemoi0WRf2uNqrh7Xq
FsttWcXB5axwd8NYbPcQ9CWsz/CslO1oNP2q3Z7OP6d6HiSXuORoPUGh/8qNIftR
Cf6e7C3ZeujHVbJscenMwsiD0XV3olvXSd5B9zhrd7tj6Q6Cbm5WMmUQPcyHmQXs
DJUtdBmkM+jCfdBCHY/cu+Tuyj110irUAmO+n4WDYoojp/bacrYJ+TI1T2T3iT/P
tav4Qh1R1fUsaQVUpSRCdQSU8A0VRKKgeBUc2NkmtweKTRXm14r1qxeQOqjxJc7q
kch1eeY7c+/THcbD4xVhV67m0mS1FeMH3v2WM37FZ2r2Hc0pk2PwFRqh53M6y3sh
AF+vcINK+niFHUR5DP66ljmt1P/Im6xJ53tU2dczu6TNiTlFkMX7xhL7a0Zbw5jz
iCwvjehLoPlDO91ADZkxSAojqLBWmop2b/4LSTKVRVWV1glHh9ekVzFohXLKRSU+
UgfRYvAPyqMGH8NiwTavij70teOvCRbJ8wT/s7vuCtbUfWY0bSxLa+QMK5hzDrMB
MMQ8SY86EkS3Hu0WgPR1PbLj/6ttr628isbhD6q9+cOFezpYJOmGlZA20VM2NCvj
MEI57m7aUSh9Dizin9YG7WtQUaHMTPP7f67aClojNbTVlnhnLmPN+QVqG+IOIonQ
7VX4SOmrApRAJk/FO3z2y125mmIkgblvYi+0nbOEGM7tGX4krf8zD5YIKCKHJlXu
CKhZCn0PG0kmRcafnf/B31QwKiTgx3t1hHmqmS90YNE+QjDGUxGackusH/AfiGF0
xjaH6dyibOm/9YUPfcLO0kGLYJOtBB1pd9uPY3e4yPHOLdKaXnfeNAeGcx6KPZPL
XrtZIeEKxwCGPernP47EtfTQCJmEvL5q5glhZLgZtDnkf85n3sPy6cC8Lo8O996B
Z/TnPZcj/dLRa7yOgzix+PV8ZZhxaZ2lSfxYtHEpXYnIlJzto+2RBpys+ftuIzgk
GST7JjtoQdEJW7uHd85YaTB3Us9cuf9SUHF57U8YjkrMwqQTsvoyVbrmBH4+vWZ+
otPleOfc4uq4toPdGEinxu+lvsQvadLKE1lmMuxzblU7I8kSVNF8PSRdB8uPNqtu
U3PoZBcnHaWndo5fI7HiwGP6AHw2y0q8ZltxtOP8KQacB/DRcHbHk5tOuTKjwN83
LZYWnB+O3SRSSFIJrEhmCOu1bvfsugDgNoI50J7vjoFAeYBc7F2ogR1J+eExU9zA
fGInmU29WujPVLd3/Jr7vFXGUX5maTe9TGIBSppOUQ/gJiUOYaZJIwtvetonw0I/
9UjdYtbTHwdPRm+DCAvvSCjVXHIoi2jwIrxH7P4+uM0xuhjhSX/gIYvjxFbuOdyp
KKLDsjWa7xPpqg7bCAjsTGbsbOpA1b+a213Q+gLihg3Eq7ALr6akEy0jP/GPaqaM
MYAXe1hPhzat48Jdnth9sZTeBIb6PY0/wy3GRW9poZQDOMjvIourY7GpghGgZYZk
f3KCOZk+pKPYYQfoVTMVeLLeJO8+E93L9l5YfMYQT8E0eluy/qzzmNNEfcZUACfB
4N6BXXN2z86mw/e2dyCLea5fVhtFy0lye5WQt9Yez54HYwanGhA3MJrwdk9VOhfW
fG+KJsScDPQHRYTBtHOjx/8LsaX64NP37OGC5XKf0/uv7YCVs41SREntmqWwK1OA
77yN4nemdQP976UWhu5c0t8BKY/CnmYIEWjcthtNHWaXdQ/3iKBjl56bbcvbeitI
3oIg8WVDSdueyiG7HX1BtVy8mVVG+eD6o09wiLuxlWhe0hue5epjsXyaFr6HzaLu
jCzX40ppcnKormVqAJrwFRVvrT5f44vuHJ95V2n/Z9DUgnMvX8zY0aHK885Ea9lM
RFcu3g96JGVb4WqIprvcJSsrGhh0az69bKXYYQK2O8Y2dvjuFInD9+N2PnIPnUUI
Slv+Skjp3l8wkMiedNt/Go51mOIWf4+RUG8Xd2EYmvJhVGDsBhbjTOHh5+0AXWI5
rpZI0cPYHdezqH4Rs76cKYhyYjKTp7Yf7kWsmXwftCi+ZD18PZNzvYgQg7kaNOm7
xfzh22ckrsuv/m1N9WJuATimPPT6TLoa34aE2nu3GMbMVMB7kdRvXzie+CPWUZnK
Fh4Gc4F/HNb14eqxB4xjvfbu9/2swuiI5zB8E6krOQJFsV/Wso3tMmIwUInrHxZL
gHnbf23nU4DH63TZQdIThVshXaruj+ufJZRuWxkk1WIy+cdVJl9PLJj0Z4I8Sxg7
+G3QWcUsJTEibJ5Rc9G8KMZyjjmulm8+OKtzUxSiFxgysxh6Ed/iZLMBrLhThw/R
K3AftQz3HyPLMVINO7JgHDvlSL8FKrzDWJvvw59PmQGJ3mBRAOO8+6wWykNItVsT
OenI6nW4zeLJk0vsmGyAyUioBG8KrVY0V9n8pAwlah+98+OPPs67tG2btoPEMwM+
Y1VM00r7h3aN8XGltDpu+hEIJn9dKurh0ah5TwN5thTEVOJsg/hp4JCrwBAnOT0y
fTUzQ8j67LFCCCv9PhabZkK+QYZ/+UmvHbKV6za7XxisoUL98xWEp6PXuil3MupN
iMaBty13p90NeUO0agWVpiywdcnqhrR73HVPzbS6XYYOtUFbsrnXcZqQEyTkWO3a
C1OYQc1xmbn13O1scIFAdQxzxOjhr1tAT/NX/ErpWCyOSWvx4eRGjYC/xm3pMuqB
GuOflo3g1dJO4sAER9BurBVlVdG6zdHhGEfZinGf4awPvrXbw9bw5UN9l78YQhLU
5l1Dmlm6CPaa3w64h87MTe6fuQwZwiQyoQ//OayHX33K5QKYUROz4X2kmnc6hW4a
b3mAeapE1ioU5LQ9A9RnJ/eGMZbZUqaaTdCP/eXCBBTgkgGdod9lMkNF/tOBYmKC
YnuFYSztQhuDQ4NwugTkD9gDm0ENLpeRliAEpmQYpBCPVo+zUGeS56zy1CJ7N2iv
B+8NTmUtQA6IyO1PoZ3D3LmFZzNuTIMlqEbh6Dopc3rz+rPO5Xb4MW3J4btknYLY
MGEjbLHEPDUb6IHUgJgV3s3/DqD263/XsY7yKkq9Rcn0OiyCa3P46jBvJ+YnTUaD
ksoADZOlkHv1SdHLI2MIRWXVIl5xFjcT+dt/voJ+mZGx+f4dUIEtHcPLoBub7+q0
6FjPiKb0/m6aQkFhDuXCOqnW4RXuwMpUmM2MrXl7tbSjVFRHHolV4cBPxz7+4bWF
0kZeby50qVvpf8uJ+xMBddLMLsYoA5+TuBKXECzXQwsKAb5lMHyqqMLn0KLrvsGE
Hs9HAaY/T6ZP6Gvuw0DE59iFxyLY0PQHx8NWkbcd0w015LrzqALOfPJYK7UHWtpS
igNDPIPnu+RkujrJxxBpcDdzj/2bhUCWpylxKLrevFsejZwjUZog20K9g+/NhNSK
UHeG0YyarcWHhL1tD2ktr9XXXIZQ6dLjZIAK34nZaOz2YJDIkCjlt4PeJGrc78Ij
FjH7cowgdPxbV+c6t3FxzmePZKny05DEVGa8MWraNRcDaePMvGbbkn1GbSIhiPDo
b3bsnLFzuaTiz00YpkjpSxVemeDWsRVUD2NARnGa+ZTCbWKQ4kqzKgPyw9iXozZi
26K3fHhtlZ/tDtAyzZErvqE9LTLWyMK9G+WD0kZqI96c4YwwpJdp3HV1SCMeEChk
kjKwWXnRJnlt4NONJ+zKm7Szir529ZaSUD3dMX22ZvHAFR6Cssh5EfOdLwkUDTWU
zK1yXGY7TWs+UgnqwOrThTFKKT8eiCvosibYL+A0MkGE2ZRmHq7E1N1FDsKU0WpU
5qKUeTzh6Luy6pv/tHevGJYW4BqWsa+JdTRRB4aChnwMYqXDoMw/IwyRLV8L7nLk
7s+EmHSDjUcry44x1zwqBN0Ck6LPhF02VMAcSK3xfkrWufvPhVqzJzfDvN6Vtb+t
D8iEG/UnH1fouz3sTFg5Q2KQ5IU17mV5KF/KUTVcywbHburl63c5OAohUSWm0fc9
vKqoWh3JOwKcMYlh2yJN+AnLAE9/MoXlfLvVaZPTaP8pzrn277T9zN6qkQqM52Ww
OoSZkMznnMUUh6b9oPqqAXH18ZmF30E4C5FNLlLM97v3YpMF7imNyXrMRLHtra+R
ASh1D9xl0X+nbdapiVOQNJyOwCWB9wCaTArooYySGZU3sFVlPCdJEzjEaviJLMgF
EmWWWN7rqmgQdlcZ9ZNmzF4e7ML22aqU+X7uWUukXllQ6JAk7pQI3dEWBmoUJLkQ
mFTmzWNLcKe6fjicl9MsYJIYXemgarH0eQ3Opx3NhGUWK0drHksrHVrma1xq2SkE
JoXLHFhbcsZIe1HBLfSxj6Y9cw2cz7yyLaimnqKO1gVW2Mq1nniB91ky0OibOJLG
HqOzooNlmmMfBfybzBwvXrk2EnzkWXyKgS9grxV2Ijqo3vy/z0T8o96Xn0Pa9Lrq
gEFMgT0AnnYPxuFv08vvlcUHrGKc+aJXIM5Hfm4323GNtCywwjeUKNxvFaHeq41C
NoMv2ZEdw/bwKQq0CuNzHwpV9fmM/yHGe8WRGKmKIXul1uqNkQo39gSSePiA5jLs
p/83VH/23p0FbKHjfRVnLUOV0qNX+jH3PAmEx6dSYy8w1fXE+bt6WvbMq4c6mZG0
maiJO8DoeTeKiANiNRMVqHhZTfhEYIgzjcglksVSCr8M3E6JgaLSISMECfZE8APt
iUPcU00xBroZnB1YsSy2v83Izj86mo+tFAKUyVS0lz9EMOwocq7mlVe7IRIXrdIR
uXFIIe3KXHiHipHzXxc2TpJniimvrFmUh6vIvlcwyJdH9j7FWLwZWeQV6+agLzbZ
mSs8o7bn1J/gPsWK5ybxaJPHYbY3CaejvSdcK4Vns5Sgn7GGnWhK8pk8rvD1HL9G
hXk2YEnBT0m8zX1lYq2b1OYJMuJHjwa7RtPWrlb2Ik5y49VLwpybfQDwI6U3B53X
E3lYZZaMENhtFTCLj3JiqRrAYiQva5Po6WjG0avTreILj6nZbIgPcn92rlkFCt2E
5whcieJI6JO94jdAHtBwyWsnYC3EqatF88KWwEihLMgev+fFdzdlKJCEiW+4HIN0
yKQ6Zk2ti2r7URGzxaDzanOGk/sxGC/aPLKPp7KKj72JozM+HatAMLcY0dInKdNv
bSKxVfxY8f3lzCLKw32+dTxdpUsWEFsJtASPvgYtMnQp77fBBSyvuFN3ym4nUB9p
/rGg1W453dVA1WRnYqagGpiPEEtBoSBePvzQL7SITgBQOjloF2egQ7cT8ijIfjb/
+oN/6ukblSaXcjDE3k9a6L8YItjTkvGBFpSyIPe93U+TMvPkJRGOqApZhDexpCCF
lTou0TZz86ODbE3zOMMtlgXA4QFP4lX6t5Pbyh2LPjPnyYHHKV6dhCgKRTOMGBTX
2y1D5ox2km8MvQxhmKr0M/4aQjJCDY/Yc5JNrO27vG/AnhneX6g1LaLh4y8ZHrnh
d1lzV65TBPFZs9kzojvHgiUwi75nSXDVc43nBE/bDb11fQhbdoHn/bnBYbmtUL9/
K1fYrbM8f69oYqDNPAhwl008uADrJmneDt9J+Xo9LjGKuk2KyheJKrzqv7STm8Dz
NMnLqYxz8W4WDM+Nw4k/m/FwT98ynjW/VfvYJ76YDKg9INB53/btBXs20Ae9f8XV
NLzjqKiw34RdiXjQ5wwcLbZMwQw49db4p7Nqk4mSpM9AIDcwHnWGx8aa/82461Is
5ZH663LR5j3uVUv3Ioc5qUL+WIlA5gKaBGjMDno+zm0I7sSsT/2MsK81a0bJy6vU
uQKmlF2AIrx/ysyay6XT4vI4vXWZcqUxcI0oAGqdU5m7H5F6mWfD9q1lVzTw9PZy
RinBR3IpBkFbyToY2xC/kd9x7xUa+jtBnjZVnRLULY02BA7DpAsewdkUtcU+WGjl
DHtXSEAXdFZGeCbNMCL8Dk7JECgBNthi/F7Ut0AsPQrymSq217gfPhIJLn5df0fW
HmqfRjg1m2qEnTkSCgDJTf1Z8n2mP32aS7D21KymRh04frYu3oYY5UGclODo87g3
nb4Nw2O7TgJKwLUdRX29Q+cfOPGWzV/gHZ2SlPXu38uJvkPZanNGYkITJyZQIcZz
1DzrbkwXMgzIyHB3xoAW7OdoO+Cm75a0JhUsSsmwCnWu/13m1Z2ouyfELTJmmNW6
4lfIwonIipy+8Esrq4kiDkdP5jzzM8Zl+fzi3dJvG3cCAySF0j3v79UF+NdMw/Nf
JSrjwcwTxajzDhzt+Vwfz+LWms5WFZob3xVHGtukkLyPMMTWrpETBa/Sax0dBVOx
0TcxMKJxUHrI9NhqSFdouiAghhUozdaoAI1My/IYAr8ATL1xe9SGhVd+1DI4rUkB
yTPVaccWfycjzq//eubjfSgScV6TyFlrRWoauDk+pBZLZlTNjlfqyM0Snd8QfNUf
MrFzb9PMu4r3v+tJWM6Wtm+RSn0WyFBXc0Hyq0nYc8lrHgH6NgrERuthcpWBqs4N
KoS5MurEnxlrivRG8Ufq0k/6torjusMTcp6kYPSO4MOrJWvUVTXsd0MljoQp+kBq
sGejj1MlJvOXjKUCfnqZsgScFfipZ6iObRGrr3pwi14iBJcoM9QJjnubdcO3ZSNW
FWVL5rydB2THVenKgJCN9KSk1TTGAjgt7p67w+TUq6buUA97AiCkOSn7KPZNLQNS
9DZOEZCxRF2VqH7wyRTP2ybAT12iyXwa2VzANHl0CItmfDUrO7Ila7g/03JBkBSG
vRvdJ3xs+RrT1jYSYaNdL/WNjVz/H0ke0n4u5I0kXZ7QlpiwOaIcB8DIXzZzaGsa
EaoRduBcxju3OhZJzyszNNvKzZoWXuzb3q+mqJp8AfxC6CJn7E2LENb0WTAnM3Fr
L2ubaduYmFuuROqo1OtHb7KfeAIr3jjztB1LptrCpEACqpAJPz3IVQKlt4Vu4ojY
piVUUUgZn0boWgNY4Bz4KnkRawnpPICTXtsoSSnB3jPGLU+qvS/iDWEv9u853wnW
/LQUolIa1ruRKcn32izj0jGXyriR9FYDP7cK8KWmlwD7ZJwSb9yFhH/ZxiASDNps
XYAuKIGkY4ZHI/PB+d+ncxO0VF2NfnHGR/vdLFviPi728NTnwDw6SROtilqfeZSo
FhNJfPaFCV1f0u/5AY3KAG0g5FOMoeo79VMkqLTHrqDuEXg1aluIfzKrGI7jjyNu
49C8E5HQoRnjktme8jfdKNHROZ2a/wQFX7n0Mivyjg2hj4vFWbni0/XW8eVhPoYx
+GitOxeyDBSFhBf+10Nrv4p8Bx79B5ugH7F+uQxulHa3Fceo8uf13LkD7rx+7TGj
zcToYDq2WpGdQHC/gEy2z/qCFegbiypbnEicrKVZFWvTCLx/if3w1TAS46edawUa
cgYiuLgYpXO8z/GWnVZTLJXJ2q672GnLgh0cTsD8DPoD4uz3KOpPEvhbM+RdBDh7
L3Uc9vADatofJca47hiCPlcLneRxhjU6gddBPXKJ0YmlBLBqcGRu5EkE9SxCzXGp
C9AguuiH7z04mzTYcsQoQNGz4i2hjj4LMpa/2z/hXg2XsgrqUu5mVSMwvKCHnIrW
xiA3VDkd+vnT0NWbKxrtrVgoQt3Egv+9dVzWcwOjauxXRiAu1kK/cwKFPl/JGdtu
1DhTDelLEUKmXvPrnnjJ7p8jwOstNF0SqZ/6W/TRuzmBchZ5VbhWQYefJuu/oo/G
OdsIK/TTP6UGkv7n9UIlORmS5moqnTGj6tbZ3kzaUvhQc4J6N45v0O7UtJXBMQau
UifV/byeJULVrLPoUF1yjel7ClJvhzRV5GOlcny+qinYdt8kM/6fN4Eknzk7s86M
ZBCQpRUpdObPgzhAafqBY5ZHOU9pILREh8eRxXntvVWGgKokcmD4g67uPVxkWQOd
GSKS7Do3MquhIp0yM+bzYRABGYCqR4ef9mCeVRzl/T22BPtDPqJYyI5ESEYfUnxK
XXniL+/y9G9GrrIOWfACeqWEewcEvvH57FzXfVc8q64mn7Gphdd8P+HdAcvuRJBl
WZ58uXlbDy1Lj/4Gfc1+U993ElrZVfiNe5T1inRyTunHaVnUgmuHfd+m+Q7tNemN
Gr8tdwq38UnKhStkTPxQb3YlePbsRaZnNLPbQLIBx8/0eilqvdBjESaAOSPriKAH
McYYL9ZODpRahNEpVqzLqEl9WhyA0BDaOa0dOHOuHDDSZWpmbqtTBqoiEWMJV5qr
XRNDoOTYrSYt1d6zbhpYAFaLyQbfaqBsTilwpg2sB78t0k41C3tBOmzitBAQkE1v
obGSa26pZ9PwhEZaEmbR1gD3cMh47qlsfCKDPSUOAhxtO/RMKxCRKRvoFy3gIE5H
ES6TySZi7DiHbK5BQqRKyapl2ghO1T+MwrcJ0NXLv+bXaSXnFAaw+1H4bOy6bQgu
79CQVyJGMQ86m2VfCdtGx194VOJ3Ihdm9UfcxKjNHDApJPDEMRa/5t2Dw51VH5qf
yQmEuVM2+19ZtQk3ILnwNC6942Y0PEA5cleGNVKu1pdm7l3wzwoysfEHoa5WWBty
EEksLXm0nane55WEIP20ZHyY2Y8AVKVasGoN52RPTe+gTItbJ21+8SRevLds8mX7
xsJnjbW80qmRK3mSj8je4PB6PqoBJ7SdbU87dvUV0fE9wahdJ03vhI+Mous6dUYk
00acyJ3zTHGepAGaV/pdDS2iRBqXxbPC3B8C5prZQriVVcBd0j6aMv+5d/grTNTW
qkYPoa257t15Nbyr/5RXeAfdz+MXZAJHCortP/E6s78ThYQ1+trqySFa73wY2CPP
gsz4ISsuqplg30jOiSeT5Ls2bb1+rK0Z3mN4iI/ZYxBo3lYB/ejeYLbNDce5KFS1
ggtZFGVIlH6dnyKKLWQp074UoeIHGVfyoXT/ZFwBxPbZr3VSeP7+xay5PaQySpnB
LW9qFa6Ygg6wf8pYJI9iy83UJVqxeuu1oft8GQku2XyV28yIzTpcHXHtn80mOqb5
A4X8fcD6c+BKLjiIHQLmnn35sBSsE9F0kopYiJZJoLEp1cgbvV4dsYcIoR8uksEF
hGpgbROGLPz7SH2jGUymRXIenZiJtJwNt5lw3AVNgQCTbtlej11o2GvsWb9RQKhg
J2et5gHUXlDQ6h8QGy6Kv9xhOkUaDGpxKWpzRLuB8d1c2zC7A2N+k4kwsG9Fc4qM
XZEbdT4fwxywZo3EAY+EgTb9Gt8Lq07hoBmvJGO8UjxtlyglhZ+LQh0IlDXPxIgf
GoNJ+FDNvYMZbgbcPBe3YicfqdMOY1LaveyHzEwl6+QAZUbHv03imJDK0DkdHDSi
qil8+YNX/WcWMLqscHyvUseQzEPQC8/TjmuAQfowsOkubwLdsc9ohbXxwOj11TPm
PKXUIQ9dbZirz01i7VAlp0BTqOLH/H5MchXltuGJIUobFv+vlXHscctasfUfFZLj
kZDfsvVrYhKZ9Fd/8u6XJVVkqmnDbPX6ct0DpDttuhzHZvfsdNExz3R3XBDR0qhU
BmEnSjj2h+IBqQY+bGcMnyj7tokNIZA6CLpQXRA9Fj+Fi5gVb8JjruyZhYjOeARd
SyLgeT27P5I30ebHNB19FmIN9WbqjyoE/mQCQEUUd0Vj8D0taIvHUO6lfcWmTXh0
pxEI8r43FvIFV05QbqW7iQVZ8hLFf1xm0qAhOF7nZKgDotUjRqAGkb6VFhQlLwnw
CtDuxKgPVOjr+67z8wyhFw0DhBOVDeZGpE29JDgD/oAAXMS5H3zIBGkT2ofzCp8m
tTp9OnikSjpqtY7iZYg+LsFKygOB1GLGUMt0RNVZvIKnGSlpUJ0TXeBt1aGZzWSO
0lyoRMnYF6bX3e1zQoxHa6xDmBFWSpCHtWAUfCT6aijJZUDixk3akchgDQDj+/P5
AbCOtqt8iP4H3R6qO7yfFkEqKzO3QvH+sEcofJbHKXt21sGOeWb5v9wtinaOaGd8
TH5Mznkx5QLVtWQzFAub+8NrW4fZ64myeg7qvzyMTKz/4k7XQOaGzAAKNEqI6MEm
/1X8P1pBsEZueIyuxEb+Q8n/8MV3SP+uEDIPIPEpZ1EybNbsErfjak5v5ghsGVNv
5+V9kh6Ptu0EZeHyt/aceNwHnZBAdjAhl0J2wJFtzmotZKbvH8cojjAcwr75bVMT
iLyM0XgQCmYUONKCPvkd5d1abkpLo0tYEmxVjPSoNcLyqQ3vonc6guyUVqRDXcsf
36chJCGmmKax22mEL+OzkFH2tPBSDJboCzWk7rp1vMNSYCw7p3Yab3cPxes4YeaA
Q9k2lqO50MeUMjwvpWM6LUcY0YlZWglfz92Fso3BkVx5B33UPnCGKgBnCeFdvJvr
p+jMhyOTdIzUqMjpfxSHaiGMeeT1YZmKs4CAx5xF3bUAbr4d391/ssI8SxB0eqb0
eHvRmQ1M42Vl7j3+EdGtxm307H/+n9T2hWnzOt8uLNjS+ShIDrfv70jciDItCeId
m6o9fwyzC/EFDV4ES19PC9LuPdyvKs1bF4gpr5rKeR5GPCNabYwsE6WcRCAcG0v4
L1pommuSB4S3izf+H0x+ZJK9sAphWmheYHRyjFsayO+PLJ1u+8hnv9W/4H5w5Pb+
gr0cV774LPKf6CRjydLz0EEc+Ob5dOrXUB3R4xKlIguHGuDI5mnlW+5BWGK7TnBP
4zu09u7Hyt7s8VqOePcHm+3FW4ymLDr+s3pT5FWWIfevdEwUHODXVD98GhBzhvAq
2KAgAgMunrNyXq00FuOAhu2timvXoCoUVRsgneQh3CzUILAqtwdUObaAhZdnlzdY
8TcRIfLgmV4lBJPLzqaxdmRFMD3kXNcN0cHcX0RLewhDrUAfdwYuco5CRAQ0FI+5
YzbxiIHgWioLGdRI4P7zkFOpvjVt7BbgMoWRdHrO08A=
--pragma protect end_data_block
--pragma protect digest_block
ReNgQfI5QBC2i/wkVljG/qDuhhA=
--pragma protect end_digest_block
--pragma protect end_protected
