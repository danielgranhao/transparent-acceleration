-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
Q4MDTmyvxrUmiKIU6YyyfV3mNS5fbTlyLKk8ILUy82e+CIthlrGadLdP8Dgw4vWljZUc1YckPoUv
9jhBJEA8C8s5j28a8ciCtHnZAdibV2fU0LoowL9qZ5TjhiXHvuUboZ58k741B4s0kbhXmNPNHmyW
S4Fdf4w3BXZgX1u62oBLQ/dUTvNPQ5IaSRrFQM0U08ad/nw1VAivPlREakXJm9s0+ARWTfj5e2iV
2VgYNNi7V2FZTSPVYAgmXSgfS4QqwzZcSZ5U0cW707aKWKmyIZ2FySoprjooRJJZwwVocWSH+evs
KF3dflxpXtaxsYLw65+k+JD3BtacyVG5jVo/Hw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5408)
`protect data_block
hgNYiZ17C4QxisScARgZkqhvz/vGd1+wZYShzesysOcMqilyTNdIBv0Wek2iJ4uv/A6PoNFFu4wO
2vdgnoREgTTZ5A0elm2uQG0bc8HX18U6EcuqJ6CeUIhipMxjzDnYKm+3jkBQrKxaUKwPO/3AahRe
csEJTetFNEN5lYq97uLyiaOYuH47m2AV1lsvp4pq3dW5/nRdnS0VRp3/L9yXFuKfy2NUdnizmuJ6
JmZKpFgu8FTF2+gyaR80Znu8DA47RCB1MFNemVxjBAQh2Chn+Oedt5ciBJrPs0Ya8oPt+YzPD8Eb
FXxUsGG1Vp10mSnx79BzE0n95HIYDqE2/GXmpiXVj7sHf9kLFbHI3E7CDlYNG8q6JiY4BQNEn1MX
/9gIPinu9vVqK2JiXXkIk/hH1VxyeRewohTPlbMEpnow6LKC8PmP9D0eYTKksRREBByKAxVf4W2G
pcDXWoTf3sDg29WDACrEaHglk+xldZxPxj5lx7JtWgMb6Z1pLiovyyba2xX+JK44KaxGaZQ9GZSz
23LurWKTD7RkCec57zaDDAzDm8NwNVim0Z2SnHz/33TCPw9Ra650CpB5lwJhkHqna9vU7tHQX7gH
uMAEgV6iiAdEd7Jzeiz0aWjCJRlAxrN6KdJvlnEnpAa+L/sK5ko38Zaulo+GmufSlUIDZbMzAX2Y
Dkh7ZtNmWSOlhtp1ZcY/GPltB60GCc1XZAf2MJydEqZR9RdRwMgpTzaKgmE/N9ZLPZortjkVwmR6
CrSzdpaUIDkG4dmDLO2qkwK4tIDPICZLyb431/i5WwSgVF79NPMjd4bfsdE7xhbX9va4blCF/DVH
2JUMYJXwP/sYfSnRYR8HEOVMRC8vsrK2vncHFkRfVnxpwgZ8PUeMLGxfiU0IPeVAul53SKVRT62q
28N5FmF4V3ZDSm5qUqtjDTmmOFLvwY/IgWFFvBL9Id3vUDC7Oa2vvj24LOxzickQ10EkFzZMyv9P
+1utmZGyrPbjU0Ezrv80eUptOSwmUTnUKyzrjz2cHjcUEqtO5Yqb3NBoW6jBQ+c5ivTpDFcK42Uc
Ltw1G5xbAQvcJAKgvoWJMldN2Gz47uviHdQoCNTpcQ2J7nqr9ut8jap80hLP5VhfMyr94NkOIkGc
N7lXGHEfAalxV1Q1qzGnvB2rQSKajVOMh8oXVGKbs+jhLuPPQkDX9p9is5wF4LmFs3zZmDlc8dWk
lf4iAvDoXA8aPUQ+Y/0PRlIGdWILDDn72AShCW68BIfqkAtKZ4a77PBmk8KaVbFO3vZVrHp9gwWY
LJZiYeddoZZ0rJIABYmZTZceMNdGg+lQcYutxPg+vQCD+2onrJhJoPjExxaCdVyhn9ziavoNbwnh
6ySI092Wmmn4ru3/Er5sekF7p6YprTubLKUsCFYKTGrV2vUj1vH6EY4DpurMdB33rxBF3qaBWW21
aTY7P4hdFTuD3uUBZy8Er08D6EAWaPfhalfsAamRLmg9JKOUSxES3r2oe8h0i6xPXuGB91nPdtSH
WqCjhjsmq19eahhkVWf7zFBbseCRk6jjaN86oWZMhPlESrOQGqodzs53CNzTr9JhOWLdH2HSDPSy
0u42nWWavSmO63kjETUjr2TDMYvPFrFVzOfeZaPSWmSBP+q9v2ILp35e4RJXhPqOg04vwzG3PKns
oVNlDlHygwE4G8MBuGZVRIIBQsaiaMa1FF5PoBKVDjmHEXD4NGlPRGqyQ6uB+XX46rNq1VUsjU7j
J7f9MsA5Zt5/FOBfSnSnsFSUOcR8GBNd8+YSus2XGzn9tf50TJS0LlJUO1hxZGcciu3PRZ+QFnG0
wwp93lNMcWVaDegQLUBuCiyXOij1A81zcpUMkW/YzWC8eF4HBU1rCvdvGzq/TkM5aXdEdKJPfim4
6BvssOXA15XMFiD6jKhe3pO6z3CvnoOqSHA9s7+P/I4Zkt7cm67hgU6cGedLRyYwMLfmvmS/+SMG
F7A1cgWIdvtWrepfv5s9zX1zV530dhd4g4B1I/CLmiNrKbkcfn6EX4dp1AmKc+hXWG0vlEH0v9F+
Ugu8GzDj9u3foPJYR4K4rnk0KqsHaLq8UWcwgSQXNlygP8TS/dJYTbdWV86tGnSqjBHGjd+JjaWw
qW+QipuhmN2GsHm+Hwq0UNdDF1TprTzPZ3qh/BiNanah2O4KR8WKRl4e5Kw1AJHp4rhAQxP1ksd2
EiwYUJ4HQRORup9RDYJPqsYRpRYkwrVoI0Fjpw86n0so9amF0YgyzvV+x9sv0tCuShD7UVo7yt2E
s0IdWE5l0CedWwKO+JMz9tO4/Enr9Y5r6aRPONdmXBL8FsHT5WPyTSVYHNo8nyKQGmlKAOWoLFVX
xvxA3vlBUb3tNcOeoV7bxNrrcpt7YGcDgQBE8eXtTjc1Z0z+a4XxvnKl2afX/kBtI06hcUs0SO8j
Nn0aTgkkCXlTnxteqi4MGhwZWVqo6kSFx2MM/sAi7ICX0h8jPyt1F5SThZmLG0zfjGx8MJQ3NUwi
s/H3zIkcQ/0sVHYeWF53ObFdC8vq81zHcMkxrk8HgNub0t5V8iF/c7JGd0OaGqD8UD9HRofWWqUq
RZIjsgRzYg9PD6qgzYtK8JBHwrJKu5rAlIQVwKnuP6ZirCdD/kgrq2MiEilu//NsssfwdNFsP29w
77nGh4CkNDDnJw2DouEvz40VWtbsbx8kbfU2XD60l+KHTOa9td37riZh/hOcQzQm773mpGalk7Vx
g9LHRguWJeadURDnE5Bvy6s8q81kOQiuWZO3Jyi8Id4MS0/zPLw54xGizGxR5lvrA1NWP1PPkJSh
uLhPoOkt+kPeTGdeAzMZCZ2J5/pRu+il7wgHKtcuMWSwb0VyTXcwrbW8xV8vBFFZ9yk1e5JE8AYl
p/M8uyzuh8BNAn/CDm0QPBwzUlNmMeC6lxIrnul2GhKbB7Q1CBAO13vPz89bT1vOkntiIM4vRf7K
fhLpFOWwBX1YLdgHPGTTAVD6XZCyAGz3tfB3ZZDqolN84wTM5sNGM1Gyr7+0ex9mx+heTq9yZQBT
aAVPFlwsBDyTCD7IezGxiTtDAI/G6AL32NkOy92Gi2+fk05vNdN8aC65cQ506qmgLWU2CBT/loMy
XtaYOWq27maeS731UjnnRrPym4Z8GvvxV7rikfBgi1T+JgmbbPWKo08UIZEFE+KqUxs9k/qPLUTo
jewzxQxHFs5ZVE//dmYps3yzCAWwhcyTA6NmbxO9k36s15Xw5ok4nVTz4VVKRHhKNGRTf9IEcnY2
Xtz1W523sibgJKhXpEmKWTYDHxxXpYl+JSJHHq8CdTw1+Gg2IMBTYeoU1CRAi1sr0x3GR+21vEO+
2A19gZiRhO9quuPEWNaQVuXiuqzf+hgDnYJH1y7OO5JD/KH3Juit5M+62JhUyaz/IXNFKjRoQFR3
4OWQOMjVwSYacqMq2VhO3TbPxTNBWUbHNJsC+riBo0jQbc5za8zkc11NXfgzxp5QFkbk9oxaYhLB
WzLrsj+xpo8c9uoCCQZhZrEooIoIlnQ8xaPysstPuuHn4AFgPhyT24KQ6iZtxJxeCkgOJjpd3JsA
uOdpmeFiKNsANfqnk0bzgvzuEk9VjcorBzyXKeSBFX9L078qzUTICwktmIxVqWF25ByNfiqPp+GT
tjHHKG2dbJ3vgTWQEMRdYyxwemQGsnTPfX5V4D8BOW/9bMBIZn6Fkh42pom4t6JshsNjtulTTfg1
Ij4zq8ry0sHthVzlHoFWq26gh8AYlLJTQPkosApBALIVAkLwaOtQaTi8CrJROQV2bIwzNkNeecgq
ZC+JDm7u/4K5zlZVUCKtK+A0tSqbwBsbaxSVw5NH/CmoP40aMB7uTx/vWEmYZc4KWf/Sgr1SAZwk
DMn8rs36yISH8pyxqbonWCJAHbsbkTTZaqdVLTOoLs3Q/53GDAyCQqjqXSy9KYpSEANxCUqAEtbh
mFBpz3/lX2APx47uiyV77BE8NCqBOUccC/qQl497/mgWrBc5Cl5zrdCJ5jZL+B3yeJdVP9zGRto+
LSZUNqdusvdj9ZRrNvaxS3Dt1dicYUm3jQmk8vqZN4dKxh7e4veA9jlABKYm2xKRVBc5Asd6VjcF
KauAyRrDzxy0x5YvLnMQwY0ILESnZU0+nXavxeicBv9/1Zo63vUosRFbxh0MlMvuIhUN3WZj3vou
gmqP9oWZNg8Ech/synXnP/9VGGTkKa9CnGQDKTVnyOwZ6M8A5g1xHWI7ASKDkN8QupDCdhaGLtwd
paTmYyByf5qaVKZ8aohKoaNW0V5Bv/9unQqEAgGvWOC7NEz1xyBHxTT65cGxxPyt47H2LZQDklOj
u1EoOdS4mdU602Ddy7M6uhIwH2OP4aZrz/UDZtcw3KE5pvXLSwCnF7q9miFX/dM6HUDowECsD4ur
MNe0LRgmn9q3V+7F+vRpNSWM33iNifvlABdcwzpk9K9ZcBOKZ1ZhkKdcVaxeY3I1g63ZEz4JnFB3
z9ryF22Qd74HxKqQGEa8Z5+6TdPEHwhC+NjJM2At/LB2mRwW/hvQVaWbmPoY4ReIQJNmR49rWJSa
CWseiidxp9iBcL8ngKPkN4mHewlRHBQ3NTm1dKD+f5f99N0c6HvnlvjUBN6X3isOqooPIatNKJgS
cSI3UVtyKKE1i9zAZWKaSJL73bYNPx4Y6NGSpjFfhwrCfTi6zW42b5lnUMgGNRItkhApMgq5d7Gd
QJlMQ+vOHwW4tJvhD4fI9r3PTIXI5PeGUl3brZkC15AYtUDVubGRFV0MRhZpkPS4m174DfbK6coC
BL/Z/FDpcr5DNmwRlMQjCsVNpptrh/KbkB9zYbp6xeFM00tb97acom4OFn1kdPdkVfeApe/qnhpC
A5oQP85X6ltGjs6M4fpU//yOxjVzQDdN6JM2A2S1cwPoUMSS8GhnJdvmrPcoDJs7zJIZfJOqZjQb
tWspVwBMjBWzEmo/3zINYS6yv0H/bEQR3rdOCjZm7Kep1qGsbGPvo4qYnrAWZhMMEGkY4bwrx1oM
FrUo+p6ak5nJD2gn3ZC6ViOY7y+5R7NpV/NQvYlQEi6z5PgoCDHP52N8KxxudLZtE6kw6jJNeOCJ
KvS5MeuxvUHHnwNabyj1DzZ8qeWkGE8OJcue4ymFI2WuuFNzN8LCsmyPULthYFjeoUre0lozOPU+
boxS+eHEUXCywe9PJudnChByqb/IOMSQOpGNdKhanhmFZ4wf6l+LF4gp99/VTRWXGqENgQGLfmYo
UDHIc8qUuQliMMSkfks1zPEXKBEDUegPi7bhHYiaQs58J2TqM26ILG8eQFKinnQR3lvTpx0SMxB0
ozu0Sn/DrSsGsl4D3KrSbwdMTDN2Lm0MKLRldH+MH2Z0DxZWtFE9A9Onjrn6GRG5pRCkDA/UHpBl
TX3kgYHwIlEFKQ0u7EDfejU+vBnRpc/BDnfY8gewMkDK9rkkLLQhRv3wRn3wWHajjQeqf+22xOz0
I4UnWmyEnsOb62uymx/t0fetawpY4dXEb6mt1Uflf4IWuphHYjHg5QiMsW85sKftrmzMq83Uzp6n
2oDLcqG4tQt4FX3Lpn/AoCMW+2rqjuEveDbVCMD4+f/dhFJfhLRIDbjWV6oMxzpD8RCgF7w7KTRy
uqNW3Wup03VbZi0g94x9+0BAGPB0E5NnkKWp+F7aCKVLCU1uNsZqex1HVFRQ9cSu5cL5M+MerAY1
qngA/GxJQ8suJRCfaldYS3WFotk4wSA+skdWnVlICZvf+Il2rkDNCqrIgxYkcuZdcPSPCwKWsmy6
TvQt8erXOeFLOFZybWjaFJ7N8qKoL1fh9FBN5K4W+OY0v+ifnG/nPKrRfDkEwfMfv7bLl/+5Uvvs
Gjl+W7XRPmZeEpE0DjSDsmbb9xGcs30ulOxwHui6pt+3Btj+ca1z7Us91gkL065uQrggUHTF3HnN
aKXI0qXKgLGxyrFGg7k6LYgdxESTcRR4kIOq1ESHzDpLTgzpsPI1YHdapPnXssnA0KxTg18TN592
6fyOBLJxJTr3GjupGQcSEKYvvdJGqt6UDplJVMtxNSNWXZB4LbdUDYMvd8/YcbyfoWRdfv1DlHdI
F7Zp70PGQLnVE/MOhx+LZn9y/Nk1dqCzrdv5xa9eudqUcJ6x6j3hXo6rPLHQIPVTg1F2JtLIogVz
fRd/eVELnFbN3SWCrnWVNsdqIac/nb1y814JUzW+5eIobTHDx4VoP/Vu+kPnP1X6+JbePw2D6wdN
S0TkWqCWx56gh83/H8oH7EGT8SmyhY7/su8LfQPCuE4+95ZKeXsxZ7rnTUiBnPPTZrixefQr9B38
Mkky8tBQ6FKJFX0dgWAJGNbzu7P6KrNv1xH4v1rHhWiQQdVMgt5Ug8p8yCkVO+yzEsH5RVJxJJcx
wM7hQ+CHpdWQpdhDpnLAuB8Hx6PBhZMp8u2ZOspMSJe5V2nDWCW/U1XVSu/R1HT5pwfJpP4iigAy
L9TtwOB/ROt3VOhmjofuirvn9lVXFdrDt2yINwqDfNY/MiR8+bPYhhyOrGJbhkHbA6xMm3KeI1GQ
hamVOvs0qpVQ0+HYKN5rS6EeOf1mNGxtLgCgzkm5MrqR86+ARUwOhHzOdczt70utOydgVeNT7kno
iCDQtKqHYU7bAIVUyfkQB1aL1O2uN9JVL5oBuCbvkJBlm+XYhvuDFlStoMeOjPHF4G2kGTB3LiVv
8lR3v5M12sj4/3S0QSggF4s/NFKb2zV/wByRnTXCJV2qiDiprQai5g1v4STZWCEhaTlu+/KoOeFt
wjReJfq/5+wYTkk3YBAM+D2M4iHDdCV91KQivXnPeZ3lY66/E8rOYEgYLsb9kXdSe0cXog7GtIAf
kGy7pa3ejYNWy9KPtyKpkGkUPzuf2skOzkHW6qn0yhUfvICJ1Deb1kIzw2AAV1Zl9lSjfZ96JmyX
nrWDszqvIQgbRnlPUqETCyu7Vw/SgqW1OplcpW3wHXlIuZsoKsV+pgaLAcBNBuhhvfcH3c0eQmDN
Osdh39KlSpIB03tjblVHXgHuoyHuKK1e2JUzpDQe7mgzms45CHXQRhbGHTtDM0xicjA5NkgVzxQE
mhFh3E8G7WePMcbml75sjCq9wm4qAHHOYMLAMIcFPR/v40Qni7iL/E5SvezWtHJWKmBiVjMdMi4w
Cv/jENOXiqPZUt2mlwHdNmIlyGoL3Oi77nNB5lnJUVde97OqTJlYJpKgXJLdo1+smNE=
`protect end_protected
