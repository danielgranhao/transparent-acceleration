// (C) 2001-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, Altera MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
`pragma protect begin_protected
`pragma protect author="Altera"
`pragma protect key_keyowner="VCS"
`pragma protect key_keyname="VCS001"
`pragma protect key_method="VCS003"
`pragma protect encoding=(enctype="uuencode",bytes=200         )
`pragma protect key_block
HFW]FHF^%C^(ZNG(&[9$'0+374BV*KWA)M4GHLW]'@QEHNUL$?HR] 0  
H.T7\&%ZJ@M!P38+.D)*D+5Z:XN^+K!#T)"L+V\4:,6=X!<-H,V _O@  
HSG$F_&-L_IK0QL0?7N!0!99OYMY#.P(UL_P,TSE0Y_&HN7O*QV7A%P  
HW[SI$_E;%HW<9#9:*QT<2$S5.HT8AT'5P.ZD[S/(]'G8A?>(5%0'M@  
HA:6+)&#R&$6R8/RR>"W=-I,2>'W15=N%JW'E?'&GP^:;.:$J4,J- @  
`pragma protect encoding=(enctype="uuencode",bytes=7680        )
`pragma protect data_method="aes128-cbc"
`pragma protect data_block
@PG+37OY]B>=Z7#/3^I$VB@^EM^!F4UGM-)N=@]G5R)  
@@:W#)46J4>CYXD/S<V?YV)>+X8O_(V +#2[=4)HDXIP 
@WFS2!H$#QUZ8T!&[53 Y\U551_/$F] OHZ#>^?E0,0X 
@%B_FP*^/K<'WZW!\S)E_(+*8<ZHQD ADT7HYVA C,J@ 
@*3CPO6O[S+/Z$*P#PJ\IYH*PE.-?)%NTNV!__+JG)WT 
@X6**_/N@67"+,&8OQYT6%H.K=^^ 4JWT8#T+U0H3%-  
@5RA_^1J0Z\76.%GM=J/+@Y@T#H&N:.T2BY(/>:]BO 4 
@\QVM#PX^;/_IAO.YP8R%%N+&3YK)DG+9O@HKW-6PY4H 
@WA4424*"Z0;;)C+/',SSECKHO'(Y679;7RWQ7,__W?D 
@Q4'@$N_Y-'%;NR\=8 ;3RY"FEFPN/E@3Q)=416$3,E8 
@==)8;@=09JM6.*>_>B::Z(2U=<_K.>E*92R:N3Y9=A\ 
@-:[#M69KDI5QOD@Z6/':J;#>N08]OS<R42>IOY#A4<8 
@L"/5 DZ,5O+PK/VM#CV.#6)7GDO=O=/]47BHBQ"UT"D 
@1P@?SN:,.&_0#L:'_8ZNQD:7;OY/1&:U&/M#]/F")/\ 
@QJ82WA!Z+A=W9^QNA8C4<NFU'BV0XQ1_,PK>D6A!.*8 
@?#&AQWY')&&*ZK1>UA'6L?IZ6Y5CGY)MK7&J5-0?+E< 
@<I)%T[$<U%<%LZF,#DOM[)<Q/K[;UM_:-8FRB#Q3+ED 
@Q1H!-K^UFC2H'?831 J@-4Y&*\M^[@0Q,%9&UQI7K"X 
@:4^3NE+_%&%M3%/Q;5;&=/7SE\]XD7,JNZH1!,?1P0P 
@=/@S6TARFKZS,@PNSZ!N+M9*.T(B86]XG0]4T.SC!,H 
@_Y5N5&6Y)UE,7" IG=6H0*P/<K,3D"_=E$W+;.T/O$H 
@[_4**0$M[5(_1Q4_I6DA24(]5BVUJWE9.P8,#]]]P7T 
@^2V..1V\ZPA)L[AZ5X#[5+6MI,'APZOH]A!*-9C8\GD 
@PAJ8J?&D8B/9&V3RK#= *!M?+*&KQZ\Z5),Z"+^?>28 
@39JV Z7US+L.<H^K[6+<R*^/LS,OD<6XCHHXBD7)#N$ 
@9N $9[)9LR"*R%9^B88 WD[<Q9&,'^S%NY7#EL*UYTL 
@5JQ___R2GPH#(U6DIMYH>D1!W\J3>.7E6FG)O*(=BTL 
@KXP2AW(/,2P1=R!N[ (;QT ;G2("P/[5!OUO0&!0$6P 
@5Z6[S#^H1 ),C9];9+EG32_N<Y.<5R1:*_KW+A6XZCT 
@TS5FD/= ,2DQ^ F8,[7VMU\-"2_ODLGYLYS52E3(KF0 
@5>!G-=_^S(:&4L_&*#?TH@S*:L>U@S69$ %^M44GE4< 
@0<_ 6O NQ648E= P_&.70$OV)+Z&&D"I$CE;6W^L_4  
@*DA^KL#@8_HD_!\N,F_WF#K)[-K59Y1<0Z'^X*0KI)0 
@)UIO=-Z00F&@D!UH=W6(*P':"U&Y),R@(S\J#JL0K[\ 
@_[GOR;9.,%\D9>\F=3&8Z-@-^%QFG]1] I0/:5\0C<  
@*9#BT=0ROPHZXA -(8+4J'.:@56S$ <X1:'0O+7U>#< 
@Y9?%Q/%FLNQW7@,%_&>N2;6<NF>P?YE@+@'GP5$0<T( 
@G80PR5C&SS6W3++HLJ/;OI?)2)JJXPC+7,-')/!OIY4 
@1L*'6IHO3*P>):(7,=X2L.ZGN2/I31T<OF=2CK"GS4D 
@1(%GLJHKN-F?/X22OO_1GT; 03> 38NZ3?2@7OLE><T 
@\</Y[AHH/1<4LX#Q7\&8M-+!0\7R4W[ 9JY FRR,1U, 
@<;<WQ83YA_/'U%U1X>_\7S01^JYGA1Z=U66=HW&Z!*0 
@:C9K!N2X.A *6^"],\4_E ENP\IJ8H6CDA1['XU-$^\ 
@(->$[#'UQH,,7G>%?@%=Z[-UHP)=$3V\^#>T@:\,5D\ 
@.U4_;V3]$XM"$8$KC0=PW=F-UMU7"O(%/3=QKM;#H]X 
@=4+M;FIV4.$Y-5M8ELC3%5><B;^^=JA#U%0T-ZXHCQ, 
@=N?M P4'K-R[O-YH3(H68N"CVK)*!D(?E,"68ZA8^U\ 
@^FXPZ4$/E3M_"M[W6H0@@F5HEK;Y'2ZJ&YFGHJHD'0L 
@*?]_8K9E:\/.4Q9U*R4%;=NJD),G4Q/LZLZB]G?FR), 
@27@-,T7O8(C(9X^5"P+F,R/HHU#4VJ0(H@7L<O0MP(8 
@"A=_S(\22!?0S>+4-7&DMBA*I@D%L\-$@X'\2^$ENND 
@_*@ /54?14T=L-$3?ZR(VJ?255#1EG<*;WIP#8A0"5$ 
@;$RH%#;&6#:[OJ;T\EJ$#8>"_/@JSO\<A7 T9!HS-&D 
@LP/4HE5FRYJ@%?6?4O410U1+^J=[U[ZH+) QITP*$JH 
@)>ZHPZK"N,GE/\&+V0^3)D]QJIS[^!W1S$H)]8*!_., 
@H$]0 _G?])7*<32@W?H$R\#J)Q1.RC=4]JI6MS!VB2X 
@W(<A\NO[[U+0]*\>OQ.^\0?1(Z9. 3A *.P;#4&6><X 
@@E&?,J)G!%QD3=2@)+CL1'!\M"3!=6:?H;RN1KV+WA$ 
@?J[YEN.:=I(&UP(!=] -)?XR87B-/-$BSI:"_\^'QB  
@Q=T#KL\*M!"WG5*\]BL3V? "!M,$:'((E]@L-\4E$D< 
@4L+5$X=.#P@@<-?M^>^OSNTF]/#5GZ>Q1\LCQF<$H8  
@73.!]?@K@&-%'4KOFF*ZT;T<6N_VF;,Z[G2JVCL=Y6@ 
@#EXF'90)+T@=42#GU]WJP3B,ALIB2PRO=#=2$GBB1/X 
@GF3'C"=^. \\AYDKZ0%>I;,G\;$&SL?4684R^52LU_@ 
@!IU[4I3-/F@@XA)#9@:.<1!NWU4">]U&5>BD/J>P?+4 
@E=&H@!2?26++EARN_CW7L?O3W539=?:+QGEN#["ON;0 
@6!E+"55;FW<P4#SUYZP(N^)8[-0L,?F.B^CI:V?>,6\ 
@GFTE1RN (HC>\O(WJ]L+"1:T* N[COO);'HJ$A'[SE8 
@[36)*233>2IH77P$M?R%87G-E-*"?FC-H_RA(7ZNC%8 
@NY<9Q$[S57:\6<Q /5VTM[PGP+@C"IH($S6WV. &HM< 
@'VW&KJ*+T,"VXQ)T4,P0*4R"O0N=]Q!5R@EVV53N2=H 
@S5K;FV+09S[GRL?Y3X0]$'\=A*HXRWYX+>R)],/3-,D 
@":7'=4?1BFS-'<IUPQ>KH:/,B-+HB8.02::/- YMP"\ 
@ RMP$Y:Y6<VFK 4020@E*OJ4G:0-.F)YC'2M?Q!+$3D 
@!S.V5&;3J<&).H8OH5@D-&4Y ]BB <RDW!'"./D,R8$ 
@)DYMF;RVS)=_@61I6.\ARIR \I6EG9X:Q4!,,FH.LM@ 
@,:].FV^8Q? J4A$4!7!/E'04^EKO8>0#YXZ\DUQ,6W4 
@BJA\;G6EN[/(IF G+<!L\+1W1BHO9)A4AG"F/6KW)R0 
@A5$3)ZMM0$H$NP&E'/FO G"Z1SI&_9&LGFJ(O6 )\K$ 
@IB:F7-Y*E,+:6M1.:QD[F*?I?P*(1=YRA8P7R:*J/D< 
@AW#4^6,4&$!DA-X<4HZ77<H97?MR_7NW%?(6S,:%YL$ 
@O>V[.1P"4@*!M33YGL1^9.9FD*6+9ON!E5>$MDN)'6< 
@ K7XR@51.1R/LQE Z??6Q *8AJZ!C+&'ZGX2Z3B/==H 
@N(CRZM '1T<,0V+6#\TN=2-$^[.^/2H\'UP?"GS1I:$ 
@[P@A#A4X\X'S#0JXUIS2)[%"_9M?SA$VL)]0WCZWU2@ 
@%W1]A42Z:BA2:"POC%Y^K]Y4O]JZ+095_&<BS5ASYH8 
@AUCS_+TLZI*)KW$X'7%O%8JS*)PZ97&.Z"V$L]!G'B\ 
@9E!46)#K-JD<E>/#)SAA85!?Z:0XZ:TFF&_STG)KY'< 
@6$)(M]8@ZI["O;0_Q^I%M ZD%FW.DT+]K">\I$-/\MT 
@*UH8,$4II\L^U+2]$6,B-%QJYA-6U V6HKP>W.M#,VP 
@"D.)NR,6 >%(L9L0.C)3R+UW-2!HG-J%L7=D.B^[ZA8 
@FIYXO.Z":\A#B*/?8@8.$3R["FK%VF@+#RI,O]@+\UP 
@>M,\D\5G*IZD]U*$+F*5%UA8MI]XJTY>TEY_6"9G',P 
@.)8RW#'XKXD%@?Z[0):B$A V%>]Q96X7XX \W% 3G;@ 
@']R?T[N=?FR0S0[\7F@P5J?*E?=7Y6Z;(#LE#-[#HA  
@_$AL((^7D@K5)&)K>L@OKZ]IN+$-A86T9C55V&DUD(0 
@XY4&\BNTLV%]CM?GDLO\L.BKS?W<"N[;.0L226!W_<( 
@V /F45Z"KP;CIQ7*#B_/"JF//'<7+%"IRSO:O@(A?L\ 
@=)EFD[:T5(S7A7#=M0<=.:Z;I/N5[3Y(!HID:%B S@H 
@<D[+T('Q$_"@R/8)*ACC(;"SK33%C@N)G&G/Y,1M#M( 
@>^FB\1[?\^G-EUVE&.C6?F9("GRT$-J97=DB 618.;8 
@,A"U2B=BW_?H=W&!9\CB?_M->D=J&-2$+-<$_N?U46D 
@6LTPU1X6&[MVKVPZLL/7-U[ Z50V+DVGU9L*NC\0V%$ 
@,0(XXIN>(XLY*IRV7?EQOE!_5B=AD#]$QE08P_F4/Q< 
@=?;2"/04/PK=Z&</0!$A&/#I#5$!&WB*.,7Z&&Y";?T 
@AQ*&+W;[\M)(%+)KGA@.!-B72K$])Q"Y]@K6JAF:'-X 
@;'%9J=*:KR.FS'DLHTQZR1)]BWB9+0J9FZ&5Y8P!V38 
@K(O7*0#+):KT0?*],;]\704G_A _8*R&&E8Z1ML6S&$ 
@(6C&Q$KPVI$UY2,*]:$3;!FYS&S3W@5V6CI8M+&M<+0 
@8]$S[QD2*>$(FJL=!I\.$@ZWL"W3FXS<HIC;TD:QUJX 
@,X=;Z"MLI_E8*<4XN\#?G"R6I+5B^[FL73)2^22N&+< 
@%5"9NG^9R-="YZQD,_>:1U1TZ#,L'NYR4RW''1*MC$L 
@"';_&E0*D?BE?$3O(*&PQT.6F7-@&7<AZ=FKNZ25DV( 
@/OL&WWVX7)FME?4UBQ(0CYBJ3B4Y/)B8QDB_[RIF?W\ 
@NLQ56Z85TGH]-)A+LDX-A]QJ(\X@.ZOW;T-BC>0<: P 
@H$N<5H"8SF,@J62$1E?#1,%PV+X-_!(I8ZECCX%Q(:0 
@.+.[TEF0^P8BMEQA02^HW!@\MD"Y9Q'QTH>KD[PZG74 
@4;?T:]U.1F1@3BK_1KM?7 8\HP\NY^E2-N%+BN2R#%D 
@_KQM!)OIQ>!16'W[.2($=8+7.-N>\W<@G@>,KMT:]L( 
@5]0O0.?!@"P!D*WS6V?WO23MS3-925BEDL0*FJ)E@8, 
@+9^0BGFB[W_N>A93/P'MLX&H^Z130:_)8>9+<?;$<@L 
@A,8HX92O/S 4X >-ZD,89@O$CK&M D>(4I?2-0B=$MD 
@?"CCB$=9J@K"DQ7@L$2A]\OX6Q/)0@)H>_ PT.K:;]4 
@T<]O^ S+&<%3@]<];5P9Q5!1.+]1CY?[U2M+=W^V(CH 
@[KGSJLIT QIIJ>SXBQ/4J;R=+U.KG"FI:QO](V#$+9L 
@Y#(4)9MSL)_>=^*G!!$:*Q&[</1%:<@QT^SI7:MGZQ  
@"B/)\M8X0/\#S'!YV\-!I7[E),(U.'E\7\PS[NO8\!$ 
@9@ZVQ"2+K*-;9\]>K9HUW>\*V)"M:E_X;4\A"7*_+M4 
@RL#"_D7.5<U ?4[N;Z#I!K!9?3]FTE[5(HP/23JD9^@ 
@>?J!V^:>87/!*R75M9U\(3JX>Y_-[1H7N5 5F,>4!9X 
@\)&OG>^1LLN7-WIX*Q'7]-<<4WAY6VT4:!5LCT#ZA1T 
@D?HQR[A.*4^1WH=XPH3H^KHUWC_8([A.256>C=AHM4$ 
@:NPP/T9):GZ"731U5I$+;2Z&1:EC:(?=6(J/:034I%  
@>&-[PSJ[ERRV7:TAT&R>*R1X:R909-,2D-1XBT8;RN8 
@" B=2;W'<RCB0<&4)"?D<^..X<2#Z3B!R3]N"9"K=P, 
@.N^*6<-4V@T];$H0GKW%K!=O*!@R2ZC7P,O>+U0@;+H 
@^M]C&(D\192$OGU'@B=XS2M;%\^H9VG&R#<#8\)9@1$ 
@JQPS0\GR@7B5^+>#F,H3;FZ!*C45\/P!>A1+I%>L.#  
@8"<3X-3EKK+$\O7CLOAWB%;/>!8P>7<=SV;N5*Q.B40 
@MF8"JXT141#O(CSD><3GKR\KTDQ#\H^R;@Q3]\^HH2X 
@W*ZC)+&4U>>545IVJ&RY';(),A2_:.9(DWC9<!]3YQ$ 
@J*,N$!%C5GRB!LMCY[#G2>*@Y<K0AQ.RGJ[H'!D71'0 
@#R8N,&SLLS_WOO2A<TUVFN46!M#%S%F!UE]RAA::#]@ 
@AGSF]6C#?,PS*6YB,[+*O0]S,%,$@=>Q$!'7"S[_%"0 
@\Q#;@XK&'/A[DU^U^49&@B7<-:M%M=20W?^21-Z[NJ$ 
@BT4.]2@#*%M-VOEJRWH@Z# 1Q:S'"RVJ7KC*IHW-2/@ 
@,CWS/;4Y$&PK;XB=\\3NF;\R77P_SR+9OM86(R43P;< 
@^DHZX)*]F8Z7JPV>+X8K!:RO?'.$CR7E<1M*Y2WOML( 
@(A6;.#YLLBR/$BL5><@"S-IQ9MK5(B;VQ0@MLJL#+'( 
@4_[?.,8[%I':2J32A#-%D2"OKK@.")"B(.SSX0=)F[D 
@I[D??),T#B>="TW;S5SBHJFI@N>DUH=(9W97#(^DL', 
@EF_1*#]EFO!DE 5ET5SZ#6$;Y'_[:96]:8]":UJA[14 
@!+2^0_/2VYZ?.Z+"RLPQP9$H2X3[N2(Y \K-D X%JQ\ 
@X-<A/XV#[0!*?=CPY>P33MNL#A!W!X:6]8F3PE.&W?  
@M1\QTU0*,2(\3#M;:_,5/C9+;.T9%B[U P[U$/Z"N'X 
@BE[4'RH6MLVJ-N.!NO?Q'G-H<%,AQ6,WE:<\V"$DT&< 
@@X61R9&!Z&8V&&Z@5'J4U9:%[$7O<C,S94,M%\+WYT( 
@*(P+3KSC7ZKF /:0@'H6K1H_SQVC*]+NZ.:XE+AL$Y4 
@HCY:WWL_$SD#MQ;%B.%"<\%"](#="$(_[D1XP_"RY)0 
@7*2VA)P_K)[;4U-XYSIO!"8]@DTJAQ 7D<')G2$$4?< 
@U"Q+@E%X>D&HX.VUET8IPF&[G6#>I:VOL3VP')OYXW, 
@Z'^1#VVRDQ_=99&M+FM7']I%DJ)#.;]XL8=2HD$"X@( 
@33(@\8]V&=>XFMX^QHBA>=T-.K_9!\4:QFURFO2?:/$ 
@^B!F9"% [@*L1 /'3]U.NZ3LD<]A2Y"1G%EJ,+>T(D$ 
@F=RP7WP$K^T0%H% /:?I1,RTG9K&JMNW7=*M>VAA0B0 
@+@$4-9Y9:=31V,FJ$:_['/Z]C3_-JM\^I+)E[#0:O,, 
@=TXPFOFO*:K75(Z/&DK9"GE6'T@,<C//2TU'=$9=TTT 
@,2>"8.#ACF?!6H>,G;8,RP 5AH8AC%@*I(+G/>F\NLH 
@U\H?GNJDNIV<6UGY(19\^)()#@:N^FC_,YXHY"^L5.  
@G.I5I0U .O_*TC@(7/0"=-J!?@!\U2-<G@YW5D@\#C< 
@<<PM'PA:&H4E7G\1(AI^_U7K"QA#VFHO@]/G&!.EHO8 
@7O%TP-5D6X4]]TH[' ()8]_I7M+=^^Q-$YVIE06G!BD 
@1'8C,W0"%=]Z>UX6)>B.IY+':O3Y%(:W-_RT*G C37( 
@*[$U_JN(,(TWEWP'P,_IIFGWQISHP![>,Q3%T).RZ/< 
@C7R&\+7;IVM(*HJ3X#6/W<,7(9'9D"@%Q#V^!T(N@\( 
@,WH7I40XOHI&KZ*-D@)D0='V+CN!_B*J$+)2&QZWA^T 
@)Z_F)"FNGH-(WF2DN8&A4DE9QQ9_5)-F*.8\IIZ4O=( 
@Y:?$XR<UNW:99KTT\GY).>DRAFL-Q@? XG?S3)8LOTD 
@OOSJK;]K Q& _SB+1Q_# J6SII+I_;A7--).'^V80Q, 
@P,5G$5\V@8'W'.!C;'R6[./+0WKY9O(E-@(3DIU11Y  
@3,=&*GLII.3Q?(4/WYMHGLR20<5>='XLDL>AWS.-UQL 
@K("\/)%FH=FT\6Q^51!&M>3]LFKW6)XO#\<RAH>-=>T 
@_I"[ 5)4E$:7Z$LT'/'V<:KQ(;PTNI;0M-8+H&2V'5$ 
@T]&.ZT1( +(CIS_A:/LNZM DM U3IH3\Y/91 ]"8A.( 
@)1Z"[8/,J45*SE,@ F<\L*P95LWS[%JKK7..KU>4-<( 
@I&IF0UN7!_JL&:Q.^)[^9?M(5VB9Z<<+L;D@(5744<@ 
@TN#9S[)#=>SR 0C!U2O!='54^C-WPLPG,6R_?<CS<D8 
@FWG/,J+E%'9RXR=.P>4\K+0G0.XIRI3V.26"^Z&=R(< 
@-]M48B&--4G$SB'D?!/553O4Z12.$%*\?39MG3?5HP, 
@O9<"R>3#$6))%PM20W$TS=#7(3N^%.4T-H?_*4>'UUP 
@@N[V>AGC[B5D4G^2 ^>0%!F!324*5W4S79U_ICB"\H( 
@#3=E$].XXGD@L (0FA^#J_D*1] MI,^>H%Z WHC^MT8 
@\LY/>,80W2!.#HJ$,R_P,O3+.+MMB.:_U3RV<VD4N<( 
@?V&V+9 B=])"+]_%>"%U0/_GJK8$[=' _6#*2QL*QJ$ 
@E6;?9K-L44F&>RPKIO$IQ=M.CNX9$?$\^K8TUE!E>F@ 
@+C4ZA24PUF,R$T;3#$48+)R?I+KJ7!1M;G_"Q.=-R#$ 
@H([68=XZTN9Y=NG)X-Q8OVS(:1$1Z+]1AV:;E=>$0(< 
@+WQ2"BI_YXC.^<MN\#"+&5\D5O@(^3+_&K!*^^I=[!, 
@Q^7KMK XXH00O2L(R^=6\JCO# L$8";RL\+5!8AWM_\ 
@,O3, 18ZT3MKRG1 VWS4@.R*(Z@^:"% :%P*H(UL3AH 
@7(OCE5YI57/B5^5?N3M,CEFA;E*W:51MMYR;.QB\VHT 
@KQ?R?;1#1@GH?]\D_N@*\_A@MHBU)KG#Y52D_PER!P0 
@M.@8>H$!D'="%:F O>?!#';D!:J3W074 SE6<?3"J#T 
@R.]YQ^2HT;*J/<]%?8!4<_-8$\>TMGD8(RAN90YRCA@ 
@X\.E?D,R01$@Y.P]N;:$%U+*4KGLP3HU",F#U<)L.<T 
@R9(:AO:HQFL6/)A#<A,JB)54<G%$.!ACV6LX76KDG$8 
@OPTF<(+=?:%\26YV[N$ZU2OBT'B2;M<UR$1@;EUJMT$ 
@!CC#CG^TX7N)-''0_FT7;V$6M&V[IP=-G=GGUJQQ4E( 
@3G1EA43WI3V435S"BY+)4 )X(;>:B/U[Y8<\5J2^35P 
@\QE'BKXER]?F&=DMT%LS8\BJ/><3I,<1-GO2<6B94V, 
@C@1=VR/YO31BA#28*@;30S$O,UJ1=5J_-_I'TS-BLJ\ 
@$[A.5CR-<!;<WL*(D"0"0NG=.B!43#HFD67XQ2'>Y70 
@,+ 3=R0MT <SXNO3@E$'79Q/7US_ #9D5PCB!F>*CH$ 
@PG X&)X&!+(+<TQ_OG C*#H</F(@@K:=DH2QP-1>#I0 
@*S;H<D+Y&=0Y+(IPLCG%K0.UF561%US^$;34[?C*XW8 
@G+!BD:T<]0Z>7KE/N\P)'MQYH,WI'()^NSW:,Y*'<[@ 
@^N4[9!PNOO:=QAL[Y)8JC<!_BSL11O'G\\@E<%SYST( 
@F)_5TJ<.U4E%+,N?F-\WO<XMU%Y((U:D3DYY /][T<0 
@[-$[PVV-G\U&\NG$[[T S4&Q).MKZS4+1#Y$\,^VN\, 
@AA=15M'?\DI&4Q7.)2F'BYSVFRCOX*$^Y_37U9+R@>@ 
@^Z!=<1F3N%VL@K1"64&X!AV;.$WK=]MW6S73VDI%MF@ 
@8.F?:LO,;=X92,!:5 H *Y<J;Y/LU0*GEM\"4&:>Y.\ 
@Y&QGNL:S9/'&G63I.Z&Y##:CYSL#+K-\-SV0;;M:?WP 
@.@BAB2Z ]R5BT&R=$+<TJ<)SIP?W\;Q@U66!\A=-'64 
@PI!?&%G,OEG4?*:7ER/OUR#,^S=@*]D02H/UOAU ;.D 
@M%-QQ*2E'*KDP0M63!HIE2RR.M;_!IK&UQSH8CWT0#$ 
@X&H20H%^E8PL,7VF$ C+X4B7R-%9Q/IM$'"GP_9'&;$ 
@8?$-(W>INT+B.E.R FBHR37#)EP=D&F%._V<#]$Q7S< 
@-F[?M!G#H8]_RG/GD6FSW)+D>?$R21R/DG>26U.>,)T 
@@:R-</8HCET?_X<C0)HF<(1V];.%>C&O/%;I"?9RI60 
@%VW(,(H>9+KA _-[(V8IH&@W#.'\26Y7-8B70'+\5S8 
@Y\M,6CFW?I7D4Z+(&UFQBL[1(EVX@#_MJ0^$2</14'P 
@&=5S6K+3SZ;KL8!]Y,ZA=(09:;=&1])[##'RPX5'EZ4 
@:3<?E?LAES(M%!ZSN.-.^ICJ&(AL*^_%V6AUIHT#M;H 
@I_!FP5XMI22R=K,AX=/ I8_\[_DE]FD.]N"\H_=Z(NP 
@#WC:^I_SN&5M0=C#PVFJWF3N9L)_Z$Q+ (:DK,Y [+P 
@TCJ7'GWM((R$/<V/8VR:MDG2?PN;%25)-Y)4),X, @$ 
@QD5EK-V=+2<YTVR+UQ&U;R4W<!21XK9&*= 5%'S6]C4 
@VM9^] JV7GZ3X_OP6S[HYR_F4#H#<Q$PV+H%U)<>PE\ 
0.0URR_[-_#&U8IA.P%ZCS@  
03=@M"2].T]\=%07"1-'Z$P  
`pragma protect end_protected
