-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
Wz2xyf/xKAgy518IlorS0OPBUupzPrvTAVwecJLnCM+jJtWgpQjHjMH6T/0o8hwW
KMrVM/8FAjuwbG0WIOK7x2Sq1NlGA4F/cYytlmi/LsxRhjMqX8J/95wld42m0H6t
NC7YhnWAk2Ql0N0lmSPqxxvlrGokSE4k4ESu0IfFLo4=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 6848)
`protect data_block
61ZdMbjLhHMJ32Pk/2W8hkxcaTy3FbuWRZ5CaogktqWk8aA6TXgDI4f5yFumofPZ
Kdf5tajubDwXNSXlURGmOJWkyYDuG3IYw5Mi2LzTtqSVX36zvRW30VJOnTzzrHQT
DjIrkttd2CKxn7TTtAbqqjmMp3l3gsAHCxD+oQT/s5hQnwB30BKUUri4QBwukTFF
H8CmgGnOPWEcxdc0lWmiJZnnkmLLBf1Oak9geJ5jOWB5fb8AaSNbqiCSfmwbjZf9
RPcykWSpLB+OzsDjUkieToIz+u40mIxRKGCUgHzRxWGahTaHGw+CZ37QK0d/erzq
HOTG4JkO4ltVYb/l7diZiGQ4EARUeBnG4U2OJRHQVGsvHFVZmkXmnk0/m5rp/AZ4
H0yBRs/8Yr5pOmFnMrISe8kq7rY6XoLTQlTL3v9YSm/meaeEwZ+99Qe69o11Lex+
mNEekBrorwHi9UG54TUE1f6k3V8mCElQA2JWWerDedO7OMYi4oU65y4DNZE+zbJS
2KLFqr9txe1WjogkPdP4C/mmf5YWl82xnKe8ECUj6fligMvna6KeWMeuyIKvPNL8
yclI/L3bB3xZACAZpXVa41IbY9ehXCJsBMitOCZ/SWVpjzW8fO0jraEf+bq8RHm0
6AxjsSLPBfL8N2isI8FZQIkJruJqoGGVHdynOqN2/o3Y65/3Usu1d2MmILCv5iid
ahPdSRwP/PLI+VsaXuy602CrUAE5m912gC8AXZDsYIBbyny7zwsTKMTBG1l74/CI
whDaAqpq77j5Ytb5AohHCQ4u3G4eTajFs8nS7Z3lV2BDXfzPeyQu6Uj/+biCCd4r
Nsej3pz5dsT5ZhfM+at8delLpGkIkfBS01Kk/jvx8QTUoUrsIhN5UEaEMYlbK2T0
1r7KdQC/rl5LeQ9IhRjp4CTrbeqCpEtB7uww7rmCIxXVTiGFXi9eGyk7oKuq2OyW
Vb9JQFtyClnAtZKoI9biPpriBunHhcm0ihDFJwmzP5ZN+aKVe9C2Dchwx6Yl+bFH
md2/VefrCvR2JA3Eyl+NWAHDZcmVfqeokfWgfV57pSfH0EsuneeOfYLBS2Tuw/7+
g2woLuOJyY9mw9vfmudkauXnacWC0ypuDSluxDycSqkrnTGxX9J8eyuT3fKwm6y8
/iTPr+nECvraijorFvGTS4uKfS3lfBY+0HmC8DOdo6fi6Zy828wKtJEBn7k7loY8
gU1GzYvztJrcsYSe6YbQBlYI0gY45nqMvMsQPjyGK/pB8DEl7PrD1ayP3t76IEeQ
r2VfqA1QZVhp7/xS/qHCY6FIvG1H8zPVWOtaQg3RDW/EcgxlfEPiVjEuzkpzr22I
PAm49PW6O+Ph2A+UzwYKZYl9vT4GyGmbiTFQMLSH24ZwkajmEKQNjMMwPSarB1x6
laqGcK7PP1X2gR/oGBzwbkZnm87/QQ9bWOmauDOQ349tiUa25vMaDyFfA4Af4WMA
5+BB9QLHjJa6c6+ILCpDgR6RQVEskFplffFrvuf0ErJxvuD9/0OQVcS50ES9NPK5
CHUYUUwTfMTHAzrL2OP6AoaSeB2upRBtmnsag8la/jtGQMo64ig6iS3oJM/mV5jt
W/Zv3lNtIj2mVQUCNFqeea8JC2gd7Yv/Jn9JT2B+qmes8UXt09+XgsPUcpd8CIIG
W9jLWOZPjiWQtRI/COjTM30NAH138effaVWgEWEsDnAS6kFBcfsautkq3SEl5Key
MJ7KdQLZd9R0jNs40TZFaIBG8OfxdSLun/l85mw4IzVYrcsB+yIRWiAUgL9Hr1ky
f2MVYfEh0K0mKghwGczUOdqrBnhQ14gqiyiG8a1aHW2qtMFXX1bnD44nb4V/G65S
TtnsMagH7sKJu33nSfWZFo2p+31rGH5OO3MJ3LY241phN55431kL9spCi677BSXI
oCn1n6cFheySPTK2iyVzhTlWqd/KnJSPEvFoqBqwaRxbcqiTQP02gPms0k3wgdko
1Jvmn5GU5Rs0FbMgW6cPa7N95g/lwupzIiw3zmHGZniXyVQ6nLZEz1BUgGshrIID
X7rLro98X7LT0UrqrBK6pkKcltNjXs3CcBFZdhMXhbIolLWIIVmZAlnf6XcN+JzE
XpLfUSgIHWu51UitoJ5IueeByQ0mANHwcDT3NUwxHD1eG89iD+x5NkqFX008RG5N
75CesHDDT2IynmkbBGbC6WyDdr3K52f3GjbA/WJmjKZHvog63TCss4Rc6tapZq0B
AJcmoD1skr8pf81iUCf4Ou4wfx3mmC+TEW+XTb1HGMaY4CxKZTpVsMFBN5P3lLTt
BqclqC8Bh08KkUQ8ckdVzWTpz8akCPwBdDGRwmSrUIRVu9fSUO+EjtuUu/g12530
urj8OAzWYOqvOO8AIXSivvZJaBdLWOPIsTDFKiUoi7d145zhMpMG3CypV/Gvnh96
flwzOFGCf98P8XIQXkPT0THrJN3PzIHIcWnZ6pObdifOhVbbOGGdVRq+jVTplGSk
gS6XWWur8Fmz7R0GnfJGAVs7IIANoUjpXtN90X+PH5TeR2D8Q/96E+FdksnPF3oH
cN6VrhG13Dg7jEQ8IeFket/vR8kjLl3Vt4fDjAj6mjN+irp6rmJwI2atF7aq83Tl
wZwlMiOIvEuzzTi3mnVISPEWUPYUPnYRE0ydYI7J8eTKPpjXqlM5JEPenopibxqI
584OKVdtgc+1JEuSVtoWh3j8NfMtwvEgY4e9tJSoFta5Eq1RApWyZ+kLxDyxX9gF
UR8CON4OEeB/jwcEg7FHPJV2+sOMrTobMksQPCY3LWwbH2DjmqJ4InMxqU95KZ30
KkYdLCzrIwqegCkz8+GVT9qOL+Kwj7NgaZz4MpOB8BxZxYIQj3WX8KYvn9Z5bGHx
EXX/Tu95r8yJucd0oZdo6hdgGV1NF+gEk9BEz/lVbg96oDWl/p0s9twl8tX6/nLI
asecRVfm++DSzF5E82rilysOGmcSVGIiEv5URyMNJQOGvebKucFSeJUjf7WrCdVF
zMgVNQZgbIA0jJZkAg5sqYjDWO674M1CdUcs/0fvU64uXWa8gkoDedvKIcXahwwO
tJZAKOzys4gP7lGlqBEPxKKbuwO2b6c3HRRUY+3PglV5CJnkB+GT5819dCS2uXmN
GLrjdsnxWSweY6IH5gJrM0Dm9ReOi89133l7ckx7G5wEyeeaud82EHcG9gi8Johv
ncFJgzyyRdYUNan9TrW0SupOeVlSl/otzDIjBXzmuAa2EisreZ+aj8abtgaXVthj
o4KLHMD3+1taGni9PY9wl/va9ClHeMAc9xiTdDq3saAUNT+If6A5jSLb5WdveXeQ
sI9+KqiTMeDS9oCtzhsQI4e2QtxUnIBaMrLnEKvMJ3QYcN3aB1v4It6UiMi2aExO
hhmpClSPHOcJe5KOGwvubx2dORO6w5XeTjs5zMOZMuMdoe71/Dhz/32uaqwVtBL7
BudGfZrQynBM6Vxe/DlIWM6uOfeekfufXy0GlrkLQxHQOpsTD00BTBt0b7Zzl1Bl
ovWufCwjoD4BDwx6f/FevBfkDeyfrF8LrtpR7NuKUmjga6LyR5onRQ6ojXuQrvmB
Ns4jW4sV7+GN7iGs5quQR49Mra8mS5DQfykziYcVn89RmfMCD9W+lDRqSeA4t26m
zo6YdgRRYaURnir1gxYd9uj0xzO4UqdHmCj3haH8l09+25vX9I7z/fabGGCsyH+m
JTbmIKnSCnTOILfDzknoHFOt11j/9N93AK5tmX7bi7PRNlAhyJxz1BajvZ6C11g+
xO/nscsGEYcjzcw3RvDy052plVVXJdnlyl2E+Jvgu/ysLgqWES108yY81zSOL39T
M2EF8ceWqTogd3NXJGlYQW8qmzV+IUKgqT8CJJi2HJYB72tPcRWvOuPb0L+Fx5nY
TnNGGkuxMkZHOs/fJL5qd9H/uR814RcMhyWICO5MaqEldVV4L8NN6KxRckiMb68a
5hbPB8k4yxXUC7TG/7t23L1e/5IWXeu32E1QaHJ75GDio9+N6yc3AwkjRWMzSb7f
y1tEPe6LciBXTW/IcYUXQxQS7KNGe4p0qWPz4NAknJ5CXLfZD85WoW9ulEMLnB1O
7RMUgcYE+03Z6sFKYr2oxl7hg2UKlJWGEZc4g0A4JVFpcwiH/Ie/1Z+y85cVyNqo
BxO3ij25rLtkSt4pbgytoHg/ctVvnB9MTmDFepb6rvDe/pH1gPvllCBhOPwUDPAn
zV9xXVsthBYMHLY3S+rOc6q6Tp1sIDenhoy3lJLoX3INMVO4n36+m5yDXV/D5wTc
FPVH4LNTdOX5jGItnYWRMQkrU3dQ/sYYqIONnaUDfH2IGdqDvxeuj42jNiIEal7p
jWuKjsjmkZkJNu1skSAc5k+dGFnO+IiqGFgFqcT7ia/NJHJamJx8FSNNIn4ENkUs
JlMqkYkWo/ouj1pslhadYg39E7p0W7psepwWEWhdSSUniCCTglFn5WghJrEZG71X
aQ0nUAX9t88HGBasZNgu0D4Ikfqpza5MrmerOKqNKjRR1m6d+caiGdLOUAWs7Rkk
51re/easajEx5bUNCUyUwXhTKOEupm3lpCgS3tEnLmzZrJ2sTGyaDTr7KqLPdHLG
aLuvV3l3WGCyuiurTWsAGIUsN2Lo0JG8pP8mT7KXIIGAuWlzVJf4Gs8AW75JDLmf
Uv4QOKNXfrvFtISaZFg124hXXGMcTGM35FqLH/zt0MRk+kFBa7ifiqm9yxeP30sX
UKJoAAD2LP3mUyikXrWpWZ3joYVwG6HddjL5lBCGI9yLfb++s/zQPZc/zBmJzeTO
Av0WXEiA5X2DM6p9gP2MIikHBFB8IEMNuwcJPBSgptYkr/Sje1xA4MVKU9F31JWJ
w2gJPT2HMg7IauYxlecQdjifMmC540gCQacIoFWEF45PEP+a0lWth1lhIBjc0F/o
tqSM9hfvpZFvm1oAzkm0Tjo3pSFGTDuzre+YroF7qSyoUCOKRDQzvvtaiu0/bYt7
pwSkxXfwRpbtY81lpx9ZCtrxty9ePFHN2jcFsA6vGklltc8wzt/Y7CWtdmPOJRHK
yQeWzCPqMVkLopVHZ8HbIx2bozRZv47ygX2TjLsxvz2YfGdAejQZqfwlfPZ1HN0/
4L7zX+ChetVLopeg1L/jP5q78tpNYhI0bnh7vq3IT1htOJ+zarz4BjcBpQ3JrolN
JLCkK+9KfLQNDvKgIc1AGaP+6xlw0aNoxwL5idIoNkmvLuVLER2xu41xNGH9E9zB
P4drTKldNrnwC+Rvni9K4d8LpGRXxsjIk3i2hNSvDHUqYFUN/kDu1Hj2U5+ygDRB
eyscXJS1kFNUdvxGbLG/xkLxfNMk2X9v5ntou4OOXbHWcqE/NxXJnBRIJlmUIe4W
TSa4cHABKsa+sUWt91x5SUH4u4wkrAv3b+dfK7fGTefm5bBpoij0b+BxBrXcM3gk
fnCHZrmBgeoLN+V90TEnbGJlgcR8qWUUVcnYf6Y0zMO9gtGSlfk8Xx/hjqdI7MFS
PkgEHaDlVkQg27kP66C2LSLF49Gpua9+/ZtEuhJR4ZNVIfFxpLZmgn7dObi7CZMh
Tfaw3iBA3h1mUJ2B++0RzAdpHuZnTq7OMSZmY6e2eJZFhX8TfgdaKgRx2XS/cq7m
YXsP/rWPuiIE/gd3qFZenNruvqpEllKC3XjDVrlRvKNmiI4VjOCZ43XA7jserfTJ
cPRZoPiDxRKEHFJZGjS2KuDr0g7pn9N1hb7lARJq3HTytYIKbf/yEMyrYtAxPEvP
8Ck8T9wlsoh+f8lCid1snzimQmEQ/rJjTFPCRbVXeLaGf1E4U10O2yZ02EBFXIxt
fkXElgwGEQ2RnJ25WRdgZTVxu8r6IxzICpMFycKPUQ8MwCQ0Z6gEUqnjJqNMF4DK
MQSbnbC66z0BJaWJ91Z6Yh9xX2hrrk5CpJxpKPIKmq/Dz86+CW8Jk3iBMrRA91Oz
LVmHzCU7gNv6X5kPhIswQDVDQb34k9fCIWwOmd3+FlUEzM/dqSuXtylTpSrg0Jvb
ZVgQ3StaMEDLulWOgIS5OsLjgIa2SZ09aW15dvm0V87NzSKzLIa72HOmil73n3VS
VJlhRD1XEnGwcfyHo/9peCNuHDG+BlPPuKtZAn9D75prpKOeLw6rlTG2VOPCNn+0
JxwKnrRoQh/gYvPEccowvf4CD6QocSxpX+jRjHoKclbX/PZM7NeJTljZMKfXMij8
MsdsQUk6QrCfAaD/uT7yEsx6KtxGk4svClKQDjRwLn2A39MZQl85/IgLnXAbLiyQ
Ddl2ue9zb0wRpJrwq8KuBDlvP/pXyvPZfu6QwAT82UYMEnwvK1VHw/VwxKpqhBd/
vNKDI7CEhVvgi+1ul8fHBALa7olV4cedGqbXkMQYfVgAiIzvn6ATSjDYrgoh/gWa
tqTQ/ba72C+sIhgQhIauv5sqD3UXKz9tQuLb5bKKUJcBZ0tC+grNPOPONcXjcom3
mp53jXIR5C3r2GlvIAOUzKoGser2w/yHH6o0rw+fCbBdT0V3LxTUf/rCzhUpCkHR
zFd7Hj6fMStZx83WedxythyvQ6/3Qb+zj6TP3lkMvDIFrT5WYiPzUuRG5sOnvbfA
kZczXwxB0WD9MOxZhFbPeirUEGdZzA3yIREtqhNwbPIA97Gs2bhaMkyum5HczRqd
m72jQinwZV550ZcE/SFv20b9qGU2dJQ3RMzIjLwmagTNrDjSU2X+OjO9yNE2HP8s
CfMDtRzgJ7kQ1LwWCwCQOT35sYlskmJDNsG7gm14AFSvBlgTymxlkWOEnF6X+k3g
3lokLp1BUQ8bwneQHq12k+3MHNMRPe5iq3KB/FSx37tdQxAdBXKX+zSjoFULNGch
/XzjVjvSVg58BzdCcPMo096cekPcA0wvGddcUYtkkEJcjlo5pVvQzgtQo603sr9T
736CUsmonpbOZdFSXtTsZWo222A0JWHmX8029QKWe2bUnZ2BYKYQOyCQdC7osg4L
x1UY79CF9nbWgO5GaIFWhzbgTWaqMaSaIeESrI10rQg2dHie7/Kb4EgVh+BKf1g6
KULcYHw8p/Ckh2RC3Ez4vJUeX4zccSh/zNk94BKzzU2av0QYAL2myaP0RN6esXnc
CSbGTjDd0jksGzvwyh+IPs38kD5Vrf9ULfVLdA2uvIT5Go4tvc/IuLDh5vdL3p1C
bVLltx+MU/TtYG5YlozYB4LsyfYDn5wUv1b+it+uD2/mSXgXxnHcwzQzeeKdRoYI
T59ZWAK3Is56h4TwNEsMLB0PM8STnAjAcy23dOOx/FhuoJ2P6/uU6bYH0c9JJcS3
ewVedckO0Gm5IkH0946J3zX9OfJ5/qYuEFr/rwSxTwA9Ba20sFvMyd0aZtoxlZEo
Ja6HdDrPn6yctMaYI6EEYfhgqUMYl4l9bxbBRmqkODOrp/uEilzCvn9KGVzvzTBX
AOzSWA6ccWvx9+uXHB1FNose+ykf/zynzgv+DZylPS9GjU3ldHKSdYnpY6xwMXMp
pqZZ51SYEpyMvoYMAzQHePX34U4xhVAQDBKqi0fb4B2ROp+9VBS/xPFdXXog+JXJ
vGScIfCwUcp0aTspYSFymOahtgOBlqmWPkgkcYUgyUaVxTUe26IiXiPjN/RB4KNj
KdU25bRyAucFoMKz33CMDwLbugpNQ2tUuPG0MedwQht6uEvPPsQ9QoPu4vFXAOTx
6IkRIIixMU0lDCb0Z76RrsbGb7spgSOLvit0Sovuw008oiu/qBEPJm2Hgo7YNm1U
kvMjR5iwyt7lSpOtniojwecCgYaAUrM1EJEgwZ1HgRE1pq+shKqkbfF7TrnLvtxR
ptjWLSYPnW+1jBZCUeSIll4gFdadMX44Mv4NpBrnk5E/VOhNMOcveAvYZ9Qvp7Xo
Jt9klIp4+amCZUaDa3sU0tzgKvxoVO+3CQErALkbONIPMFWjcG5tXFYSmKheVDAJ
g19VwFoOd88C9u/7K2PVX6Ap82ciJ4KHv8o9JTftsF+o9XdcjNNlTMb0UFPIfhxK
VP+YQxrjz7ea3GoAnJVIMrQ3CGsiKXddjtAFEQ4Gv9ONO5L/LVl2ytpAJdCBKCyV
jvOJQtmOcJ7EToJgUpz37HgevktgtEUfYEMvAFw7wq8K2NTvJFvS+dTRYKQ7Yp+p
85XSad5ej4KdHsb1jrISdJh3MyAsheoX8os424KDpeZ8cQTtdHU0MfrrxY0zido3
zJupnhk9eFhVzY6wuQRLWwKxUH/0XPMjQEPtQMU2ZPZ3ee3JHpQm80UrRuphS2Cr
dkShmXNpl+JzIlQxRIhefBolmC/T5Itzpnk7uWvYIaKhKzQVo7r7nb82poYNpNA5
GymjiMa+xdKTdPMeK2bHRZ11P2B4puxv97Mbp6KkgR0yFG1+j1B8BX1vtxoFyZ5K
3AfUZQGS+sJfaTZoijWzFZ/u79nZm2LLWyT1SbxL2KTIT+BSLmNPy7xM8Vnq4zb4
q4iOi7v8u66xy72VDOpfSAN04H8S8EtgAFZZy7mufiMBIvVmjS/cfladXaeoxQt+
yE6pgl09mXHD7QMiIl9KH8rFsyn86l/Dn3It7pGypdKNLGqy0vZWL8CTlHVFcEeB
nwogboV5oCuDridaHnz2In7bo0Lk0VvBE7XnBZRDcFdTmoV+y4JUGCswH08EwEZB
mnnGm7VvWyZsXqNQ/n18e0nNQ5eSO0lXa3Zlyoc9AZnuW/PlHGKt9TpBFHNF14q1
YR+CRbKnuMMQOHONSMuHUUaGCnhk0l7j+o41IJkzl2NwFX0byqxUyqsSO1lR0q/L
YiZHTY6KdwcOyfVSikarNja2jXja3ITmz4OUo1T7IaJsc4ff1FBRu6gK8h21U5ua
KWa7qpHvph1WGYXLDEHUQ0TQU/Ki2B4KI9QuwLz24ojZxgetmfhbgfAAnzr9B6x9
nTzPQP1wT0ITOd3JxZdMC22/Ms0XuTiI4soCnwXTDW3x3EdehM+9sL4bfU/chMiV
520aaiC/1xOZ4+kRSlDolUCCqhbBo1gQ6tN6QUJPk1sFuJUj0aiUV8R0lMPYcTiN
ICt9B3dyHBKPhdgoT/JgdbRKf4Nk1ddW1CB6UjfmkKPdH37MYaQjg37tyxOGbwVQ
WSLIW/q8uQfj9F8MVDmvWvF5fplPnhKCgoEOmi4980Q=
`protect end_protected
