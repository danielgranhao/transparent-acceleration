-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
o4cBG1xKqZdq83ZWlMftnkI6f+/LooHzv0nziVFSXvLerwC+fZYBgW/qfXeXRs0B
2+0Uw3W5F7AIjiRG1FvxRxJNIB5ImO2lpUk9WF9K0514twDPLrwOs441mpyVmWlF
pweILz6nZ5Sn8BZmjBpTpAK+2xpy+Gy3bNmDAW8CkioLiJRZlmGQUg==
--pragma protect end_key_block
--pragma protect digest_block
EC2EESYrNDb10rLyDVOZ9kD/nig=
--pragma protect end_digest_block
--pragma protect data_block
eFyi5qrMN3i3rio//hi+u1OlXSDDYEnmH/dXshcUmPh+r+KFyJ2sEDlpM90AtV8B
yg+VQJGf0EEYlpvt3Y5hv5j0OItKH4J4RCH8ExRi9r4a5zDdp4YLlfYJTyreaA0f
Dncsz9bQsN8KWnMv2pqICU5E9CigU7etJiBMlZWaYD63Up0ArMUQgF2h/ydlVqdl
DsLMvsYnHPej1NmXsQ2uQ6KtkvHNI7LAutD302zkEbbcWOutv6v5syxhwRUgTdLJ
9smmk5kBJIjCWBKP5/0kh92WMPBVAiQRt5Y165ttXnvMIpdljW9epyWXvAr+q8rt
VEnHBkBMntYDsup4Qp4n9BpZ9uoCl5PDxrdZ0r0nZ8xy5DpKhm7gGZroll2sryUN
5iNhI3PO/H17yXlkisXUghBdcxLetPNXVKO1eSe1YSzvamsP/s6/+YoCcLYGh9UR
NeLj4ELjt2qMPrkpVQzTKQQ7MJ/E7XWEdseP0+hVjlnGOzAeH8E/PA5flOlgLl9b
0uk4CDr5KYLphZl30aDYWIWUrSvwj5y4u+OM/kG4xSVFNPG55S2v9cGok3nzZu3f
iqr19VsHo8XK0So38lF/7zbtF1hw4UVG0YGZNMUYkCn96aWjH8Knw7DQ1TtaBR6U
eNV3r8Q57nknCtu3cO0HNMDOy4svskfcNVhl/d1QJTsmj/CACspR2J8UBXW314+Y
i1W0cfch6337wFEmLpTAJrIZkJQC/R4yPihMXd3/fG2H/mBJJ1axPd8AxszTiw+n
ebrnac1nq+EBdWV0ImLjcG5tgS0Bs+v1IPXWWXrV9ZrWE1eHzx9qfaWX52gRDtOM
7OU6K01XfNNoT8zchX5oTdyc2Tj9IyNiChms4sJpWdGEgvfC+Etz6vTUNtQqxZvs
5+E3fXRoo9RVS7MzYBcIFzJjTk+PATCYkZPd2NxUh+ZOM8be+GdqbClLc1hGFNW3
IEZxp2UV68OdrMBb1wRlME0ijTPK3UA/7qriz+AeHBTgDgMrba4Npck5O43D4xHq
lVGIWz1aHwPQkmNFCmRIkxMOzOUhpM6q9pQWqd1O3y73gFVyMg9Vj8bni5GqDxsh
eifHd90iGJf9YsFO61xTsmVO8b2jsZEeuSp2CE8+3LLjpwYnTT3zLG51jnYu9T3u
/GYOt6UTeYmk+KugNKDKaQjib577ztqcrz6gJ+NtI22HfoITqiAwHjFFYpBozXiU
bEdW9RDsPGCGdwT44ATV8fclH/IRGFTIYfCCcA7yqAVWpw1qcmTIDKMGQLOAwLTb
LjOdhz/j2EfAPHCVG6Vi0kcylzb2deJKUqohUZt9y6JdYM3wv6ImpsHe2QxXgxR2
VJGG2jRyDBFaralzufan4nz2wDGhlSFqi4Dz/nE0aU3yzJPrBqVoEyMuwqqlj4l5
bwhh/GxP5ecaU+hfgzkDWDtvnqMHNgLQ90Chb8TZJPz2eMavs/YbqeuLwq8lf3f2
cBGyvYKKMFIJ/+reR/8AuVQAtDjfEyXyh4Ji6MjkitxPu+wcA5fsSy3njw4aAn/7
qsyV9OcVA1VgbumvdL1YG1va0em+v4lN/JVo1QevpslXu4NtoJRV0lO9R2PdpgBh
+/o9R/0PinWs4bsy/77SbX6/oAHrPj22CTdMsykiIykM34yQ9FgS7+CL+BU+XKg2
a99Kk5c/Q0SEO2wLnfhUGQ67uMTgi56CALN5kV4MW4RKGidbFXB4RV/osRevifDp
ET/pFjXQZnFtgqVbDX6htiyPgloPUJ/kzRjuTDhzkdD6GlmxltKNRd/pkpgZ/UMN
yPa6/PxI7zvO372JMHzea92RnizAC9KnXNakUDiziqyZ6DGs1TTQNH4Dy3vJ6vXd
8+vTr6RvM6Ha3GYZARgRjl5pN7GA63q2ttKKEeG/Lf+DphuWh9cBJvhK6nKK0fen
UOHivlPEdwnUQY0BjOG3ch6vKPBFFm+5yB33Aj6KEfNSQVir+tpZyIVtdqNX6Ftt
LRFJa1PCHkbajyqBApaRy4RGTK7XmdVYo9/7PoVGwW4+TA+tswELUP1RMF3qmk1d
N7pYLtsLS8MAGe+O23xjwiFXrEkBwSw7mDS/Pke4mpEfN58qYgiYWaCvC9G8B5Pu
8C1Ksf+OL6Ne/cRhXYY2gs8fyfXG8YWkowHNUxYMlYbnvHIcLeS2QJ0jXYIbTTCB
uorIY7JYkwPOq1dNN5ZMM8AhpW9WjUWMDRfkraR89hXcQqhjzZEqiDHJZ80632Jt
u5haQk6PlS2LaUNpUmT2vLbM404huIECzom3w/gHAN7o9molbXqipmn10RISK7sa
ra4w9KNmLtDYoOCdd90Ctdv0/s2sA5zjfQ52pZObQNcpVgYTxpq2kLHUR7IvELsY
6JTz15eq9O42sK3OV7N1axxlRIX8wIetqMziGoGCniluSFhyGkcPYGngWYI8B6rY
E+KI2BdXoqB9/i7CjdV7u+iCTlujz+EsDfzOw3R2v7OyNMvN/oICCxqktxDsrL3J
j/ydaA9uzpYi6nErbE83xixlLw+yXa8n1LY///OUdowLHgmze6r7V3y8x0oepyKE
ymo5rhohXUqWLdUXBxd28nvm3a/AvHWef3ITE+sAiiMyIXyWo2m/mFjaRMTubW/h
kHLbrSa+QOnsMYN2XS3VGvPLQRMVYezyUqgpKEmMBcYDr3LuVNZhhvNR35ek91UM
kThddxINiZhTFatDyjQp6GiwZDVHsBizm6rmjfVkuqF9zShVVtd8NQgbPX+nXbgI
5fCmU+w6y618eWz7yBx1V9ZB7NsMoDGj0R0LxeyvQJhHd3tWMV8ZHG0gmA6boHcm
J5+6UKwSdZvZDRxfiXEu+1yIWStNyZqlun+NNwPwakI9U5zjfHANMAXCgg79EPUe
grODH54+tvTZErDMPOudnwzlDTOCLwxwD9mZWrA5zYbTKeAd5BURfD8PCpHEojP6
B6nosbgejOSLz1d3KApuex9niF1oQUnOUopkMoOqSZssNe/P4ddoRRP0iDJusBc5
gwRsgv8b+VtSYn0yaI2zes8DoIm9e2+syOpbFVd2zJ6c4EnZtftNXqdIqbCiN+K0
IMIPWnaq1+GMQHKJfmP+WLvCopi0cMqt9UmwwStB58zoAECXGOWqg72kHeat+JwU
pWcModMBa75v0zhwk0loChE9lUM52AgRBlHiB294Ui6D+jEkPnR/srp6cHZuAOAC
vPpz2wL4+1sECGd1SXFkhJDXlDU5I7IAnIbN7+eII0BNx396S6z58Opc+rNgy7bx
LErsFXy3RoyRWN8ZvR/3m/fOatt0FSm4qH9qMTXybq3qPxQIPGHFOybTewTcdWiz
j5x7u3YjvPIk173ywuN3BfmeuKhP5UA6VypOOJCqxAOIYOib0llWzrSVBxFoFPzc
AeJF2JyoxnqZLcWa6Idmj7eTMsGWeTANmhjDsIPEzWAJvJiOe/23kcGIAT0fMPCk
/8Biay6XLnSv7+LSmEUCbtef/gW9C6kxRGF+6FrK/0U2nB4ez+u6jX3wEmFewnDJ
XxVmEBRRswcrs2Sb5ujXvDnfNz6uh7KKL2P1532DWpZ7G/9NyhEUv1flw+jvD50x
yuf1MHE1XvIusMcXwqtiFiQzwhPDd6XnUldd/9Da3oG+Z0I2ELqqtoXGvcvwTiBM
XqngpUL+50j8SJ1tZzlS6ClrWln+PVBiVi/87+ss++l+8YQ+n/QTIB50dcLHlHD7
/Wk1SLcDBkVadDhDA70wVhvNvJxIw8Xytv4csKwWs1JNLLX/MlffS4edW2fJ8Kdq
K3hYV1vpT/wu40vlF+2gMDbQJft06jso/KkGg4EqdvVCdlDijH+AhOX4Mpiu1eAf
2AgtIJ18Jog05/p3QpcVrDmSOXnrgmxIJhlmsnELjDAI1IySuG0Jcn9POU2rQ4mx
H788kh7hhk1eBNXEGyl+RajoIGaFbnviUIE4FmEUb8W9p58yQUfbJIXe1SR/uq3D
7eFDKd01FmgW9XrmWfcufWXs/8jYKYQ9NycqKk2uuF5qbKHkfhrWm3gnMfbOOHxP
ffGL8oCq9YVLtlk3PVNGGEuuJNj93jspI7jq32Z6vBLLa5updVeO/PM1CJapoJDy
VsrxFQldqUQvMEmsy69LOyYNz0P78jJY7zsEUS9cXrHP7dAyBcMuYivCzqNiMNHf
2yIusk3v+F/gJerMWEcVPn1nm3/Zbyh5CEBOYkjWCOHyEbiAdIEEiQ1vIfGXp2R4
NY9hniiLIPPzZFMT7NRDuB68xxBqkfMlHTftBXoFLfVUyrUnxPADLCNlKOPi3xLG
RyKR4zMjZ1KK7KAsOCdMhnfrioRbDgm2f8kOM8bge/8y4wss4ZyVUQFFRsda2UNf
EbJLRql3Ybz9Mc0cPIGlbTatVDDAp1XRr1R4dRXcUu+UdSOMIEciFdmf24RFCpgF
2U4M/oreGDy3gaWNN5Sj7IcUucobaReRPz9T7qVCf+T8HqQA/Y6CA2lvI/2OvK+s
XSJnN1eMHRb8ajB0Ij+qqg3g1zMkBz668N466okKHYI+lM/0t0QFzuqdclREVhHm
9xUkRIWXOkQY9n5XZrvROKMlm9bfArfT46cE3ft1/f42JC5BkhyGFZ7YdxxWPGiO
Z2JKivq7RzZYnq4bcAK+bBCTEYvpllj/hUM9zxLJ5Zi4cEFACXRgmzdHy+cEUkxe
L43uUkdVxOyur+Sv7E6w6JhTgORgZSCOl3mhBdR7irSwLAR2nV9hVrScCBwdgfk8
5UlHJgW3zufSr8VxLWbD2kV4mc+guuqyLAFajF//XmBdqnnyfFCBxFP6JadM64nu
hpUazmlVg1qzA1EIE+tSY1l6tUYwXbIMZ8gFR/3NowXytyvvwhExJ+cQ5uXnR3PI
mGDXna4ZrNuhpGvOXtJ1hJbzRdvTfIN0bJqETShKFm7hL27Po9bmifzEHsyLF+Mw
4XQJ9dTN+B7Ayvwd/YK1mAAXA00A0HBr/wxZEuxWY8e2D3YqU3UYV85s18TceIwN
NiWN4AMfGPaa2xYZkFFGv8HsFUwCS62A3KPY6HVqLvQ562bSc35PYdlkudCBmcxG
eH0xCqPiI2O68fI9QHjIaV2ETcvar5U8Kq27yRkuXiRWJ9ayPRUb1xr4Dzthxep3
red3PxxFgwymzP3JHoUw8bjNebTU0W2mcJ0lHTEdO8K3R8c8UToO3A6XfcrOgvJO
B8TVOsIVqCTC3TXZZmad3wIzVx7fRIpzQRPD+oRsmMKBtNa9Iiz+qvzYY8spL05C
ZMx56EKxBTRul8mAVZbYyAMtiaYnfNZ9tncHQzJxYRP6SjX7jcAxE3qfP4nVpo0X
w4fPWrZEZzrG0NlQhSAyjZS1/8/FntZejnjhGWatBoexHFPdGBT/dKb4PwwlPXJ8
Vq4rAt1tji5JT1G6VNk0fuWcT7HRNnzfPYL0Fmk7Mb3jXxNHt8dGu5ydgs6iZhuq
cuanNDL9pI2Fi4rM0RiZ3BdLN5Hgtdtw+WYqrIBLQUZxOH2tIecERvWzCkP671eK
HYUjOaXAIJPgfDzdU1Jjg3GhGYUYAxpQ4FxY/wrtFsC2S5Ovib0C7BUkyiSsZmBL
DCAIYjaJc9ixjT+Hb1Z8h9fT18ehLLyQWH9VHXxDA3SHE+B5D7Q/YdLdhP7AI/VV
IwRMdVB51cP5gwy2zVfAXrMntR7KWAyG7CCiJrfD51xiYHGTCB72xz4p1X7OY+cO
bULVhV43Izlpu/CEiX8OIG+7/JUx1rfbKCsCWl3yFI8KwEiE+3o63nm/y9vSg28a
ZHy/fr50wNMphp/BXJBzyT6dDgBnV4BMksbUeHdgvw7rwLvGIpcDEMncdPYGJ0AF
uMe7thQvan5uPTbMFPVOMdBxuQTEud0s4HqmcIaqnv13Pfek6aHMci9F21+87xSD
nvEbx0uqDZrLDkY+cB1aL1ZiLbwJkbrENeo8uYEiY6Xlg99zp+HLUDyv6uRTykSx
BtjaQMlniVTCcxUMVOfNLfWZkKGnPv5bJbrZVGAi77nDg+641qMnuOQPDN0UvAoB
zRvFLDIZLVzfDazbsnjVTqX2nb/GeQjg939wdCpWiDD5ubgiA3GBqhACGEViOsjW
HozFJA9HX2XOxOgnOIOWJ+G5BJafViAR/jWVq0a3fPYsk+016BldhCmyZ1M+uZs3
cU3xkc8KPWxiR7mnouN6XZ30TzL2yaaBmVASYDzvdQJwBql5hVQaKLPzVw2UlPOK
2M48XUH4Q+bylUDIKJOR/jhQ6pepUm8XanlDwpl4sVfVzbJ0GYOgEs06od97FDqI
otuktl946xLeSTtz5YcCKRqjko5wS5XOr9sVWx+fOZFGWzbDZ2xAfITbzO55Vj8M
lARsyR1J/S2abKFYW891D1JhO1cnq7x6ED2Tk41O3thd3gyv35ITewRevOYAaxe3
MVJtNFIkZutgCbO8+XBDc3Gz6V4LCzfQn5eEUwE1/BZeouwAoT9F3/fWdrkpdLJn
5/bOrB3kfXCXyOHfdlX1KhDYLoxon+YRNcch4w5oS2qjbx6D8j8tT3lOUyjA4o9n
NRpb4pCRNn6Ww1wyl4pcZfGNWfx2stp7yV9kEbfbFxprsxERxMuGI5qDLrAGDvgD
seG76Lik5EgJjXaeGdkgLII1vpk7Swvx7/tBDRSZUXg/YO1RZb7u0CXRE5FWKby5
JnhaVY9jJdTv0FK4yHjx398FkaJfia04hWVUYFGBporegKE4r241Iv3LMU8pe/RW
LRcoq8U+JjgecP2NI86T00NtYi3Y+PPUT5GTCzedQIN8a9qdTitywOlm7uLSNT7r
GpPBZkxcP1GvsrlUqiFRKpSunCnjp/tWI0KOBDRufvVe5PuouktAN/fZAnU5CgR0
PPVNZOBMkYEi+1JKVmErd1bsQLY1FPKX62wPl8NeNKPTHGyEYfYOHVebXn/OGV38
mAOoV2uCXFAsXSU7c+vZR5tMvIfKaiGQpi+JNY3LCleBG6Z9AjUR4knUIdJMD5W6
XT5/BqbvblfZtigPIFoxqHhjrBjdLw6YhTzF9ulwZ99aaDciydg3e0r7SSWFBZ5/
lYw0Yiz3Bhm7nB05Ahlwk5jAn9iiaGnM0ETf0qDJAq3H36w8AOJFxTztKnVHti6r
8DVGcVz75B3vQZntHHUeIXzaljZiZSHHKC25fnawi8qz+ruqIwvp4ZmufGbpJpAH
BpLLBlWaxVtwsfSj8PxgFJePnYQEzGuAuYkLQW0uqmLWmHd+7lB5D/+4fsxUznlV
mj7Jz+5gTEj+ioLd1yBvZ4XI6ECt0oPd94CR+BNPYqwP5Ln8AwTt7m4uH80t3OXR
XGwETwUWD89cX5oiEwP+GQHxp1zOTltlWSM+rMJ3XHGustQTesnKq5xUh8Lvr0IH
328L8IrRPdzkNrnBrakmOEjVvVIP2dlJPpVZb7NkRD0bV+C0kV5Dl2DFHR8Hi4cY
48NTzjXxKcBWMSZ5b/ObzLPmOG9tBdBVY5kSlDZ9v95IE6GKo2Y1TB/d3VI8wSVg
sxoHmVNWF4ZZeC3Kk5WqBdcfMWaMlnuDXf36RhXyuxoa57eEqFZPvjWDM7phLupk
AXse25D0L0PDTE/DdlIDfj3T2PuzL57tMJaEJ5mQW3+je1eIHT3QJLeJWZJ7KwZk
TG+w9QeNi7LIEmf162lCqFdLMw9PhefTbDgrsPupWLZPfRzN+16Hoy0gRtnjPOm+
kK/K5dnlaut7Bczz4qu0qtaL4l9sYBWsHnN9hM6oX5JW0IIEiuCGv8i5LC25XSOZ
b7h291DZgy6V0TE8al7sqVEBXxIHBEqr5koV5m5unYIbnTivt5YGDivTiaaA4eH2
AJjebVKN4wd00YAxfrwCqfDteiySHPovOzZIs5yjlIrira1zTcYKUrCitxmDj03Z
gUfjvmH6RNT1ycD23q5u+YpMvevKxOEypDne8nPqd5NyI3EL38Cw0buPdyAJZysC
bhtXvuHScqqCsqbbYLMEbotBr7WO7SwHFV++x0OvHTM/lwqQYjJ83A8exhdhxUu6
BarzW9jaVqVFl3/xhxzJ8SnWa9DYFsH66Nwm2ILE5yL3XsD8INOLEpwcpu9EIhhn
xVs8ptTuC9+7ZV5AEVL4iRHhxAwnSX6jS60OCg44LTuqNLN0wrJfl7Mf+RKQPf4j
h/sGxej8ifCIg6jQw9HA/ii8aytrwx1A8sVGhC4e7zO7LN9QiS86FUeEfBax1cHX
KqVStgXNJU97hfYwYGaw2uoElP7f9aIJjr3qcHFajOLJexf0TLOudTfFFFPP85/9
DqRPjY3kH9jrT3V6aYxrFCud18jyXDO1nJMJSqf7xzw3GqeH3Zl+6Vj2k32VFi0y
Q47ILeCnXCy7EuM2brVmVDWBrrDkJoX3POllCflwOsgXaSQjH9TCLk7gyR52u6VL
tSsAOhfoIb2GlcLP9wYEoUsVQ/OM9A/UZw+0Uggc8v359LzF5qDH6uKQMgUJqtYG
r1GvsiCtDu6uaiKkrfD3atpNXt7GtB/cwUClIug3qtSb0opYI7CGrztiGpDp9Udd
9qtf/ooyLOEBmeSDbAfukK2oEIfgq/iWhEGEofriSyDSPu8oL1ekqXt3uYy+iKpC
24RLh7rEmzEI0ltj5aD+b7So2iNASCesRFhscLEZAJQnTfgXKDd0Z4YuESoL/G0o
ANmXtju48RX8wE8t+0c6dZvHYrl5ySnGNycJlyatGmPBQyWpVhvPKCrXPDn3Y33E
kqzEZ8/K7NmkUroqFSkhkN0pv+4TWqCmDnOqCsVlZoE/PlqGCbJbKxlRlmfqpJqA
uaElojswxTdrGnTzf1X9HE9vGeuKUewvSAfJhiwadKEaq9m+TZikUuUOoSRgP5Rs
670QvHe/TkO9Ds4FiNzv7gZiw0yyjIrd2bEcy1OVmMQZDekXvJnCNSdtfWecP2wk
cqnLp3nTJ4Ej74zRfaf0tSOLN10qxpE6GZlJXmj+lCfjIUq3yBKTJ5ar134knqt1
SClOVunzkcHA/zB7e5ZJMirDRpbpR3FCzQARcmB2yoimq7U6a6Q8rXT82lwKDEAl
b1/7Ni8nxD3++OJ/lnF1+qENk9vrpsrAwZWDIVQy7tkfelQ9KF0YHa8vcecSwJjT
/dO062YInFpEIdkDgWTX0jQI+ZOeK/CbGYYi9YvL4P1fRaxOzVkiTClmAmyUt490
lvs7WXhe+rOenQ/6aNBc1mM0vKATPitpzimfd6yUk5cL6PW33y1gn8PA4fVYVOX9
KsTWZPZUi3YGi8EHEllmXef2uUuTTYjMtjauuz7bT/5PwGi4x7klIhMv5/N//ulc
VNCTcfAXYZFcg0s+UDV0LaAcVbrxYTjzApHYK/L1Txeidtx6SqUvNk56leD6hXwc
4RV/PbFJtXYfVtOQp/V11WvR3PKHeqru6l5vRL+iRmEZ5M+p11+iJIdPBoETWywO
HEgH41x15jcDEdw+aX6+3znrXBAR7VRj6R3F/JS9ungFSxewDxmUYiMV4JNPjQ/n
iZLG87WuWg6itguYbsOHyJ9AYC/C/kTYIl0ndGBxjGqhLeQVMotak9OgPY3IHVbS
2pxvLHmRdUb7b73yHB81/N6JvgHZ7b9eWEiVm0kSUUdeSPzy/Zo3cKt8JZN/zaqn
OOXbtSa4DQa1CnUD6bFAccKrnnG9S8KVPmqzSAY+f6RRUqbmiwfpZREfjSYoCwyJ
aWYRFh935rBaUx+T8sJ0BQEHlmU4qbOy7y38ZE6GTB1Wm2vtIg/MRciCQv8I3EHs
aWfGVit++0DGLqU7f1seJBom3MzihWckYSridkJfz7iImMrJaeDxRnuGvAL8cxPp
uRxDD9V2JRYBrxs8nml12tvkI+ZTD/owHVZgsBLydsSnkAoXhafQmqoBHn3h3KIP
8V63X1wgdr9KH8dg0gJUVc6jwfl80RX9G+yjPD46zMENwjMyj0iB4dVYAv4PP/Ci
wpFkJCv2IFnXedCZlHAqMAE68xMHko0upshwK1dydr6f1LxP4WEuVXbzK0DiBOuI
jOG/XjodkawY5UazNwUU5/4+k07wscqTIXFKqXrmslJa+gdfRF5rRSlaoDB/exFj
kLFfuwQNlx50FlVyBhDe/Od/5MFrqtFs0J/x0qvTvQBALXQHP4RwdghjYZz29m6X
bQfkY4KEo4Nz2b0yRQ4PHG65xcvPn13Cg20iSo1+oUrYX6UmBmNMUdB/HEptuFm8
iR7DF92Hn4H+7KAPXdNTMExnl4v8SxrMZkbMYHNFLAkJJOs68gjBsHwrzPnJdsNW
32yFRlrGLXx9RH8X1PiYRyMp2JjH5Ij/QmLxI2bKUKg6s+TYlbrgAwrkaKDqOW6a
jOBUvTYXwKBxQfU77iZCArmtWjt2CTC69y1pl+7cZWDirsA+aNmhFVY/PvZ6uBIH
PG/oTlM8MldZBnuKZAjDRv+J9wn3pdAd8ufHldS4Jq4Y2LmaN6USJ6mrChhR1fEL
EQWTsvXUEjAmi2Ov+OaEBCZliH22jY8z5msGDPKDxCeM1xxlr8ium3jDQAAY4j3M
m8Kt3zG+eRznBiooCw2uIpSRYLSToaFxoW61MdE4ZQCSk0kKkND+6eR/CBPi4lZU
qgnYKGevnNyrr3krhUBuEnfH1/gyicPaakxL+z1d7MQgaL2SBhaiO/MJ/XMaegyJ
QMCqRTiLx6EtKkAwf3jhhmTxJS//dhBoEE6B3LqDQf4kq7kPkT9MriMEOeyqLTRa
8Sruhs0NalaObiKj1kzZzLBkofvdjAb1/2ZNZxwOrxbbdBYOZ0xLj59JTWCZ8x6x
HJwyQTSUa34m+qlZwkQqD1+b+HqcOG+lBeTjRpfr6LJ5PsJKd/ZTAefQZlFhIQ/J
UkV5dNefZGTtFcOfngbSMrQtYgvn6bpAhMa7C1Yf12Mq1EECeipF2sJE7P8ecNgN
hIGWfZwsqTbF9Jr8JTLrZX0HuJQFQ0a6yN1S/VXyEnegIYkahNpLBHgNRkmBwXT4
33iwBg0BEvRQLHvT/7jasMudf9hjg3GjtNVnij8PHOweGA3sW4p6M4yU6eYBNueU
N7bWRwdC5guyHxIu/B+/uD1RBQas+htB/syX4Zj0Qx0dwelaY9nZ4IugxZBOGHaz
FRGHollUJiJ5OrKixsAp4L+Ow2KKWviwr8mVjQBF3NjYLkoZBo+ovpABv9X9UpjZ
rZrMUg7huNlSY00ZPgY5jp7WeIifl6bXenW85g/tXy7UkQnKuTd/bApuF+2GndXk
c7L58PFVQeNuuYFfgs1UA/byptt9DvffvuxjKyDVw1LCTE4BcySNEs2bjUCOCsgc
6jTZPLSpSk4HoC0WPAe84poSpq5uSa5Ri2sU5My7W25fdza3TWIQoy/Zm529WAKK
4wUR38cp7Fidj75AAnU3h90DgKfQLCS6gklUPMuuelAnFrBM/pq3JV9u9+0o2PVi
3XDqYLa18pFRvNL8J6+3cPZGAiXaLleJYUvKw7JVcnXgGbhreAi0dLL0UqAkZlHx
+pu3nebo6ti0V5vytZDBnRbOEFpzQfoXT5Vlm8u0B4UUzhhDAt5NSUxX7F8Y8hi9
+iTtoDPS3Esby8JpyEF7QJ1MZh9+oQds69fRp9wfkEwhj9+vjuTlU6Hk0+LrErtX
AbzcCWqnXlbsTIi3j58R3hcjSrADzq0hQM2ky8ggp62SBe9a7n7aPQmNBeeCBEDu
u66BoeTY8qkndvdst1fMNwfw53QscJbhIQDC4RIr2AJVCAAkOnxQbTorsiGMicqX
o5XVVurO6Y28Sc8rSeZ+GIxcSbe+7LjTolXyh79NcY+M3W3WdeGecS0iqGX7tsnB
Z3X61eszNFmEp6T5vDvlUFdCXkZlj2jbVRdSejOaIq3BxWVLyB5mqWCFywS4Z4EE
+tGFVwmlP1W4u25cCvztTRxfLSzc4dakbeOm1dX3UmAiQq+qtUNTOLkCNPxsnoQB
mCnWd+ej4NE4cOqs65GnwdC082YlvZf5uEvDIxxVKcFzJQE5TtNrx+VptMmRfR8L
/Knqj0fn+jGkIAb5wB+/SBnhoj7ueW7F6kO5JdbHzog/P9AJStqWJKSmoUnzb7nc
biCqqT71wxm4F+ZsV50KucMW8Kz/OZqcZpEWOdG0CP9xcax1UGkVwRhBtojliFEB
cBD2S74lcrRnYT8uM0C7+iUOroU1YLLrIHu0E3C1HW6YZK6IFKvOfpi1TJRpDE8R
zhGj793TMc3i18JFXeDbtGrtVe6fF/m4kQQ/mFMG/DRuNDlQZdnwACNOCO2YHl48
2xxovhcdFR3MebNF55tSVU8q1Ugp+lLC5kXmhsZePelyPm5ekNfb23cGo33SsUnI
pJFo3FNsDmigq4FHHJQacAavfANJCEKviNiFA2iDUUZnwRzCMiB+tZYKCifFpv8l
P1ULOPMyPsCUluG0gMGRLDCqzcdctwcidN8lxvu+MRayNdJscVQa2o0WJ9PJbR40
vbcpkxHuP4cWEEJ00YE3RvKfxGYcKO8AK6JWrkmlWhKY/6ohVyHCrtiH3Lq6SW8h
g9NNAQjBfFLLRtIArvhEyjG6dT8TRgIY5SdedMPaKsEA4A4WH6kyesBbdgv29vQg
LxvBilO456nFI8zPLWaEXiil3T5/s8RtdSk/aatw2CzN+k4Nf0s1qFjUXT2X9ofb
LyRaOOWAMSK6ZWdo+jYh5TdoEpFeFAGq4e/LTXTRHdckkZtO6sk+w5cP0yPkWRp2
S0JmOFZTX0Ji223TFqmrUMyqIV1sY1CAjuwal7ceU4xc9XRAqqAYZBzyAZDYKngN
I6z2tFx8efl88LdYHGzOdHHYHKOZXuLOOn/jaAlxCPe6EF1kq2s5+lHUTgQ+1851
aavkWHraLrTNVTcRGQmMdyNEZPomt8zmOT6UGuW9D51JKv8nv+WP0UFRRLexsSIi
0x0rO3LjF2BdfgEpwZli1RcfRtHwq1HZyDdFMArdnUsK3BF939jDUZBacXOc/8iQ
r0+0pdU4p9/ATPdU+3s/QboLrtHTBCepeet8qAKKKPbTfLtHysqMmCudSZnM6Pwp
9vW1qxasSOh3fD+M2RVuRTDVRfRRKPq+9//ZuiY2MJFKXpR9ucJtBgs9glDnFg4a
W1azsKtfM+A/xh+ZFxkUaTkj7OSelkwcfHtc7CuJdZZ1jM3hges5RMKJ+ULOPgGK
aSajN2ABEtHt6Dw5pqYUKkFld0P9jr13xs/bwquLK2r0TWuKRG0s5hahtEkB3XEW
RhDqUOAm4AWTDYU4EDCOaeP/9MV+DPntwSVBxtNK58vadR7Z1/ngjvrfybrWn2tz
zPWs+GKiX2yEi2MErn1psSTEpw69sklND0oHBJZkXEAAS+1OTglxekIu3n4775mh
vG8Rju6JbJ4NKlZzlnTBIqC2WF0dL348IGyOZJdDEYl2iGfrNTZ9MXz0zf/pnOEv
tHXuJZuFKdFsVGLlv0d4hw7PHih3bVL7jQ+0hBZLp13gn+NM8QDlEj6GSrHGq1mL
cGVwsTHFT7nNkhNzq1odqFUGsZH/EuKcxKjzj0XyLudcr1Pvau6qQ/t0gvnyJRkt
vQlwpSOBWzosbQ7n1XlTxg04HpTRInq2OGx/pynxGg4A3NnCJJIAfWqz3ZuoO1sT
Pci4gGQqH/jxHfZrtWrAISeBDRalt0EoBngZ4umrV/OqTmtS5MOpk7QyCdBaf89/
4KAJju/HovvRcR6b4oPpPe1oEOahglmUhHarzzxH4XDG25ci+FuzclV4RVemDR8C
+nKHxx4soy83So5qcSBziaww0cgkHB2yLDlPQPoa/eiKDABqGubqr5yQsx6Ap0+g
h1i/yIenCRtc+OSamXNOQiMa6nAuld6TIC6lqe54LRxEjqpJqD70lXqMenydqOfS
UuysEnnBMl/akiXoRkHVtpWCthJmHpn3NUOJ8mKicvKNz5t7fioeXB4KAip5Gc93
biChy0KQg7DpI4dHWn2/2kUhXN9heUQ09I0tq+lzR2n7rxz4AG7iCs0pMxahFMb/
XKW3oFEYmnq0GmpqDhWxQFRGrDpH2tUrpKGbnUnkHuf4Yigzkpd4q3/X8JBLD+0v
mQVtF2V+kU7pQ+5JZhWcT0TBPuNi8Ke8YhqYrfZWpO4vBTJSQFloZWzqn+1KvKKS
0Op//0s53YHcaIdaBGS8k4KPG1YoQpl6kTky1hzIxRb+9sgcveKGRvzIudkKuVDv
HkLnEfezHRaFZHqCK5U2vbor0Q3+0PNTOSTNPCHb6fYuSf+ZPz3FLBYwx4eENnEf
eAlDm29CfsEBR8pm5a4RMhL5RAbzc25kv3hnju7ATLt0UUFXX4/6XoeL92QWgPW3
A60+ESnT6i+Sl90k5mHtv50aK3yN6uqfyCcBan2BEfnCqpDgaUBneYYrZOtw41c7
nXrpmVjwNiJe8ni5LL4YsbALHlY4F/0l1zjVm7h3v5RPdQVq3QeFLRrG1DTdkhMH
if1Zw8OpHvAAHykXzgvFRho+uUVf24xfv1MS8ROZhhOLV6RNQAxcrjLI+nXgl1cj
TiSwqYNm5qttzN64aGE1An5NDX50QnqaSTnjUe4mbhWu3eJH1FrDJG9t3fPEBtIb
NZQ4uDmy+LlAMRvcwfNOZY5u40nq6brq/1gdz+7S/r/2Qh0xDBRxBFQPWOWcMHjo
S0VvXEIy8eMQxUjVzVL5q9WRyvKTi9NFgI154P7CHjLfaOCTn4Quj4SIJch+SnB2
Walk6A+7bbdECq2bv2tuIOLqokM1XEfhyK5Be1dDvGzc5vANUlejqTB7H8U1nNhv
4cV0OT/vwDt2MVftB7D23HdCLr4j2oMMIPUDy3m2Kj82j2mGgTAZZ0+tLACM77Zh
wyuKF8+Wsd40+TT1ZJwEk3yVzUeU8fv23tGKIH/SdxgaqhAF0Qi+DZTRuxedKjpj
COM0hCGubqCluHas+k/x+g9646DnJQZ5xd1eNm3g8oZe1XW/L8q0C4IG03JdDkll
gZskLjOaap1c/Q6A7qSgp4iLXB8gIZkhVOYxZoZDzca3TQhGT5QBLW7UY9TEUIEI
E43kKCprPuFnSm6G+CLViyG5JawfZ9zSSUIrDYqQ9sbXNnCW+Ch0flRvOu12D7U0
53JSsxM10wAIbtV0vKQdSYl9KzbTlkKlenRQqBvMTELf23C98Gzm1hKfAtRh/qD8
qJY1UR0SB+eEyzZoCORdr0fzZnPJOiog3UrLp2cb9HNdAHstxUOvpUFiGNxUTopa
1MS9lb2ERSOGXf3aKIuZsYXDWuUAElfIHRuSgbhBZZM66SAAvMAMvgzyIUwFofoQ
ASYQ8FyrVVLPxRzOs/6PaxMGTRojY1/tkPwq4hBC9b2K/UJyr0aCQN69TUSR+P7P
PH6yDWBaDXIW+ha4x2Z7tuBQbMiuRd170cIgK2+ARJk4aGctobBhQJqSzd0t8GOM
YGDV7XFKgFqo6723kSEJvKXOxgxhiwF42rBJK345gUvV2V3zsauDqoqhmfV/UNmB
QyuCI0Lefjpkzn6wLNvFBBiUsUCCuVHrlrBuO/gJvNI1In0qGFzOs6qErUufxtTY
Jvat3rcx0BH0fNyOAMwTMr6itDytATuMTpeqCbH70cSm+hhGkaKw+qkO9vo1T/dv
lEeMAuGU/oeXVHSdu+/J4ixfj3Vw/mXwukR89sCs1Cj2La+KU+oPOgYyh4SHKK1b
oSBNlZIPrYYlZvu+x1x3ZFPuFd9pxqOahYJYOZKM2VPQfyMHrn6RQawAwzHaKNBF
OZOLTBClH4r9Jgn7hhnayCpFWuJ6E0aAIq4w3MHpeCbPehRZsxwszNzVhUIgjBDH
AuebVz6hP1JZ1DYgbR5IAbaY8NDjw/1LsDhIeJhUp/i06BtGzy6/5Vy1S8QKqJdS
KFdF7+g+pa8CVHs/uTyJ8ZXXcL6C6FGRW1U/7ierZnc11TrM8mqlkFcEeYn9/0Ax
A0rMRhtqP7gKVkFnru2+Le2uRMowyeJKnPh7PvLlvcmQpRLDr0fQI0aXrIwAn5Fu
TE8p7CjDgVmIPBvdkbSG7kF5MTjCMfzprbRY/BwolEfYBfoh7BxjgTwe7uYyxsQu
gwEfwi3+R4zZxrFz/LeDoWKOsEyaljqGI8uNjUIIswUf2bP1v0ZICQgLPwgdbjbn
P2uYlqBEtFZBDFUc1pSl4xJKGEx+B+FcAv/E0lPs9s9sDXlJ4l8ZupOCcRlNVoEn
wXZW/+80xX4lWFPjEY5YeHi7lT311duNOzNTJoW116n9IW5jaXIPhq8Up0kRIVHf
DnWJG/JfNWkxzQKvr5UD+2Rb5rpHihxiG9l7wSODOX55ntwMET1Q6F5qj9h+PlrY
pmOuKEXrUa39dG2CbisI7y9gbs3O5tlBjXQYRELeLz2R03p3c9vbSDuj4Crs12XK
Kxh/ThihBcW0gajdWOm9BzcXV6el1fGvb2AFLt5cwOTjAmRlKGowcUspdtllWcS2
iZkxSDYTydpGgcVtI535G/fgRMtoj7ACxLo8smJLk+Mv8jLmtOSEOvkQ9nlcUqGV
fYEb7px+XX9S8stB4ayXIcbdHopzkvpDgnFAVjsO+29qmF6tua/bvSiI13HUvxxk
60LBuyoUnS3QUoHo9XSRhyProtiOfnmUnU5DUtchY4KlchWpoCe7xUxFDtKWwAkU
8II/QGIU5iIRubPYsqwkg3bwiDzmwDejPHEQKLltkkx8n5wUzIKt4hNmU/I9hLhy
J3EHCjIBxP6Yvd+edXYEd2yTeE2YnE8fz+T9J7fgN7IFr9WjL3Thn4IdQ17DzEqv
sDRrBk/EiTCBPlHYG8GBVEaWwEYVBliIrYP+pwwMIsPqhedigpbBJWL+mKp4IblL
XLHVUOQ+oKGZwe7XfrBxA/Un2udClZiScztpW7xfEPLIjULj0g5aPKAcfOTPL6FN
NaAjyG2NEgmngZ7khreq3L5ysajlbIdaqfBn4WZSxxdWplicrammTsXzNtJYOMfJ
54Tb5S8itbWQVXBh1rVXz1ntaPQpBUkhPVrZN8SrIAXYkQtJLWtZWmwoYeo7u/6Y
5KLAo9LewirC8GBQYckQK6EYCa5IT1rxPmd/dEkLJwhceluQS/OhW1CDzt/TQg1l
sK3jNVClq+3Qj2tZguxeGL5hm//kjGnDRjcB18M7ZBfOnWmXtDvkUYHGC8DnZOgm
r6ZS8ohLEMOftwmZ5JA4a2tlluIox+OAPQL/TTuqPGP9+tb5JlWF50LRzeIJnPhz
uRRwXk/qImScem3I1ydgZXkYkBgz2Id+obGM0Tc42Sxj6NiikDAv+EmVAZtzg7Eo
q6hpCcR7LNswy37piVWrOzsIZbCUfDuJGlyucxlsCsn+PUc2IymGpnyQnhmS2yBf
QwD3NGfjU1cBhNQlJ8gL6x4vC+DiIyggw1lDheAQ3t2sukF1kgwjM8IqOj/ZjuSd
nwHGJ1SEXUKrSeABQPNQBpu1lS3TZsfy9lRwY+jhT43KdvyjI/sNFr9vhO4+zgqx
UEptZuk2cTvxeYaT3uTf6j537xrXizktf97kUv0P4lDpi1EzZll1VKHMZr6RlCsp
ThAuEGFQfvN5NvEeNzmwrdKpmy7saLBiAAzStsOWBBZyTheJf0so4qns665fw8iQ
gojiAL3cTGqbee8KUI9Y9pM8mIdzv2dFq/CfU7zmuvsTAdQs9BUXubnoSfipKPFg
fgI9ezuE0PkTJss0H3+7k+6toBRCwdSVGwlmViygQUzR+4+PDBxWrVnxwsmkADnN
1sLGc8gd3Fk/4O0rO6BaLBHCa1NTv2Qv1ZelBTT1uddOVGcDJ2icODAwmS2TNrZB
mJ9Cs07f0NBqPu7qOHEwTtYlk/1Bcb0adNzkJAIbzfO5ADy4az54Ne0vaudJmV5y
aGvWzjttPEyLoTgoxMbSJYQJANtv0rQFGYeECel9zLNs+DkIOxshULdKLfSZjSZC
vu5cFrD0zTy9ubmhNxRCtTXtoTflP3Ip7jg6bwQx57/Gz/+t611QfwP5AdMaGJbp
GEJqSCBCYJ1u2gs3uwWQFmNpiWGG4eOGWYacybUOxNaltgKvaI0m4xVVsCnNYOmX
PY0MlcGqQkoL905MYfYC8v+soVWz6UylrGd6u/jZ6fmmVNdyfLM4q3HJ1jUGAI5g
eiiUI03RWq/yAuo3G/lOh0UVKaqZJvJGIU8wu9fyOOZC4fhgGjgWv4fxNEXTN4Mf
j0ALhw3ZVS6pr9yAN0GMseXUipaOtdhPtE4UeUB7uKIOlKLGmzxURz5M7Gb53YuE
M1EfGBo31JIdlpxHh8mDS8tjL/r2yEaVy5k7bF5Qp57ae0YiXozEtaOniq9HyhHH
jJiuehmuG3LK50OHcymKes1PfVjEAaqZQ1eVmVKBCgFb2IOKpUsibloi5aku3zYK
S3eEZFJg5nsF177iW75ze+enwHwQ5JnmFtMk92+KtcerrfvsrGad0SzVpAj8hyhP
XTO4gslsPStt4V8mcG74B3Xz/EMHgXZSHWCeVylJbcmnz2NHa7JyJyxJfnVX4Vm0
W1j49IzdU8ilRhHWz4GXiOHdtLRGDKEWqvwGL5p5NWAHXmQ00IRlyler7zMuw2Xw
duqCJiATQO74oL9J0voOFGVhffg0g6Xqer402UPlEWnSqrGm/oCM/t4LQa6peaco
XYw+BlufwHUlJ+ZJb5MUFRqpUN/TXKLXbmqCwln4NS+gPLYRYgKbtCtEhOrQy6Av
jhlpgOVZjfmYdq6TO4/IhTTWBdWh/6/HM/GB/jiq9gfRrXmbB7aUxi7zEXk/Wtw+
kI7Gvb7rvc4ncPtfabHmjUPAh3r4c7h6i0jFt7Vo88/gu1fK/giW4AlCUKmhzqws
xuSeCjp6issJ0KY9gd1kl9XUavLJcpEJJrAeTubwtxYgY86ru3oEK+bcSEv/S3Ec
kFHOZnGB6LSoZL++lD0ge3/OiFJ/OtIgpE26xVlUZ3MdA1eBRetP+bpbJmtohQbN
43sAzHaWLrTnNSktecd8CmIfNSjFiamm5XeaY+9VX+gWbKLg6LsIZdtlirJNyP9p
cmwVv8MSDOMclaj4k3whMwzQSsRRVCUKb6G1sDX5sWVokCwo7R2nFvGb0Yy9Cew+
wfOX30VMXk7aymKcyYs5tzqDiwoSpvkC9V5tCgzO2fRlgoQK+TBVwC5CAE11n83/
AOYfN62ULKAGLoeYf5tHDzsVv6+Fa43L0Vsx7eMeNq+wkc9v/pxlVy1bdv93xzfA
1GKS6Ex6QqAK89hvpd7M1rKN8Jp/b3ZL01BiAf4CL+gmRdtEi78ApOwYNY4rvoww
Dl6Fb1bU7rzzi0GusJH9h25W5SJHRyUy9I2ekKtc9msNJMUQa5x9bqDH1U6XCH9B
Rf5KbbbKeM8+LrWi6cT+/KhtEf40pDZEI72v29nuFdToz6eh7ozJVZEyv4CPe54c
vlmoV/xllzmwrKn+n9TK7qIX9d2psKIoP5h33vJipCnRDHEmUHrgAlnN9H7XgRU4
q2gPmeBX+18rS+4llMfICE3S1YIJtjmlnEsur1srKPB5l/M3PqSirnzMPZdFz30f
drDVpzAzoT+DHcjI9jV93qWHPxO/37wYQ1PTtxixGjXPn0iS/PacvYu8kMscbRjI
TGbaQRiI6B9RNTo0RODMwNZuNfWKFr63Zwc4gJP4IwoayzQunu26bC9/SLqmwljs
kbQojrkxJcsqZroWUWlVIjtOwQlyVT3ZcTEVp5bWsN4OHdeIPijUkBOEwFg5nhop
mxi3xbsltgn6tenJEPNwljptJzqi1o9c53cplr3pkG4e8nQvVbQN4NCnrIXQ1c7+
HEUq9XxjMP1ipFnV0ArOp8G66f8qEM6FV6DKeZIdD+VuBT3XSp7q+S0tdAQxxek7
LNpg1MJvrZxaha3kXRQ0C+uAGriHZY7jN7NLedzWL12h2vzq42gQzFSpk/EQCT4s
VSx4qwGYlhzTQRCvJJcvohvH3l/PtExtAYuJbsOPWTBmyx5FKDsS2m3H4mhSy2xP
l5WSgeTTNlTW3ozlOoCvg2CPMD4TvrNDZUOJNFON0cVmBPNwoO/dpUf7yO9bRUnz
u8O0CAajN3HRqw2u7e6gL6JUVgF05+dfkDJIpZ60Axd0h6/hGaJOhPL/HgWu/hWZ
1EmUQeyOGHhzk/EJjZmXHFgqEsrQywuUtOubU1DNhoBk+/6xLxlWo0Jxz68Hcrj4
mI9yuV8RIPmqacctbIOUxnspBHt6/VJdoMJYY6Ksv5wJWaCFDXmYlCFlr+vSi52l
XV/noX3TYVo93NIggw4g/52y9UM8+YkPkrZLTYXhalGAfS8WXrurpqQv692ihXaH
dMCSxl7DJHCdRbGe1a9fW+CqZfF5j9KlwMVdoT2hTCkEP8Oz6RdBX6ZNkm8D6Bhr
AxdJm1CijyK0sDx8yuTZsgKyIa6S9QXeHl6LamkLEk3YQH8GFM463OOyOEKO7D6E
6zfRiTSW/FnfzFk/vGmlWmEDL0uQLInndE71Xd3lmr+1vKbE1or5puxj/WnXMqsn
st/2Q2BIYGxXUYYu7XvmwKpn4TxXLTqz4aeSNXdHJmYpjiB7KApCjx5OA4IcozoA
EOmUrepKyG2z0I04bo+avj4ED2TDVHMu1pR0bFc7E4V8joKd51nG8kH1LF9LCw6n
G0x79qWfd9xrfkfwBSnjQOZstnKVBgnuRLjioeIqTEm4T8bSy1+XVqgnBvly4PAd
hBtajPAqenODarZIrpprhEjIuFAPvhICVkzQmiFZH6zDlwVYLyD8ESduOS1EkfcF
OOX0jsmpbbz/bB80dpwAf/C91wca0Exj1U56SghCsYH1kns4vJ2YfIRAGABSgsfO
wIQKF83wu7Cm1W5NJFUqVYoWwHc6aGmZvcoQD95+UR638XiBO0L/WCBaGpx9gQZ6
SZV40ZDeouO1bXwZpsxxQ0n82b2Jq4YCHmVLlNeCNFV8lt+FK5UKwhkLgeJ70TRo
yYweGdbiBEfYqshCTCfRt4/oTaQSKSc2tmOiYZa0yneVH0papoOfBv8SekcTOKIO
OLr8NP3xfr2Ilnc0fRqR1KKmZ2cTUa5LzLO8MWrAMR7tv9vbPTwInkIssYq7m6pW
DQOpnYOfhf9P7erRIrlIOyP44CywKHjZCzx8bmr/u1RiIRqhhUGoLiT5vhlzgSry
UsBmKZgXSGNmvgV0PAax5Kg7ruGwqaPTi0qMviqPEG4iWCXL+iiPbPK0pjP2Rmk3
1moyvSP5DbpkNHax7/zVocMKlpK4E/JCruDHYJO2xAf6uLsO0ZHiOb5rfDMayMDo
4t6DAKj12TarL9kAoHppU8G11vRrsROfi7RRBhtWNTW8F6eGnJhvBiuFJyvFqc5m
QOBY7/HgdtJlr6k56lRyU7RomO5+XtoG2AFAaOjUSPTM95qcdj4bMM/6YksiJdxU
EJhA/zLZv6tG5hyClHX3czQ7QH60WBHhiPvNf12StvhX2DwmAkJfZkCnGsFqsULT
FOp7k+xu21MDUq/ETtJANLMuG5kD93CjPsLh/ADmy7+2vR8WbYL4Rt/E1nWxf2ix
Mr+55oy8/fURsadundf0mvD9rignTxTLylZZboeZyUSWsfDgbkGCC+Gv/9ee+lFk
NzMoXlRvM9CjHoYpnEHDjdbM00lp4GQ4GOmhi1LHGZL8aUJx3O0sxWyi7tuZ2A8F
ylAPiYaY2mebwNMCRSru3QBBpAns4KvOJstjw+c/aB6GH1CH3z+2A9aBt0r+JRaD
qijuNZZ9jBVybS9lBQPwMPIjUiX1aOT1A2nAvLxCSCQY2EuzRhVnTNgnLKBiVzB9
hDO1yr+Z9KXZQrihU2QGEzbEZf387tQnbSx3tfSKxK1BstcHWZAFI/hfrBAEYSp/
dyB27BKFvfr7z6iAjDpEZ7KeVkGGtjzsFpWVUzK1o5w95SE1BxeiLZJ+t9q1eDKH
F2bOFgeOKv8MJ2lk19MLrtve6NJd2EBh5d8Yj9sGGUfJvRJ96QE0x4wHsQ+Rkn0W
B+otbF1pR5Aoh5z1I9PSs5rPp5KCFGfpnpvg4fZ/+RoHUkmpkW9YSwmizYsmwyC+
6ixhwUNbugfdw6r/CuUfe+gwLNSoXLKFCUvI9CNQM57mnREOsitOYHgcly+KzS88
t9bEQ2wakBT+BLMtWvqAYVJt2yJZUvgbjuUfG22Xhw5EhD7MICNloaUqEZBPMCVr
tDD4Wqs/UogtYSFC9UZDS494wa+LCObepqSbLj+vte8xQPHMCmhZiinMB2qYrhs4
vbWTfOCpRsbTNBS/uW1ytisvp40FjUbZ6DdmHUl6IkfrhXYPeEaixwL0VBwLrLOr
pXeoOg8URg+e+/WTQmT2F5Qhvt6MDczLGxKiHulFx8n5e5K6ulRhRCxx2OGw0AQe
BtDnwXTUwPvnIJFh+SccLqaP09v8B7ldUQ+cuHHeHGQrrtDiSDFVVKLvTE+mdSZn
RJOQydNPdl9Y/a62mUa9SajawDtja1YMT3TAK9A1acPGdKSxMahouEK2drr6YSyY
GobhZz6MYxT+31ErqVsdf8pMz1CBeT09cJULSHuu45oizZT9wLDCfuAaTva0yzNE
gFqpfK9F9jZYCWT7kZNXmgsXXHAulbZTW30CRnNzFHsz5afZhF4tcWuib8d64IMK
LLLXcdPLG/dk0ISfq//CiYKJk6BNxoCWYlaFIk+iGxhbqWpRNk8jowUHW9GzC0o2
5zBliwQuQSfKS/8gdxZ+qCCSHS/oGBnIg/iuKPcgiTO/nXGxlEHcFBuCak5Yp+Rd
PTjNKHd/x7z381pIyaUpakV2O+FXgdAzba2nQtiokVSx3n7ulkNPYVroOptZ4s3R
UouZ9pnPB+RsOt3YvftS7Fj8KVgSMF53k3HwfZ/xnYJTHooanPZkW/79gmlAtaEj
YTy3PYDmfV9+CB+Fhmz/UYDDcsPnp5v542gefT6dkcspCohmD+S4CqJaZGRMBrT2
j1adHZ7LB17IB+DA8cOyxUYkI0p3SlIWj/VgrO8i5RrIQRD5JQNaDDwsGOp6oh4v
F/K7Pv0ngYrfHFCYt81kcviqP2uWUBWIb1WXOd4lXPfh9xIt0P0y6xlWTW3RZ5EA
lscKdll//B2T+EfrfKvM079bmHREXEoOUytyszuYqr6R59rlMTZPVAmI3cE3kk3o
gBpDpdQ0KUdfCqEa4BKH0RZ7tSj8yML5FCb9knPmxT9VLQHwIxbN/xvJSnEc0r8D
GK/OoqYBD2xMrA9iYtDoJ37p5CwOqXAF5FmepGGuSx4QqTogmZF7kzTzNsvLOwiS
Q5Jz81aa/ZRJsTTZ9oavfuQVZyoKAFghJ0ntrp69o+543UF0WONwsTrp8FKoS/FC
1MjJ7sUf31kLvHZWJUpz8AJLxqO+Y97vVSzmrQGXpW+673jD/1hTzIUvRBkc7yQU
iowmRwAixJ2/EvuOaSvHNofHmsrqT/eB7GjTEbifcMQYYu0620euTgDZT2G8WYDV
WbnTs0u42oH96E8+Tgc0b0STHfldR190jrEEdE8fzDmbii7N1cs2GFvMKO8ht304
yZt83KxBS/q4VNZOzveoAmuS78z45bukCE54Kq0XqNNuLUuCinkDVRD4IsCGncAw
OBGVW5Wcr3IqdzbhRlYcc20YugEKB89DyzeycA0LOzH9SQYCX9bEx8DentE5l5A+
f1uiqbEMtNzZWfQl9svRV22axQg+royxtWklsmoRWcP6fPEN5c1H2gAqHfYtPJqm
ThS6Mi+iItf2eFUcQeHIrCPNPP5Jgs9wtZb5MGtntlx13yjkrsQtYWJjY2Ml2qZr
sYg9ABt++8kxzRpCAKv7sheLYIlMyPoccQ8+R1r/ZbEHfTYEO2oziMXJ5eFDR01s
6eqcVSnvl+0BYepk9f26Pc3P96Jp2Voq0s5mKwf82eZRES/hw7WLAxG8hOWUvlGR
0s83nTwfFCw44BzNDkTXJqOBmV7sAxvJTU/a8phmtX45kwLblqwim2ydbD17aHAx
DuEnZq/N6O4uIPHD5t+e8ExHN256+dcXI/tcgvJY9ty0X6AvELUpS6EtL5NvNV2T
uehiRvZepfL7etJf4zpzZZRnH/SrfziIwcEbyGKhyJ5oY3H4VXbBGcKEfcxJDIez
LKWRo9kzcVCRgb4JQ7FYbiGDkrKGnIusHShmTwHbMvRL4Dy+duyDaZM+MML98Srf
JKvVfcOCYLavSnsMk67Rd1lV5N74SLntZGVWUQDmDlfDdDjsdbtQY4dzTQymkQJp
zqne61eCKWVbQv6Oi56C4zlHJJUX5H/VU/xTTBBRIF3nc9EKMMXcwq8KxlAMzM25
1oI7Ra6b2H7rrL1vf/IdRhie2VIqNHyUfnOwSr9QXf8SSC6ZKkN7da7ZRP+ucbHv
g7HZpUSohMZyBlbuwrsqOPjBG2O2cK6YK1ZmPoxh56zbujMCpCaSOkb++2pFmY5+
vPqWTpyePM5m0cnSgyGgMr3sWIvZp+Vi1klE9AHxqH+PAXinx2YLgVmJITxdaE3d
FS4jrwAN02TqGUEBJ0iYpOug6jo76FfYonnoxbTJExQBRu2Wk/aWE6FwRHMQFnnr
bHhU+rfVE8VjTru/Uf9R6QOQ6f7qkJW/QBTW8IG2tnGnTYllQ/uppgies/wGYJqH
PVblWUQegA9Raaf/AxmuSav9rrQe1HuYMH9aWY7dtYt3hGYdswGZhIbg8tilWZ3w
9z2XTDzuUnoOSONqMauA2nGWI3TpRPRasgqnlkwaWdMyoC65s8KKqu37xkLgTlTA
WZ/JhrMJkk0N2lyKkdFRWyabcvgbAVAm/crtQv1w9CnmRlTIxCUV7vepTRSV8aY/
WJbnNTuKjhb6+pi1TOI/LynQEOSJkhoR9VjRW25RAqZYodeTgss16zRyhWVvejpz
3pr7gxQuSdZ4wod8+uy6FgrioCgxKf3OQGwuBLuP3WXcZY3O2cqUj76QtzVKXSm9
nMqk2Y+6MeRjq5V82jE2IoCKTeHRmLyDCw0Khq0HOwwP7UOeBz2YIhYISi8DxTjJ
24OlDvqWOOcMSElabQMyn6g24JZqivT92lknU+2Ild+SfDEB1RKdZafp4VEdU4Sv
mHzhCu1r6fCA+p38UQOtP/W36D9q9tzxI0oIJwcCV927cupIbN7ZPt2rLDoL6HvK
f3i14u5R6rtZL9Cwjyv7nJejIDKOzfZQA/PnxzsDrjVjpBPWqFp/O3a/Sevu8I2S
109tnMioJqpbL7RZ5TvsJK3mOoHMHO7TJktFIANckeyEb44PqF0CMnekAxMOYi6P
+ZrhC56X0YkQFYQqod6WuXDOH6VOtxObPayC1nXUjpux5XZvRQegCv/B3Y55l/lr
27gmvzfQrdSXhARRNoKzoIMy1dCyw4TRkyScmJgtjY4eg3eBJq3abeSw1WKwdfBN
oyGJoPEVpx84T8MsX8HMtl0S5Q8TB4bBelob/G3UdhYWKiw4yrAWLykmhFS24Dt1
ESSFvkq+68nLCjmtxNcP/WU8z8zIMb8G3GAi0jYzLTjuQDSdJX/GWu779ZKjhXS7
KRHeWUYD2TlNHrG+w9rliLOb0XWHvv6wTr2YfKVIYEOv3sNm2r1OMHt7wS/ZOhzU
7WVslDDKmDQ8BjsOnyKIRJEtz5YiTMOZgfPydw7XUFB1VhdD+3VxEOe/HGqOEK/Q
46dL4JqKKB3/9jsgQBH8VjGDHkc/daxnUS1FxlLUW0k5rbD8HKUaaYTs7SkUow5k
TpzuCA1E22ylkIjGMXiGIynIkY8RvF8gFeT1BuIkDnEJfgPR6TTI69aGBl918Cff
pfkfkEriv8UU/nlwWNyV5wWY98/uJ9K0yVdXUftqu6d7xMX/RvYjBcDqZOu0aPJc
fAlLsD9LEFD3YK6lSl+B66JccWUvuXeJtTNDuPnwnzZvO2R7Y8D1ewjBy24Z3JJQ
7NoeXGUMtn5Nhak+dXIrismVyf1zJ/aifqtdk5bPWr/wCeOlwdPtw9Pus8ulU6Ni
V8B0y9aLpA3lMwFqrDvYS6AJDm9PFZaaQlEc0VxuHIHb4bwNkOJ6Z01BXj1icwzN
N8Dw/17swQjI9z7tHQs9tajxPr1IAGjM89LuITu01BJwOTzNo/AxA+3K1KTQwTTD
PsPBANE0C2l7kLjPQgxPQgHTlfVuANc6wjzYHH6c7Da+4WjOyKtgVUIfqNtNlCz5
gN840zNaTdiwNnZKysOcO83ntCHC75aqjL9lDouo/kyASQmUSK7dQTXGPVMUY54J
MhvDY3zECi7EpPVZO4ruGIxr6Tw3gNjHIPRscdnvN7FUVTmEKhUCkpK74NjfbjU+
CphG0xr1DAPtQ/B18zTB9eL9whNpWfM3W4qR+RiyaV5TbIWeAP1lV7V2MCj83L+0
9su1HEvgtOGDJK4XhnqnnGtC8HJI9rHjUiI6qg0CWurI3GYHEBAnmM6LjanHpWo5
oJ+YJIsOc09b3z1FICY8cuOt7Yz5S392dV/N7I6whfcBqAJM5/PcAmFu7rC0Z1Rk
cNahq0h+70eH1AN/bU1aT3qu9jR402wy9idTtMkejVhp32Em6Ecw4mY45ODM5EVs
vS0E9SLRtWMK4rG1JjN4gMl4j/WPygz74DSHQwQv0Bba6LCQod3YaeEvQ8DWu4h1
SKHyUr9KnskMVNkikIJvSCFlB2aU668ybUrbeDiFxWlsw+l9WLdhGrxcfrBU97kH
leKI3J1AJRN1LNoZX9bLFTB/yUpwwUc+vZUMbcJP/E+dAO8cqPTV0T4MRMVlTTPP
hm81Wu6dQATSjK96c9IC86U9jYhUFK4nEKl3k8O0qNu9cU14mWCaevUOJgJOBw0n
K0IkqpMuUys47NQfsLniKtMLCXzCYws/vp0R0ZQcqZuBsvZ0PJsWS7dXP8qeGHMf
9FkbuLfWFoyNslsV1Q6GekUWy6e/hQcUqQEf8hrzTTZKeAd0/NfDBi56YHicGHn7
Hj85jTajAkFRDGJ779WpIGi2KUvtTeAIxq0uJGHimt2kj3Tuev6DPF6GPGH0rJvy
VXHkU1j85zfUbKbdiYchK6+E/Dt77Rw5lxe9837Clj5OJvbhwVT3q7+6f+KGCZ8u
1RebVfoEzBE3ikLUm+Qk+jJADltFu0QDp70pyheN2+kyNCpNDenJPf0A/WaadER2
9tA6sX2h6u7B5uSCIQLva+mtpY+zWPxTUxqRjIu+m6yynh1JKFQfobp0DEz+idSz
6gdw3tAGy2SbZrmjxB48RwVMTJ2478KADbE/8+z8PM2q18AlDxztyACZ9NXwU/5F
YuS1J+H3OqJauXvsJ1vM2044smkdb7bVc2vrZDzVL1MGCEQqkU69YdYTIQ1ftXWH
hbxYCt5AmsRpaWjGJLbRjjUxJn8taVTFaE4qc6tHxeeCInXFnfau+lpdRGQpRYmy
4fwp3exRPccbQKiIgKpjP+uTvfHCfyKg7kWQdQd0mDQQrPc7qpYa2j3Aeh1MOk4w
aSKPkEN1UeG5u7tuebSX7wHN9SLxospx8DlOhE0YYqhdrc3nRVuRI2auuMSIb0k6
rHn0UoS10waE6rw8lFxDY8ypKgl+P8riIxR2nq6EQrJHYtyv9Vo5CTL9KfmCpRPW
/Lio6LinEwLj+iVjhaTJ74A7K0EFpvEcFj0BhwWMUSIEgDPbxLv+eVoFpVg2vCE+
ZPwwUxuK5XptBE9q7VUWXo6u4RylwhVpwtM2LfU6ukNYHwoEM+ip5PxCGsXgG8uk
uZMt+Ee6U0OkndUFzXGJp/g/FMmoD2ZOnmzZkTQIQajx4802mtlEGfptc+bwmOgB
KgGNVwPvGeVT2pEE9JNSfUSOOZM2X25nSlmbyZfkXP3IYeOw3AH1y7Sx9w520vkk
ec7ijlFBnE4a/fAPMIh967BshRm+EJgM0X4pkvqpn+fhuOIkGHoF3TcfeYkMznHt
bjdVz1Qjh3bKszm3eVUEXTKE4mC8KI1G0fR9KcdOQZRIE+kiiyiNk60Rt+o2Ekrb
0mern6/YmV+tQ30MWBD4oi9XpDMwMgnfAwOIS5jUfWWqdFwagou0Wp95+eBjLGgy
/iuTtpd4F9/G0NbF32P7MBjWYnned7PHVCqBacFOXMrorXdUNEEUoWccNS/5Rnow
p8a+0gXTUhBxThA7dPaLGFoA6cgiNqWsU6udKl//I4PiEyVxKAc7k4eECvPicugD
CMfCz9q9+y9wHg0OWkbckgWOuGAkIxAxcDwqDVoz/yntSjYBPKYVirowaYctjVXk
o0dDzr723r+qBpc+jgyWxwxrwB2BdqYd2SBw2B2LxbMmwnbeBHzu19XoJz3W+CTW
+MiaAElVDZ8A1p8qsv59uN1lmnHeL+kvMwh8pTYLF5LwtYHDbJw4OTbgS6NKX/nc
pw4NDCSCvg9jBWpUK6tKoLD7Jbc3G0QO2aJEdu9km8oaybpFgxtYrP8TgKYPdmj7
pelN4BR8wkQtusOFoLcsZvuFghu7RbZgFq6HuOtthhlq76Szg0CJwo+Rlc9b+/Be
3O1WS9Jw2F/MsrDsuSBMqHK2Q6qVuAn7YlPMNOP0dkQWOjfnwyJGa4oESOLdyLLy
FMsb6+eKyNX7CvKVepullXUGWLt9MAqhYTPY5LXCeXPKVuC76D9YqaG6XOkkAyFC
Qf/dXJ1PrkV/IwAU2bS+nRfMy6txuarTGb+GBIWd+IaFaGaslPrwucyHeKGMua9A
ehsFJ/8YbN9fdDKhjTfnOquFSI0nFhhgr4YTohs0Dme3xn8S+n3fLOtZC5GqaGzP
rXI3LVulxeu7zuL9tU8WRzPWyj0FxysKXP/m35/Mer3E6EELWtv2ZhiphGsrHEge
dGR7mtFhnwqdD2i/Ughaflby/BBg2H82iRs6FFy96M4K/a0EUhhuuDyofTBuneu8
QUEatQ6Y7+0dlqhtGlgnbwPlTtEHNqTkW92qAbGXFB1DzEZIu42NczNGelqKC+ex
UMSRtYLnmgq/F4L4ewLZZzKDwHzLkyf3qatG/A8pqAYPTa/bFX3wTF5BQlHQqEjr
69sqyMfFLSI2KtNAI3TvoaBN47rL5d3uJgxJb+imGsKhAyf4FFsFgIrsxPtBLwhA
7UcCcTshzGN/BEzMrNPT4hX6R9weCB7idGP779SgxH86IitASorJqkQ1hfolApv5
ke9csqWEX+9vpENXLOWUnHjwV30iOn32jsWO+J0wwsPpMwbA3jUEoM0QuNLrDYJ7
BhfzPIhRdtLK5Ux2hac/AdLncQbkKzlagBwGxZYtHcOdvI/JsRJ9k1HQBXWqy128
7cagI/Lp2G3GNWawZJ4INAVPGdYyd4r3rOZLEiHMuTgauGgitjvbw2JH1Y/RGsDa
mSjCn4Qm8svooh0pr241f0eBJqoc2dnkxFWcEuoggyRESdHSynXYISJlqFyyG9Cx
CfWuvOUkF7zPVqZZsEc8UTHWoKtwB+VTSq+0qo/eNJnugwTPjPFvdxeFD4dxkx5E
vpWXQMYa3hj77BIZRQZLw0/5eMwGenba5HBXpa1CbqYl8KKVVSV/jDzbtjIdsbaD
wvMcroBXB5PZ6C/kQWuvPhyWle2v1xwj3MOETQm0Oka9Lq7/OWxZymRc2GPL/cwm
z/qTA7+9pkcQ31Lqbet6dMSCguXno1i9zrS6Cn1Xngg+9AxsUcOUEAHk0MkEcjMf
w1HQcwodwN/spyXbnlFkmWslkwC8xu6CbTtOmRV8iqiKXmFmnT9y5h7tnpkJGTIM
Jmkw4XNhHEoJ0S5k1VledbsdjybESJMC3o+m8IFP8Omy2eJwMcZGc8VJusygsUSQ
+L1A4DAfrfCvfnnLWP7fRTRhc+fwi6LBmUCZB5+d09muhRv1d0NFp5nMxsjNWjtL
2vSfzkG+hcjzIuOxqiu5JsUKCwm7z5FqJeZ959CwvtT5jCh760uJ3cDyKPhdcMQE
r5DPaqiTDor/bytps582p4qoshfEfTRl7T93i1btXlePzy1FcMMVsUYUnf6c9PqS
CD3Ada3L+PrMBPlMyl6Al6hB5x37V9tId2wRBjKzqoQqX9OsWktUtITC9Iw/YNZY
dH/kNTJpIBpv8L8wmf5ZbgbZhFB/Ow9uaxubO5k8vyFz8qF8Al45GnyIoqTArDB1
QGwMXFR8D2/C7h4zg10J95qzMgwC2NZjMXZckqNRouXwTCEZBWJkw1MvQ5pfq8P1
KLDv91v0gLAbkZ3DB0HnulYy3y+VnuMFEVKx0iZy2xWAxz+aoZz/J8+VqqPo1Ezs
wYccwSje2aSdAwpWNGUa5PlIK2R9vMjt4kNbli3B52KK81wAyaqZ8YB5tF0NkhdR
aYYoRqOPQEecog/gGWCKyIvi56X8fKc7/oIt+KALaI6kOslBZ81UlC1xV916AK4S
PZsvvv8eiTnD8TYqoLEf04xZwcyKdvZQijVH0Uqia69EnwXdMnN6qEAjf64YOogx
QxJb9LazUbCtpK1og6LY6ZlKsPF5IXwjKZlwFruXTfjjUEpKVL+Lq+qMQnpK+GhX
dkrVOYPXRCEiZ9qP/uJqIQ+2QcIyTSmeElArynGddMhTlTH+oGLPZLaxkDse83sx
MU7ri9lStGxhJFDE/V3zUYG87ooAWeq6ugJCaOTmt4OJ+kPcaAcPecwtlE3I5Ww5
DIg5X1THHaLuV1YlttFjdWASMiHO9PB5gRStHBsp7VmBLb6KuBqRtqJehIfh8qCR
59eU8j47BuwwHXKBaFTK+07oqKBRuRGa7KRAeKnbC1m5KOod+pd4hlsrhyaNEln9
bDdQAoDvs0LVLSdM25OSuBWH+xwxIEa/lBC3yOtlNXbuir4YfJ07rvq0PJ1FU6C0
rKbeRyRWGuyXt551g5LKXX0B2k8VFABGX/x2bdVKVo3VxNWdgn+r/UtcxzI975Ca
/QXXSAU7JUWil5caem/B2FT163M1BBFDpsN53WHlBF8Uqfj3Jya1X6S30wH/geVB
QyYc/AvTg3YU4P0zaW8IOQujUUeqcp1lQo25v1OidVkYtqD4n+08QMFnXneoNSRZ
vdCsWsI6qimb/GJC+d4vOjdhoEkwHfxV84CHbZEOuzsOVWVOhVZnNHUHqx6REbUa
LS0Kye5l8E3uCHlBEOVVVG8tBbEm8X1Ra0gP8kSoO/C8ivs8rkEzulaOLjVH3LL4
XDJiH8C6CQNmljQz37KvXHMrTXsYzcT54H2nJrWy11UiPDbeaRy7P6wnsbEg9hfY
yqwXruYQnKXBka8RoJ+v8uOAof1IztfI1qzC23DEHqIY3ynda8tK4/FCq7WToJTh
7guhsIMC2B5FmfVISQ0FPpRcROlcFUclQ1CPO4UvBF/VqXSCLcnjRH3HA7dmlPcj
tFy0K824Xlcivn1IVd7agXQ8z+HbOR1CthCBSu/SvjheazBszN2X8sQMImckys7W
/WxrN6yMmMjUEEhhhi4xQNwDg5I2KBGdFtBey6G4LldJ+Eph2iBu3KnLunemGhNV
Bv9Wt/bQ+hBBmQGzhu/0dwfNwTPTTi2xCobNPlB3Fjwz/P2mSZAcgLx8FIuRMFrO
1l2M8zv20RQPeyNNvqQnchnzWee5sxKNOnmTsi3U627/M3CvPsnQsqCFTLnXyX5X
HQ+6qXdH0U5r+Yx9YA88wXlCX+6kVIQ1I81P631zpc5Ni0jDNcTF4Fg5WL2DE2wb
DMaPDdmVVgadZRClQa+e+7qFgN1BM9xIaHJfC3yovycbBFg5FOXZdImzhOQBVkdG
P5W2UXMYqTMpQui3jsdfAggbelagXG5KbR/jnAQ3nidH87RRXjSofU0+JLzPBCjy
9q6XHpBNN9pMOvmCsxuVoI79n/7T/Icz7KgGUrBpVkLwmGQBksk3YFapLG0wr2cE
VAQMqcJBt3AqFesaIcLBt/GUugFg2kU+UJTusUBpI17oDr3o8qpiUQrquQ+OwjAZ
yGcKhgBlXJMSZMTbvAfR3ub8nkAfWBRE9uL8DNTpOhi58+joAvaerDKzMzUWrtuF
YlGPUQ234ARNVLGRudmKbwtrj+CuMGRETC/RjEoFXTsyxMu9FVwQXtZgwbsv6iuq
YB/TlVdPVLvWEnz3M/uU2+WWmI/Z/aXwVChSWpnO0ydQ++x5bKk28YyWrRJTBjUa
UcTOw6G5xwTVX0QB+YHW/od09ZtzenxmrYiPRk92T3WsQn71VNtz7EivxjhF4wGW
JBoynf8edGfJzTsVLqbD5bBuUzdTgWSnVzFvZEiuu46ewmlHNvGx7EnmISscRsHN
f/Pdq/bwFtSw9W3tBAps6Fl/tnbjgz/Y3buRbXJfBo6OAi0RnFYKcPyIUCM15gnM
f99AkhrP22qMPRLcqC9+zo68IbUCKsT2uB1NiPYZt7jplCFQInQ8c0PdCXhHupvH
NhW4iaTW9T0WKR0VQe4azVRlucnWDYbkQT5e1rwX5uLkxJxu+8wQmMUzj/Swf9DG
TB9nEGMWZx068qzXhICn1gUOyTQkNOnzkZC6o2pu0qiWVJ++X895o3L4BuA6smJb
KEyhxkl26bOJ1u8YvfxCU7+Cakqnsfy7w73R1ALQxUlCA8FXoN8PbkUMUyPMPbYB
hubA3klAeUruc4e2eRIqZsSH5KmRIbRBnfoiPT8X/XApH3zzkG1xjXt9YBm9ZKN9
hc8ls/PX6TASqACfZXIg38/W7VS8JKx+SxXboSWE88ef9KBHIMn8mESoltXxOKuk
MMwyxpwEn/RUYn01IJH1A5s7u/89ksidQZMXWmlz9N2+24HPdA6BCdlIVvkuvlS5
OP4cq/nca0HyAyeasXMeN6Uc4S7SSDEQ8nNb2ftMbxr/YHXbhDOgs0pJaebGCG/i
gZVDriyOPEX0gcyfy4KjClMQdy9uQi1v+hJSk2C6yfLby9wSQ3E8zqUuB1uHEYns
nEFtSKeW3Hx0vqQqsXPRDneTfV819pqZ27zGmLON5i2BlYa/ANgULg89APaoApxc
S3xo1081fwwoQyzg9CTvSsj88qfzU9GHE0eT9yo52nLQo2Fzn0jtXzC0p33t4tIJ
v1X7xtAZwUxxSXZ5xLPmcw6yxZ2EpIAgqdH07TwOfYfhMUfDF8fiavHQXrFCaWu+
byGDogxzDXXfF68K/ZmNYUvktQ+oMVCv1VqS4mkXi7dW5xKlymJYJJu/JG6LBHmB
GugY5oCpG+f3yglJmADRNIC62pE1EeKvCpXPoJSOCMn4bCfpOBt67dqVfHwAHiWs
CydrNjvqoOcMZNgVE/IHidG1GpzIQininOf+KcbVXQvamTu/q/WUwTqtrjspQzwd
mn7hKQDRcrj7YIp4bj2eLRYa9RX5YiX0KoNmMje5FhD/N/mb98zUqsimzusj1Tx3
ictGulcqh1uWCv+kJEiW39Hjkc0C64nhXhhs5fO5v3te6QO1r2LHwc4q/bkmtLhW
M1ZH6poBSsE4Xk392BQrqbKSCFw/MliW5o7omiHmninnz1KgRSqvIo3yVCF+jN5X
oK+f8jk/uf8xum0TvRaNuu4mb3EmUpyWZGRC/KzzqnMVvdkx2aEkGoSkAHegYr5a
lBrr7Cx6r4aurVMxaZW2qQY3bhaM0SEg+HcznyQ06q3awsOJSfHMrcVh/SLMHLzO
Jrc4HAbWOBRkHjWSwJbIoWvaLQLI58yMqZ8HJpxbxLzXnlM9zagwWoZN3FY+2JEP
yLUuR7vj+lL3uVbwX1CeqhffdsLC8fED/mVYVstQEokev0gepMM7IqLUwIojcL2d
MepokJCLI+si09MRf6947w==
--pragma protect end_data_block
--pragma protect digest_block
8Oo78LKcLa5K1o+HxS6y4Gge3RI=
--pragma protect end_digest_block
--pragma protect end_protected
