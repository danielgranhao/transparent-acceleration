-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
dmTQEqquCDkYqMIoGbrIkKAtAnsCZyxgu5+jBkIoFJhHkjlX6+TE/vfrcBYBvQTH
lC+RowMnCbZs8EyFF3aGxYRTzFgpSKD5G0QBlP7Yz5BemXQG2zsMEVByJz80OgIq
GpRBHyhwuqqz1nZ4MP3aeGt39eT0XbGy4Y4XUmnE+QOpZ/16eKy8gA==
--pragma protect end_key_block
--pragma protect digest_block
ZrLM2u2eIXqltI/JrY2f1TTnR4E=
--pragma protect end_digest_block
--pragma protect data_block
0ekShtorLhdv2ONOrid0cV0KJ/3mT/UWSiXP1uB0/ics4Vl9oEb0sLgbi0w/ARhN
fF3F5DC0ACIAzJt7sqnRlauxSPSC29YZHqycW5VYaDCTTwbtjT1uGkjFLF/OW3GU
lf9BJhuk9zdMeZj4QDcyU/EbQ1J3XMCwCAi6+Lp8XvEInAcDCcpM4xmkm8ktr3ME
oZK2QJsr/ipIsSNZjjUpwzaoVdImSgA4LVHBJqOaP0N+u5PO/avyw5+VMcPCMy13
pYldM+tcWr0NVNlSn88Nkw3bFfUqZ9/juNgXy9HmNeD6SnwosRHCMbBUSZ2lGlRk
7Igx8b86uzlFJykjWXURC3dKGR4u1dhuPbG1jzhP2zI8vJyqPa15ZXMYiUYzwNNs
sOlnhL3mZFiBXM4Vx/o1Fv4PP7gKO56II7plZglaS/niVcbXVc4mYq7FpZVuu6vq
s9mV6jDZ/wAYn0e4jBCVuepBEccbKXuDf80dvtI1kyVItmM3mNHVvFA/Bdm15SF3
jfTjiMCHaxlxKqQpk5Nzxgr+Xd/cr0ULBw8Ltze5nl2Ea4sbQawgwv5Mj9s9ua22
AWeatKdna1MT6Z5e5KfnBXyi1pHyQTR8ShL7rlGFjSZu5o/OwbTJmQ5rEekmXOA5
MFsyYl1GkYqOWpAgJXdLkXt+QUZYIiEaqUVXJ6LFV7hO7DzOP0usPKOf/KnG9FYu
OupQQvixwdChfRphta+Z9J0OkTMbZoYdpRh6wFlRL/KplxUmNOL74h6J0IpLXkq7
rKpr38/DdUIwq4D2P8+bCLBU5/4ntXEXzTl5Lf1Ss8wXhskeyVBEAr2R86/kaQeU
Ull3cJ09/b8vQa/B6b4NdYq61ry1g2qnMBWlAZu3AMUa94A10FLYy6OxMgzLH0cm
CxeaokEKZkla98lB8817Hxvqkwcxtrkyb8ChvieO1SMcobAYu6faK2cfH6/HIzY2
XtSkw0y9D84DkeepoHIyuzcLlIiZx4oHHshq1/WJPvUG4y50UfkGLzrng2d8nO3R
wk299BDl5u9eAe4F7vc73WBxA8mSmMdI/yqs6FUgZG9Gz311oQXcxGXqdSNZl8Ur
VWhL/uYXzKDJ8ZaQTkteuZPBFQKileY8GhtjDNmqBOwN9ER52QeFvy/csRarXeRa
WlLnLE22wCxQbAImnRFVVOrUpkNqxvDpGtLnsS+fRpwqJiScrAGUqLtneW6mL+sm
VaNOVOS6Z4XE79t7eiYvRxPulronatCwy2NODFwsZhtm+xXk6NH0x14ii7gFyg6Z
Q9UTGgpQqNIsjx27FH4DsmUJELOo+iIiWPk+0U0I4dqbBF1tp3Fi/Q9JoUZp+YPZ
txpKdzc88oJOlSmnLTS7jyUGkaXKPFcqY17nZKGNVQ+02dgiSydhQh8/gDfGc51I
OnS0yJ4QBiFa+tLKnDlvmVMyqiPRTYv5njyCdzpZrBbfAJ2j7Iuoqk8bmkVZZbuN
Voj/gLvSiNSNz/gDMAAzfH/+7/Kqe2F2V/mFAFzRyGIQkdU/VtH4yXBJjrt9l+aW
Ko6B3awkh8QtIjoRcDMURYTbWY41puaPc79PCxrn+v6dH3JXzY0bhedpcmqTMFAY
HRBIMFUcgs9BGbiPHS+TuIJJuKPlUXBmvMxAGAjuAV5K2OUfQRz3Rb8DIoIzJ/eb
rPRA/6GvpwkethyVVTrWU2vuy5nPcNM0mxe2XpOyos7T7PxXRofxe5V2NdhWX7+a
ZXd1WKSDJ2iby0TZbUdKPYiaDrdKwXMHcRWssQyT/dP305B0kuMTXsWq5fA1jkA9
lloaZuwzmep2keIGEU6QAW5WVXP60qqFaLYO9OF7MNioDX2+QRQfOdnSBXEoQtH5
6KfQSKFBI26cGV+7g812lOH477DEVPFRezzLrWT9ssThjW8YGIBlM6v4uOBFWRmP
wc0SK3Ei07C4UPfDEeSplWNY/6KE5YcuR6eztkk6gsHQVQhcXcMLHoCwbL9gYLKg
JptvVrT05CZXwPQNFLccJgqaQGYxu7snNDJ1ZeMS/PlfnJWwa6hBZxgcQAVdlX26
Y7IweIO7TZt3Qe//LbhUHgc2XQE/u8vb/Dj6z0RxYqK4meosMxINNxiwHTWmUHCA
eHHou5UvAUjTMk13/2roQy0d0vcnlhZv0MA62fPhYDyurw1uCgy6g8JfXTZeWG9N
jGMDj0ILRHFoeaqrE0a5W9GTEW7YaF65ZiJ8ek1MF4nV/XyFmGcAz+mf4zWW6rLA
I7auKIaMe6iKN0BUHIzRvR1lWDtowCfRV/iUdu9+AmtVxEEXZHhwUbp1BGpTuXT0
benuPPy5wGzZvfVq/IiE0T/0gYjbIcvKUFfzGU7wluB39nCG2TMYXgM0P5VnQ8zp
eI5xV4AxWKr3McSCv4vVs9g3pkidNzisDHPhS7nxhvt4uSWFuoFdc9cLs/fWMl99
baKa+GSRHyz5EuDV3Ct2m90PIa/LZE0QbOUDiC5svvM9IoKll/1brpFAwUpG7w4t
CgMpw2IyQI2p0RfnbmmTyBVvPjMWRNM/yoxJzmC4umLPmcP6BrE9Q0xYnEUAYS4b
/pBu+H2YgzVk7MG42qT5IKtRNkCKo2ub/vvDfzEKbgyg9YwWnya0nTmgH1xXUVMF
X5adwUJL1b5+jUUvwL7gUu/UknjpFN1MMWrAQMfnRG0nHWi2Zakg9JInAslayc6W
zgSOtp6RdgpBDjDsOIX9FNae+0y2cs6hpmfEbLVAjkHUl6qkDIeTHMzZGSP9Xo8D
rban+xIg1i/fw5Py4PfGq9usKfayKzenibSfjqQgToFmJ2GAnnkIuPsW8Cnhzk4s
cjPShT//pIVdPGM1ilmM90EiP4ZVBI30xi6nOzV8lBwlIYDzf5utCIDf5DzCLIu7
TCxsKGSlcqLUudaxdeZIf9AIxbTnJT+nAeg0G25HUbVCpAslWoUoI0vhP+wJarRx
y94AC1oYmJGQMLBMArxxu0JCoJG4y3w7k02b+3XceMmxSEQMkFlmXkvwI4uuAwju
64puX3+SFxWDhb2ppNVHQDy9ytUIjqfq2821cnfxRDc2WzyOKX+Pi/IRu9RGfaBm
/Uo5v6+XVzNqWACD216ygb6NH073JC8kL7Nm6Fcm87xNOo9d3VPteI0vJJ79Rpw7
Rm8zSEHDzBl/vIA5+aaYGXPUVWnKnKBKLZfNYrv2lex4j0l5eKxwTtdmAxtklzio
YJ4tH8vMqlvVdCCSjwuZpm4nSkUKauH+ItLjgE1D/+rPzkzXRu6jjc5luG42fGTQ
O1Y1Jg1IL5ZNfclIH2aZh8OuVm9SDrkGJs7RcjoR/PRTlKvdhoXH1P1IwTlTuvUQ
/+wxVljbCVnfVX2OD37j9NP+yMmg070hnWe2aa01Spa2fGscEi611JzlTeApQlLw
pEta8HzJHsY9/RtRVztWtsU04H3Jd4kjxZlWq9wGaA+5F1H0rhbJJCh/80PiNIZS
J1dGMoM5a+RBMsnlro2TikFljU+kRzHVDx0HFh/tpjslPcrFi0F3qizHCNeDjgLF
UqkrJtxVUETYRIBdw/LNGHY1DA3zjoGmWcSClX9NNyzu99nKKmBA+rc7ULwbq+bj
oAp7YXFQyH2eU8GYj+IkCo7vBMsxusp2XdUJcLZ81xZKMJ1ibjBpIph5xePS/Lve
9Abll7t449N8VJ8lyupzcOLPDZJG1pr11u+/Ty2Wud6H/p8PCTqGlaXBnYjuGFf+
qmq+/edS00Xnwid+6EzV/VEgDkfx4fvOuOoruuYahY0nr0Djj7/JnzBmfDxJk7p2
TcSGc7zE1BBWaXLCitbo/GvyFPOSciw2RUZaYQrNm0JCHhFLEmP4oCOcK/uu6UDR
CYz4SYPpgAK7X0UsMOIzFRv0Z1JHd3dXTWNAoENWkEsL+eJumbekfHM26cJIowuD
Hv77O78NPhoo/fwV/p3cPB9F83E4TLRIEhJzRLRCDim85B4rGsg7zGaDJG97WK3/
XNmlwJWLiYBJhtPNfqSUKLTefHsv8VISQvrHuGVyfJcaXEGpGruCXHp0Kqo7J95v
Vc8kEVLDt9IlPAEH5i2vF1fqiAkebibud6kH6ST/XLwm5BjIglO0hbCPdvsl8UDG
KCwynYh2e5PY9qxIUOZ3q7GXVGCysuCQllvHygr1+rP+ixyCpRQJ5hPsLp4K4IS6
Pkvjv0jqxMnB0/NAVqrT/uf04SzmcX+Y61n6WttVY1B6RSSSAAlXsG6fI/PBQaz3
aX60IAmkVUy2AQDjM9a6KYvO2bwVhgc8gluPHFhQouHu2OZPR5kLzTAS10vHdzBo
98Svjas5mjiUHz5SoihkyjUeUPwz5CMl41LQPAxiSHwr3B0wGvIFubDMYhfX/ucF
KPLWgYGU9Un2kzSb8ikI7utBmJW4sj0LKJrhJDDTHWeW6eQ8Ktz4aNoX+M5Gs7lC
w/355yW8XBLqIjwT5c0e5BLbqiTNFY2n8HIszybZpTmhmGD6MOITPQUIdTQvVsiC
tllushT3eioNygG+8auhL8QaxijPwmZpfB+WFGet7iA57HtdLA5wJLi7+6qc8eLx
EQErsNcwa2jnk+seOCeUtkv0FBFnHMFUnIPUOI4yWMuEtdsjA2vz+NjJmvmtJ3rw
1UCpwZdroe0ZivZJtvMbcPIBJU8cDIr1EHtTyoaxxTd9PdtwQqp2F2FJYKG0XZDt
B1dTbxx3K/0kVlEcpaPPldIeUOlo40TLkaVYe5Hnj/fT1VFctX3MnZGSDZ+dx5yJ
bh4BScZfExAus2IRh0tMlR6H60MTRrIG3ppTDXqstj7advi/HNdwnMd556MQ82jK
jtXwbWvBWxz49JWE7sH47pEy1fnzUzbZa4hy+580ocQtP1sysiKaC3FmUaQmpnIY
wIFo5RdJsNrZtZ/zSW5Zdc0iBQ6gIqVSCSfVu4Wy2rtIi9+SmOpPCKRcVLOzNjUD
tCNqlh174JPm7fWPrVSo47ucFMD8Cn1CDakAouzVy3NmiCxJ150pc+wl5budR7bi
1Al+Aj/DtKim8Eo1B5Ub2vwFJTcc2UEChF0G/CBGnKkPmJ1kOHn3E1niA3XWkrhy
FXuTJoIdKXEInlYpO6a4T9308iZaq0ZetjKMCWcoaNeHCyHRvSeVwZpCVOS/T6lY
cSTuHIs9ccQV4cx6jJKkKDa08RWjm8HNwDrvfQ6me2J+B6q+fDqQSjse9MnDw4K5
1Jb+55QWYQceQE5oFhXFeODc7xmryh3i+iRUqGyX/46aMuUs+f9NmwpWgV4VzfrE
fnLhBJiW49MoEq8I6ahMy6ZsG9W+vvBBfWv04iAu+0+LexRZ21dnQCXrQ8n5u8PC
8m3xoEffK/VnuW2c1CyrqREZp96m3hACbOuIHV1HdMkJz8FD/4nmg34tJtH/40Oc
lDdeYgD269U/0HWmegrOrvr+WWCFxJvjM8U4Z61UHtK831+YuSvHoF6YBniv2nT1
k0yXM7nBFh0admBYnmLexR1pvOy77IV67x5kMAEoAWej2TMFFeRM488q4zEkjtrR
nR7yFnrAvZk1lF2rZPczeQcFkfYX/VEx/BaddArf4LdIQtsguAw/DJR84S/RFc0R
A4XwJeQmPl6xxtmn6E48SbkRZet8CVVs2k0uVY7TCAZ5eUXT9fudieA0iA8MB0Pu
635SnSeOLMULUh/ZY68QA3n/b6+7IriAgXtm0SJO34h1nUaXv7K6KUpbqoA8nNcN
8xLB4Jedv4G1XM5CzLzIak83Si9ANw9C01+ddaepDDXO6SoZWn7ygu7hWOi2mrVQ
k4KguS3YOtjQAqe8vrku3+o54wJOohCxMuL36AuUyIFnqogCtb+c35H7IBWm9N+6
pXHM7r3yJNDtiJwDzxVF0HRUb4vkoHZi8hA8BDkZv5zGWnKTdwcPHdxziulzzYSA
lEbJstTLp7SGfPrWYgZIq59dhs+TkkuQVPnjUL6lU/1dOVAxfTggCasCaNwG+cjq
4hUA5sZKpVt1FvdjEtEmn+XL9YULsK9kGredwalW+WKFfXYSdsfO8DRfEZMXeE4z
Ivpqc8Ia5kTY+9uV47TNd7xish4wguIA1YslBcNsVix+y47dzla4WzWl9tht6GBZ
+UUcwGxAfLbFvq1aqHbfcroKagjgzk/U4TC4Wxnzsl+qylpv/YN4JZEWzXSpq3Q4
dIYcyj0CLcgHBdYlJjnKahcvaWfssux0zF4iqbEPJ6Y2i9szgypH7rQ1gST14CgI
Mu7tJM43AMcJTfSBpL2XwnZq80fbuVija6v5MgVys45feYDRksQZXdiW3ewmVCX/
GHETq03sERUWpurWP1mHEcvKjssJDyLwV6luAULhrogr4CSWUFgUHmglA7d5jQY0
34m739Y894sLzpfwbNugTHKffe6WTevjMT+APMcd7wKSQg4IpvcTcjy6H8/pAoep
Ug66IZCgyHnh+pYphpGHvCzs4gogaowQIHfMKJ7+0lMrV2qNahL4wvraI7H4SrmP
yfbwZAApZ5m+/aRNGLb4mwumcwzWNvi25egm0p9csDc9Cc+cHJpnEQKkZJnTfI4z
RUJvC7LP+BQW5UaV7rg2aHhwLJnBMjrp+Dfzd0qMY65Nq0jnfcESNYgquI21MgJ6
ZDk/kDe2IKU6FeC6E1a0vhlguPrQnQGcf/vqBYzG5b7jtjwZpOoQzOdTCwu8E2ze
ON6O42b/CxSRl6+cT1NdHwdIjroANtF20SHqRHzTLh3rfd6NGufwGoTgdZQc2/GZ
QvClsruAeNBXhUcjWwc9N/MNeUIfwjSTKn4t4mxIA7p7eDPqa9toFdgrY6n80BM6
ZVbZ8FdyKcrarvR3cg+MHp+hzBeOdlnhDaAMJ1PbllaEiUYWUNT8cxeacb6uAK1G
C895h8x3c1ZWAPh1Fkq2Dtg2x0ru9/418/mtZU+N/NoUnMk+C3hP8e82ZDfYqvHT
MNoBGR8HkNkRjizrOXZrwUzvceg5vZ6svx3IcccgalDiYlKOkXzG76HLdqEDV08c
MSBfRWAkbXe3eSE8dQSjjGBDaAHnN1teTZxLuIPNQc38/9Kg9yZ+zu+IPutDlIit
uo22AEDD8MZzqbFH/Wp9NBD472OOUrtdd0/RvbXJm/CWdytkcjLBwZSMMHwVeQ/U
tQY1ekLmmqRf1yZdNWHycmvtQNOoW7Y9kw5uYxfPC6Unap+sunfEN2Y1j9p6/YAL
T536pOWJua4XpFcjsCdXFI5IbrBD9JuWqx9HP5b0snmTExqWyjeA02mJPwzmzh58
V4a+gLfkRxQspDBLzKqDMIEKhcYNI1WU0GFHjawhnjs17ONHRLYQkRsC+7iQ7U/z
J7EaMCcjWbifGZ7t122c1JkiP5pESNwtsg81RScuNRGMqqfnRvUd49PcZJQHy3Z2
kjnBl2oA2X+Zkvbuv9iVUIigqY/UJIEe97IWzA4SLRVCI/BwwdWzQICWfalKsMRT
VffK4xnSRjIbmZIlC8cWF0skyBcgVHP/SIsdBTZkUxPQG8XFIusxyBDU6YE5LPdU
7PUfzFXMbo3k+7sGzy5i2ohZ3XLjUZ1NJz9qVjfZyIdDYuxYz2U06B+4FquKcB8e
SUA54jbgGD2GwR+bV4WL3jmnTvAwiHKbXCJMsw4tVykTLKlHfLSOUxLG8Yg1M3PW
75skIoXaBCacRFuUXLmltWbI2OaL0FwMyh9Rjxo4cF02Meaz+kLQ+WOIWnBL4Pqk
fZ9iNvV8edTjj1GE72tHw3KVYe03wKhmiEEjCvdH8PFHTPCufhWajEIDcPdkrVeP
5BlL4qKmcYShrahCzHNeQ51ZwyOPV5xkWNNt55fNbcI0xv7qU8va7oTyruWcsn1T
U5jeVsPweOMKk6RjuwZSFVje1+6rS5MDLKuBrjegb684YzHZDGf2I75ZCTwRDVbE
yuru/C6Kp+nyUshCfZ4Xe/ps7sT/HKFwQVLzQ9VTA+DfpLB1U9QnLvncYkfkWw1y
RYVQk3bjtVEO9n1bIqJKDY1Tkzf6pHdFS15FsSXtcf/cO98gcSjfuwe6Gs8oAjaQ
klx9z3rAkCeS2Qn0hnHKCBFysYeeuHy+yDkQoWiK5TMIGqAtyUhFRkFfzPcTiow7
UIVLSfXlOzwwD3LBkg25eYERf0yXuJ6w2LBLlgnYe4R+ex8VS8Xaoukf2Xx3kzHU
40e+SM9K3bAc55v8xKhtQ15q8I5X41UTEy22n3rYc/TyLKJ5OIXgjXFsgVtJN5x+
5wr0LHBRHrD6WICfu0AaTKwI/Z6xqbolzrXS7GyHYeufvidaAov2JmHK51+pE+7L
6UoKxzGaW0x9CIAg06IrfShb/PzjVDvuGrhECQhbC0zOnTtenQhO95V+3Azbbs3f
/KSk1kgdIAYkmGtgJNHpBYSVh5o5iiK1V0OaVDBU1rK9V/MQ1kH0DskvlnlI3dkC
nmMZLne4p8QRJI33P9h+USW6JuIpEgBNb14J9XIe+vvNuxA/AXFTDnKZmXkEIIgm
plbVjs8tTvJXcxpBjYroI0+gof7KhrrA+BAKx4ya/OVZXNf8WecwCA08TpDzG28N
EwCgTkNSUMCWwOUIQ6qSeKqY67iBndR+8mQ7jlxpgkug60qI42fZhqPZs2phOYkg
FegOaz3Cbtmj4i2pek7ZKNda9I1ng0V+SZmlnyt3XsU46AdrH8bsHoz3zWT9Qyjp
uQr4KRFvSwrqMzoTp05M9f66K3VxH/x5QWr3n8A0jtzHgWDq2Hm5vx6+FBJGpFZI
n6fOb1IknOhanxSMx+KdzYfSfxyA5XHz4mKT/mgbQ5nqG2YRV/rG8X0iBNu4MZLh
mGA4O8JxaJT5K+8k7oLA7QqtTNzjw+ngpHsEv1O/OPp4djtzblSFNw+VvEMY4nGp
ViodqG6h8PKvhoZWOELfGpLAWk/sSI5hF1lzOgorOKU6rPsvfpX/YXSB89/y2xX+
cxgxMdW7zxFZlsJIQ1MYmfhbcUQg9iJYiC+p/bEutCDi/uMeNai5ooi7V8sWzMWJ
pAn+XANQlc1jN7B4k63O1tmNfwW+2IyoHgDJHVnhylE4HpJ3GKz5CiLT9IddVCpv
PPF55FzjBkPojrmsPMGiGD/LricXoBjplXunapWAnfszk7RaleM/i5W4vPWB+FD9
zHAqg7ChWkj42DAMY5Q73KEPQU1zSSid/iSfg8YSzqFgTtrSQDcnRm8DwNO2EfaN
zpv2k8ARzlEtAKwdpbwt3CtFrZiyjFzz1nU8I/sXri9jI/qwRofgMuaf9Hw+J2GZ
tCU+qljQwx/bmQiDXObP1lkjgX2/PRMWE8LCzzqkaNKY4qU+kq15loTp1PF0JYXU
u/cPiLyUg4hc5zMkTkj05RU6ze1vY5F7A+XeJ9XJMq0tK4J8omoiG5tMjkHC93dQ
JcEChZ7tT7NTtDjQJNN4AT/6l1rOJdTWF+7gaHeOCHjsS69kjWxg3aa9rHsOF7AQ
Vr7uVTsbojTs4h176zKQmvCnnWUjY29Seo/4f/7u5IIaFmwZLYIBcwAG53xJrLMd
qm6CcuV7G+/OESZ+hH6tYCn0fNvEG+EFq6fbhIlEfreiKPha8P4/2CmTQbnN4LwO
McGvM9jrnu7JWzJxgPYPLabN3ODeA2kloZEjKuJaOTgPn8Uf+BBhzRZCEJbhZa5Y
TVAMgI+0QEiA4K3yW3sJkPaQvhBHrKKwMhXPZGHA5cX57RbmxwUKoErIGJ5EMx86
BV+ccImjA6KQ26SEbh7UJGGUf4tmgIvnstjD7G2rA6hq+41/m05giTEUE9FnfEz5
Ti+SkHYLmd89voWJPJATemXTyALRa6B5cBeOi2ThaS+hUgYkgSd+7P8dqadl/jlX
MzXoAdGMK1jU3W27Zl2NeTFxLMs/a4RhoeoY/A7AFB7kviVPnbXm6c6i+bjoY53/
66tOK/9jVixDQIT9gaVzljTdojUsxR41dqK4QQ5DW9VwxVuolcqAYiMLOZcYeYou
JiM0+wJBpy7ql4kobw1xuS3RwhTjrjkgQ5/JiDB9GJ2hIAvh7xWJCZaEuVjOFcXM
SspQMRNfCkvfcE6uo8c1fKUcKsr3gcnkzllcRJuajFDEE8UDWFSqrUHr9cCi+aaf
OoM5S+aNxHV+bBf0wwtDI6/fews8H3R2BiAeMMvOY6ehwOYjHTKbVAAyLrJ+AQmG
NkY55aRFjcQ6RAyCvULDrBsTvmhK1ydXANZpdJicgyPQAsoHBjNQaiZxU9idP9MQ
M6IZkiZHrVOZg+EBgW6tiXf1axFNEAcosRPiAPiOKRXXR4PknoElHY1cZ7CeUkQ8
0zWGftxDN9LAwdu2KF3VGPyB0OP1a3PqbOlda76qUC773FjUua7Sa/6W5HF2NHgU
0bdtf82VYX7zF7JpiRrood/sCO53c+fXaKELSiqpE+YLIL9dKdLGa22LDzLqo2U2
/mHAN6+wyADecLXRhuyb+CrOObTBW+8w0E4MvweSfnWB/f07rUSzPpC1fv1NJE68
PQW/xI995bF2sDetFhX6tiSljkTxoazzafYIJTqmM7P7bvJh6jKTlJcH00FYG4lp
MVAbwzYtef5UtKz0o9FtFQI0BkqmU0UFtG0Lp8SIgfeJEobK9b3eqbG78bxcNJcf
Dlgdvbf9Of2U/plzMukDGDU0r4C0E5CNgNN9DyjpGgfvtvn3kkP7P0xFWcjCRI2T
HxaDARoc5hD1HJlbqkIv3S+odoGbOoJYI2W3GupmmoNNQMTfFhOprXzcogYONBip
LY25jbxX/HfGWitIEZaZDA4ZrETbjaSI2P4iRvwOM79o6RNDLwP+YQls9Q1V9y/0
eFu55JO6jnZV1RScml2FOnaATeF/V+/vP/o/J5u8/5tgM9omHBja07dFxTHwqO0j
rGYx7+7OdlRND+DYgID9u9tXrboPal2YmR2HVjtQ4lhjvTWmzmqMzxezgSLhbHQs
ewdEXyHwoEG6e1FJaQaoaQUtDZPqtIRGYN7K/rSm5NQ11RE7HwsrGJRD5UW9Yoj+
x2seg+CPrQZJgNrUw8iYHSw1FuMLI6dEPhWiBiy9z0BIBBURE6fjlEUjFRVLGrJY
5SKtAaVuYgOfxhpZQMIVHHSDd/gEw/whxeiSlKthE7UkLgaAvQlMhHlIDm82RKl1
v6b5qvbak+VdtNysWTYC3hSTZhlTjmZaBkTu15wLVrYkb4CiS8jpKzRQ2wubxHec
AQEfLVBHWmJ7xYA15LD9HiwIVuLr/rdGN9U7eJUvUMxIsPFJdmFYTV3V8nS34Cy1
ktM30kBzIpYnWtXl7s5l5JCLjHkaPSVhD03KT6pAvj5EvwBUFxnFV095JnRXZlCQ
uKyWrB96z6LjKRAEbfmheYlE2Lia8wmwAoLqKCeWtWg+rRNwxa5j5E1l/A29LsHg
VlikstZIHcr8rbQu+HJifnKGTWBB7bvZc1678tN5c8GNFtfBurEbbF/wFxvs2rBj
cCIrX6RI184bHu7VUlthJnjsDMLTE+Nz8r5S1bAyHP9m8QVNHxj5xERBiIatSMo9
uw/ZbLKggRuwivnYkP7Pxsnn//+lAy0rFGLcb58bS5nDktij8yPaFFZXTuj7mjws
caLMbNCb6S+/kK5aQKIsC6iZdqtMKH0QpibRwQXKMYY+qSrLeRtSEvxlpFy7Mnb2
3YnXxnuCBhI+FZDDD6xQ5caOURAiw8XK79qm2ti6WODtnVOLRZ5Az6WptotZPakA
AL/pSA3Yb0jgYWmEpUaq81RnKYHuw6+G9nvSOsnyXGhKHRQIZywgDW4Cy9srJZ2X
rwFlGDmk+i3AAaWSG7WEi1ZIxegMO/uRN6ZxBUqibUJ9KiwVyKWLjSgmQB4nM7mo
GfZjnkmjmG47ZC6+DKOWW05o/9bApJ7GwJ1esrB5JC+/IXehNp9yrIMBMyNeJpcp
5SRysuXAyIsFwXh5fnW2Y8lvDL4cb84nekn1T3eqOgHg+gIyzXu+Mb9MtwKBmW1A
Brjx1yWe8ZPcizsYMcFe4njCWgH7Bc3fQZbmI8UI1twsWhTalH7693QJi/crGzQx
LNF9033jPC60pMg5CtoCOf77peGR1gNX5ns3JYgVPO5PM74jDedEuKb3APHCW+8t
0rkbmd6GRuXpiVGbz9p3zVBq0wXSNXwIGy4Rq4fM8YllS4GWPkfZCaVVooNVzJMA
/fapxPUgzf2At17GV6jTnp1fdwQ2Gn7P+U9uBZYvBLYvL9mSW8EOc++ZqShNjJt1
CdMPeQCMRHseRhKh11Tn+2A8ncZbhxcnPPMJsPnMA3iKXjw01lTstmGXgCbnQy9w
cpINOoFG/8xzjLpvfLJEX2vEKgTMaRU1zV46yfTJXVAyTHSJj99Z8yBbyadvr3tl
5KaynCrxCfEyYdz8z7fJAwbUMUxY1aOy7dZeCbonHBclYU5DK7/RG2YP7J8JbBax
jTHDrv6DsREil/H+j2Ie4HDxGB+7SIkGh9AYP2QaGU/PGeZodSwIA0W2V2nfM9cw
JLh653a3yRqMrracqTGIYwQxjHlJbgyyVTkytOAq2yCkYXmAvkNEAkYgBJtEPsqt
SwtxZx2p0RfQ1h8cs0NpJSLVO8xE4HHv0HnfFvr08srz+aWJEtaNMU9yqOVwv1V0
8/sJJBSti8yhCImZjjpKQvJ3OAdL9M5qgL+fY5FAqrwhH47DlzZ/jECDxszAjx66
idIaDtWR2QGYRvyPG13gABCnEGblhho3ZyCoBbG7TuFXl/2sVPu9ol8+dTcnktuX
VA1bYbtl7AWuByOuSO5o2F78PsZru3+IbyDOUd20QIbmiVrmjp2sgMY4H3w3BZRe
3JAV2ju1qDOeq+acRsD7+7qQt6a3oicB8eDZzt0m8muO+qqvZZ0xtsp1I90YiygX
oHjNolnMD1TNiK7RarP5KVw2B+PRvt2I/cU4QkAiDD+FfuWu3LFeD0T8hPBcQcIW
qyooX/jwebVvrgJXQNGx9g70xCpXYNCE6h9AiBQbEetri8jFOL/xkGLYTt0H4vy+
bsWfxIWkptL0f2AnzHUd/e9giaCx6FRdinmrrvWLG2FLKoq2JmY1SyoT1BRHclCC
6OM7xTIMwvkiDDiN1dJWfxS3HNOXL2SZ0IuyNKVRB3b7XDkB3EhGVQQRtrU/Zejj
BXPnCybunv9N0umKKvbrtJyswa0W3JWtqdmTX3lUHUh324Tfh0W6os4w1swRJHOl
5LxaPSxl5nVimz0TNlerhtTyUsO7W8pSO7ATVhwJd6vn1TQNNDBDzW3551vagf8O
Wdrh7WshaLDIkSQHVOVeTzkGZg/ma6PRGowu383lCNzp9jFcx4OfFNY4Za5tNWid
wAyfD4i2E1hNp5mQAIxnofySnw7gPjmXovFWtaDsxsP3Vh3HrbVvdxu2soPz8FYO
fIjgXn04hfXuZ960BeTMrr3lISv76QU3lgkCNhLSDk9nB4D/kLJfZtyuvVJccWxw
L0GgsYhL+xRQoGLSpAt3DNe5+Uhkp+YFaNwSlN3Ge6EIRjgZfKxZup5TKKHOHtk8
p2VOdZD0QeZTufBVd0q288/tsLDhxObWwivvphKOxp8XZVjkRxYlj8gjJSK/BjFI
2jy1esoeuq/adPGwoXDmhgNvUCfpQp0Q8i3QEE/g0RtlaVA7gca20Hxo2A2ILubq
Vix8BE/tWHTdpQ9BxS39AUlwVrlQbX+8gVIZ5Qynqlq9F13tse1tqviMGsTS9ZKR
7E/3yHCHJI1AngWhQeXg1eMt7pkLHuCZA5TVNhAoCE+zAJE5XRDG9xlsbSq7Kr9c
JDBKB9HKT7EFTeTWNiYIZ6S3jKfeROUlzE9qLsp8/vAlBLdP2JXd1zJ9HOaesDt3
FGf/EyPUoNK4nFxX2ei6litU5sc7y6Xoorm0XMiUjewEIFAbIwsgqP31Yec6oZvs
EwICatVOXJLki7TLIHGzCPaxlmRemUzQ0ExA5LM8d+EMQKFSVEUZ+ADJBLlxB0B3
EjqA0jT7GcJhlRB+2PgE5vECmrQvdfEboWFCw0NVxd7mWD62YdmJhVOdeSTGYJwB
Uw33AXAPFS+UgI+UQGHn0amvPVZKMKjY4h2QdSA1vksH69unEiGE4iWXCyi6jQBn
7jT0VslclqjwzG6FSd0X8tX1K1C/Ss4Mvun0XZDmf2qm0fXZbkcR7TxbyTr8cdWD
DcVh+9ibn1O+m9gXfhoqiDoqu45lE8uucawDl1tcv1jIpw/9/iZgGeCA/41vNxFB
/gXTIgxcx6iinW1CHT23OFfr2EI5QEy7DCD7beRMEX1IatiEcwgEz7jL2oXAC1qO
CxsaWtvIo69QJ1fL91oK996zaQuNNXwISLrq0/i6uTF7SbBSD6KYaN1H9FYkAfCh
ZfKC7NtPSMa7MKCuR2WQlQjpLaNvbN83Tb/tjH2nkMtIDO0jSfPUFWemZY7S4Z8Y
QX3BwKSXpbWle+HEEGJnOR596Jqey6Bouc3pCEW9Ya0YeMtGVPNBWMJBoQfwxtM6
2C8JOQdlBW8tiGJnfhQn+xcoHk3+zb0Yg8mgVcC2qNXjjmCA+WuafOPtrsdBkX63
5PTDls34ljMroaSgo/fjfP0YdPuOWiVpjIzNWzUPDajIPN0406XDjl3fIzpWk1We
ucBRAOpCxonQip0umnpxUujAFV0USt05IwQYGep3MlgQTs1Wa561c7irzsA3fncG
ggUe/WMwU/ZSwBLECLfFp2RQyfV6gPm9D7M4ggU9TFfYGvPHYXwqKFijcDXXvVCa
B/bHsxZo9uKkS8aaYyaBTqKejrXUOqaRFm6O/Ri1ChyESl3S4f6kbdG7+A/xSHns
Q3c3IVxGN7Fvsd4lHu/SzDXokVDsLoOoHQ6IsRlB10UJtow9P6WCjGmPvdRWK19w
jzSbHb5Q44E3N+DHoo+jg+vnTWxgSTnyIyYtb6jTVFziibFTU95v6Q4EcligYFT2
OaH2eckxgG4KpWH24SGH446k1K/fuvU9f93z8M3icj/uqh9xJy9/VFmdpSoiLfB3
+LNd/j0WlqCPpQXGwfoyWJrIkZ8d4HH8UyhiTiJPM/b4zQNgnq5q7M86deBrIrvk
SplSoOakJwrX+qfjKBfmluPEDquYl8HhEQdAF38hOuIubXUBMG8vElLzS8OggWiJ
5vvur07eCNR9kCdym03mkbJeq/vtA9Si8Hxd+xTzDJ14VHU+w4ouu4RziLVeexm0
L3aS8jp3gxa/pVivG77ZtiXNt1QtX9+cNZLklbD/GhXBxD+nVsysi+mcs1zKxf7j
TEIT1qPHm5tw9SnkpBdTBKUL2FlUcIB9CNMYfwcaN3oBid6l9GY+I9GGx8EVWcVm
Ihch1Egy5/PWrLk9WYWUKaWwL4oM+SSX4UYGPEpHAGYjogKBsDh8Xezb83/qVYR7
kWGwN6/w5Z7grHPyHl0rwzzXCMALc0VIu/Yna8WPTJUrPaa0+UI9ctEiwG4foz06
/MYesrDefOhkU298R5Fr4y7G6QU6+4OZ+xeNm39r4VD4lm9rYpkIq+u9GMRj4T7s
eG6oVv+lBhdufj7XCFzxl6YZ5hywqdEN1Ix4x7QhZLYON3rsvPKzjQNad1pf2g2s
eOH5XFushTxTLdfW2b3vXTDuaBeSbhV4mD3M7WbMG8dEgc9i+0vfyqqZd9BcsKNu
NLktyNyS9+Y6xvVZGBqjxqDVYl7j8e1OQ1zeDR4GftBnVmLXCmywd8wB06t2dTEv
DpDa9wU4BT+/QBK72t1CEL71pgHR/3Ou3RhCJeigxD514HAUV4WXYXrY6mfT3gZ1
r0o7i3STvb/6XI0QrcMzVeOJ7xGRpqintgq1/jPLXUDhz2lAhQ9RuAKgkJxqU+Ra
xcNLybzdQY8hltXNX5rVPZtrhP3BNl7TJIz6X4EJFZBbRbyuqBZK4NNpemGMruZG
hDFVqkTVOYTCjiFLQaGKxrzg9xeiok+qOaUmfmXwJJVTVTYUP3Pz/Cnn6xFmLkMW
xCV+5zVYqgwSl6a/vhsZwogMynuEuTSwdhQ0yM8ZSVamTH55S0cs8bgupX9rdtEU
DQdYZdfaIzrXwaW6Kkl8rKddP7VPK7pUaTVqtSUJoh0uzQcwSiqt8qpFR5K8svQ1
Y6dhK3Is2JFRQZmlVneoN8pHtyYlpG2IjxLW/Xq1qZSfTszkeC2NIIANlASA4jUw
DyQlUFzYEX4I0H+/Jr1E3dBsEsPTVuLUeALPmn+T16sME6FGBS3tfhGgvmdYwjVN
Nx3EJZccdrGj2qM00WLGgrVmvrikP71mKrVsftshjLySJKyXDqxXixvxacRsMDV9
SMEMVLxD2DqcBwUWUV0P9mUNhCitIkvzk51LshSdjdJ/OdFC+yUomoig/rYX4ABm
T5EQsddv18bEf97DsM1dshaBYTjwJhuJRgEWRZB9OoZVE+S8CbD4dzHs2FghZcHh
TbAzx7qJqAzn+1K6JfbhEyTkwFNaM5oKYiZU1U3WNsBJBBPaT8+js6V0PN0f+xJR
UdP0ZgiBv1Z6L5kegwLpXNuNLo8oRF9blY4qz2TRgo8lMC/GjjxC1Pt5f0J+urcD
6h6vSB6tl6pha38T7s66/BfdxBrY/vN25I9S+v151N3yQZwV5bTIxvUwRygYAcUG
lJmxL8ErOtrFxcf+kVb4/yDEQkWNMlVMOPWD6bYlNTF17X+d08TJ60tMIaAYTm1B
jdfkhJI6C25rs7uLXrm++dgUUIr36cGNqkbTjFYxIb9Scq4kwz0yaupbZaawaXKP
RluJAnGMbn9bp19RH47ES52f+CsnNCq9XEKhxZSh6qKlx2yyFh5fP9KPEECGcT1k
4Nxo2NU0X6KDs43+OGA4UAzhARKD0KYOEz7eNRGgqfnHMwlEQUjC7eG5Ad1l7uQS
7MFmvWV8avUfSHl6GoSW5vBu1sDG77XQh/NcXsOEf4qgYX3NqwrbRyj9Ffu6vTss
hokZTdM3aCoG2a9y86uP8nOBRXuoeLkmav+Vy14QhyYfRb7Lvhb8oBSATLhJdQV1
p+B3LrMruQqFaxzqCqJGzvQCXb9po3e6RNNkpIeyRBtjWpN83FPACK1YvEPTh4DI
NQISzhRHE8haAI5RXH+VDkJKzUTq46NoJAAWbccOHa0Zl9GgQWmUid/jw2p0Y32y
K4uo+1Gmsu/+Q83l3zrupYRc6ygsXR5X8pv9s+n7jnSXiMIy1HRzT90h5DsR3wpv
Z8hvPvT1Q8saQhR4DgNrolJTkYSjGPz0WNhlO12nAEHej2beJztAGfobBGZhoOAy
tvkMZtAG/v6PpcpS6On7Ca7Ph/KT3f9MgBH+cMdoPqrw8RberrOVNxJ85Vnj2u9v
ZngnzFgVmOZZ6eRvgMuAM4oa3Pdp6gJSSWGFM8kP6ZSYp/AJhhnnC+DPWPa9Q01u
GsXmbaURjiujL+ZadseduzL++GZQaL97yjJv730ZYHdq96Xqyj27ZpEZY04e8n96
tuunOBIunOOLi21GD5LcyrL75sUlrbsVDtpBvCUqZKSWwl9t7ea7tPOe3uAqBp4g
rs9Nx/5KEFC2mAvxME5RkWFj89IlnLarDEkK9T1YrWHidN+f6pVIoKYaBwfjIxg0
4/zQsimE8SKJ+w7Aqvhq+QGoZtzQQgHDbYmYY/9th0kflagnL946E5kkSchS9LHn
ZEUWDmWambG7JQoik4A8W8bM+1phgxjvzVEVKvDNVHyOMBEg7MBOHOLyK3COT01m
vowXHtdKm4qA851wE5CQB+5HnxcE3HvpZTkrEfc5Ivn6PTA8uk8cVTGylLcn6aA3
KqZEn1qKtZI7GpiJdopfmBJioobohxzTQsdRAMHQAn7pAbtl0tk5UXr9CfQ9hMnL
2rxvhvyNxOeqNHoo/F4cISSrDTOuqiQzl1PoS+F7VKzx4GiNHBWdSFOTFIh/0hMv
3iSJqAGLarGIWXNf5+pys4ngcpyn/zS18gRArgVwNndMK2Vn4D8aVK717EvVwGtK
docaL83Chf9rZnzG3RF1bceUln2McibQJtpUKPE5DUgD6rRoj4ee7b+JnMJFNc6k
RTWUQwdbxkJYvwjjbToQSyxFUV5yxliBIuNbTeQvZ33puZD52MX/VnIff4CmYOlg
gFBar3CQg7Y4zSflzzxE5QNf4avLApZJ+5EZRpLjpLiRbRTr/jGOS7mQBh27Jgge
uD9hU+jg0p9LrBElQUOUNAzURLtRvUVNd1/WG/ZLGi8+mrV5w0koSaghem+1Zk4e
lDrQ4BO3jlskKTG7ihzpyK/4Qw7jYABeyQSgnHy6smBj+cW6QlfexSveiPcbyDoP
96Dxu4jLlujweLIIhw+CmZiEVDg8yNE+X/sewjQvsuU/R64StSX1lq4PHkKRKXbe
aI8DtPzdTaq/Om4nMaWB8QP+IYp4Q+ndC5k+mfuY9FnUUN2oKAC2Dutlr2v+DH+X
5RZY7d/vYqUqUAFh+qnMTgZgRD4uoD8v05o8OlnfUN+78mj5Jc5Tv61Vy2RirPVS
purVXV5LL7UeVlHxGH7jWLfbHdGZqwl2Ht/Fi27O/JtRKD6/2T/j/swkzCjY9yF1
ce9gQJ76yzN/wirMLULmr9teEIZrwDPWGWDznHHnXikx81fBYWniPE9s2G+9UZUq
6N48/cZdNAQjSHBCxLQG/MRpbjV4y0o1ZADfTiu+bgMLVa1e00CLAQfEuvTIhapp
ECnTPot9bqdezvj+DFN4FFFv1xt0396AAS+3+GxGNu5uofZUP5o19c/ArqXMzSjR
iDVydZ3WO/n8nB4a9/gBLGYSMoOrdI1nEs0E8upd5NgWM6WE+5jHiaOlMakbcVeq
0nfZ6hLqsCKiB3dNBakYle/Q2ps5G+uqZLyXt8lhojejLEbved74H+yk5ew82Qtd
+Xb+VVFYU5SpP+9p27N4ljTZCJsKu36aTtZ+P8mZi26gTQU5TMgoMzLxEsgSo2An
2TTbsKgrMyGrTP64cdQvBRL4l7gwpPOtaNzeRfImybKJvRgCR1w3YlJpDtMtd27R
K2RuDuCbL/JS0VMAcb7qRxV6BbIq1tavGkHClDAzAIezIai5xg9/CmOpJYzhAwhy
pWgEww8nP87vvyDb39ksoKmG3+hrm45ZLs5oK9fPXzClvkSVXqPb4d93o75AEiO2
ZFKa9kp2U2alNE+Cn0rl7ftwVbB1X0bqQ5Cdo03QW2TOce7XmUCgJfARbwJSRTPn
6G/nQ4HalY2exEclYXQUH4C6uNDbvvlkudvfYXA34LYy3VwY80wogisV5dV5woYz
Y3Go6/VeyskdjpSmP6/go0e4i7aEdgqcF7WiyohPNPmLo8MDUOGam5CQvhT4VjeZ
oMl++M3vaAbA4sQGWhJn8iCF7lbvNcIlR75k+YzNHAXxXkbmrPkJdvtDQK3WWeXp
tCJ/qblpU/7nVqscfNGm4Oqb745pngaxaqVM90EVnSn/RqhSLrTdBEx/yRr0gR1o
5c61b5jdF4aa63irzdYwivEYeyk4yqJRdQsbpeDG2zjhpmFLDpONxLkBk5NsD4N3
nEs5lEwC5gK67fjxIY7m9rs980+G6CXR6+LEgvaf0s/NrtI/92oQgqqWxNBpUQvT
SbTAlRU7xevr9SbgJTaeSzfjqts7VmHyC5V1BrwuDmjeYGFBtKZPTp6GWbPquZHr
sxoGsRuZK18pfCnQK+bL52OIzKSMo3d1DusAqhKwml9mXZ5C/0Z8VUwS/QFskT1x
iF24+FsrBQ3pQzc0VLrxoB4jDY3CFi0jOPW17dLNRzK0RpkfLA9f3pnfQlhwyDRR
+4dfrsy3HIYowB9zivG1eQFe3NhIYocKKLauF+Or57IF/IrL5uVEY7tZowq/2xWw
dDvSXmSbTgwyrS9VAYwFdjFdQXJuTm9QFnUnLtouRIWbfYXuas4nJvIYoMsIOEpy
OIXoHNSpOsfI/zVF1V0aPKo4jltgwumgZDE8KHTuY0DJSBBosuJV9J6MnLrocSOG
IB+rcJwYNLBbPgGnIilvfVctANXnNvNPcEwzpGUJST8Zq7niwlcKMZxpOqJABCoO
InABe2aAdideomK26AfHs1ksjUsX3x6HPxt+q2JSLK+d3RUuwVedaXibqTRn3Xpg
ONOokHePsfjgs4YOmclq0lOU8K4HgDq6MfF8eOvq7BeVUa/PtAlnyOq4jlvqbUjm
TOjh2SdCCV0lR7saDNi+bVqvMEE5SMLSKpyZ2ziWOPhoiANLlPvrWCbOiUrL87oV
EBjBe3Sl/URwUSo0/9OmiU6xQOtuxfV9y+O6nahkKR+j80P9Lm7skHQQw6sFQn/7
dtXHD++5x8kEb1OpNXEldaQYoY2CxL9RPpYfnp8E3Lk+uX8tG3ZLjq5ofS5KGzU2
vz2AkPReFRN3ZljPag3Mhkm84xhRXesEgjGnwLxBzi2aD+nVzGt+YpspaVIYgbkP
6nNbE1XJGVi2i9yw/DrNTv8h18cPPqsV4DGmaSdKk/lmF72KmjUdkjoUamm72BsW
SWfyrCNU1OmRi0AzvaQHO6THphLGlc2EEn7D9rVVY3EFBu8wca3fVp4Kmt4jKFdv
li7KADdS8xb89iseDIR9uahjTCBIsgcCIaH8Rj47Ihamzm35P+xYUCGG+S+efwYV
JEFtT0kikKM3n4HVYExBx6cqJ0IzIQ4N5r5vQcowc5lfA++EdHFYcVv2r0OgIDPq
Jwb/GS85oUKtjTR4R08VYg1gmuvKcmkQ1CqOvrDnN7XNo3l9Cx/4wUr5zPCpQjWG
4m3xyNpW0yhqg8coW8zAvZtn6GkIWZaycf4MJZDXy9+SrNXYlKVYRhJGas4pGuNL
ppdCviw0U4CdUL2u2mHnITZqTHbMvqJLwXCJ/gmFqXT8YZAUKBkRv76J5byB1Le+
X4EC0ZDjQqfsgGmmDLfNsyNhtBkS7MKMrMX8RrnLhwaByNs0VtKZsbLYxpftbIaL
pYfVM6isqrNovCeQJJjhnPep9+80MZHyc93lDXASW5Fjw3zQdzBrVBCN05qNSDSh
1YDezdL61JeBNiX0shbUW710gvf4P89jAUBPyLFuu2V3VOkp6sBW4U2TN92yRo0W
K3yPnppQDj9FhHhP1ABrfOICN1V/+dMbKhMXKnczc5jVhw57WmUAbpmhADpgSP8e
KoTMhTPez+mQkjWfaOaJnOHV9yoNrLbtGHuVcF6Kh9E7S8gMyTKJBeQK+ZD6xMkk
HLWRgyUnwoT7r59KzGRKtX9HBzgy6aO22Htii6wW+y5Ele+dJb+tG99jt8QWDxlj
7BbqBP23Dwtcs5Hl/2QBPokd2qScCTWlgwW2AiOuWUjDbRgC1kdUsMA5QJOXLGNT
zhnN2VSUkBpbfwoF06K88eiLZbQ4+210qToX2eaVtqViue4QMr3fNJAk/HiB20p/
NfPGM8103ufNtCHXF789sBhQ9SmwWIAbVZdENFL5QQUNJEQ8W6wrGa+epWRM2H02
xVX/vWOIP8rPjFb72U/Af+uXGFNQnxqtTjhA4BrWtpt7ncO4e/w24/ZHtjUilynE
gTOL+maRqoDN7XCBa2PpAauZr2n4rs6KrOAwyQnHPDMOdSSOwBlegGa2z2q5sbQf
n0mCs9+r+G4UidfS4L4NgIIO63jAb5UlbPb6b0Rd2UbMgvoA6193ZMnl0XpHIHfX
WU39wYIJ+Kj0yobBTW3Z5R8HOOSAmXD0XYbv2CpQf7yF6ejSF6A6LipkgjDlzOPl
4MKwjBKGrtdluaguR1Co9S8Rhf7KlcC+X8jkCJc5ncNW3pfcKVoi2Iv88RSW8vDE
ipzPvggfIQoscoRaGh9T69b2PT9YkXTtsl1qf63rqVYG2STPPCfscZbGFkPOYOj7
HwU2+ydDjTbFPXYJb7Kv45D2ZrnuBr/rAY4Z4bfFNoqObYiZAMkT/mo7rijuVI2x
sThQmXLmh++vsPYYgUdJSN5k9Zs6AK1qj9CEuJJc/KNt5onbh747iuYPGoFIMTf1
fU3lVrBNMaVUm2DgoVjGn9jPDGsPW+8jIPUiXzyhUUrSNNCQ/GrDff2BOuIiIDGO
tmSNxX0Jm9vEgrj1hSIjSaGgJyfaiAeDuAJZ5rt+G8T8+V0AhVYlFyobKsd7G/FF
8KttUwKZMIHSVtD6Rm/MGSNFVWlPKB1UnVkqEs0uV9gwxWEZZkSOEVNX4tw5xrho
nteiRrMkiiErlVek22sMPfVuiOqlv3VIJDqG4IUR6vReRr7ShlbveWPcHio2xG3Y
4F9rJQnpyA7IKIxxHeJ6Otz3BE8aysOrVUsMCP7N9r/C6GkBxQwn3rT4AwO9UpTJ
nCT5GeJAIO6ngwqrkbSHE6SWP1RgeJIY21LYdVnEReizlUB0AH1FODrJSlAijAwk
BetxgatR600OWqtv0NIcKrpIQmN90jXDEyej0BcIZxuR+9F6B5cNdGH6f4n7/FNf
fIpQmR60KVL+neOtifbPH7tdRB28OoQMwzSqK/QPF+sRdROQCSC1Ml6SBDc0yTmt
Sje25pxiJFxSK86TRs/jja1ZBxhXSjOVqAXj6C5EwN/fHxfyF2pblmYABEi7rRc7
e4pdewQEDzVYVdItqdRdr3sF6fcWTCJuhI2UBRF4eBPr64TZmS2SSRCI6606jcnu
W7xJIjlylR2PddKemcGfWd1FJlEmEPdHdbLkVIE8T5AoGoSFoB8DadnZ9KLui0at
/yUMm0DZVxgPmdSortziDDdjrThjliqZplKz97I0qsYGaFMcLFG7sXeYyS8lMLdL
FtMeiKPgNbfQ1bvm18bxuJw1+c/ho2A/rEoXKy7ZrTKNdsMSYTcz/OiLXeJW1FWU
s9gcWbxTC4OjtmKnQowZ9AOW9OF1OWfRE75WeWtR9t/0IV4cCKVby8JJuy7v+/4s
rD8JJIBSxJOU1W4hGbq9jjI6HbzG+fjsJ24wF1ZL8Igis8FksCW9VLqLnKJttBp2
mI2dpjwjgQpPH106jqtb8WJP6Uk505JRIlrQVFjcIw/U2FBJE/mzNbpxOQU4wpCq
uyTnpcbwJi0d7RvrSnuO9Z+Mr118RwQ9Os2ODgMp+50BUrAg+B1uih2NyFFkWC6C
PHkmNLnTrAxmR1n/mFyI8AVq/UCay51VrhvDmlj+Rdgk5GaAEHqZbIBHLUgaqAQL
otG69XlMROCiJMHo6LdA29uZXRFPlBSsbDccaHO9b6G7U04BUpO30xTQ7C+5bg2C
dIdY4T87pVzMxRJvDe1g1tyqN33c+r8g/CxcJ4ABNhti/qfF0GlQGj2T1CcO311n
7XXOU4kgJtVxSNdeYls3CZ5itcL5JEr3TvxgF5OmiY6CsBU6pq2FDhoQYpgnhKzQ
eCHlm4bLvNh45sw4nI1M1QniY1T1uIBoO4KpgUahWGBnng7vIzJcc3zq8O0f5/7W
Ahy9oAGewdxYs6w8Kz911NKjiRncK762Nypbo/sVyYliCaNo2WwQK84pgdieu7FY
3CFCmFbtjGQAgEsJDRHnNL67NJXYRMIt+f1vZsN3hVj2zhP7+7O94N2gKCksCjXm
uPHtrT44KPLyKQfFPz5QD6F4BzFRkQUu/freHAkNooLWx6a48EUWaKksUFF5b0NI
mWz2N0popZDkC0bOPhcfg38HagkLLCEq36js5xeExInEc7snl68FHxAv66z3HOVh
wPirkUpz+e2L4RDR5hvds35OZYKIQsiqYQf1hXcdBjq/9EJ0zLWIJhVEHsStp/Cp
8QCLizbBeTfke7QqYjbwQcDfzuobNPu/o6Y+roeTnkvIrfJyXP07kL8QXfe5daTQ
kVJBbTWYQJ7lvYVrcVrn0LFWmMppUinwOnDCd6puediZhugTXbrnDV8ZpPiux32l
pkWfXxRgUrWZjZJfjneymFvo1Vg3Tu3dND/E5LvXXLC35Q/tBQ7CKrL1NdICp/8l
7FrQGqv1L7DOLYskFIrPbqjlDLdXAuF+wZ/yFFEnxVxQi7k+OTSFHr7+A/3/RALI
8EXQQs581QGaT3G46YOI5lFBzmu0sCEmZdwcAI+V+8HxBzW74gbe9Cr/lfMWFFcX
qLK8YIkxOiTvxj0VV4/2c39koJVqyQD4bV3tVGXuHNRCVW6KCUup7Gb779XtcIMk
np+y1U01JOrvdyHG0Ddh+WB9DerCrYi0bkjZgRzzckYRQMQgAdUMLPyD6ffwNoaZ
FU93/NC2XNb3N7LH3zS+85N3Rprl4oXKB/nBuk35f9klpzOn3oR8aoEgOHdGEPfx
6x6jI/qruoUpEWOZmX6KljhmaeJRMp5i0YFguW0eRKrCWsEVK3WoNjVI7eOFs2Hp
NVgv2+/bvUoBPat3l/Vw5SkGEuz59B5+wOcebLFfpOMsxVtDwCXWV30lTh15Q4jS
klob5Ntt8fTsUGlRpBDX5kalHXQz9wKtRbO6GHXDWdga4OyTSNI+L2XgXSnVkBr8
qkdrmtnVlQCqBxUg3IJP2KLPyS1+JBXBH9WyNTB6+isOp0yg9uV3G4AowsBHTvO1
5ZBOiW3eziNRwRDznXHYHbWrlZPdZnWoWKKRU90YEMpAIe/XDGJ9y2KoVJNMi4oV
H720UD1FaM7dGDoNNp76BVqRnRWYBFhAdUhbm0sX7xWM4LaHRGfER84430cpm+43
c7+W9PLz+m8gE/G/pqrjQEnIel3Lvs3I/GTMk82agraGD24DNCKzWyx6Z0czUTqL
67WCZSYYeK7agRqnvlaGdiFy6mKubt3/0z89NV5P+00MTfglPGzZKzyTHJQwqvHx
CDxNP2yQbIqSBS/ByvfPEx+K5UsCR1y+WdSJa2NfthypYKSkFKrQw9WuUb8KkR5z
Xv0Kr8wA8L3b45ir0zItA64sbSKlOQJtqOS8WlNRZq42BjAYTEB4lXmh9K6NlFYx
uu5VFoqZeru9XWuW3LefsC+YjmgbXoS042MfM1FUIUoIhRokDEu3lwiPpZTFcgsx
bo4NissmbR7+agTDS/d6IITyZK1PeuGrOiyLfYywGunob5mHZCVZnKXf8i0Go1UW
m/u+eZlAKZXmV1PFTMyepNtBO01Mkp6uBm/S585SRnG+ThTTZzSqsV4PsH4ffHcb
dNFnAX8MC5lrPQwmmgrNfGaF0a7RgBgR8jobJzU/cZ1Xx8XWXDTG0Iwpyv7z1XHq
X+063XN0+UvIZhOfuYMCYR4rDxfpyGJbODyJe4S997qJQ5saj1Wrwpfoj1Kfb/ks
NGg5YUmJ5lejTgTsRUQMWcIYBc+8cZGeXWNU6TMHjRkxEw575FsO8OhtlZiCp6gZ
H/JXa2rmERQnBGouUCFi5pRvW38p6Jm9rqApKzP/bfvwLeQg4JLELJLPX6rzszaq
soP20anXhesD1JaojV/9BIYTKdVjmB9wsreCHWa2P7iLqv0K6nGapdy0ei8VA6y/
Iem5jbKQcYd9YmC0qYcZ1Y6eUJ8ZRTKPkGFeG4luT6afYMJ2n4LZxN+TqsBGlHVJ
wHnO0ThCI+nUsnoCT7d4zR43fWI0Rc2q3UMltxqXfQG1bTIiLG+VIAvI6S9Or10W
Y3id6/1jFcQLdWrkJUHC7BLiBg4sTWWn7KI1Gf3mbndo/J6v1pMEIFCo3MF6LmU3
gdoGdTv/iKCRoGdA1adiGE+rMp3vkoRXAIuNJoU73fFFhqiWSxo9/46XQqNUHUAv
97W16xlkgTvB73doh2DDZw1MgoiSBGHDb9t6Hira3zx1Br1YDlRJSrHI6May/Iqq
hOwx7Dr8zat4YhLM72WK8uZhJNnlpDb9ctCTsnGD10ZoymJW4UzhIc3E9XWaH7yD
no0d1KvtbhrMYdkIyt+0++YKnntJ0fDLwbbBvM+kCsHenri1F02qfXi7F+X5Ptl0
/uNpfiXxa9UHXPbC+iduByKv0N+0EaY20TzjoUr5Uw1529QxSAvfbvqi7rAt7iEF
GADMazNmO1RvLqGrYpjuzM8xsjkf4L0AeAzMko3nXY9L9quHEFYEQWbrAC405MPB
CwR7/vj0ozVjMIuqIlbb8+HeiUJ5fC9tDnJ0N3iXMm87q/1yuTvOvhTMLAbRBhnG
PUWse1K81K5GGgVLCi0cg4pDSZYvrm3HbR9w54nAMFB8PioZ3zbV3bZOLnXWCkHk
kG9lERZY8ClNuAFJSVcgth7/Nb6eV6pJAMpNrkdi0VdrIh4vqEqNcEUaYqDngohr
3cwZZWQBWSwF/swC/1M8/bYPtnaoyiUlOuSxS9oOwJsxityty16cU5AhNg+Wm9mo
x9taOX+UvkTGPIwLJY9PogSV23CxSWqgemfv92Ax4B72pl4L8g6H3M5fyqp/I93Y
8nkEdb9Nxi0TdYNqFHbmmyWHHgEXpRl8pLnxBGZf9r0t+qTtPN51XzewvU3Ecgm3
HzqihgvmXb1ARDWL9owLoL3BpiClsxGERiVbMjmdm1gqnbh2Heo/OGMmSWXO+gLI
bbrQbshVzNiHIR3g8TL3B/n9kUDKU/2/J86/bYeblrHuTykQJDt2Xjs+p/filVbL
KJWNXqIjtepM0fj/qgZkOpEyzl+xmHafZ+qcroRzXixJF9eLmnriWRQkmLGFXOmL
K35h0Kx8B9A07QUT7FcCM/IhWPIl1wCShDcFr+5Hbsvgqsc7Bk1UjF495nPn6UI4
azGbhlB9xLeANIZ6eCzZ0nPVCKgH19MGz+DYv6OAYjxr9q7ElYJ++F8o+73vT/jP
VBjfhGqDOxLdhemKOFFTTy00JBRwykB0quVjiewa4V/9Jle/0JXGdpneS8bTFu+0
2IzJgBD/uIQALEiPRXq7Vm5JXTucotmOTsgFTQTnCJYPXr0Ou8GPHYr4JX5ktshG
+31wRiLnxJ5Fckgeju3RgGBPEPp+ePI8LILUdaB8DS9mZsHgff7wffN8i4wbZZGA
2nrRlpL0yINN/mM2XWLA4KEnxN0aQBPg2g+vZGZSCGQhea6TTDCvggyoBUyPPRGE
/qEjd6Nsn+RrCbsb3d0wWJv+Un1/Tq7NogYsd3BPD46oARkJeThMPt63LNcLcJ37
B3r0j/1ggRKOfa9+5jh1e0vfomIDb8YH5jjtwX7Jx1POjHXi8HVs5TGcMGFXSSYn
okVCMXXy/cf9DUDNTnC2VhFJ9bmTIX7BNbqzSnQiTWTH3k2t5bz7hhF7G38mYiyw
y+0xKlvLdMXeOdNeI0vcZbACklRR9Yq/3Fpg2jQMfojDj7BQ4VEbFxHQTNpTlVKW
mmagk6XaTWi0MRGqX+pIJZQPQYzsVRngk5vxOaBr3i0s31hdBFoGVwCkwaAaP9Ik
k2cEkMTwjX4NAxQ3aKVRxhmX+1f4r04YDfz2vpr28YWBwuhUNvJutNZWhWXwZSYj
Qak1jfuyS1x6yUyv5Fcj+J++srnTGDkU7KXp09vPP2B1DCKLY8esHEJKyFiHq8PS
+UTiGl4dOiLmMHyeYLpDHjw5OlAxiCQXwX+B0+C3xDpn/Z9DyeRNaR2soXn38AfG
LHvnvAScCNX+bBm4CCl4W/sPYusqhLp179NM1cBV+mHCbllRAI2MxJxy/1/dhvW3
DHHCMgSJoD1KTj+NEoiJC9ntAe+3Of/eX7pDgQxhdaKclShLOd6MC2UwHXGq1v6i
EkpB2hXTXQBI+svsa2KsJ6GH4GD8XJWBXGpFceBTosjTvDqIBhqKE9/LlXLH7LmZ
DK40wLlSEprpL4393hwlqLCoBrq0n3QegCR6yAfNRsE+W4jU6RdnLm4pzeWcol/w
nubMK3JNp+O8i4ykrhMReZ+X6+DdTbzW/1+bxxxc/uq+i/8kIBeVpEgq2MFbqgMo
NQs7Ph33+0gvCsvpXgQ9Cxoil7HdgbeiO2Sd+SdTEDQ5O4XaMW+w1N6rbuOWK6cx
8icULVfL/obW3BGTSYVSKCw1hNLHibvJrchcZJiRDsaQ6/KE9z5mg+HQcABns4Xn
gyxNitCrsBkipGSfn4KNpRqzdiq3p6lKnaeJUsZNO5TiZ5nJLx5gxAstwWaiYJMY
5sm/fewTRQ/8yshEHwfm7FzhjKyTRNrSZz2SDuMbMkOvpZzhGK8XfbBKu3fvnpYk
aBtDiAIjNSsF62zkkpKqPKmIGAKp3sh/dyRP2u1/LkNRz6/vHGZT+2SXuURpgqua
o78M58JOl/vUKBsy66qqWfYzoM/pL6Wg0/ghSp6rc6+b8TO4FExRqfKHVLqHVaKP
PLeJ0Bs0Kxh6A6o336PZDR/bUQWi7brrE3q92WLQBc1ZTYkzSgjBDBQBefS0FCb9
mFiNB7XD1oUiuEDB1ulDBrNoLocWeZ3uJykPXgoiR0EXYeUmGZ9zwpbVJIEc0uJj
M6VeUpCeQoOAUqg1EelU3fXoHykNzIG/QvxUAhRqdpByqAnsqXt/t/OH/gKXvHr3
9VWhPpVAHJzzd8u5mGMEdEINxd1Qx/mkJv+8Ho6EWeqQAj8WwY5FRcnQ+4fuc+rm
D2+Tf32S4UsohfG/MNWIRfOnak+C8A9wJLpzP/9tWhyuWk1BH3biWvP/e4W5Ik9l
JDj8vNEFUA+U3C+w9VQ7r53MMI5XRBFyRt2SXryHUyyg6oNkUx9O+F1J8AILJswC
hghe44ShxiEtrAhKBbvXR3upgz/hZSYoE+o+071VcStNkXbXoD8vmD0HY1dE4Vvf
O3aOO4uPqO23by27JuZ5pbDkMpW3IOEbeKF9btGuTR60YaWsj0RPtUtC9jh06lJR
U0rWI7+95PQzunjmphQKikkHlvorrMPMBwefRojUhf31/M0mHnp5jbpKvawoNcII
8fWip99ZXLx9KJ7YGf6H8cdbG5kJlOY7UftvNJKkVoib8OJSmoxaRxnRFU1nPm58
GOQ0XYopOQIMTuUuWp//N7Ct8z64zy2K4vyzWjTj1nOhZmgxqQFYSGgeyi1kPeUV
E2jxXeBDU8GsxhF5K5m7/dLCU/gtaTcIsdVohLzBikoIz2GshTWPebF9sSxf6gIE
K79/LHd0bIhX4onIRfNzRDnfdITKazVfFRbHVmzlDWKt/8ELBUbDvDHRodCxdJ65
yGnYsD6+UcGZPeTn0YOdFArjVx9cisorwdaU34Y3v0utZMAv6r4KKL7YfUJjyEXB
bv8dvZ9i1V6Qo4lOYf044DeHni0lNOEHVZLWOEUG0yZv0zlFGJlxhSuWaVJp6jHX
KazPn5yiUSiQROjkeGrrvMm6og81ga/4yV2Elsj5MfUk7xElywpdOcB//exwmgND
RiBDfxv1cQenGpf4HTP27N8HQJweQlHqfxDwyyvBZ2RhzS9prtrcvDNrgzlT0sAw
51nutLKJ9f3vXaLdXtKZaQOvz0WKhbKnLfOvkKnNOu1SuOx1haieWgabXPyTSboJ
qvwCjDFynoSxmZmEmXl1X/zsTF6ZqVfG8mwOiOX+07V06L+jWPhnfkppIUXKDa2W
5I0YtHjNAVqVxePHu8XHENK8mKQ0x0pLdKe6ZJ0iaqRlYp2jrZE27vC0Qk+E8YwR
vQkKRxj3hrdu66Uc9CidUAuDtm5jSn41+Rt7HFwH9CbGvOL2jwKSB+q49gy0PRiL
buvdCkxKy0hLNDo09S3NOMlQ7IcosLG3F7asl/GuHok+4yKo+rc+ZetHYEufFCDf
K6/sOyZ777+VJFJyN6HmfM258ipWpWPP/GVPWlA41CsT0/TL7zOgRfohfk1bO9k+
y9E63E/TWP/nIJKj/HNU27s0RuqrQadchmZTyGopRWcenZuIYqLBwOtyT/Es3AeU
sEWdGBbGZVVF6LFgU9xjFXOChl9SBPid4QC4/JGbcc5Llu6ongfJOv5keFfmeTPk
4KSnXFiQBjSpNJcde98hC9LIhcNSoZODcrSIG3CjMhI8dHMqqAB8NLDc62X/cahB
S1ZWNvC/NWjPMtR9pLFRHGMIOFRWjENIRjxVuUuaDkBvfyqDmB6ldWHy7eBLN0gi
wg3oP0lh6IIJq8nlslkentgyIReWzniJuXUlMBgsOjrpAb6Bu3Pd/8EvLA44cjLL
j4zx85noTML3WffNkAgfS8TVPB/8znyqqF8hf2Pl8Sb7ir6nkYc55uQEoRNdxwPy
pHX/xGfdvexfi9gCn5adIkhRAQ4YriEL2LH0YzG9H7GBlJhMNszvhsQHRoRnO7ZR
WQx6EbTuFyXtgVBrS4s2KpLE+vL2oV60P4iC2WuFGPkDFHMpS+NrooQK40jecbP/
uXBK8ff9OsD1qb12kVgCc3t+w9YXTWBOqEO3zYmGxyuVuu+pXOKVEA8hsIk5sbBC
bW42WQ8XoZFjVxh4nNSFcWqLPIyCQnYb9ELyrxHD/hN7FXRlx6xCSQKwVlUvPyuR
CS8yO3pEZzFibewkQp4MmLSatb1oHW9DtjbS3NLgRs8q6cTPpTq1gA4rxOuFCIa4
qBGq80/e7QnD6Wu+YFfQx5nDbzIBbz+QepjRkBUc6TMURXQhP/cNro9nuaGHlYY/
XvJJ/+ktA6m4nOK8f/t+Y0cL7N6RkflnI+dBw7fxloVBdGRMud0AMp17YcuEpELX
Cev4nEVFa3CV7qBzMpDiLaQS8KBybG/GPwPZQslm4TBOMGqf2y35VJ6p5l8Fx6ct
TJTPDjbu4ZhexBvMWXNcv+F/eyXApNYh9G8Geo4aZiSeYLdjwOa6anGojktIcPNz
Jfh4dda2dZloJVYqgPOUC7LqtRAyHn6u6kC1xBJINA3PpVxKg4nc/ued1aEK1w+P
UtTiNetLITdZdSFmsD5jpHjXKDGKhNZzgSbnQRZPayOiuPEfWFrmBLeCftrnrCOC
9lBphgtnZNQ8P27aAAZPMzvJm3b/9zco2ms8KKGpu5oZYMTJSJ6zD+tQ/jB+kfAs
ekIquhCp5fyeexXGVCm7lRuSCjLf6FyU0C9gnzClYtPjrn7ps/5U5iUVmp2qxtXq
RdD03KeG9eMg162Ireqthf2dWieCPfd2wseWkX7Z3MUIjWm7DP2sBX5bFsZFYCH6
VsmMJx8KIhtuCEyoH8RuzkLflL6aGpqEj2EwgwgJxzqH4XTw/0DSubz7h3ieTJnr
5UuFpOzpBbi88bASIaRuRQhGa12RaLKup8rEQODl7idP4CoV67A6N6V37dOQ2yYs
+uduuwmBJzuYwu859HU7jCpezVOelweTxxLam490G/DF8OlyyfHPpFP5Zoo7l1P8
qeUrD2VvqNpsQ+B0Zfi98gMTQtnn7YVh9l7cPZmMTzxeRqGiFpz2E8mhb3FnFkf6
6sXV0cduLtfQSg/3uKAeZvJd53P5z26MLfgYoo9EdBwtwaavHD8gS44u7REwPNyg
3ld2jJdQPzM0MWRqT88r+iuksxG44bZXZzAeatQVsZLtXnJlUrKStuTq61maVc2u
4oY2xkb0PponFLEzNSvWMwfnGsqIc92rifSg0fa2B6Zz5HsEoMYrv84W5XBOWbgY
qaq09PSAabXsY7AuaY0mYBkqZ6JxZol4DtGWlaBBXijbSWA8Bb/mP2yIpafGyLb8
BEbcNj22Lwf8KSqd0bED91iA25jSOv/HYvQobQVm6Y3wx53NVmGXTQl4zolAhUuF
YnRLweWM+7LJexzBwHLd5GLkw6teDZdGRTdTXX2vJv6jufKuSkLKf6l1Z2ITJB1q
VFobB5fcM6aNqA5TFkpuIRi78G7sAQFk4/hufb9hpNeX8hBcumNqVfcRbWRuGW3X
IpwTV+Ms2GBvCDX4LLpmKsqmqZ83gZZjQ7j5W0j8/SWxoUL4CLBIQYeXFH6qn13m
W5BULDub06tusVQWq/fHcIN3bSXorJdsWopcaGriyKYpdcYcfJtgvHSL81l7MyiR
mg9dzVp43lNgMdkLg8TFA+JXhqExVCKBax8h5b47sX+318RNUgvXyLbDPflvT3i+
OitLjD+3zIEcHZ3lO1Y1BR6pw40LoDE9cVDpFG6j/yylUBwAbo9Xy4SRel6fjhS/
o0lnQmSxKlj6fs8cqoiMt7uT9A03xtmUkzdjcNUz3/Zl5BsoHc7HVJgY3g5KE3Xn
eZ5WOciFQ+AQKm38pTfrFCo+mYElAqDQuhYNrf318dQidXZ4gxBzq4kipn3KHFtL
URJArHHLoB12msK13DdZDTrAUg6vNa5b420AQHHbI9Xv5xFAq5lzxt3jDy2aetfR
Ii//xMqymVsmt/jVr8iEXa9vRmW1zKr1BWD87MUq5sHKdxoGkp2T0j3qy5UCxxHL
yqwCJpkmaJgVrqS8bol9Oyl9nfp44zEpTnIjkDl7TgfxSPDYHEfivCNBaLHaDnhl
vxw00bSsjUzQdo58v7cNUJuDT3R5E2XWhKESdA+csWgoqfDFZ4xqrIxSFRIoeDK2
p3+Cg532f3TBxFijL6N3n9csFX6jxIfao2OZXw7h5s2Roax1twb+4da3ElcgB+rd
Fzfrgd7b1bVFiHJXrXThicEfyaVDo+SFCrwPrK4nreiktGMSN2Jb5zAX3TWwRVXV
weFgVASWSa2XAjZTgXgWTThHs0QlqHmvwfjAx60jM/NhFHv3V2QG/bCcHsbnCHVq
kMLlbEg6DENWO+af5skSVK04/68RydtP4Xb0qwDGgSxy70pPbfSjNkvXbpMQpBbx
QI8V3tZG9TMvmVqRCpvQNqrd7UkbB+XclHWS6l6ZEuofWx5kEWaheVKSJ1U4SXC9
awE4uzXvCM57TWaQ8zST4eTRpqNx5H1qTxf+UrxqSgCRG5IZsbNCnsPD2nNwHNIv
MyxLfzdCCoh4wSgEspBTes3dTCUYgh0YAwDDqZJdYLEvAOHkm3FWcA2IeAXqn4Qi
FiJe1UQB/kq+l4XuTLOmUZ1+0MiaFayQB50a8HpbC0TdfUQL+fjb0O+hXhMDx7xg
+6J5Z1T1gwETArRxVHNG/K2Lmrr9fPfXTDX+j0RyQLgvTPhg5NaoGOVWZj7YnDeQ
iUKAkpIauRUxjJgIEeKZUHiTcme2s/65ibvie/4MXVHkPJBT5HfUPpa9CjxLkPFU
I/fWHZZ3lGwM4fNL9AH/YJgzu+fSUkNQXwSPj5pD53e+QRPuuiQnAblULSeqRBfC
OEXgjrvVgsatuWinR0qYaB1Oe551iayGTCKdF2JGP6fAv77YbiuSoIoOy4LTejQA
seD/nNNs80GZPBUCEmzHWQxnSDCuiePTOhDgkANYF6R05uBEw2yil8R710jJe/7v
9LFA/2f8VfWFBvj6fiiNSGNrKnFcQnum0tcLZaa8XyiCBU3xqpjrYQSAgLJNxa9K
S91X9udJGeeFXoU2tDrojjz3i9ra4/zA/9BIarX3fmY4fIJC2FCkc+fKl3XTaxSb
BRcTKXy09/uUMPcRzwpHnEZZsEJOmojxO1m0+Z8Pg9Z8p4JUCZcOV/CJ8Hx046m/
ZlGqaIu/gnldzjU68LronItzH+jJO6fqQ70ghpXc99oReJzKvf6hH/wlP9L1I+9K
qz+ca4HZaNraX0ChP8a71WftP3TkcvmbxvnwmJD5OzwFiTJjtdGG9BsZgB1fri3M
4n5dkCq/ElHR4gdsjQUQy8P9WElz6IFRHbK6vR1Swv6LK2FLUmbc5vvKfKkBEvo5
aR5q/KUpY+UiBh708oB8UMu7unLQI5onOXatp3+dUe+H656YppqgrmVx+dG7/ZWq
X8Tr+EwjQs6rcDyENeW8j2n1qqgJFFWPn0Aleeu6XC6cpmV/Dkl3GkfBbSX3h50H
in15/rwlOhgrGE7R1wKJTBdfZVahLRiZTYVIOTtJlCnxgnrQHqs1Uu0NJI5bIXsU
JiqpK7hNWGm3hCBbj6vd+cxDTpRiRRtHap2iRodtwKMxc/hknMpq3xVkOxap95xK
Hf+3+qHiz9VDI/viVwyAFTy7U7Ptyptiktc+Ix5VHLBT7UBZr3JXzAtxGzdvqzWb
25jMVNsXl/a7FAWvcIseH3FNEwU3IjPchDBjVwv5q+5qGnWKQyoJ9V73h3qSzgmV
hq2ULjlzaDOy3OZMS3q/NCMUGfsvgCGeJmzA4aeV1GANrjxaL2jm1DqS85kiPA1l
wPvrLyaO3xMtoirz+bM5SiY7K1FSqo/gmtrYV2GQ0heipQbLeWM4tFI0Jo1kz5Wo
ukU4Z35sEPqwLLywBl/nWhwA2RaprMnXhJOJwiwquB1d2u0dgb+j0/2sl0aJAWef
2ffZzw2beBRMndxRs8sh3ogNVGKRlbz75gIO86lSqzAT5CuygN9gUKSmSggM+SdV
QZxRDL3oYLFOhmGqIiVtThrTWbHYSCINn1yYGk2/pKqv0JqXP7gvet2S/b9CGpNo
jP4Di9ZW4gXbIiGWA7Q6TZVO1befe0vdToBkafamnTapLv/afBrGFRcNMFlYoJ21
Uczf0UcrYGg5Jsc4hzDHQmOSJZ5xBf+bXRw9BaB8F3YbLaHtsKD9b+jwIkZG+CQP
uF54L9JA6ZrBLp4bceSDFN1JzULWpJsvwSLzkVCpTDX5OYPwSU3fYU/QkBqRu0/q
xHKcng9TttFqcNBrWMJWXBq8TQvtHKC9m9SZLVbG0nxZUpoa2PWbDtmGt7neUEzM
p4xnc4VcPcTzQQgz6aUmxQF50H3pgH/XxYpoOrjmwYiKpg/SDd9DpZ10YPGNj+Ty
VogdFitStvPl6HhqzJp8++k59zvHdEpIOPXIKQiSC8Chbzl713umHiGIMTRcxyyR
JGD44M9JAqNVt8XCaUHzcx/GD3jWjTA2RZMggEve6NIq6hh7v93K5+DXywRrXOAU
zNqYjCj6UbXRtWJYu5122CmbzaKWDm0yqqf07jhTLJHXMuO2D/C96NgRgZHm96mD
9m4BGZRuQgvy12NBYq/EwqpSVjj7/F6ZaT8hoBleyRYOl7jClO0IkhTsIMii+qVI
yVWJki1SX8a1alkSxJLLWOGihc0mwSsmK6BlD1OZ8TeZnjhtyUnTgrvsDTUgxmUE
veVxz2nglLYmBogRKfZjQkjDxC4gDkhXJhACfWyKOKsMSInO+dhqus8Bgr7G2nJ1
Uq7i56kcUlXrBkUE432iQ8JoLC7oSrJbRWQPt0YWbgI/XE0vnHmrC78Ui3zZhOFI
1CpZAl+QO3cEBy07275ir5ARbLa6dd0U/8T6rvf/yPDeDayLaOi3oaSqG/iAPtuj
9FEKF1Zq6sb0Pd8rq9FHD8LpYLN+Uhbyex5O8JcVrwIPuAaBJaFSnMG3L48CSRys
OdwarRJEse/nnbvwHVwZY/R4NklWoE5e5CPlmgK8rJPkzYE4pHCAiAXEpqNDPph+
KRmoXp7mU7R35bkb/8k9MbMDDGugY0Erd1+TNJSRHksk0I9sPBhdr3RrJiGQEDto
ZgmkF+4rYtIoLjJ8VnpFiC4tepq/6muvfp87izy7wyihpa9OZM+Aa8VPn0pmkHeF
L4PKOD7Q4InZdzQZQQUlz18awbxeBrn+23FkEBeVCKMz0uAKu8gniZgCrgjvTE9N
K3+RJfWy8wBnIlEnK22qgXUPKEDqAoOWFV9608a+krdQImBNQ5NsyJqIfFKKvWuN
zjqrT1sWUonPX3x/nOwgH16GshkE/D1Xvr+5Swin6le0qHmytyP1RGAiSfijpDoB
N7PnfsgOtnBlEaYe+ryVYo633w3xAneSwMxEbw0JdnHPG2p7zquBKq1mo2yL63zb
GIs/0pos0yNMi096Z1LA59eSVTfJ6rGh5cPb/sMcIb7CRZx837Ff3FWVL1podtda
TCkp1Vlwwc4P1BEgZ/1CeMm7B7O+aZUvmCqxb3S18aEaLU/IZQsc+n1N+YCwBvS1
YmjVErOIXEBU9YYRsMqOTpSNs3PxZXVpMEEdQie4nAs8vjyd76DlLY65LocoIfwB
MYbOk97phkYmTCniHWSiuYy2JZWoNgLn86F/gaZ7xnt+mov3PXZAemdcGmyEHyJG
42fXl4lKmbzs4ezyMckQLFcz1CWQ3BnmH43Mqvz5Ogwt4m8a2Q5bo2IrFaNTYTrt
uo4HJvr9fLZQTZPqLwMMsjQj6tT2bSWYF6/FTiTBzx0Iw8cgTE2gpN25y425U1Ki
KWg1qb6Tey3Z2lrXAd5vPvzliC0fwncNACcLsNEdGzhHz/lXagQK9Vi3chv8OAgm
mOKS0yTz1U5OPfj3YG3ogU0FVbD94Vk2bKdkbSVY7RB6LpR8LZyi6MtU+ZwgP1Ij
ll3c/Wze3Y523yqKhkObF/OH29F3Rq0NTHdFziQmHqOB24vngP/FA0zvIr2I6edP
dQiZot3GSq46pVClJ2nbzQpDfmb5cTbbRMC/7mo2GFfMq5ftJPcYQBF9kHgv7JNi
h6+X+hIjoiHR+dORutw0R1cwDhZ4ry4fdCZqq8DyrTjkW02cmDXGirTudY4eKKtp
+1r8+GGAfmTi61phlb0/E4qth0d89dc7egF1fJxZpmVMfGHJMjsvRg8ymTP3iKvD
I36Waf+ORINdRG7//IliEs7UZNtMILabSo7QdKG9kd0yCofJZGtP08zW94OORBj5
mhUlB0VFdBx3SE31+0vBU/QpuSd8v4UugweURcJetkRvBCQ2BHVK4Z9W7I4Z3HJG
5BkNyhxAG3dVFfrQvQPVPtUh5aGbVx3A4PJwZCsaSREM/NaOonFkPxwW0w2bWBrP
l0DPO8PZjU2UONfuIFjeQ7xagpZawVFhvxS50vB9kBJ833M+unqu3Y6JITI4Xe4v
e7Q8M+c9fEOc4ZcGfoCqCz7WziqIvdX8+q+xwSivXailjH/jCodgXiSyZxAFiR5z
4KlqKLrBfvxbtKhLAxryBpsC4Cxj5t+5/9B8mCPh+ZtadA/Q5E4e5nHVJHA77Od/
19jhzSGAwR13KguweSBID1LtcIXnTT6j1+WgX7aDD6dQT1HoVwt/nTvguPkpQAaE
u1gbH5zGuAiAkNsXOCkwGexOoBzTT4FC3cdBi9q3zh2nS1k1AN5hv0pxsNsJ8sWL
jxWrAdehVsXfy348qcgXvjjOceX1LfQoRkjwqd1PHvpRSnDiQxMXg+PMmqNfng8y
fNHIz3/oWyhc81Dn2LLkiWQizhDemoAiz4XrxjpcfS6bvkUtC6Hm2Q+D+Gc+e7Ve
Ep+cmySDnz0rVb7zjT0UCBGiM9GcQCJS9TQE9OY6P4URKCS8srU0G6DkFJnvWKf/
SeSlRwFqa3hxAQ8d6qD/Rankc9h/c0E+bZU8YJR6qWhuVr+maVNSh0XVvGoD4w50
vYRmyxOqoEf6uqkg+J4jecRQA1UrgQZ8dmjtXrLu4R9ipg/Ff09ck1plmb9V/kLV
rg5JPV2iOb+iIvQ9y+On+Ap2nvA0exZxzZ6F9FvuI3zNf0/OJ9eLzQLLs8dUY8kl
ISLoVHFWTldbULHaErSy7faFS/12nxdJ9QlCWgMV4W0BQiuzfqEVer/G26BuuI7s
gI5U31ELtg6c8lpOdaUoK3IH1DmOqpfdbRonR6rBswfT4AXA9wjwMxvdVVD+PEe6
tSi9atgtWUlySZg/+OQHA1YmqFOCXGPnhOZVcF1mTE7+KbC8aYkSHuebX9tlRYjw
IuWhKIaMTMw/tm62DxgZ+lv/iPhisEEebg5nShIolxth6vA3732m+nVQf/LUMgI6
IyIar00clOlsa09Aum0qykknvpTdMHvgHu7/NVI0moocKdwhZkbMO1ezyW+QzrKN
bTDsaBctdrH0inMKnGmXyFf1mUNc+WObGgd3Xribwy+JRo0FBzmrwvGyhrnc11YB
Rsjs5E/SMnfVUciJ6ZowLHZL/nPPWr+SmP9BSWeZMsv5Wj2gX7zO3lnyBNuYhsJB
ROxtB1JMrgex721FpRb2JllTUzRATtL5Jo4LNf89So0FIi5GvxfSuXKql9rds/VB
h1+GVlIjdymD5loA7do9iRDfWGheYn9otFOkti6KSTsge9XN6Hmhw8tGLjobCzzD
tHTjfuV3B2+F+HZ64KGOeX3rRClPykT4UXIfSUmf61BOM2jec9Zl9R8bXA0RvSry
6k++UC9Ptwkv7ZftTWChDGfh22aNNaB0M9ecGAj7GqwoKIvJwc17HZnNI52ye6iX
kdFGtI3rrO3vWZlMO6ZGQ+Imxmgy8BcqwQ2KtIAp9I1/Z2RK4PzO+NFVnB9zSPJO
zPnZLkuMX2+G4zbjmdZi2vNltFw9bxHrLyupnk7Kqe0KqGZmRf+pP6j/GgG4lsuD
AfIqG0VntHnbKCOcLcmVqO2YlCa3Zl5aIZjNFn6PsBd6q+xJmksIqiT1VE5lYOM6
BvlxcphMPpmDfvzX+Jwrr9Lsp86dWvcvvX5jRB0K1zy06OB/9fNgV55191NN8vxs
D3iaAmCSitCVTWI5ECj01L4CiQBrAx7H8zkh1FNa7TYERTXKlmOAa5Ug34NgQzbH
0ta+wmF4b9fb0i+ztLuKBpaNEpDz6lFhZ6QIwcCym5q1UKieb5buqxorKaUmH7t6
5xWCXKWiitSXt97ILJE63HpZWiUsZnmkp/vuYx9Cs4YdcM799dsa9bebCn+6EoUB
wU5zRX8MPWBgFKpxMHWvzbuVomQ3NSzppeFzy7MyBenfac9ozHMh+AejBvRABQiy
7qSk+SUdPLfDXbjUh3iSQnwN895tB8a/WEm+hioY4rOzORchHpXra0CF9S5PJFTW
Nn/SzETy+ki5faCkWqei5gsvjh1GlsHbDU4gIn3QdXCZplPG3FghXg/rFQOTTR4A
kmpU74c14GonKjo6bYw3UiG8lG241YGthOw4uCg21jOUDv7azn1FZbT1eYPud8kx
HvGWbJjBzmWr3P/iI5uXRYOOwWKe45sBo6l1c8g8q0qwE+tJWejG+H+KaaheiFmu
mRoomZ6CfGwyPmf/MLfKwIuQ6b8nnHdvSCKPN1MH2KRj/zoYYxcNdvL3E2N1XsEZ
Ku26/6SPaNMHvZ/DyI6c/GEt+lGEDXsA2mu/mnsmwcIFprNouYXuu1ObdMNCK30r
KNFF7D/9f7OzsWuQtj5KBb8yKpCMzBg2vN6SNY9951fYBooELB4lyzhA0ah9JSnW
oTGpES2LRMR0yn8ExFpPfEJ7xPeQw31QgL1mLo1ZZzwHGQDaZEfTrka4em1sY04r
UymGMiYGiKIQ++cxeMMD/yTUEfd+pfUuz7fPDXFhKFZ29BntiQAC4JgpDzyBDyLr
GveTwvyW1WrC9/J672BlBLpE/ywb+WqjWs+gawb9atrEZhA4tcFgeYJxojdOcAup
kDJPU95ldjtsHLJduvYCGDzTGWQOEaUIqz8PJ7smCZekhTkhWCNzJsOBFcie03Tz
HDHMoWMaK0V2troa8ESkbnhKqK6SVrMKIXs6HDEjAU+DdMy8ECCWOCmfZ5A8TyqO
LDbWEnASGa06htCR23OJgqcplyy7+qU1ooT3jvlVTXf51+twZNPLvzeI11mDgFH+
meordH0alygKheXzTMcEIus9b4drB/RMiG45b6QGs1T6SzyxUa0NXT7pDQ8SWPeE
tENAHXIWqfC1P7p7NHrZNuAaAvPnMQHhxYGk2V3Lh7AO18bF9dQZCQFFuGpSWw0R
PMOsJwKO+HKR+sG1KZN4osAYvQoP9F03GfHcLGQh01fFuRb43oJcqUVHnPCZ+jGn
c/X7usRexZtanibeBwNBBTe/ZJXwP2eOlnlRsE/30IZVR/XBsdrBABiSixKu4VOr
ED2OXNbHHNjN+CDBUVNUGypIuf7C/kU9+6i/Rcfqp8zC0Rt5yAbRUphV2TxTh4fx
S8VE1G0cTRC5ENIeYy9/r82Yb7l1Jml5m7A2oFQBcvwHLadyGjohmRXmkjgO8xyr
EN8DMiwQJERWUzKP0LoiJ5zTAkpV7fNToCVFViTP/dv0LiDn0QLE78z3xk2uueOS
QmJoDBujp06mS+voA8o7O1A2pxvSRI+tejJT1Wz1/9mlB1SOvjEJ740cEouZCWdw
SFzOvL5Isdzf/TbjkXIHh+LrzGOIIhVoLKmn+6pPxSRj778C1nxjxCT5OL/4FGtz
lYIx1FrfSOeDB0hlzDovH9Z9nSw0bQDxmLjDYjlK/TnSms9zZvcKWbLLSnDI4seZ
XxQ6uN1xnUD0WH2PHYMc4nFJ9F8+YQ4ketu2LfMrFxG3ZKUcxeDHGAbMPWzfk8nd
vT2ugxDK3knIZBE3Rp8hd5sbrtn3T00uKxIGJLYti8g938fBWzIovzvny/XSxGPp
i2kckOrgbPRe7YAf4syzn6hzOWlX45R2mB8A8iKDoy2tND5tTq6XwAL011/5RFtz
zkCsacvKSmoB4dt5yWQNVQMTWNaLNVFkdVd+hd0k2M3X7jhXTfHQBQcJAtyRHikA
OkI+xfJ/A0QR5WN3x6HPQZR3gLgxX5MGtCJayoVkNQK8Oo8tKFduz+veVm7kpMgC
fQFYjs1JiLNHTV0WW6EDLuaGMFs0MnSzcYPmi5+iC6qtq6OlXpkoHGbCMOuEFDig
IE7kncrNUdCy7k2w3h1lG7uzCXQJzgiyqBf4nH3nSrI4aU6KbpR3YBFl1Qat+pUV
reS5M3qBQRQvx8Gp7XwJeLH80zBjewV4tCSbaSRGtTJUbPC9+S2Inna8mbQeW1L8
KJNAw+JTtTDpBQ8avPPKw0jZE9zSX5HyYNq9RXuDolk6AETHXYSllhnlPaHihI7r
Hx1oYSa/qAh2Ph/ehTIleUOwd+M20bvlaUNi/HGlK9CFJkl5XxUqJ7cjzQu6GHFS
Dh6gkb9alJmYZaOpQCXum6kh4S8TC/N674kNBVjihbEJwHACflQvAt88tHovMbLe
LgYKR2UXWU/cWGuHmuiUMwZ9Ybkot+zJjfHtlFBOMk9+2YegzIqb/eN3Vo2zVtSQ
3hr0HZZUtvVzQD+5OkEgXTUV0srapdGeHNifCp1FIWhyTgvDicFLbaX6lFoTKAzb
vZLWCcp+BkGfRV80JVbpC7Jr8XVbQrgffC0l/TMgPecZBnSPVdVK2byoc7ENKA/t
3PkJqA9aebvR0ctLmN9Vwq31NTJyUKnmLdInsK/pqMxb1+zU4zdsn1e42csbo5dH
miS03ElgxlEZTblqb0G2FSdT+CD6aK/PVDW0mkXhPg85aMnItCPD28lbbRqqC+t7
zxLzw+tq6/UbJeKdBy2A2jkw+/e0ZrQ4BpvXj4ZGe19WCKZ7ojl1laI+ldFSVWX1
5hFSCMLkAYDxByM3F7mUT7kph16ow9Ddr1yOGDpTlYzfKjOgnlue+OhpurdeUG9N
YIUINEvffxJqDPaWzVnyvXZFnOIUS4S61HMmvog6eNW8NgE7gWfZpwQnoyN45z8E
B3u8+u9qtMzNIh5LuBOxeXoiFNPPI53zK1XoELb4bwLITg00Ld9bf2i3r+XiUPxJ
YxrroJ8KbU7+6E7yELNYToBui5jYtbWthAGwXvtYAZyCk3Yy0X+4IVlIq7RlNPAH
Fxi6UiocYhDcFv+CVskgPwb46jI3ZPAyKZintn4vSTfh0NrS6uvFQ6wxwOWp2+Sj
8BQIM/c9z6uZlxkV6oMcXQ3hn39WpNhYn9WWVBNb75CjB2/FlZRKBki1u5pbA4hY
c4KpRqR/tdCxnMhtPGJ0pFUxsVOelPfrDlZHXJG9NHYFWaboxlYpRuaTDKrq+Rvq
5+KhAmfygKuZPqrq453b69+Bs0M+bO3O54ZFuTyOjEcepEUVnOoknK/hQknIIhIs
HIVAoOjRXgSxA5izXK1xUYbcMeaTSSU9Mp2ru1u7gEToIJ6AJ1fdV0P2icTR+nUo
oNdtaAeyEOHEx9PSHC9oxv+HAdDo3iBJHUWkHVOHKTVeKgjm1l5fOdgYAeFZsEya
sLZ2cYul/v+4yFJNivf/7/pQuNTsWuI+TRUO5SibJ/KhREH8sVlLg+tW6KlnY6rq
i7F2kxzAHiWZ84w3vJ3oeT83k8vRnc4V9BPK5z/86n998hE6TaZfporIvxhd2vFe
e7MJ0dH+OUKbfQg50IYLONxno1W22NWGdJ5pi18PSMACO5FrvHFEMZESvVDjQ8CZ
XPC43xp6uLZ8JVVQB2pe9oT9TRuTjDuK3BX4WjDNp3hlwWrEPBmMLVufEkxDmeMS
+HuCeyPSnBmNTublujwq8S6Rg0o6cbvfBI6zFnVHyDe+zpWaD7i2fEkJNNIgwfYl
tfRbANV0nf4Qpz9HRONl/DcY4l/SbfKgCXyZp9fmBOT9oUpl9pGw+JuxhsQ6lYnu
41y5Gh7QEwA6kS86bcPMQT9e/QmQk9hH1G1s2wNWNwup3/z68+VngiDi4oZq1Hwc
IULy+5Jeanlbgc+Egz/bEeNHuqV4nKeAzJACLqmZMOQE83NHqP8PmJutP9zERGdp
N6aC49PHeGBNvoNxIFcABzJmOYAlGzL/CVHDdMAZwHrZmFPcG/PLxrXbsZU3o7yy
QWzo9BLIwxsgIeLruIMVKf+QsYUXPbckOkt5vSG+WKT+K1YfV5lfIz1gLAuueXSA
/BOuGfVDEfiExE18D0LjdGmMhINtXOOl6jYYq6jOAcqWFnrGmHjg8M/95+78qagw
8Y0sOsZGL7gwPISjFuTLTw442CzBnIDm4MGCdD746E7OX7WafwUZHeuTnkIqbtKn
TNa+1d2nhGPlTRqy9d2nEzeuRA/E6JKpEasX7YqcMqR/bOwy4SUkfRYQc98txNQS
LX5Ua8CyDr/B/T93/fY75GDxE7HfSJazoitRATU0Re4PLdzOzf1bJ5s3FXaIbnIt
Pn736SfCdVM6F3FXU3JxcnyYKEwoRLbBEpkvcLvfoYwh+gSXL9pAnzcs0BSiSMu7
NpK384doqArxuWOBsAypH7MUjCWYVkDWW3RUWmr7AXDqdr/iNKdyB7zGkojGDvkT
d4hKFJWABuROCMyQWYMZDufzviAFPm+XINuZPfjsaPv8qQzEkvrQjmi4hC4SM1LZ
SXHQ9DDgAaduefh9k43LQTzf5S0neR1eRrKD/FXyNslf2PuyGIJrCrmFv9VWp6BL
Rxm5VouoIGtmXht/jGItygb6hS8HWCe4OUMiTzNLGG+JFIMRyTTRU462K9nEmMM0
5uVYi9N7Rphki8k6CQevgQJ8qYAvtfhv/ljNpIdvqZNXyHfzZLDi5OMwvCzLZzUZ
Si7pxaGjAzsAkEPKT0joMffbjeYZazEXD0jb1SmsjHEqu8qX8wEYJgVZefKoWuPC
veetXTXqorgUCgnXqtFV0aMijXG7BddKMiRS1MiU2IMOwKg9A0oDdQNVK+UazOCE
deS+VWo7wSLbjojH8GYl+dR+R1oYlA7JqWRhNaK+jNVVicSNWaT5zB/K455kzsfc
zWFyx/8XevAiTNNcFz7QJkU/2TNkTzrInO5y1cJLeR4L0D8o9gUq5S+crT0ckK9X
J0d4qfcgCWVlfGl89HXY6iY2iNqRRwWyLZj7Ltp8aIAHyP7PBOD2tPGE5pdv1GwZ
djXH017Ru2/KFhBfQwfBUXPvD617o+bdYdeGy0HzCxJbnk+GxSAbE31fEv6UfLZq
bcBPHjjj96pZCmNigvqwBV7e2H7IIwLUJFpK+F5D6VLVoqNZP9bhSaEcMWnkEG1x
yxWBGdr7+53U0MC8D/HXaTlwG0dWO8UxxJSHCrcSC0LogwEKh1Ij31ZFjiL+l/u8
MRzcgBl0n2QkLPW+4278zfMUFZlGvbZLgD2ptJ9uqqqoidTpnpEDHJg6Z1nfRa7W
5pi+0FC/gMG0oy+2MKCv5UfP2zWzizeu57x/yzUI6ntU8y7Ih0Wdo62NaUYpQwEm
RuWG9IxYIHiW4WmRlTEi0TkqKwenDv9PI52pF24oPjTxan/X19137LKF4q+HhICL
GPY+M4UKnhteBMN+nAKRNYcWKpyLjuZXUywTP/rXPe/1tcxyYE/KYAWkSC+0y3eB
slFTfOGlpx9Xb0youXslDrD5Ku01ZGhugcjBz1MlPscMYkuC9PBBt1DJVJWTjO7E
LW+/Q1lotdo8RNHutsdZgShwhqCMM4ehY9mobvS9gZwLqXFRdgqqb06NnAz4WC0D
lomIzeKBdwtpQDjUxTYQXy/IyRFkEpa6f176z7BCj4KebSoPrHMXeaM2Hifdinsp
OWVFDHKqvQGSwH32L6/ZbeENNwjXkt1vKyHexNb74K1f2Hbt8QuxW0h22giJeTsl
Cd3Y5M0EdJc0Zw4RFlhkamtvtBc0HtdNldenV8Ut6KU1jdy4ayiuxZqjJiQwOxiA
27YaVKHM/vYXIivclyL4xkDWgwOFMtj+8s5KRzIiEiGepWPnzRmnz3+qMYnf+Pjl
GFyPHESfrxQvq15PMKEN46DEmCQasAvRH5ogrbHu0KPeysWSH5TJNivwH/Zf6bdo
yBbXVI+xi35RdEwsXclGtQNzRjv/VO5EDrhEKOyZ2Beo2T0P5B5iCfxe4KGOjlzH
BguJo/YfwhQNkFIz1b4HXSPAbLNvCKF3mBGdfLFx5zpzVMlfq3W1+UnItLjIdbYw
BOZFfG85swxM6F55MhvPqegs9dQCu/cJtjjGBvr5t+UlRt9DUO+1gTri737OopQL
5VzN49I0AUVh7+W3XtRpS+LgU8ilj3X+q80VKuObsqMY8lmQo+Z5hc3W9G9OHU9N
PgGcJI0Du8OQ7iLBCINCNIWigT1X9EDXBIRu8oi3IBqpVrVznihD81LEdtDWhWab
z15bg3BTv3umIM7ynNvFZkatWfXMWWFDXb+Hhtpi1BEzkKLRG03u/H7KvH8wS6x6
mBAfP7rFZXmzf8Fhpcwhqvv3RJRHr3NisTKHmQrmC3nsLkR8iQbiRvDbXPMuKsiK
OqyYaSpxiaHoE3k/5wvnifCO+qqlp0y5wFdEKABALQ3fOy5xhBNXECExcHO8qxrO
1mS1WXRfgLfaz7KUnWk+/GMjG/QhrmoW0U3ddSdluGOx59/U/fD567zn/a3+Mlie
tUBwjyoxXmzdLmPn7KoCd7gvhLpwoZoaf3GAdIRpdoIyR3AVw+uyzb682D1iKtQL
0TXdQjokypd40apK9yXi2cKlxtQHN/7MMbtmLgteSQKsDvHpsSC05p8D38uvpq7s
pmQP/CqF4TA9U1PfLXUMs41REBxC4HXIMiG+f66sAi+R/ndR9URP3Up3Gn2sTUyO
TwDk3BrSLTXygjT5ZSK0D863rO+ksFTYp4u+7FuoIYhkpsSPMFfdOH648HaydBC8
PDLgM5383nJ2PeyYaQC9SLduqREqmRI1p5nuHqn74GgpoBOKp4KP6IXGQxK85whP
cpTOgYNp9nOYx15/O5XZiTZTMbTgTUYnMe4YIrqOPdCVK0XPH6+/JASJVnUg2tF5
B4OR3p4EkfPPQ37EPpDDKybyQ/Wzt30J9n+R1CINo9R1lbLkflG8EOPA2xE9ohk7
RYxU5NtoOFufm79aCjPuD88ZA7fmQ+WjRnTJT5St8sdtvAvlwz3GFj7N3bRKQy0D
XzEKHuVNZJnLsR34bItGTtwXdmSeyvDW3HrFt4Jg/7PhJ5fOjb0exsb+1HBr3h0V
giMHgUFHKK1HiIDWiYUhf6qz7Ny9NLDdhuiT0kiP8CwVuWZxh8qbBjFeKO+T0JrN
kg75Kpb/s5awSC3moiZ5iqJ5ueCq6nt4jXN4CRvWVD+tfmwG2QepRPZ1IsZe3+Vj
4QopnZxPVG7TTo38ldhyVy0vcmPekH+lrHSh+2JKxKi8qCqZTPf8HJtazom0ku9M
q3AkKxvVJnSr2TJL1y98GjQbFMFohxTB3bHxX0wiIckjOKCbfUujyg0WYZzx3xqH
tYWE1U/xIFrgMuL53mVz0x6sFQpIopMTQMoqWF5tiqWgqNRSovV9xuIm/LSH2eM+
mxA/E3IKaqGIX2dKpmPZ7StsYJVianwfGf5nYcsZDhlAkkcjb+mkU+SmTbzRi6kf
n768b6D4rGZNTzMbIWXvfDud3HBHFTXXTZlejV8+fKs9PEfh2KvPpy8+Y+Ia6FBS
ndON15cNpZUjr0Un84F3I5GxsWD1jU4VLKflXNki8dx5kFwdIwWzZMTOIayt+5Il
hxyR45gxCbpyLVUziMRLHZsZbFmUi2l1Pwqn55N++IiG7vR2JT7/0dmJhD4Jv9xw
wzKecXFdwQP0hyUD4XBv7udqZ2dEBx9ACckZvpFXii9gVBxrdR4s9eOjoVeguG9Q
ya1s7ddbC/Ldb3FE6fmJ9lssjoxXRz1PQNcQorp/Bn+rt2OdyevlOT0UAQJhDDcf
8AKcc305O/4R++SI1gC2frkt8WaPFgs5NNpjSluHh5S0f5IoMStKb5tGVedMPocM
TsbbyXDDODi4C2esWAdKoSh9Kh7BnXxwbp7sovhrPcjvIIsvBKKaaYxRNWuzcj+f
XeDazMd4kbifsov1iAZpSVttdAChXfe/SnrEkWx6Q5RnA1W09hbIS7soyUv43SD/
aZtUrkWHFQlObOaZX3J/KYEbhOlcKIVe9Uwc4cdi8U19cGe7NvkAHK4YWiJkpQZ7
ls1RQ6ly+m+KNmQ5BvZJBsYxRe9G9Rqh9Ri+lFTrGInCVEAqAXriEdTFIegQTF10
8TlmykkJyOhl/5fpWE3iNsMHwe2ZNcTSikpamvQr2XpZqfuQ6kvRuSv+78zJ7YfA
qo4P44YPtj9zVl1XoowVJmrBt+I8Zgp6gU3qsyWKElp/MNWk5toNk8h7WZAC3DwL
1N46xyWF6mqVZAJ78POr8yHaBhB6T9asgvGqsT4raB6j7vsC44vVN+JtvpXQNSBP
NShGyzWeNe0jRaz5bZcCMQLbqfoT+WGEsQ2f3vkv0JqGq1NA3xC9qAR+veaguRCL
DWMwOiC0tpprHJ6tscHss+aiM874utgOOCSEMngvO+d4SoR7xexskvuzmmy3xEbx
VTgMNxAxtW10KJrOyn8GdZe19PEaJvNZvDp8mR/xoFx/AY+KtyOR3y09nbSUoxuA
zJ6boR0KCkDXBD3CPkV+PVcG9AJRuVNjqA1KHbU0cseDdi+9Ub8AY/vB4wmBVw5X
re4CS9DoeVRGBITWS4X0AuLLb910Th6vn6R2At/CNFWn7KK52ONUsmsNcATU7dLh
fggboW9QcBAglYlyg8CBJTpcy5wTGZKpHTGmStmiD91nvnOlGNfxeL2RdKHFG3rh
lhfxh3P70qACtmdu1sdvWfLm83f19yiW6Hdh6d/wNOb8b5+gFuSwWyAiczXvF+GR
s297lSOFBs4TPf4CiLLS+5HqNpOApTk2MjulrBYLNaJoTWQiwUR8nn4f2HCgMHAh
0gHAKMyw5CPkPr1s3GOFGrUQBFI9a8hqw5gH0I2mEqsxALkClfCKiQwnSdDbPCUn
fz/tEpwm+jrvuBRl6zKTLm6y0g9X0iII8g1nCVAX5HhmpxgHE8Ax1X5Sl4h8q+RX
peKRo+0XY46QzvTnFM9gguyNc85eGGHxplUR4GAmnWFiesVdCpQ1RL5R+lWDDP5S
kqC5ROsKtRDaWJYtZluJIpfxQjzeNF3tIahYCjujYaVQ1lGvvAdypOsBh52DGGjd
ADeusfW8L15H5WTOa2yTjbs/XdtSe+zNXdXoALrzUDRzgfbOIAivHyGeJV7TK5IP
VbrEcxtU6ZKqgCEUXU6EbzPBUd54h36eHJxc8sqBGwxnGsFRZlLYVc4ff5LNvltc
Y42msED41DTYJnKkmY5OXWpJ+v8WqHi2bMVVtFiuhS/ps/Ssbo89HT6FezTf5vkT
de6Ig8TexAFEjsHXDkMTQxf1DJpuvqs2zyY7JJIaOpH7oFs4C8Q9IBfadUA6WT0E
znFe8E6vij8+hspKXYBcDzjlemCeg/l9QhUENw85sSOy9/BYszjWgHBqEJQbEI/S
zONGOarowrccrjHXQDAqwkW2YKSLWIW9FUTR+mTzYM35DaGnZ2A+OCLXQVknKmAF
6z/onsd36phMAQ/xhKyB1EycNLB81YRmYmb6oPaUMbpl6IQAYZWiT2Ty/O9G3Ban
3EoB0Sp/RSfxtefr1OKaLCksCVM/dMsVr7WK0nfQXQsXpjeoEdZUtkFBDCM9uzLq
PAU4D2zFWRN4R0qcnlgCmS8qfcJCU2rlVpiFc92HQU8/12UeS9DWu4ixLGqwwfLJ
goHM/vTuqOsrz3+XF+Gf1cNKQL55m7Yawa2xcnPDfPjAeceE9IvaiV9CKAJsvd/+
bsnRqQyt/PHSXXFAHvFrMc4dcHhse7NgJxiitt4JJkg7beENwzZNEhKaAIdNfQ2G
/Pz/cClKQK7bkUeVx6x4+bc3rnXpuhXHB6ZOVuoxcchR0aE35BeWFHV9SdVJpk2x
kwrq+5JNATlHDaEP9hBLUyL07ols2PVSQEBl+cdI7U98BEqqey1WJIAM/kWnwYOe
mD6k+3ZRDTq0b60KD/39FLY8LfYRqsjHXUZzcImR7BjN1Of+2hE2JoH24CTOTShE
B0K3OCSPPssdxGlSvJDFANhVnddEgu03mPJZMUYQk3851RZi+y7UTm/LgboP3iR0
+B2K9oVkm4Yee3dU3YcDKZtYyaEyQLV3+qAQ59Z+Zm51bALU6do4E6vlBl3nPtV3
9Z5osx8k4J2Nss09PnwxbGGNyJnVFP8QzYDKUYNF/vMH+GC0vCKUXvO0Xm9RMLqI
IA6p64d93wNoTVzj45cT75ekTaSoRxsFwo+gKrkvPihDIpWz81IDzNHx1nCweqHn
+9bdSbLw5svfQF4kwK4ElCZTwqXs0Zy6H7mO+HxlP0qNvwr6sj+0ClcbGuKd+gXy
4Kv58BMHnk65OOf8gPF3TCOeDX7eehkKi1GiPYZNMX/OmXwgDOfUqcRcm0dWvg8P
kAGmWJO7InNGsOEYWu83R76yI4LRlPdfGKh5pA/YvD9yW9Q3C26sONx3RuzQTPV/
fvjQXJJGvjSytMX4huhr3LJdyAmBdnuoRJ0OF1qvWo36m6hNAX7Z22QXAnEfFl+j
3+j87t4994+mgChvJDA3UJpQsQW1SvRRIvT/O1Klp2o7/hSNtY1/JXqKAz7zhc+B
oWVYAkBzXdhl6VmFPRUZY/9V2v5fkWamv18pd57wVd0vzvfDV64J/X0IdCpaD9NW
j/aK5nUXc8/FkhKIZeyNmttZteCE1fpZ0CgrW5yaPywChMoZatlHWSqOqPKmeiRF
DwiUIYVoUMna0ngZ7EpliNwn/COUY3ClRtARwDemTXSgNq7FEIsd7JMSaO2nVAHD
W+3qY/Roi5dO+sKYZVt0lcwHTDfwdnbM3qSLHIfVZlDapC/s2gA+10+jSnqupQDF
eImF44bu1NLCSkum2cXo03Vbh1ljoTURuXOzrQL6x8OPH0prq8kWxFv+rJCI1ECq
0Blg7xGBqSd0JVRaKsWS0dabCB8N/gDkUnxrhNDbNgwmlpVGwAWbuDMumbzEPngT
h8te62sWfMCiU4GQ2C7ZIYqEddS1HDHxSwHNzwtVYuT2+TB9T28vyq6FMU5nHWNR
S1fwoEyuuaTnnRkF1JM5pyhoMehcL9H74+Dr0udxTKVPb60qUByiT22y1SnscwYO
IDVLJiQePXemoFD6/XpxCMyvhkCDdwl72Ja1EpO3UDFTRb64j3kRj4cIr4G6RX9v
YRWui70w1FSwah/f5MIuENSp6cybAsiuHXc0PXMu3zKOPz+bNJ6Y5oxZVvhUZjcT
FJHnWE0XUF+FhIwSmz88aiitGAE/h+XP0ht0zSYxNwzqLdRe2cBV+0rYTeSFPLHi
LM8cxFoZFqfXglYF78JY251mmxJTiVKMgIYTqO7QFm9r8sV5HhmfuALsmZ846kyZ
6Xnx/qjatQ2WjMbCnI77EEyn3SjE5z93gVAAoRBgCsbI9/mgAvH+geS3JcSpnCCm
ALrY27zBS9YkDHKDn7mS22H6WFkH7aB5hhpQ9pb7MfXyHSZ8rKxx5kSr1cS7g+Fr
YhSVWNymubdKgMpB3m69562uq22GVfd0+2+W73nOQJTTeRkH8OkkctsDxQnIpaS2
yA8albsFwICJ1tYhSyIhkiDEyGjpeX42ARn1ClLrc7ABx6yPJWg/0niRGXro37Ct
loUrKcpkiIC1mzmttqDdf5iwQDQBM56ducwxPOs9dAPCj9MO+IudsHtGsbbGXuI/
4Ok8jY7ZkLre96oDzzJeCuu9tKcdFoaONNsTsKF74slNXXNTw9fl3yXxBai9G5Ja
rqcSioNBkkcNaoT4Uhx5TaUhni41vL5IWeEu5TZxlwo9bLvTWIshNBoU35fw8lvn
L9wIjWAwDhCw7rvjmfXQvE0YavXSqLyw0o7GYMSAcPHdTbRkcBueD3bhdp5LQhsk
5PJ+mQOd1W/MYcuDGG2mqBNzalaaJEO/+rm9P/W/eVkp78aK21FEXkVDEOLy5Vmo
M2b8ZD4MfkdcPXtNuY/YuaoK/J0arqDA4Rdw4l1bBEqqlarMSTNObTS10HJ0iKA2
4mHDQY0sN7f8FfqkyLDPMAQR+1kqyjkZfAY0aWaWV0l8WFpsfvHzWw3s4NVX01KY
9n4+urpoWibeRJvMwyehvHOo+fv6SrGo5GZZ5elWA0Vzt9QJB0yt97BmQwRjfyLR
I+XA9fzOyJWmxnzrtgcDhI1SYlOMa80obFx2oMpro4O5921B5PWxZfBWxdZBbYrq
35CbIiIU6rlqPZ01t79q9X+oRYsisqQ0VJeBMAIjB7xZgVA9gYGTpFrc+p33YOWZ
Br0Yhp92gHU82Qc7/IALWpzpFD2fsNtiesBbi15+PiX7jkOTZr4ve1EZmuXdklf/
Y+w9LvCdtfEq+zApMs8Np5CBIlvCwmcakxEYZg/wpBqtSmXDgZD5/bUoqcMgDv7R
69NNTMOnJMke1itZBTr9AiR6KmyHs6bI1ciZTtyBoxr/XL6s+kEEC/wxaeWuEpsV
SqXBRUmn6+TW2MmQaXonAE41GUvlkJtADz17FVsaT4syuMTA+2YhDOLrCzKDXxI9
IffIMov+bp5Nm0HTJCKbIR9toJhld1q/Amu/kv+F7GGJaI9/jPvVSpWZhAuhlLDe
9deL6Va8lJLjrfQDXwlrYaGEQ7FhQ+dSR5vNaTW40qaCcWlDZr1u6y0QANXUTz4a
wsdHXDoGEG0yktqJz04VoyPh+ztEaM9HRo8gE7fAb2DnX9sfYv9EhCEDKDMSTdg3
Y07zDFQAOTKWLo3TC4nlSxtnfkhfv9ju+IwBbiiloKLMppdlw/haWQUliFstV77B
DTvmStkjMwEJVBegYxbDMj4GXrhZcr9aGKl9R4PAC9g1I84cypkpZjJdfdorZTYH
moWPXyOtUCTZvA0Z1/w0a8o8/OGVwqQOoGFVOO40qZFPZRRqRdJ7m77W0EKfWkZG
QoULw0axi1yQmSA7EDhFhn8+ISn6GouqUf+T+N1kzpnf+RMcMNsHTg32E4vgD1Ti
UKy+AsCckOzlTLlyKsxMmwFqPF8GXPKM413Zifaz09yLTp6CQwryRsvgONyi1/+l
o12AeqDQpDSVPuH6SzjIo2RjLfoyRhLxy840cf4rVmxDPhuS/UfN6EG3V/FcHjJJ
35UK8L+qbZjZXYDkIjme3R3JhXv3Su+ULzxegdueuV8TlXpkeZCSfYUecfqFiGf5
NP6zEsF1GSIW26eFAHE2lEl1NoUYvxAtR6JQCE/Mq5Cl6Or2rOOOwWpb4BGxkQx+
V1LFez+5ld1v5CFCt+efb5ExqJUAISbKLS0a8kjyZvp/vcwenQUWBwo0DktkqHWI
6av+NssPaOh/e750xGansX3U325CilXCffVDEk/FKeBXFsPBXgJNTo/9cWFg0W0Z
9BRxCcoEtHDri9L3bhibIGMib++7FlSe8y5ue7LJqe81czFLOuUr2Li3PCKCcdgI
WR3sdkM/5Bj0QqzC1PGlkFeRIV0jmQ0e0RPeZG1W7wN2ue0a3WOs9rS3Niqbx6SE
ylyX4p+QU3q20OPy186Hb47YD/eLFZiBq54U9jAyEg9DMW5Ncgh9tRxHm3zeyjwG
GCUTZMwmTyI81pfBIw3S2pQ08/xgvPCTXPiBYr3pBp1vkSG1DWSn/fCEI2Q9YhtK
c7ZaAAsyRX9HzXmA921OdbOjuldxtxiPczV7fHJ86X7kPV+nV4BWSNPMXzAxOJk/
LfLsruLeuRRvGaxytkCM+7NFBQAtiCx6Zh1UxD0qP5WEYLddrfAsEltk35K1Vuyx
sj7JUA4x2iswsPZtVrN74QUPUXL6OiNKuwDJi8HXv3bWF+hUIh39VSpyxAQzrGGE
t+SK6PpBjCe199jYlbCpUv0e1DXoV0hhRawSAq1o6AJ+gYK6odrqZaH9oMztQXez
/bbD4JL2U3Hg5nTuLcEwEhPiicz4m2e7VnNPgXihs7NsW6jTIJV8NY7DRtQ1EZSC
CtXc+mz0YZr1hlh6h/Q5r8s5HApG5LhqjoYBxXwh0iUVURa06BKOvoJKAEoD88oY
vowNnlsTfppjAaDUNGCm2mKEGdTu8b39/K8/VEA154uKz/UJh2MwXEREoClmPPQF
T06uMWbfmKzFxJFezfBYAp8Yea3w/83A+zQjj68G7/RrUSfIEusqmagGFsH+4eZ8
s8vAc8ZI4FEVz8rwu27xG2KpCAvYSz2bNiGrUnvtZwDcMjbLvCw/OffS4SaEijUy
L0ecbUOSv9YcGslABhcBYBnw3t8MsUNBxNtL36oKyjHpHiilkbvQGJcS14Le6RHw
cEnU/niMKhM0LVfvMgGOSEvBw0EYAzbZH+lpo58ecLlbVFiguWJTH5U8hwNpCrtq
+AMoulxwA/EUmo4FBXKtuPuBN2+lVvt86eFoA71DhzF9foNeP1Of8sEvKA0jy3JV
cIoU9ij/LcJJYw10vAm3Qw1LwoJ1BIf68O96A5jg2g5nqPtlf+fioNo0w02U9Kba
YHICfSheSxKLFqBMy6uVvgFs9XPc2h6UHhS8wVTVjUeflncj8c6pEVdOm00UQssp
yEodGkPFr5Uj1zVumSOQiO1hOs9uLBhJmENu6h060DtnfQJoPRn2Jgxy1GdaAO3p
nM7ud3X9V/ZTHeEbEEpce7g800XPbVkskk7DXE54fwHTX43EnZbAuULtEaFvepnG
w+hnfAAY0HKQOB2nTEX3ltF21n/dkCh5tgnqlVDcIXAsKSIIEHyYNkjFgRct9mZu
c4Z4TbIiT9SNfxBrcGtMhJTjk8i4kdUsYbSh7Y6fkOUvjxzgifGbDeZXD6yhR46k
x9eut1WGDW8mJo94uQIw24D+vPAGwNMwd7FxTOKGBbkK7qFNRVC0GJwy5Nw/t1I0
twVcVs7qFh49Ux/AVFKC8hSMBEB+wBQqnH1dTBV8dzMia0ot4qWEfFe3OlO2TEQx
lvc9hFNa5vDwvdR6d2UqnTruBEgYGoukLWxDHeVyVwaLgADnfejYqCQXsJfjasqX
+/EN4b2Fg2X+NCkv0I5bJwJFht0M3YKCEZnQVwsS/avAcRtzu7kR8nIfmjIQsmF+
DiVgbY5V4tcsHyLkMMBsZG24moSNQAP4QDmc2FL4sJAU3j1YPvktWiP/nhsWm/j1
rR+WGWABUGIFwXEkltiMarb3UYdf8Deqd4f9QJ1nBYej0GWvACpwiPeMQKM+QNxt
NpMZ8s+3S2wA/my9AZPTEK4/FKIK9HVtGoKIzTwLTvM26hlv48IJKB3s8ryh/Ay+
Q4Syw5d/96JlPK7Qp4UHiY+JMFoxaCxYMju0kBslfeN/5Hn1BFuDdE4lL3vphMEt
3mj0AiL4j3IqrEfjJbVMfaQ0AEQ4bIQpyYoslsa4wKH0OcF5ZjMMlbagWZo6Xgkp
jBtASEmYjB+KU2l1Zh4GS2U0mSVU4rYqvg8i5fHQz23vMFxw313T6CknPCamnhb7
UxVDOgDIH1CYa5Xn3VvBala7K7l3jhuQkAG9kFnZHMGVd3GbBgLOOXG3uQXxvHL9
CpeBmwNSO9tyzZd9p4EwrpaXYDRZpjxzpyqvKzUse63tqqs5qA87pqdn5B5k/E5/
DKAFYCXMvYwu/lG6ryVgSM5InLNhNyzpZu7eZInEQvLjWNuYht+hhD9mlmcy1kUQ
NIlADangSVQ4ew0qbmuI3t2gEq85F6ISd4EEz+U1mU+dCihzP0WIH5u7Naf8tSjA
vxTjqe0iWbVls3SlWoyrb+L+XZAeIW54AkqR3Gn3gRvYkvoSttGcNIQE+VTar0LC
6ePpHbC7sD4bfXjoAEN8lzLO79zHGbuRLu7z1IWGeBSScl1IRxWkdfTviPyECwOz
TT6IYXeL9B5qfMCces2RjOHW99sqkjf+dk/oxut7WFVoKlUrleDzKW0yBoD8AF1c
zEGTIefxKatO1rozk3VDYYZi3demaTijc7OB/f4MdniUPukcXX6NpwAvBH6L7cPD
ISgaizlAPjz7sEeSQr9AYWidyYbX6UJO4gyhelAFSbYczh3iWucGxjv4XagwVZy8
XVEylQnnPSDrit16UwN2HpNELMoqHBZG9GwLp3ZO5y4mgXn5ASVLL6aXfcHoAlJB
/ZXMa6UpDBfZpOKcXN9m9vT1oxsarhxcPX+JeHskQGk9Q01+ihSuM+Vk111Geih0
K3r4LoaF/INw0I392EbtaYk8JGoXWGdxwWj3AYmu1jWLWNeJDILwA0VKe3da31ti
4pDJc5y+cma9hFTlAnlIBe5FZ6TW+4RLQodDv5pwrfAZPK8vM8+/AvjQBQDiBpYC
jaFXN2BEj9RrgEXwyUG2pXrTM6q+tWKZid8y7zNZeyJLH6oYJgY42r84kSO4jAB8
hMG5WOZ05nvynwCMDKfVHGlSRqk0m1LFeQvdvIRqMBXKD7MZ8AP79EKi/7c6qU9M
jUKVCR0x8rKASndnYbldTT16x6YOJ0tRlWkbrD4bugJX/wnZ7bOimj6PmklE5GQq
J4KVKlQi+7gmJOe+t5mOLZqZ2+qlrbZ+xWB4jX5PYgnMkVXdckSbPqUUi46T64E8
2CsFIobB/3zdlolo3KFb8/nrxoTjl1dkTbnHvyWjg986o/a3m/zLCb+gObTuFBxj
vWaeC6UK3GXrm9PhK/8A38gfQihiABweE2AtrS5dH2ecB5iMT7gPDQzuxQUcxr7e
Lv7FrgSj6KUKIqvB5uhIjRDIuzmhpTWt2rImZbMSF42D8iepLWaunkqEvAwqJmYW
bV7L1LuntDOhkbZ+G14GDvCTy4dp8AkPiLYTxf8E2fxo7pzgjrY7GxUl6G3FJCoq
NZ7CKhSN5Wzd+oFy5HO3mne7eg8yaPSh7NULzYgyZJU2RYiEgK07pdIUVIyLNLuC
PjDnWPNiY6hxoQRSQ8CKLoE3Hj/mRhwt3fhnD5bWzvR2+oyPNF9yKJSYV6Txb6ks
DqJ2FECu1uiA8FcbZAZmC/lIuxghcAeOU10FLBg4mXRfO7otw0i1wVvNfVLjykEo
b0dGusWb6A0EKI+F8Bvkhrm9hS16MMKKvQxrYiWk21cbCdJW4zKW0sJrTLFkNjQd
HFvw4hv2dLVpw+F8SKM8iDDyNsSAjK6stc2i9PbQkGF9I+o2v3e37BI8cV8wehKA
fzG4ZCkvbkChtynSneSPiR2HfUaaeujiW9P1VIrlq+SiB2ucKLj1zR5KeHYGOUpa
Sd3ZP0bwEDmBB7oECqX7GAATlyYLSqhkyqifEOdgJPiomrzfnKz7iyS3xdG56Qsj
zJ6DeOI74KKAp+GdMnNcfGaDCgbRR99SA+sqq8wKNM0UNRdi+nwO/7KnJXK6wDT0
9JaXUfspBVd050zCo+S1gpxgiL8i7Xo3XtBoDhyADTWam0g6VDK+mV/Fa3DPPg5W
yPZOlhAEUnjK3yrbEk29dIxIGCwCLycMsjzu7SxQRVz7y9+V42vQpzg4+goTSoD4
U7LD+NwnNo8INPnp4/6AjT2fV8D5bI/z18U15bYrfSuvCcv1vdjYUWKW13DBit3M
T9+gxy4aKyVDj8cTXZfsyU/3ZGp2qFkchzhNYV0dAO8Occa6vxaBELTQ4qtVPDHG
1lTu0KzHbTowDfm0YW9783FuhvPdIMWgz3yZlu+MRqCqR5JFH3FVw1IquKEMicRI
uD8E06uEqIUUPoQEd8aIsAwve0eCy54qVRMhh0H+88rMPRQdptpuuIa71+I6TkjR
erFUKLwRdko+nL+HhBzdrBEdmX7V8j0WcFn6c/lxetQYnm5vlr2XMbewGoaMjzed
ZNPTsVz9xZtjh6j9qR4jR0DH6VLVtZfLH81gynsrZGKMAaL5ClEmiLgF7G44kbd7
77R+CUtYGabD6lP5hxFAwHY+JA8AXJ3n9f/DbA5ouveqA5V/BiPXv4Cxrypz+dFG
343CA8UR9H4H8qxSx8+JpKitv75SxwygR5fRbHo/uDr+d9RswH960lrz47CytyR4
R6HrkvtMpc9CUL4hzbcag7ZNY7BnzYNjc/Ycx89yT6KOLD2nPq1McaI0VWHG2h9U
XNQDy9M4fHqenZUS12bO7zllXU7GFdlgEVUxfpHHPLJp7+idx8xYTGre40fNlEyX
mfwVFjqqwiQRSEzl8Zk2iIzExHJUcb8d4V5vs5I3hrLn9PBIXQWlMP81yBmIsnm/
CQPjp/iYqhuebbVNsR605sNnhLYTIwyS7l/3WvfL3QQlE2avFPt3oGszkIna0w5d
HMvSB1ZmonbmveRL3832OxA5+dxg+4hY0eDTp3HRgQGEmQ7ttOcB/bvymcrszVxO
e+np6I4Q0Cyofza1WGFY6ykk2M/kBjYdz9a0sokchqOMlWiRREOEPNtLqVXKGljO
RT0HBEnyaV1wona7rBCXf+WOOWMr4gNDlESKmX/eW48elBWa0xf1SW4kdMgTTxic
6rwgSii0sGLOHtWmK5d39xxXlhxVyAbCTvhAs6hUecb+Ewj0nVm4UNWTE6sFP5fN
lup2MzWvfWkzivsuHak2KCv7+DrGIPUykzENLMltN/LCMd2bH/BbIZjgcO7d5Bst
s18GnCnuPBUac+aqgLsBT0ZF3vbeC8oYP626XLjVpSRJway3mxkZ6FPG7uR+/oMt
Bd8VuH/GpYsVo0xchPWmU5rGXQpUNhk2av54MMyH+MyiOEU8ScxjRATf6sPPvMxG
XH/qitUIBIdET73houKlzuc90ldWkviB+wvyhTLmKiFdG1ass86T/r3/9soWIB/7
B2k+ycm1+BVQM5bwvrOkPLHCChfkPJfhdVSkGRFBkonx8nlvkRuTFr+xifmJYfLP
tbcWW7iLTgge64QeaQRBsZPlR8eWIeI/e3ton+3ZDyEmsHyu0Ub+hw8peUtZ9ByO
N2d8T0cWqLwh92eSxTv85Q/DldaoB4FfZnf4wSduH/uCZyHYir9MmPz2yctGzZx9
qp8m21erRq3G3C0MFyl+LPDffl4NUnIW7Asu+a9wXHoZivyzLGT5xBhXQL3nwknM
XQ5xUm0ufSVYJwsUwlrrJIABCgsuy5ajc/AA8GGeGHuS/FSAMb5t5W7Ikw/jJABi
6ujJd/Hv9DfMn54+VxEtPgJOQX7JKIXWGyKemXj1zgU8SpIwCXV3x0FI5nC7a+B2
7c+UP0niwEzuG8Y4sYHQJJ+LlW5m2krIafcJ2G4tEyAg71mBJHdN2D7HsLtexdby
4nsp7NQaxA7rZ8XwrFfzwPXWZlHZ2d6ZGY0/RmGPlT3IRmp8ytZvgqMdlq5anNIz
o9oL+yKM/ClYx7aw3ONv+TGYNaHCimJUd8DunmqaurOho0oGpk6u4kYvv2/DMyru
6oUnChnQcBh+wqfz+zInNPA4Rmqjdf3Pk++nfm/aXZMQBqb5KXs1cgHnR6xlNEe0
bk5/WQA/Npv8kTHN/iTxeVLDixlhpCYgHZp3DzmH5SLlWju+9xJaEKOR+OBahdgj
2aRgpYgeOFL2klKWYCw3I5oN3qotomn4D8yg0PKHJOMMf8EFY5x/Kd8wVleLgk5l
rS2x4v/hbzLr72y4AtJVH51hwMbF+ueqBTUgNKipp7aC+RqZCBTSw6VLK2dsE1eH
r+cpB1ooN2S1lTCK9psksS/xqAE8vy0xigU6XRz1NN/xl30darjl0ldf9A7D3y55
Faxjia7uTYQhu/gRuhWVTpN5Cm+E/K3qgzMelAd6yEdk6syG3Nn46upLejaUycDU
Q8KgiNd5PiP23529vrwXhNH2I72OWQralU/VJOBS0TBpAP4PpiLQXCfRhoUkdaBO

--pragma protect end_data_block
--pragma protect digest_block
CZB5H+Ij0Jn+zSsYi+VftMz8a+A=
--pragma protect end_digest_block
--pragma protect end_protected
