-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
2Bg1DjIY3zY0vQCcrHYXCagvghz+FFmDKLrLMR14IiMyZ7t4hJpQtGpAJ3arfQHP
x23ZmVnCTV3Dhs5vnJR9GQjx7SV5mGzhuHPGIOJq0p6wtMAi5Eae2yrJENa32O9T
KduGEFKssSfncW75mpOM3I6KC786ncw1BxP9HWafMgc=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 13056)
`protect data_block
0TYgSqXecdjKrPUm4UMUgesb9upwg/0YSyIfNrzC81PBN/2suLFocir+om1gSmBE
A/67gVeHJTU8ACSjKIXv5TU7epYrS7SoBF8wMziT/WZZV/j+oXRjAXEgcxRtQjAD
94B4mGpQyswdHjLMHv6uPQ9tTW3o43xnVh/FxccYzhLrbuVNOXYC+C985RfYkRB8
pKz8yjMv3DY1WzfWI0OKPsj4WipmU5aBtImq1SEgKv2652IGU99FP/nnyIvznJ6C
B+URZkcIRqDrlDjFkaNAZVURMZ/oS8Za3zO+Phso+cQGlbDytMOBVOzDwtF94Kso
UVjMJKcUY09f72hVOPfVMgyyEgmfm2AwZ3/N4vnIWNICz6LO6m+o1RAJPZM49P26
+vjM1aHazK9J6STYDwiGntLS3Ayk99tw1i1j4eroBjESK3FoMIJK+wLj9oKMFErL
uRR4oUf5Ua2Q2117lKon+fd20dD24lp4w2FgikUl4tdveKL8WsWSkYQv+zQNn3rY
aufEeQXAI9FR2DVUXm4YvHrMd64K4pbLxnluINTHMUYxo0zOJz6ZxbNRpNHvIQRt
KUlZb/mqhymUT6e82T+KsxRFSbhpPusBMJh4wYim6jrQBkiVM450X5enUoaqJbgb
shXRlnE8RE+R9Gc2dGjXuv1dsbeYWh2WFrbzz0nrfuJpl0otOyEaLVCnFbuxOnDw
xzO2yujeo7OulSNUW4OO7TjdVG8pGU4H0ZgReqB8cq10s/3QpR/3cmClmIqivWI8
v/XX0BTpxu0OmTyeG//1lwuujqGWu+/iRnpdJEx6MPOQV9kv9GPaLH6DxGEgJPUb
KSglmI4/47mPdt7cGAhR1k+3d2zC/qajKOlm8v1fD5vId5yVxfP2LAfg2iAt3FiY
stWrVUwFNh5rRzAABAbU4DqQuQWJv+LgcWNRJgJIRjn040r5lPJypxp+YLDt4X0s
lowc8IvX93WVN71Gffy4G6zHkg297LaaWRCeqAJrijZIOE7fBh4XiNfiXA9fEC9e
xWigIvCbXKjq9Lr1wLyqcOzef6obhbsAPX3zfqjP8guGy1nt1QoyrFibfcKZH48o
5zu0dSp7BuEAZARhE68F6+6o8TG7xmBdJ8L4kH313IWZmrcG4vFz0J6qulWqPHLi
scWsME7TwS8f1kZJPKNT/b31Uo7ZUQHV4ylflWMttY6fjBgbLCzZxnIkhus5toCU
FG72JeGLsXU0e3Fh6da9u0F5hVzklo5PhVFJIpkJjjExhLqKieTAz8AtrPimend3
AUdE4wQSUII109ttXEfEGa8SpJMHgn1EpI05sqie0QqQu/yj+Slh7XSVOwCwrSwS
M+48/3o6NJlb47l3XLdNkClZnYR9LZvLR9+4moeHbr37dce41CcdyBkQ5jBgQ+UP
CFM00UPkwAH+VJGBliWOv+kDOB8UtWhwpeKy6indDyPAgGRXipZVuYPZQ0M0axri
i9H65EsgUWrvhrmlb3Lx4cuJk9cvQUF0p+6UlMvOhsiJh7GL1oKDgNn04d4Riq2g
yM/VblxgF52E1jfnpBwVFK2cOSXAeEpHOiTCNCD2OAXF1B1wFwFDCYbsw82QGZfF
wESBjhw4mfiLOugfl0gurIT07NbWo8ghaw+wHj8i2U8VjeMH6OIqeSihYSkXHKx7
jXqHthIE6yteZN8/5b8C8UksYOZQ5QMXRoYNte/TPQOCP0rY6P3S33xwgVYnRMh7
WdJhP00xwf8pPARhmL0Nfk8Vgnj2Iq9O+dsqIDCDJs5UTgjPfpUWrJs4O6b/wARv
3u3d2seBV3QPCxARvdA/EOgVBipMpqk/MnqfAjdwkiEnWdWDh8Th+7FNT3jMNvw5
8tG/zvnbIn7jTT9bTS0BRbQb5V8Qrsz1yKuMr+tpfjwjtQTtN3Vj6GVS0IKSxQD+
vWo00MpQd9Y1TGKrxlBNoKwtKDon4fSsPEE4ZkjwyBXZ03R3GpNXWhYqaNxSN0kR
KJ3WLSqX+AeW9uDa9Kz2foeOEpUgR51Qh4EGD4lqtkVfKP/SLqadGAZxNeJPJBXu
dsa9vMwqJAiD/S0DoWNhXoNoxUCX6xWCRNQ5V07lMv8NlJlInVl36gvt4KLEXJDJ
iICh8SPZ9yvPNX10Jdai4OhgBxKstx4OEREX0fUt69/D/p3Iv96KKXP8BZWpMJ4d
llfd8ZgnimnwHCVPBd5YuKZq0jTogPys7lWtJc9bJ0Rh1aDMn0OQ65Sz1lynl6F5
o9yvL9vtwVCQcWJHyRqcOjrDVwXXH3RoDOAe0WhZ1e+V+nxhkHx5MY+g046jqo4v
E/iHncGXLOo1q6eH88rgSaaYsQft2WQ2TQJLDAmXA3QdWlCbslt/agitr0gev9Yk
Ch+62bHoM13mlgzdN3m9ttHAJyPEEfhRZpvqSLB9DGAvi9ya8kj749ZhoJSILLoN
SuH9rz4Nbu0/yd9QwQf4POsyLA9ebxUOQxXka7GwMLeuBgOhKwNay6blCoTW1cAB
gtFJY163drdB3IqGQoyrAsDAC34pYIPvEmUJJmUgbgc27EXoXSun8l5sHNEBBI+n
WVpv3xxHKZtnfuC6oTC6UxBFbM/tRLhvvLcI2+IrqjY+6Q5+dBdcfErXcBJXOsxj
GoiPWR+MDN0iWyXR/0Rdz93FdBvPbaqTfY/0/DLpw1Hw2vU/XJacQQ/ky0KBEV9w
GVxCu+dgMsdThRAeaZtiZmzlWtFcS7Fkrz1oUKSoyrSWNT0HqJ0Cs4ofOO/iTs8t
SxziG9aQKVdcslQUfh3HuMunvQBVnxM+QDzApPAB56TEPJ07+HqsyxYRPg06vJI2
sIUnGJu62SIW/Yz6sZxoraMr8nZt4QVFSvNV/rskHtjrjnd9/aNG25e6/3UzYFKn
VskbXOQ+w4KzDQCAzpyadQ1u1+gIGzh11ldXcFqcPQS5JrqHz97xfpx5BobBV1j1
5eQkA5N/21iL/FZdkzt8bon3rBZQQD5P36uuTTAJUv9e29qiHtZddLsVwyBBvKIl
zDBbj1jCiLumEuqin+jgejscLQyFkqcgor4SzNU5TIRNzQRX+3uS5IKZLM9aGabS
0Ft+ur35b8BVf58dBTH73fKclRjjycK3k1FYReoAD0ExeeoFe7nyXEWbGALhT/U2
xCnyc41ctWHy1hTLlcgUt3ixvhloM6zL7qc253FWysOW3OnuMJMhJ96in33EWbj8
gtKNIn8L0IpWfoZzXS4IfR0YcG4SlGcRzFuYh5ralgwbMFV0LW0WwGjbcfSW/3IB
ZxqfI9wHtH1DGDKVrMweOlnnhpJ4C+JBysXFaniy5C8JdTFg9NzciMDhxbNk6qTE
ybmvUFnTLed+THTrMyj/a3PWwyZ3y4WFqELoJ6/QlRXHIbFFROce50EIqt87HpKN
p/fhFzJSD/tnrtUxeHidukxOA0La/5oRSRLdvKq/0k+5zRGjfc7Ss55R7uKYl9jE
8oz7V+3aoNt9taSep7lT3yAx4sGr+56HYIPo80NjJ6036RlbXA+Lo2BY4Gke+98C
elxe6XDosMy4EK/dNO9XlhMGJlAahqql+iyEy6eoB/0ZXvYY8IH7Qt5eZQsuhMxs
x2EpPU5HGxlBhtLl+BLliOs2h5WCYyczOSSopLxK4r6O8czEugI55pzwQP5XH38E
VmHRS7tqlwDLVGlzrSUcbPb3kkB3U6DznPFZ7Orjv+7zUCzih1L/PbVsFsnSpk6f
bUA/znie+EO1nagEYkanh6Jo7O+ZtAQPOcptvvCl7DLb5q3b6G7HPcjWAgQEbqPm
10O9u7KdTymIB19PRjtcivH+kkmXAMKfVPCBweNlNZ29ysyFMTjjXBERxmH2haDO
DcR3f71tk/Ic8rKtM7r/SFUOWGNf1FdGk7Y+UZjJN3J4wYaOQn1YvZ9YlvvIZ1qV
7qBxBNSjOyfHPco1t9QmTFRbW0vPKie5NoyoYQqdxhEp1rPTynF80zsr6H6wA9jG
vr+7nyF/zRBe5ibxC3YDVq4ykcPy8Stv8dNmZiRs4z9ZlUTKPy7V84zxWGS4cuPb
+lP1+yuodrWxqalL1s4tp0XUSiRNw4qEB65hB6zWmTpPwoTbzPOc/s+cQnp6ZRMV
vJSujqiyyXy1Y2XFyf+appRKDl5koFOhI0X0fnJsUb6zrPhTn0J9dlT9Ax8mq7w7
mGG94EKKnWQIlU0MZr+5aMS0eLMwCvkbvtSDU1wF5/absh5gOqzYob1QSwY8NuCe
W3vuMp62Wy2s6bK81D8QsutQ1iHblSFtauXKj317S8spQ7usA7iecTci5Do4Hx0/
89guD5/uLa+rDZYnCPafuuYiRtA+x5GTkw+Jion8BLcONGofC1lfMChyYu+v7IzE
1sVyihnOz38C2XQM3MtLvxh9D8W/htK7/p0LI/qFvYxbXhU5/nGaJuqRv+CKWLoU
iB2FA++dBEyNSlaIVZSyAZQHF2/D6VPxcJcQLolRSjJ1mAWVsJw+lwULRcxh5+2I
4dgaqhzyuupb+lH+g7htJpDgVCnPMwodBJBCAsYDBomA8tll/wrk1Rt96hlPjkyh
9/9XKRv7bs/1IwPCKL9P4ktVECZDmGo3rn+iiBYYZHTPwkMPFCBP7kSKgYUwO4cK
Mo/EuP4LQz2V5MHCI+kP/TYqS4fxcWz3N6LFxuWtLlq6ApL7nmuOQnsY1tM+sfoL
lVmlpXkXO1zv4pkb1+P5CUm8oP/+g6/E//KEyyRFiEiEvgbamA3Cm3hJc3kKR/AE
JgTCNOq9HnqPdh7z0FIQqx/x9Rtis14HLkzMcIB9ixJN/Q41jnAgCuY+hCBmtyFv
6oi2DviKCkTDFepcgkvxSxkldrTaEJgK7Y1WOgZD81hN7fINihwjf9BQHN+Sa6Ou
4V6amqJXEagW25y8b+dYV9SHP/ExFmjOsym7GMG8JgM9oOigCVXfhpyT3xlvBSEt
xp+U2jrHNN3myMfaRVXhOdwDVuK2/0OF7O9zotNIOeaXL/mgT8G5AmXO0OlzQ7C9
+NgwavjJlabQroZNH11JNUNvmXmqDBxbKEYtxAmf0qu7SD9+PDXgxYBIdPuwXciF
nJbYwM1C77UfWPtfkg+pkJMasjHNfpz5GRGN9CF57UgB4rCYSmMfIrW4PDO1Sejr
GMfbDcl9YkbX8mqQGI6y32Qu3+0oSnRYd2N7Wj2te75P8Uh71h5DRBBMjWBVHPy1
YPoGu9MJXRWcOaMZS4QjXqKrqc+tiRVOe/59p39ehJRJg9IOyyR4xfRFBcbhNAlQ
pspWrv/1DeFE8TNjJ5Jm2LVrdqmJFssZAN6aloYrQcAxX4iFYDzBQ/08ckXcEr1R
pPyyVMwGxcZMADlSwwTlObEsx2Vqz4JPhZNnuJ743zn3KOFc+Pa1jNRvL7XYvqZf
D4nZvuHMdiI+S9hQVuGm27KCjaS3WgZBggm8bUOrliid0p6eOKWZcVA+yihRVAEu
VIQFaeA4458UrEiFWKXFAnie21VNQlTPa8mYw8HFzMN9wjQ1KXFu19Tpbx/NYuZ3
y5MJD7xf6um1vDn6KU1lO1FaSCvWPhtOquPDSVM2gRjIBFZRFJwIN0rFXzWjK7x6
1dWu0RbywMBLq2JuwSjLD+qKULBTskt4DYK5LnarHx56q3noS0xECykbw9Ns5w8w
/5znd5Bz8ibYfUwBXOVNQLIHzJAmBcYzHwz+Q3xJX929Na/fUvFlhOjKMg+9zyKN
NgpDHP7/oOFRXM4doHem+x0JHdt+8dosQJT70P2H3F9VmTRoX7AFD9vX2jQX14Mh
QsAMsSjx/lBeAxTnIhnpxXGJAOWzY4E0Dk50kn73yNNz6ohYRgSi8E+A6bdG+25C
uh3UYDgI1X9hBLqqMkKshXvZH5+2j7GTy1nn9fXJ4wiBSPPKBwcrmyWxfV99Z0Ef
4nnPnYu1rFLZMJOkCoM/k1qUI/rPeOJUYhgswg8iqONFRpSJNDTWNZS1MfkM7QRg
Y19h6Kqa132Mdj7nji5cKfU0U5sGahoXQPCFcDsZkiQ8ddSkp4w3XeymFXVVpEFf
NZNY7hlJLhWD/l1/dUzEeyymuYcgF3Vwt90T7QLBOl28KYvTKt54yZsNBVZc5nlo
P161MIOh/T2yb756G0qWYzoynHLZZxQspLM+DqPnhRP01UNKbEIvhGHKjPwVnNZz
u0JkqR9ZGHaDpsWiaBhvaipWBTmt2ycXgE3jlrZ45BmWv+6ZR/EhxGiUMgOXMGb/
gNi7s9z8STyVFYLZoNyPoZUcc0a1beiP6qLcCcvXgPwhY2IaWAY6Uhyw2TktTFYV
EGDvBef8YAGkAnyA8SLCQxeqHui8z9tsO2MlgSz8LuwPGO1sIkLdbO9GYPwM2pws
gYYAw7PyJK5N+UTCH5bdJjzg1y9gThdWBvqot/V5DnmOVaXqLFRoke2akQtqO0vg
727eRRhK8mcV/aCIgMXvdZGJk/2r+kRKGCwBc5n1X3X+T6iY+C37WTF4Ni+MXojj
2sLlzyVkhGWdluQ2/OkM+c+bGPbRpzKz4W+TenJsJHB8YUtHqiNnW8cHxv5rS3Rj
SthHYPdIH4G74Zhu6pctBjD34A8dLBGx3d68VaodP4yvTrInJsq5hwDYRnKWwGlK
Li4IhB5vtgy0EoRbYaLBHIU6DPMtpGNAXPDa8AA3ruZbMCoG05CcBQ8fBDn5Y2Sb
WYLBVzcfXdrfXxo8ueqlB/IJOCeDLmeZrIxtU8rn5jv9GnRV6MpqqylQpGIEdajc
FijEluAA+9IH059GcZFM7JJe89HYo7x1Gp9qJB0rH5U+cmSzck5R1TwEpWcgtJpc
siMB+GENg8HA6TJSb/EKzUgnXtcRn7Lu3g8OtAANm805/dPXOdwrlbKXQgtAKg0b
Pm1E5GClyTjupKF9j8GcE8K+EJqr0RlJOC0AcG8RvQx5xdtboi5SiiMatvCmnkCa
yWYkOcnFeOyphGGYzqD61XKeyZoLBItJxpANfVU9fms91zWGqiNdlGO/6eMPqmpV
8SeyHTXfZma+syhfoxNpBP9LOev0TOx+91UPgQUQ4CUOy4U2+TC23KOpsbor1eQ6
RiCfu8HNHdNDX2p4kpaH2OZdSmNIUGLLMHT07FQAeMjA8i013irGl/iFfRnNLe6p
q317YZ9Woe/5nPcXjw3wPVFeMFfZfhLJ2KEevHnilgIQ6gZvctkRTlZteU8Gn3GF
k2p0rV6xE2mG2nHy3ayzD0WUXT0AvjvYQ7uDID1W0Lin3OhM84igaYJLCkqMoqk4
/iN9c8xA/1AL5Ev9bpQ66zqnkR/zrArmbosp4YrFyZx+MyIHOZY7j6JjmkBUJ6ML
HVWAs6MY4L/5cG7XgqnWzKMhiVy82w8C5Zv2q8Uct3VzEdvfv+YhIxYOi2SbLzxI
BPnzwZhM1gjp73RiAjgJNnYqrKEgkvFd5mHjlMhakHX40wnBoraFvtUpiW1VT0uA
UeUxL2P9nl5nWi/za0J+xxs3usRwLQ4vnryyiAuBTd1Vgd0M1tlxUPtkY14ZKElw
ZDYC2oAu6HStdVXv4/q5vVqUcgywkdSLsG9gfFmq0JSJsGZIquIKvDk8w2KVicBZ
gUXN9orfPH9siLbUQBwBgKUBFaXzUDUJVtofp2yFUFVewOw3dtRvRjwVtmq/qPVn
anRB/DFAF6+mNbHUar/x0BUvJp8079l2NUid0sYan9QK7LvWFgagblln9KKzmZBR
M/xwRVq4vbUQVZr7Y3+IudfJylRXVIG6zvbCGO8SnoCIAP7lJ9oTvf1/TTkmosb1
m2k32znci6fn2dGxV2sVgJPNRysEKY2Jyu1Z7hAgiXf5VAicf5CfCvfKDajyTZUZ
lbMd+rCxeBCRI5OOBAU335GLzYE0bdMXhvgkHG1sL4FSRnLonc4dcL49qeltPNJo
8cqeWRkeug1r+SWOaFYa4Mn9GRNN0oayAFwFB0DooWilKN6pe+bs9vvlGHNUnOPh
taZOsUOJ7VLYnWv1YptkC2vnlZt9O1kigKthyQmQSBqBgZhU6ZpqXXxSgCSV3SFS
jl5fTj2Jr3GxQyyO9MMrYf8JBW4j6am1UECXmy9j8I/f7G4ElE6U6oTHobYhiH2e
Dxguz85mtwmMKylvQ+IbzAGf+m9PecJT/xXqMLMNhQF9t9T2yugj6eV+K49a5KqL
PXyjto7ZmXGI0QR9j/HZSRM2JUA3q5pkhWlEpLr49A6/33yqfYWhIMmQbLBcPiwj
ZA9XBTEnYkaLDldKdeD1Dlqkzyf5WkH4xj/oF1swnh1lbpVNXkMi64vgRVRF0vXm
briLVV7KXTO5fVJ0skMa3A2gWzRgOfnn0CtHBDVhC6PUc1RW9SIKnYwW5ajlwxkB
5sszb206fLTN2N3gk9nM3gZLIm+C3wo5s/lc/0kEvqOy07UtgtepxAK8qRD+1FdI
N1jaZQTV2LWg4TkYCAf3z9eNq7Er6yjhFMM3oUSz6u/fwVjk8AJjN15GQFb9eYSw
Cgi1VrlK96BFLvCPn60Extq8WJhzPQQWMEaptZG8PLgPyiE/9LZN1vkyxHR4UCzp
zyF37HIu8WSF1DozKcOrf79vCXG0ztpcN6cc0HpnLtFtBA+B2vkTLP1pNFiV7gBq
pc6v9iGcNdUSXbnQlOMjaFrwAz2ZagXjCpIlvcnSq/vLWU0bZTY1PkhUfkbkgoTB
182odo5mh2h901blOlxURM58F6BJgK9QqoSZzlNrMBSlNRpgvLO/8zlTV5/kqjZC
S+ipYlCzk1JktAef9zYDVfqk1+PQrS2z87Q/lCf7KminZjfSaXehdzFen6Y5bTXF
qk/aQUP5RhheIyGw8mGaDYelwMz7hR0CTKfSdMLJ5J7CYtv20gLrjYZvUPI00OAH
7zzEGKin5x31RKk2B6aBrXcCDx19kcHq2uNOkCatNFa2bIZgACUI0mqmjOE1uMLR
AxO4JGMj1mFZ0PFn1Hsk3tL5MyneczG32YQGJlsaQ3bRJLopQxPjlI5cqGRMNHAK
opTPd+5SUV2Hf9fGhaQxNqGlHhbp5ESdZvvNBwB10CRDqBKDQL3Dl6P7dhXqWMe+
1yEhaNewwuEBT+eUkPnaHrfP1utFbSygNTo9UtlZr3WfD0vZfGwvSF4zuLvZcJf7
QBJKBijtX+PCmFwZo0Fl+SOYGodIODDuzlTVR8wNpCzNOtRIoEM29tAjywya/3w4
kCcfj6+Y89kGQrOjQGsFWsudsHTLSMpuaHLNUiK4umbfyP2JO59rpvcL+M+TV2aT
fOLrWn70gsDB3okDfbz3a5BZJ3Dit2zjkiJyk+iJ3LOfB1e4ONpbNhfeO0ZGXtaW
989NtZuJWO9swcbqsiGGG/9TAWEM1TbKIEIUzDXtyXuZoli3aOelcp8IwSWAY2lD
I1T9wRtCOt5YP3W6xdDqmoae1V6eyuCz5tjU5dPUhgMW1t9v3U33Crm9TqQl4xJ+
plvaF07XaX7P6Jgfwb97WOnNyEO4cJG9V1pziquWXRBSWdLkC4HqfKP9oGpSvrgz
r1EAEqw48pimuzUSu8pOp/EPeRh+OqUqR+edHn5e9yErdTr9MXd7q9j4pNCUAbd5
eJrhUPNSbnZ737UkR5vCv6Bzx3ong6bntMfQGtejdHUs5W53aWidwRdK/8MiusKf
ur7WiUXSPZvX6//KlHe9TmbQ4LeBNKkHlCmUTa2lv5uHgIgC2pVTNmNBsCg0+W03
WrZULuMnzUm1oCm8zmILDobD6kMjUKKqpoxByfZvNQgaPFTddv9899Ro6jfU8zCc
2HYJKUcGIScEJlokWxr2154H6VfHRrUAaFDEUSAPX69NK1YcODDVw1SteLJhCKHp
HnDBgP1rDrYZM5ZbVT3PMUM0e5HfD8LqbduNkQjDqiHZXCW2/UvKsSjGawhn1KJS
v59lJxkBkof7Oc//IxE8fOYMXpZpCJ3lGwX2D2L3Vs2AvO/6YbMOocIZb0DyG8kB
/vOu6ak5YdA3nWS2tnoqeJLTruSJdH6cW1+t1phhl8jzqnJnFNeQkPr/nhz/ao7O
R0WELbbKtcyjdnzmmtFSk7sk9/JVCjIQA5j52JYMcZQlIHDtTbdYU9y68tynP4To
CkseRp8EuYALdpkYw4YkgQAKYgOF18S2ESvc6RirrzqyIdnK71fKqxFtZL96h+0t
xuarAUOpbv3T6iN13Lhv+V5Hxe1ms+wz0gOXHgfKjUn4THyQo9zZK40V1ItVt5cJ
bI425AUiW6irWK23lPqYIV9ohxjr2BJit5KNtxAjSS/CRa7VgCNePzBTd72H6EMK
W0OYvmaYc/z0M66hmyd8ksa5EN82rILW+P5+G08fd2eW2nITU2GU4nluR9TvkNQV
OJ8uj/F+uij6AdlwzbmqrMbwfR4tlroKqV8tLOK0EH4fRtohipQeCGfC3OgDpU7z
ICP3GVK9TNJCw6chSH0Du/t/vpXZro7TlOZs5d6aGFhTAcIBwxVweDd07UgylfwO
/tlHH8HLefAEoal5aQnJ1Md+H6JiW+kSR5M3bGJgmONcD9mb0BIyYYaLfIEn6HUT
gfVFDZU2TeOmDOCjq5rRwk2hn8ZY5S4y1JzETExFaFIs6tsya0dzKqGGRxQvDrWL
ABkrTozVzC4aM6ybjVE/RmPjZ+pZSiZ4yMHajmzwtL04ThANlRiVrndzU3FmJPx0
eTjR12I0oZuOy/HhMXZqsrKk/NjzcHLkJqt6jpZY0qPrKGnVPE88e/Mjc0HwFVFx
kDEBT2b2IwF2SAKbVUVQz7FWRPzKltfZn4/D55UlAD/h9KLiHzlKJwCM4+qlP8nZ
h7jNUfVu1mUPa6XL1RtJkc8tHwMK/GZRmSC+9ngn6zA3f9wNqj70QttlcFwI728j
dWIm3hNIv7iA+hJ8qjQrQv+gfC11adM6Dy91vkIwQLVMjyJnO4Nie18lRBvn3x7U
smPJEFWUB5XyILPBoWuuBas42lK+wbmM7DcppzCMqA8Ow7LqbfZ+JkSciKSmrvTd
wJRab8XhcMA34PF7WAVWcmDEXOqtV8Rg9xdLvvOt7D1C8B+9j9qHIbeV6SbdSYxc
EO9098ZeTUz/dxOT46rB/DHXXeG7wIuT1v4zHp4leDlcVh3i/OfWUAn6mxFsGOUx
i9hTxrNCygWZkfQq2Vum3o4BL7GbHy2CziZMOAPU1QYjkP/c+yDE7psGO+fbKFfQ
BWbfYn6JM/By5cMDJAuPsTcao8weHwriVjziGoJ+iKQqujXdNeygs2lzYifhSgot
Vrbjr9BfrMkOMEAVmFSHxwqcwElgI0CvXhEiVCBRrrWFZp/48OL2HLPQvLnNikF7
qf95cfb+s6LThg1HBsdeGZ25ADt43ul+M5xr5/FZvGD3zs3dH7Hl9/hHTgP2YDB/
na8qMnQ12UIUJA/d2f4MIASbevuWBuqR4F1A4nXv4SFb9Ok7Ey9oKAexhQeuRYb/
CC8LIzzOs6XtjSY9S9DojDk4rqFgIZD2SYtkQysm6GuYo6QsvhxPLQBwwg7LWNkV
81ozGdDl88ALtq/1Pft9I20nqRGyO4KyJDanciq3JA6WIk707OiWLPUkjHTp8izu
hfPfdFEWUcFYWeOACMOGNoAMIqybfNizS9R9wScMdyPT7s/MTInbrexjNSj73Otp
vcybKkaYMyiqiyAa6FzDBAnE1PUSROyJIwHH5XBrpQrBCY2tjQ9/kKQ78/fp+ziD
rmzhZvvEcSR2iuki4Css1WRa3qZGuLtHsfuK04FcFlDjMAa0WcB0xJqeO0v0tloZ
oaeMe+6p3XpQWUgyNcrzIkqCzPe71693KdWp5O8dJAmjcC8dsIbYrfB61eRdxhQ3
mr4qds3DYtxaizIEAuXSX2N7mqqrBQRp2CtgKZKpZq293LkX9inZB/cMIiR62EF2
XFboRXEkEVz0EK6/Pv+eATWjkLFvtzE+oltZRfk3ZVvuBST3ITEWJyHFVCJINnLJ
n3cxS5wiwE0mq4NLrpNPygEVFh3/V3fru4IvVpRs5OgYucxjNe5Mm3lzUZmtDf8X
YOjNGXXXqudW9YESbPwGleM8PMamlOj2HCfmBCPbC8Taf2mGDxUcySUwiKVXadg6
8DdYptIRSKI/UTJQX9GoMQ6y/0aNjwYN05pBl63t5hm+1nxaERvuTMLKwAQFOH37
VGWBXWTEgqV73sHYLG+WgyacwwiRQr2aqFQqT+TL6f9jsB1MK/5O8VRh8SuTUBi8
KWCMJmHI4y10B7qntj15yMb0ekWk0dAkEGMKiM2rhfUB6edghEBwa/jzogpLjlcV
j0R3TpNqOIgyNNB1GBakS6BDRQxvUKzDPC7rtPhhWjndCURNAXp0RdXjk+6D3kpC
dcg6KOEjhYFQvgyrlQqRYGsSpVS9mKJdRuhloJ+OaJ0NeIejn0wWYKZulRHk0M34
DhmvyEAbSf2Oq+X2FqBI0mIWvTvoQnsOWrI+yAsDNFQuZ5/Fh7Bn+9v+2YglUZq7
IfOgCbjSqeO8G7l6vIZLsF7071E/q4le2JFK+0fFgSXO2Oea59gSDX9oFnFNkx6X
Vdyk2/5Xsm4Hw2HoLLRnwO1R++yTPRIiE1nhADYskTep/vI6vaOrevB8Yn18V2w0
Mdl4d4E2t5rLb5Miyw8azdmos5hEqPLSjpbqpkaTdoz2ZeoSjmovalCg1Tyc/gW4
DahrqXYf4PCaYxr/kKgE8C6100K3j3SlhjIg1WN5hOWmeD7smsx4Ra+CVYJM0p2m
WZsFY8+Y54I2jc4ng+EUFGBO6qLqXEPyJeqLUVR0ltnYuJJ5pb0MhSs1zxVdj615
EJynBfJYN4UQWXF1spDmTQ7miSv4xLaEcNqYo8cmpx3KLcfxDBN1F4oSXd5vJDpi
eldQfCbAB1tt4V1sw4N/XEgF+KSf6TekBVYboMk2pmJwd0KxvlSqAju0vlholptW
eJny/1ffp1sK2XPHZacfAwIrldbENh7vokwceMJ0y73MBqR9fQqJC6VY7nISS72e
COddfIRzMYtC93iaTU6hPU8lwkvxg0GxD61EBrTBh0pDY4cTnVw9J9S2nUJpMLXD
hM7GXP1HRY7Grt1n3sysI1Vd7aJvH8MzDct87mQ+yggW78li9OnWUZW2eG1Iu6tX
XoMtpRPaHNoxmWDT+wA+91Qce0IgkD7GLdunOyEHxyzzBQ/vIjiPgcNBDrZoBcWQ
ClOX5wVhTJWuu9v05Y1tQdJpincm7PpdEYxWGMG4bD7TuK9f242+kYEY78Ivq0ma
nyNPPF3/3xl4E5FytxE6CjZiRbi5la9prvVxcvVWZnH1gVwT+cl5DIbkqnrTZT4w
YpyVCfNWMxZ6RWEsbvnADY1VBD8FIrXLLRW8jv1LT7P40Opqe8WIqoHEfFXiOZrX
EFQ4XrW22Cf/+FJ198KPeWQem9wkHXAaL3pwosQGyVXOq3aOBUbq8eVxOnV1K8/I
ZUuH3kmSc/GMjD4wKWD6QfQZZnArRyAKB1b7OTkFZWF2nMlY7pLDz8FPuVIsE0eY
De13gkw75US7hJM3djEJmrE87Outx5pdYavPToSH/FeL164bAcrH9+l/NB1UBBZ9
GpzKlrWJTtvdBOP7FW0epAGBoWw6r9iwvyw5i8ncJ+kXwenn5KLoP/2OzVJgfnB1
4CV5E1UHNbw0gOwvetIpg0wAkgizfThU1XOWpRcD0itEKt2AYBVzHsZX1KtaSuA/
EatDQf5GPiVLN6RtCK+Vhz1ehq4UI4qBHyysZHDd5pp72r5GOFyVd3TBP+L6O46W
4Qc/PrTYzAGaRaFmGDu+dLZlnWCUMceEju3tkAmrw24BIQJ4m/kFlxpOEsFbFjZO
v+MP+3Z/JIhQ5deNMmztpc4OLEokZrwrGNrvNe+120qv6eyQDF1glormBfwtFAzI
1ISdGHxZweHnmJxHzLzb7R9IiBcgyIsNO0ZkWQdp6NlroC5ofOX1ZDvGAr7eWJVx
vLKjM5mcUNutrfPko5q01BijQqErWdjeR3d20o5TDcwlItGaZfJRKS9WA0C2MB9j
92ZPOEmGE9CnNzN/Q32MCoin0INpDXp1S0tn2gdUAse1/jD9kD1yPhTGkdpN0/LQ
33sUKpP6IYj0cldvD+Kd5NvYqDenItu0aMDG8oakMNThFtZsTYtbDP7xLyseo0Lx
daiJFnfYQlN9MygsFgj6blyF0POGat6qCLB0wBQh4j8dU+4gAxQh+mTPrWu5MPfn
ZvabrRjB+uwKCtLAFtfCyC5dHLmvMVOZuoVXEtFuEN2oqN5aOISrKqPDLdVoQ4cv
/kaMyjcqsxcJZUxCrVnCCd7oAtyrnHuladHvhKnuhHMleQEgzZ2xfMWy5N9eMWxr
u70lMDRlu6JaVMRd1JrjRPDWk7La1iQ4UQrX8sGME0ACJxe54VvkRG7DoXJtZKvD
jXDvZk8cE3vIYK4MLvrzLDxZ+wXNDXd/+u8geXO9Epu0TOjrrAutl7nG2AU1DcBk
KQkCH4hNzK6eISQ2JkezAmHXU4KHQZgH1MPdTdjZDi1e0kZDcJjRk7chHJ/TWdEV
PUQ1mgwgXQP3UOUpYC1SPeJ8S8eUAeB30j7BnS2KTnSvhmNEIpPOcByMQSP6N8D+
SoPoeakElK5aE6/domIrAUmqkfGa+owJe1xlk0+kUjbP9k9/ef6zLW6rNnICUepF
D2/AIc6dAdlKHSKQcDclRnkh7VcNxQJq5gmj9Eu+DnZgskdnvoqjyV66CSIUlxJw
k2okaPYwA5xkGf+l2NofiKxCMz+0PqpFR+7kvdfEJH48GKUlZ6g02se8EOno2u2X
NWg1pb/8zUqe2QjSKLteKOPIdRb7+gknk/wMSaq+5rzRwNE0u8NDYpieSWNGDtrq
OSbwmUOFFqtYKKwhvd8Hr9VM9dP9SfHDJFhqU478MPdjDrGz+AjNwD/unzR86tzo
SRj7Oar/Oq1QCcvqeiVx4ty9tjnKKb/fRd1tSW1UuHLIrXdg2tvC0663xM5F6I0O
Rtr7dZNZ3StTff9UDWQ++96cIS/VGjlvEEb8UEhHGQEeRx36Onb4IvC8iEN4zENw
V90xQq86UYZ0lOodv7lxNPZdX85+1x/YsytLfhMZ2GigctQTihfo1GwoOX57Xxfd
JxU077oocag/d00N/oQ1jevkbfyISSiOBzYr4OfW2gE42QdEMxe0EBmsjk+Dz3Zr
ugUAWVxFdW1y8NX9dmBOo1ZY//oW51Sdo4sD07oMT4Ufzk6xEoRq34cYNmUMWX+O
G7KJkS77j2bIAlVlzwE2eOSIhIMHKmIo+ZTS5tg/u9mKiru21MQzEVT2jwPy22Wc
6FxXp8XIB44Etx0hK5RWDCixllvpUy/1UPZfUmmnwKa9LZccfFpJwZhzdvzEpmVO
PPCTOizt0DjmDRfpaV0YQR78G6/T/v/Lt0MP7oDrpUlFxY4cSVIL3NRwAtEbyRfP
7femtZ1Vlu0IFBEDSvZL24UxfPsOaDUNZD1kJBcudz2jgUFBUmuX+9aVT/FvAeeI
EmhSaETAQDfsZQecSBFrCJH3hq8kzJs3tkWO8x5Fka8vX5Ai2DIGApjwJeXSCm0y
Hm/tEDPJnWdLymkwox6WX1+lEZW0AqDHJHsyBXgnqJShRBGqmWevD/ZfW5Qikasf
ddkilwC1dpKMmdiGoJbcc+ebakscCrFNeAeWH2THT88OnDbbc2OubVS7KoUTxdn5
bbBcpYLmDSTjnxFLzIgEr3eV4oudTSJfSvsP1HHdgFbvkQOYd/UZQHgMoZmyjLbG
xAqD4b0c8+LbJfGR7iC+/BHxsT0uj0uj+YKxMgawFs4YKt2JOCbQ6hjhhhS53Ij8
0ox1747H9bbf1pF2SI0p+23uRDCBZh7h0jHouB2Wmsl0WdHRYl/VKXO3O2fsyn9M
bmeEBuXO5BnsDkfEQw7C6JEaH2AJ+Yq4HhMZmnrJrXaTDo3QO0Zkt/aO5K6mSsej
eZOax6akkAYFlSL7FYx6ItQqrNMlTntlXlfqXZyuh5u8DRw3GhX11X+NUcKTNnEt
bHcEc+JNV1Ug9QPKtK/7stVZixeaxq0yMacgXfhMDQQd4vAZXTeLiiZP6ulySijh
O7hxgLk9ttyimDtyso/+gfPPBwKZK6vU2dGGxj9Spbyg7cnh9nJTawO41kIqjGqs
CX37nlnX9+xpNvoBbaVZEhydkXl35XBS+azejnJlrglvIUlB/o4LIK5au0SIydGK
ISEWSDV/PUikhcP3cGj0aSFiXBbUGwHa6k6crc4Cqdo0lE6wVb4IPgOSoB8mePie
T0gudkLls0s7II02W1buK2dzX0MSEnNb0Vu3543/0/SaTyTYSN4Lzd4waW/j2lrG
edWBf9kc6dZkCKQXdKaeiCzPNarEItdJ+/0sD56NgzCbl4zdujiml6amLnfCEAi1
vOLgG/H3Dkd6bTGuSP6kyeFN4E5ifYGE2tihRiaq97R+azI/NIZUl358aMpkBYPD
/easLmo/R79fWU/vCK267Z2WgfdQsIuQKfXLBbUVa5LXt5GpZMlWEjMA8p3RBVzx
sGi88Q200db8xsO6r1iGt8Y82Lr92z9PUgYaGGnugJ50FVFLQI3M2tX2I4Wa3sDY
LqWcgLN3RzLUEWS1lupUvY9++79VlN3OLfGSFuhzR9Yc1RAKjnpfQfGqzwRq9Loi
ZEqZtks6SwH/iC5B2Fav2evcOrahHwylE26RQHqq2dnIOIK+AcuczImwOIOigVIC
hdgRiYHx5YWTIzj/igu+Iox546QaWfHFL2s74LErlvHbEOfE98LxF37xXfSWsXFs
8IO4fKsIREs53TQrEl9/Qx7fB2ZPX4EH0cZ6oZKqxXkFxKog0C/JgK7wVWp1MPXR
+oEMLIxAnawYAfjJKVN7QodidaJGRH+G05R79tNzzKOyk6FuwdEAq2fNK/ccoOXN
E0YDGYw8ScvhYovgp1WAo/UsLtpYBFrAM8NrKHe1yo4T479McZT+3V+Q41fMQmXX
UU3U5Mg7mmzH0VedLPloOb4G0TKkdQ/WNNqCFLlXPcmqOtkxwhbpcW35n4QpUN1V
RTbhzCZmHGoMN5zdFOFk388zffFrCzWj+B5qnCnj+5guTbcRRl62mLu28U+cVaA3
bWNZNo1DJC+KaAeHwiHyNjYXNWablIkDVKLfPqqvS3kXMJF/l8riSKzFZKqMnNSc
0g/wSfPRjGUv2qZJfhs6//z1n1Rl+IVAHpSPat0Z9HnlwjRIbNjCTwJ9vFX0Gr7Z
/bezOdyCkARt4KjUhpnniRrYFYUybvR4i1TpuMKqwgOekkCcrmKnume1UflbFcaK
GVB+gZtTzjRcJIxcMCgRSFpyDGjJh8VJM7Kmtjev1NegSZbkbOUMEr2X2Xrqfte2
tbm29Wp2inH+bWl8LnoZgVXxzuIMVcjUgzHELfkvM0I6NY36PM63CkNd+EHTIl13
OaNycaoev1kFKJui6Y3GDP4+cKctcGoo2tAW6fpMvTvH5lFgeNerHlFS57hLjmKV
`protect end_protected
