// Copyright (C) 1991-2016 Altera Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Altera and is being provided
// in accordance with and subject to the protections of the
// applicable Altera Program License Subscription Agreement
// which governs its use and disclosure. Your use of Altera
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Altera Program License Subscription
// Agreement, the Altera Quartus Prime License Agreement, the Altera
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Altera and sold
// by Altera or its authorized distributors. Please refer to the
// applicable agreement for further details. Altera products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Altera assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.0
// ALTERA_TIMESTAMP:Thu Apr 28 03:59:44 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
lme3aImxmP8krt/08W0Ri8no3iPy5LfaS/VCx8kf9u3O7GRO/mX1QETkcO8e80Jd
ZYFlpONUQe+bY6WP0Xwy09Mz8fM7d3KKinDFwZHP/yps6e3vUWguIuHxeleEIbkR
vdIeqjRW+oZzvpciU4OsxO8wcX+DA04czBNc1/92Rmg=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 10464)
btp9+qMCknN7P0OFYX7D6IBwKWUSGigBA7abEWvLW5bKIA2b88Vzt/d9Jp+bog0Q
QBm2b4zMq1xn9bAfvUhk6q/3ixFy+OTISjodw+6RItL83ksFrfHRGQ4YQ5qj9ow6
Hc6aEkPqgnicFx1ScHvOy+vhI1cHUEM1yBacMEfA/g7Sys4L4HAr2qtViq5oz0LO
1ngeLwDl2cS3/OM5JCISNzeoZDL38acKagzL4VA6cqtXoHDcM/E7mMVMlbD28nkS
uVJV1Ra4rvSNevCmxjSdSbDVCkIEY22zxz2waOhWl0o/Kf/CTGatHuPMkShPTUl2
xc6RhZ7J8o8ZVh0k+hmDJJ/tH4QRE2TqX+AnPkt2eiwAI+zz8oy907xRr+C7w/XE
igQGEAdjE7DVu/6byigmWHY4+ULNW9fCKFZNvmX/V+RoJxM7WXmALJA3xV0hy4B2
YpR3xullmVf5C/L3evFXH+37tGL//575//Eu5yFOP/G06wDEdxSdKkznR5zPxM3S
9BfQ4PPMR/F3+Z4ZPcTcjxIAH1vb50QTndZGwi7wu/o5pF8zVBcx8P/8MIGpMqj3
j8Qnno4N7MzxXT3RcqUZg14CHxKsqlBO/J8DolSjJPA3cAUNoDutmP0VtgIc2YiP
jQf3yYaagM+c5DtLf67FYb9nx9ZYK3HZMiIwdqSF0HedL61QABz/hVZFigQ00sCK
mag531wj/wVrf7mI0P9cTqL5PcXC+fMwBqvCoLQJ3HhRpWs0N0lWTmQwhOa3lshm
t908skcWG67tx2Em7JAZm7ERVrbfWb0La6gbRpc2AuprWsrTB1Sf/HXEcFYhmwqe
MunQNZVAoPrvo9AaMon2QggfohKCviakuosMEpseKWVextaagxJqZbaM2yvA8Ept
TnX/X2gWyfclTM+8GFKfFyMLHNTCdrbyPMylo2+3uNTSmoLtgkSjHHXwT9KwB2T2
67pq5hiLplhanlZIn+eli6IqDnM7STM89KAtxwy2ElI2jPKNT3hSPAQPHDhSEk8t
2ZMLxfiipv/kF0mV4AMuuFUQNUN+Yq17ifIBDaSQNBxGrlbp9HzwCihaT9asvrd5
2IuDReu4AuPxVf6R8RZVLznRRQp9rbjop286JNoqriUNTpTqnZmG7/lxrdABRmmo
S/M7uvrDfDRGD0UMz6tidnA5j0LuiIG0ckuJzSL/yZ7Sm8/xpEb2CGVvLpFs0TIr
nRNNdsFAzvGxv9WDPc2VB0SCULuz+QCTb3+nGKSmlFQyZIofzdrCKp3f2eJyxIDz
mChirMdYiB7rrxEEX8klXApjbFzaF6IFtSYZnNk6WbVNspQfXzR+Z4hXKyl5qJn5
bhv3I/gQSdFo8Eu0Myi3uIGb0/p9nNUZ3VLRKku3WPEzjZPRW5pDvDXwPGpbDN2L
8QzGhS5J2DWJDEhs3y/vG9CUFUTUO4wP1XW3RHNvEmyufIwCAvg4T8TBfciTxLME
IsBgHr7R//f0ApVdLF+kqGxs0k1Od04ucYmWg3eaA7FveRhQ/gczyncLzQFDdoub
ueJm1XLuVL1/yp5w84xostLmSn+pHLKx/W4la+ehmO9M5FEEjrQ8Xa3q64dyzr9f
uarL9zeFe5f2wyIix3iyCOq3eQWl+70ULscegTyf3PoDQnKCSu4s7AHOH3QXiXTN
kpN7nhMkGD6r5dx1l/0P+vz8JKpCchYwKrM2WDq2iy/BO2eHw45Fa7/D5gaLXVez
+rh7ltgEPZm/WeMCvKfMrKO9kCGen4hs+P2605QaekvETDeDebg6j0pES5J9GFCQ
//lo8XX2ALbqVsL6OPo5vQuFfGglpexs4lcSsY6C5F99W015mlN13gFvT2grcC+P
eT0bWZKzXMeXh50kmMbEF23TPxXtwQ0kHYRJ8KG8tsfZuEyQHv1pnWR9zKPmnZGt
F3L2StECWOl9jcjFOmR25ANLsj/I1x1m4nWECSzIwJ6G0HaQ3OhxVYtFdzLCly2H
4HweknboBBgc0wHVtEEHKYhNZnwibBX0qMDFpxm5P43sZ0Ng046D5XKG9VZv511i
wl8F5SzbLR5xuIdUj9a8gq86qWV5GmTXRoKzQVlQvoyiJTEAAP11k389nJakPFzW
7LvgwuCAtTlzUs8IvDr49vqZjEiJMHDbHsHDWUg15sKfCT9YBChQC0Af5G04Nu49
jz43RuMHJ49HfpG27y9bvIT73zqIErNxWCysSKq7FefuH9jfIhijBN8Iat9tB4fI
nIVbtbCFfse+RU3jAVWRAsLlaLrjZpi7g1JtJ3nA1NmeqonhhLMhmyACwJCJvNRq
BzlKknvJxDu2jFDT4kvEbhMypQH4zQCeLALdsiKPndv5cn99zLfDUenYRF8keK5y
bIVuljjun/2MXu3em0vh4Bmqsx4z5vIx7RajxGAphjYoUev2ZRT7LL3Nibo7ikxT
iN79H01GjEXjC/boyGRtFF0JyD9g3OJbvnlG53Sdj2hNcvXCdBzXkIvFBK2BIvU9
57wzbDtj+xvPRioI/fkYvFsDE7yn9XzAG19cMz15ltbOQWfz30f5IV3eGIu4v1i3
67iJs3+1yrpwQJtFbcMjsub0RqPYDXzBEBY3t7cwD97FKBbG14iwgEs8UMv8fnJH
q8J0jsM++eJPWwJ53VCuCHaguER94/lt0UKHO01bkqrtaj5fUvu1qT9njSKGYPhk
dELJwY4gf/IWPTV0v/MsQXON0V5w4WvQpRnIpZQFM53uUKqNNrGR6AxyWHWBZHax
EAapSpTHs/3WbjxtYZxddzSe7mZRNyhU6lclQgjuOQahmzSCBEcrsjypRaE3Hdq6
ajkL3/fbzwkmnzwVM4BZKsLeFrGUHPCz8SM3PPXq6/2cbyB9Qpnw/Hg5WlELJtAO
JyMVPHEjSXUYytDy8ggMphWduE4D9zIXd/tVURpq9DSm7DvjIyf1B3Y69F/KWuq0
WIsIUN3jayYluhsHEL+uIr2BwdjIxD2bZqbKLP1IFKGDWQ1pXO/ceXyzwTBoByYz
xQrrbD8CjZqMvqfPx3Oc2A8VVczNdlaKteI2SWuhkiZ3ey3HzcKLOGZi4L/LasEc
G9ZAIeAZ9YLXd8V1EwWCgd1S1KXVB/IUrcdMs1mVYmCtmauBLjIYxXK29UP73+Z9
5tXqszuOWgBzPIf01M8SWxLEuU1uXpRPVeE4WbvRyFKJhpEZxFU6P2t3n4U4QbbD
1m77RjYvbs+QuIV/e+jktarXv75IMTxxUlrspRn4UJLFcx7wM+S7UKXD4MKvy84W
TbJCVKEc6X4brDndXCzME528i357zFoir21CUs2Vp+Np0MYtzqljdRQACcZaJe7N
v3qxd2s1dxKPWkDjelfNoP97aE79+aEVJ6NM6YQg0z1hRgJLVZx6AQar3n5CLU1i
eX6gzpWBvR+l0KPk4tuBMsRxFojxQAk3NChmp0CmGTP1OyqhrHHJ4z9C/C35ZJ9W
hEYgFyThADUQjWRYO8x/R9vdzTbDZ+KN8jq6JuRqcof4+22mmKvk6VlpnTfdWWai
WKY7OJfE9nP92DxFShN717q7/Jl34sVpzcYWxK9Y3f5HMn+R6bA8NmTY36Dda3Tf
YaYQ/I6CXZIRnr6tLFFR7PZeE0bXsiHhU3u/VLrU5Aghd+hRCwsKViPt8p/BUYC6
s7DaCrTpl+sejj3WsetNDYePh9dKwWePJvogDpExSNUV+tRM34nV5S5/j+wG6QUh
/sZpJm2PIWXMZqZAHM8pA1spz/dL+VsZuWppNd5bfzagbbdeH7IhR582vGWqw8E2
VIcgMVS95CSrtUZN+viJXU9tGrsjclcaj9bz5MQHtY6sryd2ROL777WbM4MstIT1
2AXVNAWDEsUpHZhWpff9mCpl1RLxVaB0B9ttq39A2lg0QOq1p/Vq0C1MDJOCiB+R
Usc9l7rXynMe55loUQDAvLw0f46qbToY3Ro2DUj01EzkDCswKVwkDsO/RqaGOSyQ
RQEA+MBxwmUFA6hpHBKWOPrd7sLi1zwPSV3bskZr27FVl+BFtUpvHWVux8bJDtiA
SPw1OkuctrnYWEneJUJOovrNILQkHEG0AYhuk77yi9gNrnvBRrMaDZtJGOlt67Op
w1aAYzwCHg1g9RtfRQnMkFdP3Fuvtzel2WDFtxaUwqr+nR0DxSfJvfuvz/GkR7Zy
CGj0BfChbKJGaRd2rjF+/wThmTedteYSoc2b2KckW9RUosRhwvAQwDoJ0RXV3tFu
dWSaVNZqb5JO7IwakqP7J75XFGsrL/81HkVLXg6hT5Gbfo3KJZ08IIG3Emb1hHuH
y0ZraVM1G6IWsz3/unNOzmFdqEZxZQl4NNqb3i2YQrQxoUok+bxARkEx4ao6IpAY
7r1QHSsr0RSXbmIAY++nZndXjAiT0W9VqYZEbAmklyEGQKEx1/CC80A9+Ear8LOI
3n5TK/kElLl8yr77baLwIqGDMM2vWHRdhx28NNBJDUW99IvP7Z/23bMqK5xLSjWn
PxEX22NUSTINejRD+/fLYP2x9dIO/AXsFDgTLQUuejiNeCRByhI2r3DuWXVtjMsT
SiuVbtE3ljbxd2/mbKWIWLPbUM1bYbvDE8guDbuZAyNImSUDeWNYrjs0jjip18N1
jk/Tt+lBtlePCCLVvmVyAt4fz9CrjrmBwUXYQB+CFAH5DZUUusBbP9DJLi2jV2FW
J5OFlo3iUW1PBIMdtM+UxtBCfJVbgoNQgaP2BDfiTCt+uag7w0Ug2RHBsLzMly/i
/VuOU96FnZWa3NIlKyfzqhKD508Qz+TkUhHNBorIAf2/TnkeaP8WSsOVlaPaEgSr
WUM8BLbiZ/m0cxDFVLQRSlEp1sSxRCeNRTtSSD5Fsk9LnsKC0TM6aU6ek+wu8ZPy
+sUpoaeoWI9UN9qJGaU2C7km9iE3jaaN8ilia8QmWd4ocCSfREq0kGxra2orBkRK
JVi/iz51NZhvL5pTCVj8sy8tOdg6j7k4mQAHnORS3WS4HcDUVNknWQd7ZhJ1zkBy
Vy28NIDCItPVI4BIJHPCqmX6UnbQkTPEAMiK9Hmk0Eh+t7CoL8eZXg7ttujpnGbG
37bcrdvrGH6yBmfNiq4Zp5F5u4k7RrbzxsnTWPN5HD4ONrLZLtyWUG3z1i0knQ8E
wYOqP/Z6i5F+zvo4U1z/TTRbKjtwo2pnbxJ1EXty1KpopBcn3SOw4KGLuOf4quw9
CPJJfm/dNMrVjWw24L7JnsSnqUk8AoWRNeyUc94QMSFySR+tSihN4eMtl6VHkvXE
CaTooDzNao4pLpelw80F1+t/7aZexI9m7dtVUFp2yShp2YLUg1d5+8ewbS5VfoMD
KfHKo0o/r30pSLDudyyH5dBrruCCMnL26I5ij1/Uk+hKKoojkMe5yznBA5Yx0q2D
yR1Qe20C+whBTzPGArr8ezF4guGXib+XzZUCnf2GB6/YaCgs4mN37N+IWEU5h7hX
s0/N919VtQIcLZmkyYhtMNAi1PMe/y4GBPRr7tes01mQQ6Nx4lVcazQim+oTW/6V
pZIa6m/mrrkKONzFxjsdKDgIm4wb9vJ1DmQ9b4k78PyPKW1ob0pWsx2a/b5KyTA+
g+y+zUIe70NuZPd3CAwMmhWcPSXZ2WorfGQTXI+T//qo43T7uWss0S0XJ49wXJgj
nxE620aDNCS3ZNfKxxn2a6GxrvYCqCk+yp6ygNoXy4SJ1yjtRUNl9NsdDfkPDiVY
Egv/Y2NyDqnVe72/mfB2S4nt6u5vfSMppswP+njv6uVGQxU+JRm4oQIqgYHXu26S
KEtU/0JgowuVIjHWX9Kaj/46g8m4jM/GY2HmIpbQDw/OaSkByoGeYrhchF/cZS94
qk/9p7RsxmCFSfid++BPsGKZefPj1pXvc9ycENHT2CPp0hfzojBO6JJKE1ZPLDHs
t6AnE7BxpWNuLupPfNXjo6Ad+WIfnVu2Yr1RxXa2GgPnBJeio/e2H4qEzUyeikp9
z2PmFoJ0TpAvz1w9TVRSZwOmSLJAtE2oJeY0jYevBvPOpE61PSI8uXcagXqtADZd
0C0GY6SHLh2VaMkyNA41XmzYiM9BJWTkhp/RJUrEKOab62rcHCDkxe1wNMuLOrQb
kFYNFnTCJW1xRCrYKPbDpgjaN2mePVihMmZicRBljEw7c7xeupMbgaMsd4vK6+bt
GkTbP+HmWhwLPlfm+VFg1a5UnrlzCIEBB4T26A6mcJBXYtExYCt9/tkZByEudwyA
BsbrlHSTTFXmCou0IthUW8fux9Sk+5nFCg8ENEZATu7tBDDztU8hlRkr0//9BE8n
UEBPU26jmg3P5pF/R1NgkQ4Py+uBo+hErIFNgVaYiD3lwfZjm1HAJ3M3BC/FBIsH
zOYdWo8qMFD8BbkmYLprVDgUGhW48Ijs85jAsP6syL18yZdsDh0g74rK+XPFCgv4
fU+jQZk4/8OwjstCC7u1p11tY+Lh6bKZTk523ra4dJ1picS+cEdJk+CX/yRghs1V
M8H0Kby8BenkXFqhnAuSU7Evsqzq2NaHdsaCb87H6WV2cEbJdb7rCqdL3UiFHhJ7
M6KX8GkmCnigd7tbVkxH6hDKyJKkzjavPucojNy1K5iPBOg/Yal+meoWxqL/zZZl
FE6+UNLnTOlinYdP0c74+Ccq/VMX9bHI9xpY5SHrbfOUpZyZUbQCH1Slang2Ng6c
oFDay86DVl9+x+Ji6AIEKtXR+uYj9vrXWJXQ24esnUVLetHYb25uFRgDXlDtSElm
jDslmucHyQxHdmwyJsDNKrBeGlp5HyA1rV4JR9+iADS4ldfnUuJnBu0hV9yRpeSj
ofbOsFCj49w4ma9zAS+lYJxGygfx6mRu3wd2+v8doqo6qVd1AutIgdguhzaI88+1
IxtYr4kRhi5gjQvuY+uvoHnIjB3RSMzl16qg04EG5uzyOCPGxYZKVHhCUoW4kiaK
V06j3BB0QnzYnFVrAFRG+yn4xoKLAHzg4p0ZSnDeUTZYIg/FyWb3zXQpJ+5+J45F
kcMuRs+JKAbMRzJbWF18H2a0gLMPTu/73UacGnspTEkYRlGFYc8URS0uIOaHGLTW
mFhQ2CXQr0w2Dtt0vg5KVbtkUoG2MPHhW6Of4YD1RNeEFpkgGodyfRz2Idh0eTE9
QDJPlCVaRBWg9Zxa1IzAy9cmqijc3KBihGkuYpMEO9TI9mESXU+6lLz/et9+Tglc
E53zdleKN99lkkciXXKVSfqhf0/Dtap0T+jAG30YaYDn+D7O7tMmSKQln0vc57Py
PLKa1WNb7DDzpLC8Zxz/WBPfjubM5QjUqiu9FqXVgOr3jVtthyXFh0lYVHpKCsk1
ot2TcOkc12OmojcUChE0kRPjXdrJ88Z/p6BMR0leR1rXw/8hXZCqzSH+uzboLSkX
mFlfTkXOBGxKt2wua7lErrHf8lErL+WHa4my7lu4p8hjCOcHp5p3UGNX1Vvd20lj
7BHwcoi0rKT1mUdkpeT0+xijGaOAagegPwhQwsO+x+BjcY747m42QJN/YpUptecr
clafBHwGa6W4ipxAYN1DFdwdl/8TtiD0YuE8smyED3/SEsCSvphGgo25xLw515mi
tTF5VO0gwpZ3yeEqiuxS1lssxsNwgn5qPp+e0O944rG/SpY0m/gWxaHvloJpG0xG
z1MQ4HHti0MIzVfZw2+6wQW1ZicrQ+0VTRgT/50SvfIJfAdjAakcq0kDDnuWf3S5
tOhqLZg97UWkyTFtLjaAGZKTFky79IaqzcFECwu3KuZqClpaeHpD4o4SzjKF8xsO
rGAlju7RmFa4fNzV95aGNF+TPAcsVUat7ess25LV92XAWMyRIC0EntS62D2R/kuX
sf77a+tXEs0MBwJIeiO2IjaK/7J+KM9LULVa6biJM7R1nOIeTyYt3bBsVBpA86xD
XSFnQOEiVa+MADJf4a5ABflDnK2cztkk0YIJhYIABb1SRAaJzhClpgXo/X1+b7I+
qxMPKKjw/IOwgpKEs+ORNCQ8dpodIUhhU3QOkFcHmfmBbqiz8LjV4noXlsuVJ20i
71senwCubgRm41ObEmsJfjhiT2mFoLjExg8ZNYhoBA8AfN8iv7Ddps1v98qHh2To
dhma5Iki8i2RWOUXAQxQiHx+0y36Iw4zBBkXrv6ls1Bs5y8uU7TksdYi3OAIGMWo
CvST1SLR+hBz6D6fKejjJsH3LINZkCq16cqCLWKp32dQcYoDW/mfFzF7NE/zWboD
J0S58NZ5BDMb4D/O2ueo2qHVtp0x9lvLfrS7TAIWS/SJMVMjjuu5AjKLQMOqj27H
hNeOoWSndtwvy3QCQj1ftqtDnfaEAsvaA3u9ignAgzBQzRVvY19jCKc2XxKYX2UY
3qkCvx1s7fGndyYHu8VVuvZnwaAChRZdhdhSCLfFUtTRDm89/EUbckXdtkuRwcbx
8lvAj5z9P+nSGvkhbUEUJzinzYMCN2E8ZvXeEFOwonX4vhP+kStAH54Hn01gvwnO
ThCPhBAxu0W3HDnCpHBxDj6HLTTY6Z0sd6juQDlZ1fOGAHRbdYhqlHoehNp1rnbU
zvVosQJPQaq8UqKlgvWWt67eFJFzmLaIwUSBh0ROgTFKeMztnDA7Nr40hl62o1gz
tGZA4LKWD1pfAVN746ZToI99Y/vU/Ps5gXaNz9Vhjz2DRgwMy/fC27YinNQao8bH
7Y7qIOazTRVNMFEFPQEtDLNRAjcJQtrmAMBqpTD3J8F82FZAXj759c1m6N+Uov5q
ZgkRQsmRXDrGW7ZihE+uHnBxcHmfN8VLXB2AwgAHPooog1uibPfWmJYFhcoCTcQd
T0j3aGuvBTlQF+5hpMaIdkAgoj7IlUZ5io/Yxejcx9Lz/RF1XQShIehCRVG+3uxt
+mTflneyDxI+3MF6xMF/R/g91Kd1Fs9/3O9Q7y4EPBePdwWqu9LNA/dHAV9B1pdF
eEx7VIV5y/WCdyKz7NaQcMl2xf8DM9wGer7WW9+bwXwPMYIW99LBzaCnHeoLRk+f
R1gTnEwchGVZu2Kygnh+Iib3f1MjpMgRBoM7sEu/ce4F2fb7LR0tspGbTjwuGoj1
eu+7bhhxc1LMkB71LYKL4KYEScx2W6PUQ2iUuCUMd+u7LD4SL/kh65gyY+QdOUCs
2BmyrOAe09W3eNoola8tkZrwU78Rk3L0+rDC6JF5Ghuhfwg4ORo1OV2d5owISTNz
FzXrhFx9XTxwS3DpECONRVSZw0UbkkCU4vguhGIw8Br+DZFMacPrbj6vUC82s7cq
B3T6idKQdOlbQzo5q3CeRh8B6b837u3J2eSxvVVRHK7UU8gCy4byhzHu30VehYcr
jsCjxuzwI18HjFYPNzYh7dloL+dCS/+wxqp47Qj51bIbVh9scSqHRm9Qd29h4LgK
TzNMJWlfgAnJBY5B6L7/uPH/NoDqUiUlDbdttum9Wq5wlTXz7LWCdVIazVf+Zeqy
foEQqdDXOXP652lWI2xAX3t6ZrmgD3y7baMeeMPGL6t5YemCSRBNd/+7/lYf8W/V
5YXRyZeLxwgrGHNSw3ib4wVBezzwMkWgdIl3g28NpS5bQJ36oQNB9wk798s1h4m8
rx+vr68H63MDYHxbG7ILQBmuXPx1k9LPb6nsRhWPJbn6qubjTBLDSALqYey7Dpdu
W0SiCgw/6+TjcV3xV5WI+9e8GHybHAiZDEhVQZDTmB8tsD07FBxqzNoUoLUVPwKW
oBE4yixKTF60jrUvMQM4KtgCPP25lOkXpJi60lkc3KO42vgCoq48NW+ANddi2ZBc
q6qbWFwfdlmz/lt5lXE2JBcKdLxUbv3mkc+1W7A9T5QJsDK4l8KV3vlL3V96WRNY
G3zTLwho4GiWRrXbZlNUR3wPvdh+TkFD3PwwJDHjq9gqa7NpEaIqVz7Sp69LwFWi
5saM3YReqbL4q1fvpCSiREQ/OJPpjFV04qmuc3JBgX1TevRaNlsB7vn6iI47g7Pw
Jog+UYzLzni7dmYst/C2f9sDcKH6I7DTuUMHqwQlCM9idlE/4Ihc1lpAwzJdEk8o
B2J+Rndm7TueC86MvnY5N7yUtuqwjm0oT0U58RS1J2yeqrpppz/1sXhntLdPRt9E
mwtO9VVM3p07LuL6itstBoY1hP6WHxYJo7ggV02zdttpN1BVe+4uZkvuZXc4xBA4
EhjYuh/kwge+zs1916V9N4x+k6Xur07xPuGideywFelD2wIpp/9DQrAyVvci9spo
VLOzO8aiGC7lAcoIh8nHa7OHuVpH8kpGjKZFXTR7y1FNTnqb3FTYJBb9c9e1XMPr
FatK9liSRmTy1F2usQDM6jsyHfkEPF4HHOCQQw1Xycp6tkY6PfFeEd03OoZOWt0P
qlUmqf2rTive/bOnII0kGBlWcAMKUAjH5FX7B6adcqNKY/997kxbQScUqWBIgmXk
LHTT+c57WdWeHactYUIMgvhP9zgFqPSfXUtTJS7WC2CL7FlrCgTviyNFicSHZmva
6v0/JelM7fN3g7l5xFcX4xG2JijLm6BtONftpAn6BTAtVsjwnlEOZhCKJ2gwe4Df
kngvXD+RU1xMrNK7Lrd6rUmaS+FZKzrC08tfDPAe9SBVfkpj8OB5sad6K4VZdl2e
Xa9/vFb0djZR3zlyfS39UtAK6O3pRHVp7I+xLHPBuI3+NM6BUHXnXaluurLCmoQI
yuWciGRcra7eX241fdB8pr212QnBT76OEgmrvmJz2MJwB7yB5Te93c3m2ONpzWMF
yyBeKbATEbHlcAtHP5xfmj9T6FLMNxY50MNL6Jxcc4STJLwbe3IM4MQHXs2EiA78
UqlELIKEafe9ruZL26BMfeGTIqpvRutjSSUFNCqVKve7fsLEZfXmfB0+8pRihmcA
5FuXFkAmgkHrier7uifxXgr6NQ8P0idsD9C5dgB3YyYz2SNKsbAiiiGSqrdAaEXr
zrd2rXYUUFfkXpbib5D3+eoHWqxn68PNcn7nm+3eCCfvg98wvp2yMdyFkDlLpLf/
AYW+RnlOnVAA2wPI6HpPFBT7sddF/4vPon+TEmDi/ZuiVUSBtUA09uOEo8VxVi8u
Nn+3s2zLwg3a1QOFhZUCQXt/Z1ixJqKIrfSx1Dq9UpnMuXbTAIxlngQyZFgGU7xT
+uGgtL59MmVfUp/ubKFNoyrWPz0IOC3OQw+zvUzocyCIQzemwxLNFKS3kywqEqs7
/bsW/BhWUHnC1AVudHMoRrP+YDMRD4Tmyq7KAnyKhPG7p+HcArBZFvsLHIzgNSV+
D+yTuteZ4OdgeR1S+RHCzzxK84a9cf8Tq7CuuXhTzbouJwYDwm3rlJwSIbWnnTM4
w+mxR2LAb+GrObK2YJhi7GmC16No2qiLxi+AnnPaNWjMjaD+MZErT8x+uRcqMGCY
daEAwCjrZN5hLPNeX2qvtbXxHRXUO2HaYyEngMJ1C1xTm1H7ExCFxSt0O6pKgtpk
3EKmcApM7d5jQH6619mmz4jnGOrTGsm2VCPySvd/yN1LM9llVLgcfiNMbRIUqSrK
yeAuNRpFggKkVwB2AkhUei/ysJEVw9eNUUkQT4FAO3xxKyoHdWrPLP0XkbaNtzxS
4NVqbyS2NnEaBvohjw6syO5KD4PSbuV1z+YtV5Xget1dK1FfxmF9ui8iLFs+5aTk
8zSPtKpIW8/UQ9gC9pgmPR0y4V71AMstSFBhzAeOkR26enipGTE4V6wV7C1B2UDS
1jQ/sZU6EyubkpLpD3ch3WHzDYMLFSHykO8J31Hy787UBnSxMVQya5SwO/WPiWNt
QKt/R/8rHrk+H0s++0zuZPnSJLdX7oECbTeY8udED+Ob4HC4qfldQT/vDTZ5f7NJ
Ta7+eOpFLq2ss4A56wzP6oxvkL8eO8b+iRUwx2EwnY+fl4gPeKyaKo70dYsXj86O
tfRPX5FCxsDgabOzz44Rb8au28HqznYW2YFXFL5ARzstDR22FPg1XUs7dzuqfbxA
l7lyLWIfmX20Xsch/0IF1z1XAtbJlYpD2IsUC8kna6/HCV1YKTAWay2zSgXoz99l
2rLI31YWJw3oQfPX5Ol7ghBNwePpW/7kgASwUGQzJE7gMQ/7bN+4o9pJ8jfrPwr+
XgzcLU8C1aij5ZyZhvtgpjhqPdqtYuglrEhxGFXH+0G3QHQnbuyC7YppQvygG2EY
frjcSGlLobQmcilphAc4yLwd2Ncht5HcdOKt4SU2AgX8JoqviMwHyrbUhHJ6Y8SJ
TYshedM5J9+G0+4LllS++inqJRp9F3JMjhnQx0A9PfymZhy3lVrzwiOLXP/DJM72
C3F8GDZGtraN7nEME76AhIhk3jTU8L54GR/bjejeD0lh2hqDh4+SBaACR8YwD9tl
dtA3p1uzT5OLi/VVpCVn0QfDy4ZvY+v/6WcTImD4jc3Jao0T/SfxGyWdtLKMEJIE
7hVmRZFTmnxKQan/vWGyG30mRFFRPIee+7nwVhs2+VwekR+Tkz1o/T94XZVR+BW/
kWXEPPLoBry+GxDmon4dwvNWczwAFuBRVgpF9eWqHWxBir4VmMae0ZZAJZETCd3c
Fn32FO/jCIeF2YnGpTxUAQ9p/eN5hmvf6M0vissJCLDP60JMYpFTzs0lzj1pE5GI
ZXc41JCzTlVwE22x3R3HestPFHYiRUWpeJgNlxMF0NVhDRr38vxLYNUtCFNY4BA+
y9kIHdvwHGW+ydZ3xIHVDzD6rZj/hBIdj5CwvEN6ZeNDu7VdblSggOl6HdVQSHzn
C7hGctoYXjLltsvYWkuk+Ug+fNT+oXjEb83oz1H854HZliuindLIGrLv0lqljsv9
YYUA0OTxLIW810yC16oxOsIS17W9A2tklOCF4R+6i8P/f2TDDLTMA1zVotIgTxRe
gTxfMXzcZOgZnS6PkBKhAXTFmoKjFTsOdPZMU2cR/J3bhkREvyRCryD6oqVVTT29
aT1F0egZm0sH7ezwA8U2fxisEwM7WzjrwPO6TmuRf1ThZmAqHasdCWEU+tgtq57W
mBpqCLf+3k8q+b1vJ3vj4OmfnBZwPOC+JRQ4zLDxiZ68+aL7+5dnU7ZuhanN0zq4
q1OesXLTKhV345V7T2NxuuKLfrVKHXbMfr3GT75Yesq08NbDu7PYF+Hi0aZgt6Bb
Actz1XVmwcUUhSsTRWPnRqRspLHZIe+ePSeBpEDG9l42MFn8shVdtJD0YfV/1Nx5
Cl7lxAZyQ/OIZKvlXvE/6vmdDanHf0zoLvPxO+e84mSygjNh+lBxGbR1Rh7SmSoc
q3Lm+olYtpVt7aPO6SJO3K7fv/dnbrSWUSwBJLA+ZD2osnc7ua6r22zLBPwtn0nv
isN8WJKYOJ/ftbxVbHHI6UoF5Es/4L56VMKRjcXk7FUbTaaueli9iVHLXtpNfHrq
dZcRzd2cwq4KL+F8sfzDuBRGLA7mo9LcCJKJyaQ7tY2/P3HYdXy/f0d6J9xu97IA
AdFNKF3b0+XWp6WafRihPlKCu+/fFW5goJQQ5kKSSxyguoRSV/yRNd6AFO2BShvF
s2yZhaHwc/f0M6X/GGlTLj5TBWs6GnGNaooP2BuWnmH9HRhoatQoEjaN6n1WFnlH
+bpdNVnP0z3Y4LgYmkU9j/ezkTxQ1TseG8s7zfRohqiM6u7gkhUFx+kx0vu/hzDf
0QCiMrf8rokyv4iQugaEnRpuEyRSl9hEA6+Wfc+YuQaVkm7/LGMTTbDxACcNvgSq
9hGCGPUjfj5RE8Cf6NXhDHCbSClaB0bqrkhcL8V4AK+Ed5A4rP1F81V59b3MnPlA
CT6typ9yF07oTUsPfbEAyy1vHWVWQZ+5MOVgV8G46J7xNam3pKUgTJ57KYRcU7Nu
NXXhbSYZYWSoVPp2p4Itbi9sKZDTYcmUOFphZU1iuPP9PcVp3Dy9FzlbffUaJTJ4
yZS8GqMTKFsuV4v/wYYxJp890k0G592W0kwboPN8iLqnyuv4+C0PSuoY+06+jnuq
NYxa7BAoG3oo+xu88epuReq/sareoWeRtCNFSdmGSS2tQIJzDJYPXl8CUjRzkwo1
`pragma protect end_protected
