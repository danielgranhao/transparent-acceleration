-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
fZKW/sddS/v7kUz3nr0ZKd0I8S/qAx5Vl42q9L2M98MbQTMLSHKAYqq4fqqap3Lh
/0xbVuWrwDI9+cH99aeXnP+N5q4ikwlhHtEP5OsXRFmNto/C5o2MLRx2bQbE/wO9
jBqyxDwZMOaLArfw5W/sYaik24bW70GHXr4CqANt4mE=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 9845)

`protect DATA_BLOCK
elk26WbduLViUn3qfMuWXus0jRieSH2QZmwFqbtMnzjQMC8O0oV1l/2eoV17laTj
fsKQrhlsAqhvpXKC7yuFGYmakw1apf07IGI2ihlKvL3vnd5XntjcD92jw/EDFCZ3
T/O4teHy9vXO8aF+8FPSBmrydwDp7Pn6/D8CvIgA8eTfeAOUBcnqNG7o1mueJ2kP
b9+4UXy601m0PGHSkZSXA7HgrNC75Z8u97+Cgu+VKIK4sw5XBWBUK/7OFg8wNlMo
vHLGbgnTRVdd0h6r2/1tzjxU1YZ6mbVFY2yLwi8jFmXaqXTNm5z3wBd+X1sY9gpS
1prMQy+AC0RmrQBjhRunCUwqwUvcaUbkLdBNJUvY6f/4YJjvwhX2AX4hKdFw8lM0
oEKsPIQWwjEqM1V/fOykWEqYKGYu1qiAfK6muqie7h1wvl1Se3K1YyNvD0y3Elck
2YKiXkWyRw21DV+lvxdoO2tpoZs801rheiQS8TSr4rFOOpLejJZVBYGxfWFgAqWA
lqwpNXSldusYbiQrqpSgb2OJHftrR01uZfcMGcNAcFujtm0RFHQeREbjRnXarOxH
lb74IvbV2bIMY/LNMJ+2B55GiEQmsreu+UKtKQ7q24Zt3qQBkjhze2OXwJY7owS1
UD7b8BS38IFfvW16zALk2eUnHos459FdPz+TPHWf8DxtTBwS1S3R0rM0A1OzR3ct
C2TGKZt4dHbXkrVYu+wgIxacY2V14brmFJHfcsiXjwsRt9HGqZAErvc1BkD3S9wz
qpUTV45pjjswYSMbSmWRv9cq1sH64ZUVasUblEIhOVr3hZrG2NzlmUlaSeHdCYvp
5Qlpl46Hm4fWo/f0qUZ4vc2+QkBU7HSDokDYe5n+XkHSS381vZjp/OfxVZFt+7wb
u0jgQXxo4wdPKb8IsX0zBdKLg4pSC6UJ/4S6tOiqj9EeDLwPyzlk9p+RJvLZ0Mpo
jtfZD0wa+eSbw9JV68mQ4fhNa86mSHAUtQdsyt2WBZA8WdP67lBgwjcKXunWjuGr
Z9njyyilQ2uC9ZsOJhpyEpYfbCci6s5bx9NS91hoMqNvJ9R5QEO/tmyvwh3SQ8lo
NBPIHS1Wy4UHzgwU2hOHTc4uzWcySVFwbpI3mwNBgFMIhh3HCfI43VJNiKCmQ6HI
1dTolXa7grwk1cjQqA5FZx089fVvw/rMVSx/8N1ZAv9BkACbmSiBDK5U2IypyuZH
4oqNtYmLiy9kWNQepLHBWMjeSqtMYkhVuvNSxTUCqkU2T3MDSJvoZYwlYU2vwiYy
l0eJQ1nDTk36SGotXHxMqDlKcIA8x0HsJ/KbYdp31Q378ssUcSlMyL6OFGLwcwIE
XPEzHQm2VC8Fju221rYHHBr9B+K1jAk0H5pf3zYSa1SxxBmAWUIp01SxB5yfG9yt
KS5JT39xetV/cSlVuegRij25nz7OdVH9I1Li8xlHa3Mb4VAxDOCNaPqXDurfxmnh
RwgGghablm9n6ZKQ3mlAABL2eqIAqUz02AdncwMCBSKFOhBc3Ph6VwZHo9bdtlC7
Fk6fMB93tsaz0Dz9XFmM/FFxPXDiofnDxC8etgjz//PdZH/4H7xiIaupguvlxEWl
TkdCXlLEmsepEqoSzx8/llNrAsesddan1sGpNp7dgXunJVBNnlMtslpugL4SjkSZ
bRfrrc3H9RspwZcLKBnRQVki5bhs4gfQveCMei1U0ZO58+FwTA3LSnyJwfQA8iC+
2sQ5/6GkR0BVYbzZqjCBbklZ3U7snI/WgSP+tcafQiPUqhNlWKoEUqhWU7quAOJK
/CPQ1JW373P4sq7MTGEiIDf2DoukphcphqZBDaYJieBZyXl6Hzx+EuJofCXv0aO1
9pAbnpkZv7Yy7fcUxqU/HZ2hW5+sAJR16bKzn4cCjyaSYV+QmgvYYk2scaZD3oZ7
A8JwbdUeVwKaUNhLVdkddrZ3bTNqD+2ZVePSCigZi7q8Y2RY6F0IHz1BknqA3QP4
1lnJ+HCraS37tgJhAMPXDlGwfGHCLBXMpb+RWh1zItcC+ZrmswsgYYlKHHsZ4rmh
MKMZkDelwGSz5825Iy3mrewIVp8HfNi8NBTKIigRV6sh1z7xY78YQR6kdZGQk3wr
2tpnlqeh85/pM4nZqtV9LsUc9c3SPOYVZP8xAW9lWq1L2cunVHu5EYdpHznfDJ2c
VGPms14d40LqADcwRfzOCYTxb9I6mCihgxA0KEe69ITKb4OmKjjMO/wB41s8nobv
4f1vJwREsYWr958FUkilIYBCe+uyvEGAtob199gG6kgsVwDamxFIYpwpMRbZW8c5
tQA7tg7KOgyLCXg1etqMr5txRZzkophOH0Luu/9486eejvCQbtWYlC+2Ozok3edt
mMMiDGF7sCr4+l0rGKKUw8xtQA0CdqLwy0Kz7NWZKbbeb00QFYl9ZBjQiQOzYG5o
IGBOqoET2fSyUQ1LHmU5mhWwuN/uk2HdI8D+ZELMpB9mDDtBvltQKhFsc8628KbQ
vomD5uAI5ytRWRWynB4Mnt3UaE5uaDG//J1qfSmlWqJ/eeprrAXmq3lC9gjsGPlm
8ybxJpUbxC83UwRH5K0vagQ6ucL6BF7YYj70tAnWzntqQukuAhWCMxGLVUHAakgO
xFJdirlxNzlEERxbWyh4LPmltZpmOVJvvldlVfcySqEduecHRx4NtJqM5tqHbWNZ
244t8HNkJqQoUtpg1NE9hHVJhwZa5Ve3+7Ch46fyU2zYfeLQBS14KpiXXwJPc4ga
hUiXUD73hhR/bZHkSNJ3hDcZcxApkChfwCKGseWrn+KLq257irBqlfjNCycXtotv
7BZmts3a4YdGqJUCfzYz8Y5Kw3Qeg6bLfCBtuA5JHK0+PNxEyaAjbrOofXn6JDIa
1QtWrHsfhht2i9/rodgH6H5lVlfK/TQKlDoXBmqPQJs/D0fhdJAk5mw0armou5ej
Wk1HuKmoQ0aDerxfbGRy32SvPwTSHuNdsXLSNf0AkME8VZh5ZMlfdchJYxsZM2ba
HR54luiFCYtQqzamSirDtP7sihktOUPj0+fbEIcFcK93mqczOgGdroBoeuTAeVl/
KM8YV1W3qxx9uYM5ivhENZXiEH339cCtKPzlmHjsNsDcMdVyuliTRG/OtIpJGVx3
OtU9nJmIRwK7FOYKMjXQ1i2zLiNxliS3aAQBqJrCHte6wh+j39LOwPNuoIbl7hE7
XjFZ4JW2N//3zL8+4KSMZ6ntbauoo0BRzFH8wmwfNNE/z3OV+JGp2zxcS2G/KCSm
LMtnXQ4BLw2jTx2Ni8UTusrcbF/kbxsUVL0zy57YhlRsgnNopbAz8Y+xpu6tHSii
CPIFoYp1hfqqiJYey04jbTmUrqcA08ILvA90n8JzefIwaz9i1osf+nsyTG99yWyg
1dLUPrmEbqafdRjCfZf5+Ey6YTdqGfLLtbbvCGZuBAYbnajFyDVvlWgw50484xmB
if+fdG9Tv196okGwUGMaqcN17C2zMWrpu7OEz3lBjkrto8M8+MYqECQ4tg9nSHW1
GaVINDRfuaZ2NdBFsdrmE+phtz/7XGJ2ADsCvY9PFUT87Zn4uP1ZjcoDxsdCYWDW
QXfmTEsHF0WgYyu2EuPMf6UYqsfKB9MEdFIr8TgWPTGfNqZHXn5fJtwWFK7vc3TA
N5rqnPIgKbQA7LUvrRlJwWsqcK2AVs1Thfkqx3MHCHhK4IDI93ugu4buRySCfDdw
hN1wBbrwRZFTsmeV5py6nnQNlO+iI6jOHZtziFIm3H+LnlDFYC2WXobVs1icjjle
ZIMMJeXseWXMabWhc86S/vvCCzX7xEZFww+Ns6NsDNKhtgD5BReD6e+wTvhqtFRG
fBtl6bNRsONGBFpJAPSxZPoUo9mtZwUw7z1i6UShSPWeuKilrKKsXf+OJWyGeBcM
kVN0MOLjfjxEqEDIvQ1DspixT/cfXzrrvXTfite6CV5gJrREQiu7NO+7uze87hjD
Rz97h2t7N692Q0XMl5w5ACELdh45+JF9pYdcKp2ALR1D3Wht+HYUrwzCqkH1EaX1
pk1u88tqLabtOb2n85vi/ykomvRSa8bCaroWoiyZfgN90/VElYbpEFkX4UUojTtF
ZYJXHgwQqjVES87qNhcT15DV/8mW0qBwMV6PuL+TIddk6a5WRhG9OnKrr+9BQWl9
cn74C4m2teUKzqaUI59mqSotMKomzaGx8Vl8Eba8MaMaUtZXDIGZOxlZwkEAW8oJ
PwBwbNzwCtBkGzlBsM2sQOldZLVJBIT33EiZlvZ/bGpTcDiF1RUG7IW5cqux8MvH
lD/d1gjmG333P4y2vGWoTr5/Ea1o6auGrYL7CFo8XYlX8x0oK2NGXx1C5uQ/Ryu8
MembIGcH2/VwpMtHKfSwpwqc9X0IcPhFSTzPb+1X+6b106LibvjW/AW/R9m3hJOA
PgPAb0WoHAHH8BRRQX2kfBpbiVDXGV6xqwDvl/YAX09WqzVOi0HL4lEj4mQFkCIl
98hlBs6/ESIlTxzgim2l6LfkTGJhpB2khMMKIX94MJ+YEDOt24QNG/3VYw7EseQY
Ugc/fX29nkMTqMQYlv6Krxwb2Voy+8V295k3hl/FwJmSfPKDfB6jRcylWuAg6W78
wMZF3yME/1bkmA+voTbROY4HrKYNi0aKjXBuu7rKfxuqaTGH8PtgRg9aMcfbJtlG
q1W1IaIvMUcuwcirA1YBr+C2Goi0AbW1ZZnYj1lY0piKMNE+gSFP8T0pw0kFj+vQ
gp2z0tBnq++mrPyvdLEUJqCFtaaPuhm2ceygpWvgYwJ5KqWM6/VFDMPhdxbBzeXy
ZJ7bohUBVQKt7V+gM1//XZqn8eMXGKP9OLIGtMlZTrfvxwXZFbeOKtBYh1fMGEm/
A4evBWd6zNKyRQdEwCdzzHwwK74TDPl0ihop/uv4ihqGDKRSGOVAtfpsEtr7iIc0
wR4tHoLDYoi3S1VVhxS8TyHHQvUT2GWiVE8UR9DsazFbjprZBi944wCgaVv1qM+g
Qf5QWSE/5p94IuKpdH2zG/9cshgioAW2qAApJX0DmMRZ6ZgAtCOGrxh6a143bhmP
dJUWh/EhYcyxGaFuQeo0DOEMuSmvg98Ws0oLxPC2ogXFDGVGSXrfxj4VQ7E+nG54
yyuWVUA8CAAx/aQvqhW5RGlWZEHvEW9xPugo/yDqVK13UcTaA7bYqBsxGVmZOUWu
8hDMJb4bwFNBW5R9BfiBdaGx/QJJ0wK5CNRZNSIckLPAsApC0dEbIJCmogFyIKXC
SAlvJh1mCd1u9bXN1Kna9UqeBGeIkwiTV967boLDow+Fkoxcg/4wnyFRr5e4fg0q
5xNciNwHgPV83OEvftwCDJpa1Em2e+S18AYNRK6iGu0ntjUf7g5hv0lDfzdu5B/a
aZc0UXhjTqxnejZGc0mqm7N3pnvQmwaitij/tPCGBJEU8oW3qYAZMWvFKOBXXbO3
MSgmdi0PExqGpzjD7ixAKQiJUPJa+uY+DQ+ZruPWvwr/JV4dgB29/QflgdtHHfl8
wZCyLzxwGXFc6FAx784aDVnUS48q4L6mw+c5ojSJuLGWBM+5EsNoPewBdttlbW0L
1v50L3B7bcZx5R7EPkALy7ujEReveqpc079imD3kts2d1nUAU3tk69kmGNmDYWd0
HV8mozLaS0Ez/BJ9taPOWaHg8E+V6z8IXVhEbkYJ6/N0x4+hJe8SP+OGTbfO6Uyn
+NJDs+7S2QmNJ0dnl6WCuJgR3E+G4q2wGgXRNwkYUxnteLO6qXPydFZ4j5TuF9LB
fQ0r36uZpvduns6pzELRknzgzK4qfWn/6uigFvvr5qOC+Wp2Qu/Sv9m7k0o7nVbI
F6N8Z9gM2aUtWw42u/yk/Z2DBZUwFaN27dc7FTqQeBEZK+bNIDkiDNRwVQLyqnlM
4/SA7dxeakyd4X2rIoIihahW7+B0VtGwttxrmfju3zdFHf+0/rvN3Bjvd8QzUD1a
ZXsCyhNhBdub594cq2EPd5n5xLKyOI6M/3X7y5RxrXD5ymQzU/a1dVtNe3iDY7cE
qfolenCf0ycADBXFDDjAmBmJcXRgQCOrCmpVINC+UyjtuB8G+AhDaX8DmCV9tgHR
BOJePAHVV+BaKcaD+VAr2yoEaux8id7dkdiwnvAq8xwwX/FGFhsUxQyGomnNR0lM
l7+sXBgwUF1wbKKLk+N1YsqQzYRWTHxm3t5KPtxqZQiQuQ8dYZQvjB2+ZLt61qVr
kee/oGo1BjoPpyuCJWJN8deI7s//tSK/wBt+OWINmUObBd4hZ+j76wmSyk5ja+qm
6MFiCIT4h069nyEi0no/r15vW4NSsvwGLfBmpjuqkPqcAg3svQmXYGOI6MUio4Vv
33nDMifoVboYPc/PDVNfCq+C8ZaUowpCLGBr+R+kiMd84B+CtT5hEuzOr0+Sn3ff
jh/S7dfBJDAIzptQ/WnMSNnMIt+qTY6HiCJLrTUI6GuyphJO36eNhIK5jRQdpLMv
y4wBaG1+nZV5rd+7d8QkX87eTnSouqWueEer/J68SRBvpeRiAoJ9uWRNddBbbCuN
DxRUouhaTen2t7IaFvofIwwbdz8Z5OkrPNfAEbJtarG4ELyxtnLIat3Gdor3Lj8H
21Qh78xVw6aCYvo2jQrF2OMuctQIXHUEQ1jlmX/PpraeYx1qzXzw6K6b8bD08siL
B3Gz3bjNUQ6fiPOopQkbxFrvEwmFqpfsWcguagWW6XDPaZmYvRHuC/J/PHLTHK3o
4meZv2gqiq8SWAXjJuqZLUNcMegdgry6Ufx2wZOP1j6TAcmR/6Wb+gcZYVzJzT9J
4Rc3cJif9sv+VfNnm69MX2u3ay0tp0Op6Cy0TIHCNIp54paadsx47ijW2cRojKIS
0zV9K1MvO7vovII6aLLS5NQWr2hCJ82nAAb/sFextNETEcLWiFmizHSCXRanJgzj
hVpGN1+xmT1IQwzKU3ogkWc8Ype2e1xEaJ9W1TatH1HjLX8rsb9Cg8eJSZZNjrjM
XrJuWwfKlt7yYD2LJMHUUxCtjqprB6iALoZoylRgRXkROBSliGUfJbBw+VVCAL4C
k9rdSnTSlSw7kGpjDdrJyaTOLNprHwO3PVdoxjSlDrLVmQGzTIMUds1vGQBTjzvQ
HYPSh0m7Umo8bboBy0n4C5kXZcup3+UvxM4X/724r/P1pqDbAptwCmIUXqfGTSsp
XcoQAJ+bhTncIcuxoLv10ICruXc73lHpRqJBdQy8Y10BUTfhCYauvyc4PlzK8i80
ORwFtJNg6V1EndG9MrRxUjN/gJ5Hr91fKFNDSF/YAHTFw226xqqXF7WKjPr+TLGy
bdhtUH5jHzS8nOTpJjeK7hpbwQ5T+vx9AwWNtHR69zCURNmOkPjihME9X/eOoECz
emB3LMhcN9tciXSUFTz7R3rT6VqiI4Fqha5zzT5NCPx54jxlOAI2DZ1trlLH90AW
3xzUSHLUodxzPG9cMOOR8wbQi2UO2fyp5NGA4jpRQHrrbuZP9o6C2NlJFxIV+VLz
VP4DATLitjqbgOsJyRt6CIRa60F1xvV3i8HsMuPqB8P4GzOjWdzJAeyPxYZqAbSa
bhGN+ZjMVjGbuxKwuDWH8d7ln5uuRlqz+a/NIIdDHTBxp3nmzyOMxMxZRfuj3vK/
CzPU7eSZ5bCIgUSA6kWRXy9NXsfDCpffkIQa0ZAZ/188FxFIR843q5TUIjt5APSc
w93k/GFquBfKcgfW7F9ukuDRyd7HCbHs3l2NT53KskRaPQXmwNUGaeIOLiMRRG9/
g0BtnthRYQNvWJd33hON+FdrObFdekmDHW3HnvYWe+LTP6QR7/3SiPlluPAOYcBN
zLbaySMHZS48A96EWn4eJF7KFv/n7Q1ecv4GcQlKVZ+fr3kzBhBD2SSMqqSGpuq2
3/ne2AR6BSIFgmSGbG8OFVO7sl9esAr301j9QSOmJqs4BmjBu3RbnlkGZZP9L6CM
cGvuXTTT2wDzKsq6Ub5MvqyBHoVYkeT+3G2R+mdLdkM/UEA8XRLN9QL9NXRKT2gD
tLX2m6OEk9/SKM5G3LT6W0YxX3sFL0c6E+t0T4ZEARQqIMWXLtfI9Hnauq7p8yK3
kHKjVfxpdnxWIBpXruo5SkOuk3j2VkLnF+FK49xTJRGlQ+R+Ca5tJPgQUKZs8QZ2
tIdc3DXyphAxLhPlDxt0T4sIlKe+7RNIzM5EFsifu9VPuATO9d8BFccl/FjOIC9I
sci7/TNyZC4Rp8m98ScVXQ/A7c+TsMpbN2F8OGioDFQwal/zcawPFVIWpIwcv1QL
FRWC8wlAf80tjnDLbZTUgie44ikSvwjkUDIkhDYcjB9aKs2E+9C3mYOGVL7USeE3
GCOSJrIGJw2umqIc2C6AhTn2LE0IM8Vp85xwSyVEYbr4EiFphSY9jfsXkZyN4xbY
Iw7USZhWPSFti1b/YbXgpy8V8tujXgU9cgyVbUsTaF6Crbte0gY92Zh78qkECv5m
fY78NzO8FlhPg8n/puyW5sqSJolB3J18m2TJS7dMmUVSujotvne1M9qMkaQflfgy
3swWXt7AN7e9f0hZf6D1A90PAaZ2L7XPZfdECPfEcPcCLqO0OJQA90mqTLlPRPiV
YR7aqVJ97t0BejNBJq//mUTDI3k64bU16qIQKXFadEu5PW7GobcgM/iZeN836H58
YYs/n9ix/R5QTIui1viVgGQT4zGg/SUZKkup2mSTmQiEF/H5UG+i5+DQ3a99ewAv
dLHizOPabi/u3PW+FxspwJg1GS1ognGpqA+NYIMoFYSmP9boepYqS3YH8Px8ljoV
tunT2FyPDMlu+Qq91QfkcuyIiR9GFF8c6RwpATtAvKEozuYRDKvVLaVysz3Hz/e6
2HiR9HUYUzeA6n9dBsyRQM5HWgPYPzn2YfOyqiJdBaEzqwIuqwbUkk5/NGgrO75S
FiARTlatfir1FFhFvAKHnnPoCD6F/cV5d4nn62RjUAHMGqYO0p+QJPEbpjnKSimJ
cdl5hxA2vU1Z2UVuQJIYtRpJC4OrysBxrM7wQA4bnf920HJjMkE5gys6ZB3t9vgP
gw1KwwHvqAdZOqx9rIWDuRvkZFuJU3XAAoQY+wEoe/AX7GLujaxiAUF8vdW+Cdgj
VNNzNca8Aj4RV7+RpEzDPy3kyE/biubukc7YG/oQ3ewuuagrPl+/kpmuoASbrZ9l
ZTWMdMdjwt/sojXr4snyGPA5cstS2BuClorVVEUvAIQ0ooEwRbohNj6LUfSn+TYm
LFL8d9ngB+W0kx9tf7xlB5wlsIB0HFLHd3ZYajp6j/nYk7TRyLmWzSwSywXwdpcb
TRDTjsAnz/6BgUEgBHoKppvKh1QjZzRuohVBo2Zsxz1tq8p51dTZ1d0nH29Vl/Ul
j3ueimoIcwhYQbYzkVS84wAqix3OtrNrnIVmlrB4+WzvdOg804DwEKradz+xErXE
KESNghpNZM65xb7IgbxSZrU2PiK/7CJYua2mKzYgAIV0JaeqPUmP22l2Y3ShEf4r
EgdZOGP37zv9snjoO/mVCcH1oIGHNfliUezLJGq97APpJtBHZ1KP/H98hwR8MSge
Rq9oHOUZ208d6kHfrHypFFrmSs28ECx82QgGqLEWpNs3V0GU/Y1F9J136ht/fdI9
jTZE9/0aQAzBZa7SITCOnEh+/KZlHuISUdb3q3QnQ/P29uIjCZp01pPdYmfqatGl
UbIySDY2L4JaCvQZdWsJ3TIw24nr4hLGgDvAEo5GXcGOxsysn+dU4v9hFaVNuuSz
/h4acFuvyNDJvSh5tFw3jfItK6qSPDZ/Hi4UKrOE1cVXdykp6rzMbbKZlKNI19kJ
YMv1i4w6LTJYaP0dj9scN2ewCZS1C7Sz9urAVixXiQFr7/LP9TH3p43dFHqowm33
hHjklYuD9ALhCcLrUwRQl5m1s/3dMQdFMpluR3yLJngCxphy2gE8YzR+EBun2P17
XfkFtFONIB4Uk3oPT76KBSJ6uKnLrfz2eRENkBlTiISUvHl/AqAwfpzH7Kyx64cG
VhS5h8C/PzhJu8iJZqH2VwvE+D/rj0LRtXdcNc29ykfzLfVZ5NzhBjx0JEXnAtaj
3fBJdlv8VLNgxrDAKqL6VRiURKSKNHYN/VkiQRq4dQUOj9tQgPV2iFrKhs2OMFNw
2oC0ELWxIXM5nx9HRtpesxR2PQy2Nk+nryR747UHWjrV3Vbqs0reZrKiH2gOJwLJ
I7E8DxyiLav9ge2/T3Fg2VSKwU+SrDXlKT/Q1FS9xhCLFVu/qxNAdNpeLfpgFAS1
XqpsboTEmRXv/U8igcTpzQAqWq8ZAFLzkmV04sECwug5PL/bEkIJOiQSt0pY1iPo
o1FqGsq4O9W+CU5CE2y+5XSGS1KqsbCJ80uLJwZ+LLtQnFObU8ZHKOHWLy2K8Z2S
Q9QQQje2BAGSaLAHyL8FyINKAiSulctJQ8fEiZsms/FsEaK+JfsNsYgAzRpXQ3uL
rfTabwBg+9+Kloh3upS9jQtU8sFrZbnl9UdErwvKEpYNgIBttvWvwCk1cpKNxJAm
YbV/3cgIbxi+h9S7RF1N3Nv+LPnELMEmRpNRmK9vm1lIn8CXuD2mkaJHARTUrRgV
7OwhRmhsS0rL8WTKZYbPrT/rqzs2L1VvGnZiLNLHiNrmZsTRvwKrOvRhcSV6h3SW
cGIXhuRMzmoYsyRSBCZV9LtjQxT/a6vanRT5QLQzKT1kH0EciTM2nfdgdpbrw2Fe
fb2Y224wWlqufNjtX0pOILih3LBtoKp9dZWzG2NTfFaH5itstG8tn0KuZRebcOB/
gycm9re0wDfV960q0I+GblTQl9DFgNCcOFglX59lVSPE3tU/+jEox6zMicLbZkeT
mpWcoJ49to8K3WbfaTjfGfWBtQuS/KMpBmfLYoek+1Jib8U2eeifToiBSHU87Zov
+Riu2ThQFxSkydmmhS4QOHaNdFlDigXZ5BqsH/HMFuOFDnG7khqD/Oau01RDlSZj
T06F1e+6NeaCRgnzpnwaP6eaRI85+FvBH73Q6UvytTPWrkVnbqPf5dNvzep7K14i
GYQseU3/tUBZ5VDDyX46JTPYo1QU891AxO8TW+8nVqH9yLbNW5bAx5U12GR+LoQy
mBB7U7UZlXn0nxdpMuOgJt1iBDfVf6RP8AWeSChUQq9gVPlJMAvtTM4AZOzXf9eV
kEIlPMh7jH5Xl2B1jnDBCu7ztLNdb2WHryhFO0iOmw8SKfVIBg3Qy+rz0xBOUqpg
+Dxs/E4h2M8ZIDHGWNVgZYT2as9l4wB0wDNqkI1h0txLr8Rp6hPpGjJ5vzwFiU2f
1tYwyPj6UyhaOU/AROoGnj33qhYteq1dpC2a5DIZDbs6AjUk8Z/t8iWtyYMTKCQu
L3GQgxilymDWbDDfBrLUzS85e1uzCOxS1cOxWG8bgHfwQDfNMaPGf2nFUAKCYIrW
U9ct5ydlF6zgA9n708LU8k0oWt12q0CB4S7wT4lXKHMIZI6CMEuaHDGgVpCwlhO2
lmVFS7wxUfqmpXVTavkJ1KePyPd/Vd7fKb0iKVRczq2ttMlsD+GzS35ncgWXTQBs
kDwx1qng3rJZ5JXLoAS+83VQ3sNdGIy8ZQlABjJze8rvd4sZvf0ozpjxgvou/+ng
qB1E4De9OXsEMIQRSqkIvOqa7k5Hks00oO3V50NdI3t8q1f0wn13zEhAB9ZhiKKu
N7qBjjAd8QBX+m9CHhX6Sw7k5t3xoyN9pGIF0I0S4YHXQLFgpq+nnGL7M0aiUQWf
SlXiKy5fNM6lKwzG/cR2eT6zVJaztPLw6aIiDLjSFtcxEmx8LZ2BBgF8pP2veojO
pJLjt8jVQ9JBAPwPl/Pq4FvUu/n1SWC2UJ9UmxiNI4Fb7TnqLBcxj260FHZMkUaR
ZKGw4TQC/qqtDJ+OSjmXSFNiIlERjgwSfEG6FZkUslAcYOkX2wCGNcpJZyIMkPsI
/PFrXPLnjOSxL5VGW1m0v6mD0QgJG69pi8QBqXlTejBGf+Vsb/ndWSwUxn/SzP3u
nGXTOPJ8kRJ8NdIJXZviRRvyBO6i8ZqaaL5dquMYR/b2DjuKquiTxFe1gfs3j2RT
OgYO+aWeRv4AjTrAniQMlQbawjf7Mv72whYb3pigcHCiMBnj9vNDXqwUZmM6bHym
p/ZtTvH+e7irSnJEVFoM1bXxFMyxPZJxzPVMbZc0+OYHAVRetwh2w3b6HJ5qsCLY
1r1KlaKWUiXeuQ9/d1vxR1l0hrWTBk8P8T0p8sDln91wGtZr8LCuFeh3xuqDuS4e
J8m4Y1WmXNaK1OIZSodNbTAf7DZ7NfibaABHcsgeCS4mf5i0n8QiuZM5Ee/NTGUK
unCSTVrem66fvAiRS9ee/SrTdrHAJlysTW3fG9wBW3gxumD9mf/tzmlPar+c3dlX
AxjrUADhIn8CgrS/h9mLKaPz5m7gfIoG04GNDzUhf8mdKyXebAF2yjWdokmrsxOc
U3aKDn4UVWdsiG9RUa8VkvqbIrhsRYDQP02ppoRpuRcU+upEEmyyHK3Tuh0/HzqC
kc2n6TjnQ9ASd4frjjbKQHtjiueWdbYDsi3me8HSA7ymP9fxSDjBvduJXuUaZx4j
b8bP2Prq55I0H9CIJF239ZTNgUcLZM7sAhdUHJEtD6LNKXr4vb4kpMjQUuPrE+Pv
8Kk3CFXKwzPGEBZRbXzX2zCKFvVE8t3zan5u+wKq7thL/q0KGzeo3fFWAOCSg35R
HVA1t/2Hgj6+pQYYo1P0IeIa8EKiYhX7//CrUhkiDcpJBcvSVK8k37fj/mk3CmKF
q5QdTLyk9f9KO5Y5DzfuoXpUXzNyStu5W5P6jYsB0W0agrLT6KsZj5ZMCKSE8QWl
z24SOeGBvIcLKcZKhGd3bv1R+jOrPYU50Uj8/dJ9MFyEMgiqUuiv7eU+gNtrULnI
uuGTJmQnvjf88udxyLXtlJFdIwzBlGu4m0v6aI8Nr0vJq3nb8Tkk8bjLFvIjwDFs
uC995Af8V657anW6XT/ShxPQDY6ks7+i/J8e81hU8RRwTBG7eQGLjZNEzWrmSWws
OSwFbOsWev8H4f9w6pmugr9Oo0DdEmILlOQRZlH4Fv53+ryNQf6aAvxw+zsWDm+0
Ul2GLIqo/6q+8DDEBRlNTk1jn9j0M5S0LKk8cNAHMpLzTsF9IPH0N+LqOwid9TkC
YsW9iyd0cveIxLH/U2rg1Fv45MXbAjog7S7k7wgJOf0=
`protect END_PROTECTED