// fp_add.v

// Generated using ACDS version 16.0 211

`timescale 1 ps / 1 ps
module fp_add (
		input  wire        aclr,   //   aclr.aclr
		input  wire [31:0] ax,     //     ax.ax
		input  wire [31:0] ay,     //     ay.ay
		input  wire        clk,    //    clk.clk
		input  wire        ena,    //    ena.ena
		output wire [31:0] result  // result.result
	);

	fp_add_altera_fpdsp_block_160_o5ob76q fpdsp_block_0 (
		.clk    (clk),    //    clk.clk
		.ena    (ena),    //    ena.ena
		.aclr   (aclr),   //   aclr.aclr
		.result (result), // result.result
		.ax     (ax),     //     ax.ax
		.ay     (ay)      //     ay.ay
	);

endmodule
