-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
eotiaC3jbVPsldfJpXXmVfIv92c3ZFBXYipM8RF85agvGd2IOZfivhlqhXc8L2Ye
3gfbREvfoi+jxYZHivuN4MgwMzc+WouT0TLtuvWSl3xtA3GviTZOG4t9d3d7WBmG
yj9BoteY81BfRCXDHkYvwJLWLvn6t/g/DO27I8ytgmtNJOQQjN3kgQ==
--pragma protect end_key_block
--pragma protect digest_block
NN2RPCScmSd4v4+ZxP4qzaLZKys=
--pragma protect end_digest_block
--pragma protect data_block
o7baLs9TjDGy2agpIDLEgSgIMORJJJLRGmgKooJfNKS1b3vbmG1sSunl/qPwzR5m
2Vuhm14PjyO8wGviM2g2S2eMqw8ITjiuwhLlwSS6h/nHaApHkhxq6PxziqpEOSE6
bCGCh30k3p+f7USBhcNoF3B9IydO32M6WXTxMgEBwaetNDbjdNMjMwnceqU/oPCE
gZMrcysWgy8umVab+akc1oZyo92Kd9gTQx0oKWz6ncazaX+kCtG1LrRABzXnyA1t
U7pwfGtENv8ve5n3o5Lxlm8SmyFpKsbWTamm8h/4bSVYC+k4gIkyhHhkYEKAb5T2
1eXGPbSwvZw58a8x6RhsD6+6kuLuMi0POmIvr0Z3A7AITPAxOCxUy4zviR938sem
IYsRteJw0mQlxz9qK60q8wmgaw636gL/7tWN2Khg0xQ1/GJ2diEp6ax9R/DR1ROy
l/HLkhSRnWzGyD7j9Hjz9nz2FG2Naqpy8CItVEjD5MraqfOLXM7O8/p/RBEy8AYi
oXL/dl35QeJH6Jop0jWCNaPv9sCxd7r60RCr3OL0isj2/mMa2URiQpyMidhfv7R1
gNoJ0izxyEHKAHL21m6e4laL7xDT6QlFCR+8FUYn8cnJiIniZI0Ffieqq3y3R3ba
F4LE4eLiTqNdzmJDdI6uT37yAilWt7a1VyafrJRsjBaIL7IYmd8UXxMISQKTPi78
p5G9F1O/ckc83sDnKJgWJ4N7AMdc6KlGpYrEgFH04VFhoG4iY2MG9Mtwdn4mjHIY
TN8gOS+sAMh42OgOdLUI+rdQGa/EEivJOtI/JON3ZNsCO/fN1M+DmkljcC0x4IZ1
K1o6T3MGgixGuztTVMz2hCjLhH5bARTh+YEk4udSlKU4T57BIo0MtoI+/NHF4H8d
iFNfQko+BbWUKqoaB7YJAA4zySd6GVrgOJrDVPIPOroWJuXTUkwIrHI+ktsYOUty
loIkEZGJrrb0D6WgTB1oRJnPQTWoKWRI9g2ultte0l24wULiOgKk6nfaAyjq9uz3
5qW5AcEJfaqx8/JUqQljd8zNfLFpkOlKerFsUU4p9+y9+j/bniI92isDbrjx9ym2
JjJh6AMDA546YggxDwvgWLWQIjpzuDYPy+BjXMVKs1b7VFyxz7TD/fR5gAJXIOOY
ZW9AQ9fqGdjGleFG49+Hvv+Ol4F943VbKyBppSEy8kHyNbLxMiPW0rExdsPocFuz
0+3JOomzCthJizts9AoRocNxHtNXqc2KV7Aol1KpmvTD7qe0IaJif83eUZn769t7
iHA6HLz7oe0y0AJDnCu0hHebu/THV6vNFsPtslBseLEjKIzuOO/PmXAWOV6Qg2fu
5yVLL8i4NmXlF/bIE+EC59/S3DH9/Gzogx9m7ISvBzt8XkSp+KiIXMcrHsNX3Yuq
OO3C3Xf3n+eWRxxCWbymwhDfACr7Q4X7QoJisxVgv1qLUS+YZpgMSqaOuUvqeDGF
ds4ELl5ylgsVTbsMTwWF671eeX674iVb03SMtkj5ctk3vGYzjxDjbgBvbj1Kah9q
2Sav/veCSyWNAIz4DwsyUcfq/GlA4j2CPkX9O8ti5aS4BhUvQEq7xmrKcNF+SeSm
PhK+OKE45CU+6+sjso2vU/WUtlhE4S/tHVY3AuKUpHhPizHfL7l4l+X48ZNURavs
4ChCQTtaILrWJtKN5832GT9bSOp+IXiz7amxw1ZzaiZdzjdcKKPONnFBDDPvYOeb
6kNpHAighDKYDN1gI2aKL4S/GL85vFn4nB1vpl53Zb9Mx0MBb6aI+CXiBAIoKojr
IKw9YOssMcuMAmMEbD5nAyUDUhA07Ukxi/r50I0ply8TO9s+OTsPMstrdpEFGTr0
KQKkc1KXc48zU8Xt7haBQfSA5j/qNAMf9WcOK2kLDgN2j+VIGQqhMdOIIfRVYOq2
DbGpwkkCOZgHV3/Ok6qUewXPxbY7o6UVqFxsC5eQEr6EWbjiEZsb9EQBr27DlJi2
FBkwDkNJ9REHkUg5/8O8oo0GEnhbOsID3JARObeUK4/dqXC0ZjUO54oqmwyCUse7
EC3AwCaLsyot2aNRNRUUIHJPqIHxuZBRoBQ77zBQqQUmpFWwEySXNddzVGvAmIYm
dj8Wr+b3XTfPhb5rqJ51l9Vyzi9L6O8DMj/YWPwvUBmwfO82ffXqvbpJZazmvsWu
V7BdTLyxfov7it7Zus7HpjX0eN8sLjYTIVGX+XZsvl5q5MZZrghOr1CL1L7NLBGD
el/e/7C/Ar9r1WfRoOzAj59YSkK4GBvMfXGhANhmA3VntM4o0ffly4k9rWvTrvTy
2NtZb0tUwiM07JRHrhaE+9imOu9y3/e+6lPbvjvN+lkZysxHhJ8z9CjLGRrab4PD
DRWb3WJoNGTUU2QOWM6E+0flwe9RI398riQaoVzUT7Nd34j+AIuNWz4+9zqnXoLP
lAcyRvmONhu/ht31pMSrgut0/crc/onZ5Mw7zZWB+KRTxtjgTuLIFY15/ScRkY5b

--pragma protect end_data_block
--pragma protect digest_block
WIg6mt72gAV30PEuCntyG7rhPWk=
--pragma protect end_digest_block
--pragma protect end_protected
