-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
TYNwXRSVPRiFo3Rcgms6pTPIkuBLODKG/y6AiBKT02X4PRG7HjCSBSJ+RcdKiSyW
cEu5lcQKq4R8DevpgizXRO/y5USfFW+y+O/I0MPf/LTlKomMtR8nCexvDbX9Kxuo
Qt00DHvxaxFaJWw/mqK3Z5Qcep1pUczYuzbUQ581yiM=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 47964)

`protect DATA_BLOCK
FcfdjQQKkgcCpgnIkzgTFCNlcu9jubvdC6K/5QFi/bM71RghXe/D4zFdczPt+WXx
e3cRhPSFlJHVBEFzoRdJLlcZxCnESJHcvKo52ROIGmojaFRNY0EKLITNF2ONZ3v3
Yi+VfpJ97wqsKHaXI2KdNWz9HsxV//yJI8MHQdMNTmgA+9khKq/buBSciH9TW9OQ
xtrzTCYmtKgLs3LfHQIBbT1aQJlX/KobTo8t7BE5eri20paUMhV7E6OgqjngIVWZ
ivCsSMOtMkI0P2lgL8CsLd0+r5wG5USJZ9/HFaC/ufVQOO+EhlZe6WYhRIPmth+D
wTVYLbp42nZpWB0UCwJSszG3nz/xHFiJkOdUsBGbCCANJbkQJc2IT70v2X4NPLrG
yN/isBB2yjk5ploWvgAK6tLvaMLSmOIgzWDTJ8I/gVn5EqfByD+v4zKJAx3Cu0FO
6hwYu14rM+bvPu4xjHD8Pb0iJJYM0K/dG7UPaxXuVJv+vxJyQLnbJDkCM7rmqw3l
7bSfmiaqf9QpBnsOUAMJlAjfx0X8zetVYCgXugwJY/Sr3Ux92LHDil+0SYlHcw7/
ubkUyma8uUCpzaOmZsYYwZCJIwz19mn9LSiYYYwuYXymUgIZcc25lkw264UJnLBh
qQ8kdPnNljjX6Hokl4MG00NOdaK3SeQJT3i2JqYBhdoutAUDBSEQf9O6CfmpkFDh
dtgwX0crQty49XTP0ll5NlsR3DzQOBu7+UyI9UzZCflY8t4XDavuCsJsUCqOzOo+
JE82xkOejRmIXWtn7aulaUQrHY3qegDiHZ/fq3RqfFAQwwud1x7cxPbdgs/DZyHF
evMMfllrp87FkZJ5rWiwAmtvKKq+jSut09W++T6UgezgbsNbibJHn5I1lJEbK1ho
VnJsMePQfyLV/0CEIHdFK+ir3VGLP+AQfC5AyGHxnqWYGhjnbuX7L2J3GstzRtxJ
7R9FxDEmxmGSEVLYuEkkAs7CQRGlL4FRz7dmzx8YFNVMltQWTyhFVyqT8OT+snrm
bldnbNAqsjzmW5Y43+IOUtjF5cfnCQt+nCYT9SYzn6AC2BRnFlCLCWb8h2VOIZPR
SDHhhQtSnTDA981+RiUycO2WwpdTozEPA/0RHrrTb42BNeoaE8Siq/Nme1TZ0NGf
nVTohhKHMaWB7UCozubIC5ClVk0cBz7/GWIqaI7z0M3LQY6iiBIEFxq8dOX7faPA
eFrbR8vJTI5tspfGQat9JI9s5VGr9zy0uzxB20mS7IJndxfh4AZPGwlEiLtFdoi/
jCFsY5e4sdjAMBPFJgfFtvFaQhkaPP4dXGFjHIiD8QcQWDRfeQX/ldcoDwNsHAwF
VOyvydf+fo/+p/8fBcYwoa4G9UQl7A1sRu1p9BmkabZV49HQvPOFrtSXhZhrC3Tx
FCAAzdixq3DwOiSrcCZOUnW+VFojFqUESKI78JX9ZaV5FI7EQF9sscgae0anxwib
+W9vmTqJl5Ogqze9IyJlpp6mnNpoC0t+CBlPHn1jnse02FR0FADts186Tlm0T7X3
8wkcdrTz7EKcu7VTKOjj2JGC79zDGWEBMFaTPEbNmBPQP+ajBs7SMImrmD4tXZjN
f9HGwnd9Z3XU06T5UDShUNAxoCLOTkhH1qAqnfEcgtfhVPiWg3MbJOHCzoYagGqQ
ZPeq9RZm7RINmaQ75OygH3upHyEoXfieQLLy0VW7KnEnF7xIArQrcs0Rm7z23z0E
tmluqdqwW1i0GqoWVTg1VOcszXD+JBDZ+uRnZI2FEKkuPkn+burnGHMGaVk3BCVc
cvW3m6RDpfAh2SVjnGbzKy8+oV9M8XMyi5Iuv6/V0Ybyd+EbydPKzDDPFzY+LxC2
nB2Um+80J9LZNG123efyRDDw5fJiKJ0GC3II5WmhKhPsWbqVnwlnHghAtvOKoerX
2FsXZF8TDEypqM8AEibbzzomVmjNhb9yfUxnRLqW/EmVRrNGaCYpvgDRktKxDxh6
aOI6GOY+jtkGvRxhF4hFDD/+dxhWkkXWLGLiVQAxV/wPlZjjSYT10XaeaCedJjg5
t+PzLJBno2vpvYaJ65fg9g65j5D1OoPWJUFDkqgrwMyvZxY9mbbCTPl3vrF54qq6
iRElaNFmM2wABb0Cipz2OZNlYSn5pTIWaMx8APEkhyyg8xXA8RamWGOncjswwcXV
wIpPRbFBCqvWHwDy6M8ECYf6HjPdXFQu9lrIVrJgG7NvfuB+HgMS6yT7E/Mn0lak
M/oeL6zWotLkwtMlnAl3U+7Yz1hHH6r0gFvN7aRrYV9vr6ykfXFCtnvRxf1IXJax
ihIrjG9Ve1glhZuhZZ2zMidAEThUSzvOlCuQuWxLLMzTxm0NNZps9AunHJoHxxjd
ExfsmjPsHy1KCecYQeH7vESXrs5gKcJNLZ6qs9VV5JOcX+M3p3Xc/9lMMvjUnSG5
OQDt+oJNb94a6rkV83dM2do3Cq7JgSlzZqVM+R5tLIqSthuCiEz/COpx/xhEd7N9
g1gGkZAXerYt+BDZMau0npeqCGu12MQXnXq0/GJ8shMaqXBlIt4WoxMftlNT1vZh
A2cXrGT3CB0U5+4PcGa4o9oJHvd0ajCySr/4AnwHE7AcHt0D69BH4xdOyRC9qq5G
DkJNFGGFPG3A3FKq41XODL+OHddLSXhV5ewrkNuPe98acqN98LMqqeIAlPVsdlu/
ldiiDLdZyaz1jYDf+Pc59P3DUlc3FCglK3CfO3vhhNyLNBuEc5K6bC19A61+eyMY
SbvaJDwiMaSHXEPKDFglXZywECfV7et8v03wqyM3w+g3QNWQq7dVLJJAGX5oT/ym
SMZlP1ZpE28f/tAvyhhPGuT3D6Y8U4VhCCiAKIj7/JVcDnslD6/5DeH8dP0VBs5C
j9Hgd2Ypl2HFNTmuZDG63fzoO6AVr2E5ZLvaTFWyI43AmlE2IVJAHDfwtHnJq4Cn
R4mWoxI2oUgC9axnYProsn5N1KCO2EBpcu186OE79E0HHeGmyFk1IIh+ppS+1H8k
UWHNRn2w1NLRP0+fCe/boPg20I1uFkIBkTQUE0A2Ag9yz41Q02+lwNGy/CLouF2r
W0I0NqBjIXlo6yxjICytvBuyQwuC6T8kuKYUWvJTpV3Ip0FCIxEnZn5t1bHVkCxx
WQkQdcn9y9YANJij0qLth3FNrpYiYJCRisubTab8UPkzxG0R3/HgOhrzUso/L/SD
Z1FA4Cr6KHlx1Ww1kZkBm2PgnrQAv5di5Ka1GKPDGMGTCmVsBI6fODl3VROaLTxb
5vbMfoZuVne9HTqQob4BCghQj78oDHp0vcBWqWzvUZnPMsE9tK8EzSwVbPY9Manq
ahq+MEsW7Cf14LlfWzgtJh9KMZiDUGyEhQ9tNCtWRNqDAmLRDqyc8ZBtz4Z2g3zB
Mkr6CitLdxdxa5I1RmBzSEvE+CznDD83sDmVbf/Tf/Fl3hv18o0wJawufPco+jZR
J9QQLPHqgzU62vVv/9CwdI52iFNjnYOLxFx3Sga15Ex+IheMEH5qbN5HKZ55+loO
j3rTgHEcfhD7aBok+irsvPMpHwB1tltWgAdaX20Eg74lwcyR76qMVv/HwubuMoQ7
8dDaxqH1ZokzbQN0qp/RvcMd0yP4zhhoGSb6JdKWBrhFp7Wpb+EbPJWhtUyc37zk
WYo9QDYTjdhq/M30R6IepAEF0sJHTykaSyVlpKineoq7l+NC6KvCPORyKrAPHkoY
9qTR5ReKsk4aMlmx7v0+BXK2MPQTRrBPRmd7eAiZmWz7w/EV1HnvfSj76enY8mGs
O4Ag0YS3F60QP5nl767lZ58xravn6yfAm8m07ark8Px0LQeUASd9O/w1w6hdVwc5
m8KukDFzX8aAGLYNh0JgCjDxzUgrAh/9KUgJUfEZIxOMabA5A89FMIoAuG3JHG1j
tzPDYLA5tLob6jG/KEtsmH/9tPwyy0znXbunk9rsekIJwnkoDM2m3X8q+idsfWUX
rT5sn/UuZnrRldcCa2GeT7+ynT9xnh8CXARx1gCanbn99MS1d3kB4LhSg0V8obtB
1LH2Xt7fTL/WhuSd5+10VbbSEUzrJDDRjA3+AxxXxQ0QSFoanPTZUCYQ6wJDIPfy
7/vHlZL6/2sp9Zem80v4lQ3REEBwy09DSP1FT+PrdsJ2cKiycTSUTXx7fmudslAb
oP4k6aAnZA3xWxMcnmBxStqO8ErlZuo5X0VShDON6U8CdVTcFbsLgp6fpeA1v5Wr
3kNPzPcUu5eNGzpBfdBxUJxur/ov/1ZkCraOmqxOM1VZez7R/0MEFMr0Jd54Syyk
fS+cKz+4lkU4JOxmbrbiimcxGnp3g41ZSN8+HcJdN/HEsueUIoMakv6HC7apMy4I
dz5gIL2C8DXVVKfBOqymxD+cH6SVyv2ARcFLheYK4gmimOYztNB1SuzdGzpSmvU3
eojaQxGJ7dpbxq69Q8cn+K76WAizOgrj+pLy0plyVS9H7HTDnpuf9Nxa4bQcETXB
JrdniyVot5+6ra3zz6yvqDx36UC9KH/R3xAwPHDz5o5O2NWZ7EFSoXRRB/X6uJuL
cHDbuv3ce2cozkR9Qr5MoWnZjwqRdsXw1p9jvXbdURQxG21yPCtXEAZZpblJNcTZ
oj+4MD9AFM/2iNs4w7HH+iyfzUwkUwV2kk1Vlz1NsVGy5+LdWd5RSqFAErEJmxyG
5w/Q/wNNO70OqcoQ7Dci3joktzIESvrLDroGEuN6TH8jx/xiWLffOGKy7i12xXxc
7kpdK/RpmqogBQ0H1BlfpffKl9kzuVVSnuwXh1ETppsXSLghl1YjIXbqZLb4agzS
jcsACSGAjqWbsCPaa1rA7TkY/HoAazxrUe8ngo1xki8SyNWftaXVjgYNOoGy6twR
rDQw2whUVCwa0oNF0jlcNVA1+D8cCeaXkv1Foa0rcmLN2Qdyscn0eFvu+L+QS0Pc
b6cYx/+Uh3sF4+fsVrH1j4fGqTf5ap/NlMFayUU7lJJ4yha0pF6jnvbBOh8AtZNU
awEh9TUgk80o/7i530cWypGRy/ZhxblZDkETP6Z36UhWBwKhaykV+8MJwtHTaKnJ
EPg1eOb6mwQoV20bruM3VqIoFppz5RjXP6yuWmXzSf/yeJ78HecTtOfgzgvjcBW2
YAFvqD7k0LigKsvEUGwtXYkudhGPtowrup2PDKADhPxZKmIIuz907j6MYIxtmWpA
G3Dvw17kgWO3EHh/g9OZhHxqHTzj6mg6LL1mhZxUDcpHC1/asgv8KW/oLTh8PQOI
mdh3kzZLPnIqlrwSo85gUZ26Dalobig7t+LOiuaEi8JbzgUnT4reECa2nMQXFY13
izO0ojw5Ek5LzL7GzlHuKgdCFnQd09aA3blMIP9Jl2YS+1D4IGji8O3iw0m5TeRX
RH5tJ1165xo/lqoUfpwiZvccDnoL7ZtTc2ARD4hDaYOjZiojXBENaf4bCe8e0c01
vnihJ5r+epF0AkTP74Lcvf1bvgV6Rw29hEyet6F2BpJuiwjeyPp9sdnYQgup1IIC
O6tG/2Dnd7yIkU/Zi3zG/jDcbk4GlIasMnF0251h9qehkSuBnqUdqNs0fPMcSbBR
FzbkyafEfSmz9C4tLs/cTPwTpzgJ3+AoUACrmv+/xPqnGYqn+aUhLkvaXyTz+Uzq
t/enfjiu2IHvF4L0Ywyua7nj2W2NN03McU7f2QVYMhz3KDy+SXL07Z2Hq4WZ50BL
bFRf4UbXj+CyWAVKhTPFSnlAeS7S6mMAc/5G5ibCaACmFJQkGA9NOJlQPH6X5Ckl
ERbBQF/itCXkFZWYxd+sXUv3f0GWoMs+3oZa6Fjj2wC9sHeSTzOEHjShKy52/gHf
Ih4yvwhWO7AsOIBP5dxXXLaHFZjzXWPUJrQeY6HgO23ao0yn+wSEUOEPG1noxtER
IJYPVP4tNR42QoOCdUcSjxYjpXpN3SPLt3G7E/OGnxkybb2i1FTtoFepGcOvNpDu
dMRzKDNdhn6L14slsYtGTSJmMeakCrYs1ts4Brp/lID8YJcz9VbhF3mOe19HODqA
dQLy+t7eu562st/TyXVhhUw/7G1YoCxt/GJw60Nb7bx4qNRQGUxmcdv9eZ/4WUCT
DbKz3aeUxMvt9VeA2Za7f21Ww5oVnXX8WJxqDbSUiXMh7TQwvuyKQhnR2SBL3qEA
XobiJS92K1NzvFqKl0L9zRCW5INROpO1sADcIKTS4LfsIAehGcn+5qs8NtPXBPRy
d4kuYNVh+ONWKEumgQaqqC1cywPbbaLp2JluYI3MYjTa6v/MbHnDGbH6YD6X6R+b
udlQbbNR2phgMJ2f+D9Cht1exUB2Hu/F77+YPzhkZHUwhh7FIMlQwHBD3rN48hpf
pmCTrv2Y4UimH6yG7o1aIQjtjNtdFmnJYkkjSKj/fgQ1vUnbXVGOBCzdUX8hfQd5
yVMKh2kWHxS4ZhybTTovJ/Rog7Cnki6InwwboyZsEfNLUGRF0lhydbaDf+K/fPOJ
W9Jg6OB0+ElrFOIdImvFNWRfPsOwlbnuv4DJiOKlqvf5+O2YTLMKtwKSFodRvykz
em2x3AyWwbx5/8TCJ9iunKEzzP5TC6xCAhlC/ngseCuTzIl7nVetfkuO/mXtlQQm
/yQBX+Hyr4M3r1LrDooJq7qz28e07rocgxt413RYlpyP7g4mLb6OMjuTiyBhq5Lh
AIPhfA/CDHhekDOc2OUYZsfHQVREG4XzscglgIMs0RbOAz/2YpyyMwWhU8psKC+W
tG4wvSLK40UYu6l8M38bFnGs+0cjdtvbTphiDLdg+Lnr9j/ZfFfJ6W6WvaCSB59e
OKc6X1YMp96uxWc/cFQ7EaN910ZPMKl2RLlIHtZOSPCrqu1QUTkHPr2GlSZ/3XPK
8c3bJ0alybIwKquTFkY38HeYzQ/Bs2ET6FuuTKwT8DxY4B6pLqWz3haEnn64nEGr
zoI00GqQtMhz5GumzgsceiNQXVtf2mb1dJKWcGpOZpYCEkMBSm+/wd5tnulfV20E
bLNiCPZaV2DPOtcqxS2fNisHvln/uzwOX2/11Ght92PS/N7BWpljkfCh/qanJlN5
qAdNjvIegbFXTDpKQIFv4mZ3g55heozKrY3nEKY5kUOEVVBXEKlECUR3W4KFmJWM
T5KZdtohy2CXJyEQxpoC7N3elPKqvRmkvHJKxVc9o65XSTKTfZcfPmSrEW7N02O8
MCwJ0GeY6SzeLd162egtm28wzyO1KbT40s5Uo8JnNxCFxbzWoloImMfagKf8L1RS
tkZ9R74F4LwW7ftgZS7ypqEJbyYknLe0zT3XI6CZhFaNPjq4toGFXQTqFiMSWScj
oEi8WHwsCfbheNoOxLqz0zWCyCgVHSaWIWjRwkdoPqL2lUCbQSu3EBp8GfJ9v3z/
B9kKd2IppuhqxpdoKOniMrSwxA/xaks2kdeKVNRB8bzruuX5/WmCxbJ3jjBNF24a
o3rXKyc4oZrvPI3AiwVfcR97Ra6hsaEbB/SBajJ8sz0xgR8Z/CsZKEdoxGI1mpgQ
FepoNb/aAkO+vEkl8cekhxpEqBon6UHAHfpXyqDv940VwqbRb4h8WEGeYdISFRpB
s9OZb/hUvtca7fbgIUp4lS5/8BLZR5vT/Yg9q1Z/yWTztGQjaS45aGO3qZF/5eVP
1pJpOl4lNpu3TPi0+KIUdd7Fi5vhXydM63iWOYnBDlE55z1ldXIJiHWxlwcwTFiA
6Ppnv4WDzW3/pilyShq02eAjmzLDijwcFZYr4M5WaFIlN4qVZU72hBYWvhcc92Z9
an/pSnrbZUxBI21HBrDPY84I2ZKXmjhk7yiWhlYSpHgzFTyzyc1oe7EY4Viv8dAl
4JBMJHQ4i6Q1bFGpYj9EOFXY+Gqv+ngnJiOD4LEcjOPRtCotl9tVMVjQdYJbb44v
DOhRDc1VqLoBKRazYQUKoH7mpYJUoV2e+KZkMZb+rqw42ryIf/SHD5BqMgFXllJ/
JeO0hMmzbJSYs97t0MmcJySvXEh/bi9xP5npvMteSMuipwItKSiFQFPZvTOO5XBr
RMLV1hKL5DZXuE6DzCwuwYPUKoD3EZZg4rPfhE6b/K8OOIpEe5HWiBckD94mzXB6
gbaBHvJOfbbUqioshiZXZs85hYI16uL3tswmx4RAViwtta9OcRtT5hJaCER2s8/Z
HcR1GIq0fCexFzRPzFSUtVIjuQMJmwtjFU+CE0Vo5dFscCqkivRwkXCluh1SQMnd
Sa0FxPQNgZLcgz1nmWQBwvuDzq/3LDIehAGUWhc2Kp4AajFV3wGRAAz0ygYDiIAK
JtMOE5jTHhmJYDTDTVPpGPqxm36jJdZOyjcKnMmRKwqP5nXVb+j4pOCkVJF3W8/k
bmzSG1mVHCZ8YRcEpamz/I4ZMpVgmEgg6TIlHQ3QnkGZ1TdkwAnQGl7cxlOoEFry
jHjpzXIOeN0pnPtvoeqISGXzFhYHQZsQ1TnzWJkNJaJ14vSyc6/kcmeawJYwFwIs
5CqH76lrXV08WSTnGCMn/4y43Nfn5xRr7VkqOvomGka+CyoJ+jBNPrWsQvpnFGW3
dx5LhQERrAcLD6z3sspMKEIu1sWM+5Kx01NxxutXxvOmrWThN2V3RIjiaIpR8d8l
0HYr6bldStRAIMeafKYwTUvpsV/kggDM/lYtWwx6JFBXVJ1dcos03Iji4/gKxeEi
lHskHUW+yInYVf6XbvK0zcIkWiGzxG03FHWw26g3bqXhiHcofTWS5rGbo2mHBfuz
qJnUjojn19su72Wd3qdvMTpREs7IPqERuVVBncQ/NH4aCpxLtPffF2x4tu47qbiQ
EMy3VcrkTaUoQhTt4nY4aVqymjXiPSL86I6mUXvaQ5S0N1hoiV+Orp47RoXTSFb3
JJ6nIwp4TgBuXHNPwRihnFml7dgxjZ8qX0QOX8VG9gho0/d19TF+MqHTZax9+55j
TiSvpBVYX1vAGzsBZzPl/frKzsUTiPONaDr6sfDBDIfmyjAe4lPOAdAmrMfQuX9s
/FoTjxoGtpobURgGzTqmGfo1sXEd/MwBdIjr8dv12CzvBlyQdHBbw0IKA8Qg0BW3
eBFWFmYmDKxjoDMtAtLtsd12YNj6CwI1yayvFW+URQsjKlhcazNSRJV6au7UqNUn
074YkWN+DqWJpvaEMlA+aL0LmLk9i9nIK1OWOWVIM+YltdnDZxbj+84bHTdzdCoD
zFcdCe1lbrLd3BQknNAuhptfnSEQZpMUTvbMQHGbBdXe3/5p38zG+6yut4ZFm3L+
6fMc+Y7mIDNbjLJ157fcSNfBlg2LLJCXdVfWuDtvs4EHD9j6pC+68jUGqmyEvw+b
xshmjv3FvwO5aIWPbuPEJoq940Ylf0KMy3TeYXtkYVJ/ZwMS7gTxzkxnaAtZV2hZ
R9gFiF0LlAue2w5PVNYYJTbEEqU2paYx10UcvMPK8YZm9t4682E3aN14c70CWLei
KLYYbHOplsjhshL/o57CYY1fgbYy/kY4fIYU/GjbB69b3l62qkjsUekmQxcDlJB+
VYsqOrFkyAWS+YAAoM44Z4BJiAJNMVm+dlTm8LFNFqaaZMjYHMvFyi8LlCo6huOb
w8dVYP1T1dXsYNaGFl7kHvSZH2U+w+JJR0Ys3N8WdQkGHGGDHhYeOVl9JhiZBYC0
rIE1B06elQKCzhFSgTR/jKK70MFtOQB8911GxHE/QFdfZ+Jd2RNGcuLc5wb/Q/za
7FXV/4s1waLaPVAwgamHbjhmnV2TcjgrdNGGJFW/EhINOwRdY25+G3b1wTW16ifA
xfwhejM5BE4hwF30jM3hQbd9TM/5TsMM+seMU5sWi01h0s+Prv/LJG2Yk9lqiqAy
zyV3LanvyLBfVeghokAUAnX7N1CD4gqvCK2ZLrvdth9XTWfcDnYmHJexodp4YZAn
1bwpXCSH6veYxMwzNDzBFBiVD4HewJn626ufq6dZPZ9Rf4atNAQ2hWD8iSuSVJKe
l+Ejj6fs3XjnqBGXUjI4oiSB2lnVqKMdFlxmTaBqY+EqtOYLYMgwAacbVfm7TQLp
/eBn+M6S0t4PYAf596v3FIJKiGrCsFzNjGGCv7cRcu9JT/eQjky46sXFIMt1e9uh
2hxT/U/XeLs4z/MpEhRNGcKLHgXmlVzRda0Xovioxx6RRwSSXory44m1AqShmT2v
B57GSp7cjTu7D2/nbWv4IS9OvjQSBOXL4sfM+HRFEda1dm2hbgeTdPMoFgeBvqUS
ILt4gLUYq3KgLvvdUKr0x+Q3Aua3Zk50PkbN4tOGW0S3Or2aK2tICO/uDYxQ6gWa
Mvx3Yp1wkt+NHSPdYY7brJ+/0eCAUXWGfYaNd1LGVeYD84kWCtZbsYclfGtTsadM
f8zkzQnXSCiDwTrIlSz/huVW6zMcZwziB96Vz+V3g8ypM5ZSQhVB5oBibgU5cPuj
O8I1f0WjqnfAO56M0Q+uBeHAENFQmQUs5sqJDn5UGePZl8Nc8mU93wPMUH6pFt+7
idHDe6MWyAII9abg4xXdYaAE7aZqDB6zJcq/X1sYvoTOTyedhKK5MaY7HSOyiEBJ
dFCnpVy8XldbKxLznbdyfECRNUooGnjM3xXmxp4iUa6TH1AS0fYH+Jsdd823YM3g
gcPruwnHA6fdZqa8uQmrb2LcPekTZPtRugTwXtrhqeS3Tyjz3Kesh1Xr1O/hD3ta
1lXYrb24FKpcNT4cUEw5u5cdm/QrImF2KWhDDfLQq153x6T/cpArzvd1vlhxZBW6
xeGlTMokd5Nj1AaM0OBoNz3HYHpVLLcYALPM0RERkwtw6F6zNHo+oaDfwBm0XUw6
Ggq5hqz5nsH6lsAfbQaQRTVdYNNw0CqH4WBIar+QhdatmP4mUqqq2s9ge4qQCj2Z
PeuOMAblm5ONqRTew5x6Ka/Dy+AiYRXDGRCSJCr3uEouArp6m9R7y8xtOzeC5cXe
tzNZpW5rBMOdYYYKO4dyBOdLys0qI/Jw8VDsuYYyNxD1S9N0/2ZC2Nw+KURaMKy7
pmAZv25vENdbmqwIskmnjWLKnSKGedBvt/hGw2jNlQsA7+z8z6yEaRZqOmDO9v5T
olL4vUxNrKXUb1K9rUq9TeNpcj5Cl4dvlJTrJa7RCZZzEb4VxrOkIzgz7VAQaP/a
/CAkqwX2KGL9ZBQp89bltIsxd4ScNsd1v0nidvR22ee09h0RbE57VckLuZfz4Boo
U/Q/BUYuW0WEH8295FXSVUS8VvVVvw8QJ+UbwmqYMNx0JCLWbp9annj1F0xWfy9B
NIqQjW4HrONDWpwIjCx5GvRuY7OUligzLKRvWpnw01YQiwvlfU9NNWzv9zTbM3kD
oSClUCTM4gaRs8UtY3Io82ibfEEftry0RtwbNFyOovztqa+kjuNAwDxZLYGJ5AvB
r3/C2O+ngw2Uk8g5wqllLNMIELe6s+ERAZYtwGDSdOq7xRjD/Vu2acbc+hsS6BC1
CO98h69N1Sysp7QcyRS1NHQMUT3lqResp5yFVVM+AAugxRJW5VRN/gw7WS9iKk+0
5uHwI36bqzCu2un3ifI2ncj0+sYXjW7mGWbKeXYZYqzRUdAmJhjfXQhgUQIKXLff
0/foNGZ5fB+RHKjOdCTUsp63+BAlh4wZUgOsRSWHCRRZ/0Fcv7rM3NVerkXsSOgq
sacTRUhzUeMiDpgOok+jrbonHJ02A4UWPCQpdtIA/eKk22/5JP+XHzRNDzYA2HmU
IFHl5up5DgQVrGnft1eghI4n2yYG0FMBDquZm5LsCUuZcoJGr4Hi5QuX29PMm7v1
C6Rkba+oX0XxefdJ4yx3Nu4yOBbU25+SLSgk1s7SdwC5HvLjstWMBVB2xrnbmMtT
9C7YvM/Rg4PK0ZLeSrCgbZ0nBpQatCHEOrNrOn/UrW33wls4rVN2+LFhUQMZWVJY
LIBRGA4NGdluKitvlRffRLOukaG0lLJCzNP19tVdAcmRuehmgoQ3zUpNgQ5djD8E
jhnMPxWr57gBpqvsMrlv2xj4sJL8IjDqapYfpDLh5/0D5jKBVhwUFx5is+7PHxlM
jKthJQJMyvLdhj4aoxkOB0Is/Dna+CpiNSZ7zqy1tQc5pMjfSrB0tPcjeENzdfo2
Lld8GN7LDrVSujX5HJsLBWKOpuc4dggDaToGlcOMuF33nrPOQPLA89u8CDqwV7Op
olnkDoAewe8dOZvuf2qPwKyJ+n5mwgqvepCqoB9Pcv8C2wmQaOr9quMI0Fu4fdMb
ULHRba/DhIwBrg5EqFzmeFsuTAzf6ep6iwtIBy8nlkS/5AXnV50AlY1xoCwNmuT/
0RGl7egxDDCk9detJK8Lr1A1jh0i0iLaEf1SoRoHDDwfUdqKzuZIt824Dm28BnUg
/1hHfQz6LkIxbkluKo533Bjrx6sKLdfTT3jHhCD83ADiKH69gS8iYwgaWWOUvW60
DIUgmhJsASgyAUtnZ/hNcuUu3JcKK+O6k7HwSX+l70j8Nl1uDr1/3hTrrqqJSeNu
uu0fXpyNoDeL0sJwkyp/vJS2T2o3+d/wWBdmmVKR+cwngZc7YaNzv6EkalbJe8/h
Omi0bVPl49zGs+V1uNxTcBsCJriNs8A2afsXrxQaKvxtQCiK7TrLt6sPB1lha8D0
VsK91/TexkJnGkc/HQiV0SRHwHkoCk9MOwA/o5sKR/XAuikth6T033Ir6zYu/OWZ
/q5HpJGYBikQ0DLEGcdboocl9zT42zBeT5TvdKBp8iPwTOzxviOkm6UgfWbsuTzL
u053keQYMJpStlFBN80seCz4Fu2UV7IHIar4hV8egNdtpL4mC5r7jjq+FXiBla2p
T1aOR0m/hOObYcLLNs24v/enMB5rx+zUjkQI+clMRP1ND78w8uUM/iGE1USz4aDh
cfE3J9gacFREBBMXDvo36xDLcyKWZIRsFBUeaH0YCLLogZoI8WxXeh2ZInTV096b
35QiLgtOv/t9vCZT60SZgf4XQMPISV2Ep0bVsypnmsVmVdGPoW0WWPilAxBsQeUH
amK/t9Yg2O+kPYUB2AZ22yKP8lTatI1xFhE0oKIOk5lPLv1e4yiteDrvE0DTAFTe
S9srUoDxte5GXaUv0FqrH4AjyYzJVggGMUzM66S9COxX5KkTVC91+uAHgg+8Tcmi
LbE+R1topn9dD/4Udz4HlrjfbvEKZIp4TzPE7UjmziT4Kk64dax1vVZ4wvDU+EbK
Jh6o6CtO03//njuFIrl1PqVQRV3Hi9UHgYho705xwK5gRItMbmVGl4eqmpmpoVyj
OKg+ge0No34X1paEcNGGSNeQ2sYmHGZLIBiogbx4MJLEelNH/Zf1SVnUzm1hDn8d
D8bHhEFI5tBACwYX8SfouX613R9oQxKKlOOPwUsDtqLHKhH75q3S4Rmy+W96knNp
mFraVXiWasEa3dKZw/FdnBcDbEQFJ3XyANcthguu4ojDA88zkS1ISe17O/cvF8Yj
zTW9/Ecyr8TIalnGyoSo1x8WO2Wqa9vaJq/A4AQiMWoR31bTH4EKf/QsUTDpjhNF
pEMW1tCNupli9dWqysQq8rFxUnzjrGF0alQ1Ywpfuq4SoG49feg76dRUBM/ZZ94q
jT2NpjkFgAlcBvCyFYHmE47OJ9otM1WZHqUtutwqLoSotro2goe01PgrfpLZMJLN
VXGlF475SDTpbS4dqQWnLY0Gf0zfO5H1nY8dZgVQIP0ocKi39LD2qolvpSLiTKmG
FcOF38r3e0Uxul4eYnVvbCR8QUy++Zb8ZKdgSZ2/Y/Ro6bLjNYhG98riscNJap88
MagOzDt85sEb19T/A5Pc1L9F9HprPLqG3y4kCOPimczQym2WRAVtX+6nfRyDDmeS
pF6niVLNutSBKaNbFx5oyGhCwJK26rgUhLcMel+EilfhxHxc0rgnryTfCiLRefzT
b5uazHFs6LAsIrnBupvtnYJ7QEjLI4paTNVGNr9tq3ld6HXTz4QSPwTyU5QA4rtq
PAdDWk9unpUSuWgx3tkB0PBOc393tXUbXS71T1CkmJH1W5bOx8A8aH3dTeVyo35H
hxCreGfMCTBWRrQUBLxkyHFqwUjqqVx1pF+OVTjMm3rMJ/55o8ySIr1tr7XbBwVJ
V0XS6JXFDu0Wq3qp//2o2ix5EEpxdnRPCE+jBkwN4/WK4CjC+MlZFOqBFwV8kkgs
E6nhe0NThpUvh3cvOzP/MXx/oqNCVwKyyzqCsiDqh0mZ3wS0qvhhEG8NFntuvC6c
GHcRbc2zeeEcTjH5EztStv9Ylgu1I9OiXNHqOtLI7XnUYme3FCx2a+wcfbWaIsy0
BT7a+d5TkGdLE4uBBw7DLlqT8+BEcwMtTqgSOL0/22CbSakbuHsptYM/MW0MZ3LD
SW7I1XdkRbXIFKTyrbJtftA19wjJQT3g21hTkuZOcHBY7p1iG+UUh8shw9/NB6y3
xb3XlgwQvDLnXHHqXnPBI/Z3pSWTWE/kCB39FxxxH2R+hJYVbvE0k1WazmctzN1u
lO3rB59I0NLSBm9zAUrgzDkMXECjcStcijqx/wH85IHwL8yNk/zJyEz684BzuqcM
/Mv7ASSJ7rvx32yM9oMJnsObB7Qp7y46VmGgI41u8NIdcaDhXLkpD3t0wHQtC8kU
CDjsrsAzZVQJJpccZH0IHzcJoZrxz/j+TR16CG8YnOQcCHG4hJDkV+VAchPs8a6Z
LzWuoyM3oSTsXLzCLEpHUfirHK3u5NV5TEL1x2OfOYEzNvf1PcaXvzQxWDtFGZWX
meHlBL63mKm6+d/C6R76phwQhQtGu5kenhcSpsBn7hFjYWeQXrzG4gTQRBYkT/1u
ES7k5GPlPSlXieZAI2vGjo+ZrzM1Bd7rHQzoV6O5QiS4KTzp5L3jHec+jfinq7tB
22IxPHCL3kEuPaJ+yNLmW2OoRNg3T9K/haOJznTaaRuypbmKm1x2sAR15smDveh4
B1PWWwK2eOCroZ6XjxKFPpaIDV+9rXDkyfT+OTOkYSH0LK0q8Ul7s/ft5KV6DAc1
B/bhWm0YUCIzEvXAPakm+xhAFudWzOST5+CH4/dST6EVwuby83hw5jZGoUZhXX4y
8+IoPHzgGdhNaKj8KzEGEjLujgtcfkXcALf973RtN4wjheMG5GEhgvi/Im6+7Zz4
vRFtdN2Md16WVERPoIpiUI4ykcyAghGJ4Zb5jddDCv6u7Gf6QQDHF2ByJbmoxogv
ReAFOYslLM7o9YoY13x5D66MH9ruj4ejhIg4wtx/Pr9S0D9X6TphPH31RKEMtXlF
Xmng4FDS3OZTnjJ105RoRCUADTSDmlRugUyItNzBwm62cKE9C2+PeXOrpmuIlrEs
1nNBpuePPuDq4o1zAV+MH0yuAmNgM+YpOZ5l44z+EFhUbLrRKPXUCJwbgWRhaXxm
4y7L5S1tYZrBoZQ4wavV+nzRXa9mni/HQZ6XbvefOpW3VXh+xXoL5SvtqVkFAn1F
BKW+169ns5fynr06McCGPe1yhBGRA3ToObzXWKqUG6LvQ+/cQaZwO+Ur/e/10ihl
v5aFeFTRxWYsi9HKNftLmvVQMAp/8i+EoUenqlElPjLTOX2/tyrWCBg/RtoBzVlV
ZbJ6x96p3IYTbG8NSb9nTlcjhFiH5mtVsA9SixoPGQKl9NvbwOVCT6ldKnjzXXnS
NKdW0n6hvHJcMOQCmcfVheCTbNb4A+yPss+t6yZ2VOVUj448zbXnO7lftAbXtg0w
RkeyaBskookdGG7Xz4/nNluFQpKFTupH10ROFlzHVYyOpSl+st4Da+Css5pLtDZ1
Frah162Vr2l8j5tFhwD51eDXu3mjbqmaxS0ZEq1yjF8BSMvFjdq9Vwek3wKIMcEP
BFea+wkMH7vlJuA4DnZFo9TTBFc01mhUPZ7KDglcYf55yKCVKkf/ZDT+ZEjZeoM6
ycH0xSLy0yYT7Sp6yej+D4E8Ja7sHszI0PXe7Rzcg+6sFSlIKAE52nrqF7KG+cNY
pTsuUo+12FpNSQG31Be/SeAkzBt+m00a875UdVmHlMAJK3eaigvnqWWKsvzYJi0r
luqBk+TxBT3U1PH4Jh1ADLYHvbkmvSmsMwWF0E/j58tCYprQPM4Vco/y+uZ+L/Ti
QGMGOyEAeMyp1Mozx3JLwL7x//ZdKYfNkcTVyx64yxZnw6asgqUIp5EaoPdlleWL
pE7oO4wm0B7OJN12GU4xrBJBx0JN00nlcMSce0poZ/ghaXZh9YNsLZ6oMtfQhvRu
Ta0pzA0otAH2Xo29oGpEmf7r8ZVmkgVbjq0Osrzrb8yv3UuQ/B4PgEm0bJYa5H+J
kp4fxNusuNs+KK+1Onuii3TQC+SSxS3JoQMKAShHPuIInCq8zK4xqXHMcCI3WwKG
8INQBMk6E0RJ2jWoZ/mE5brD2mRG+jIhaPTPvAHylTKl+FZoPxbhr7mii0q277Eq
gK/glm/kAdrJ8sY81qv4ITqOY6gEzhTbfsaMHqKns22lX7ix/3/UVo4dpt8GaMvp
MiPgOKxyA9Kir8dtJHP2mRGKra9deH8/n17ODQWV/kVMGrt2mpApXnzyYwmPLSdo
C+Ywa1JUs17mpvhO6hb6U6cUfxEJgVTkqun1S7NJwlwv9kpBGbsoBJWVEG5wa7Pt
OicwwjAkVb7fw8PSxDF+S0TFLItn/6ki5Ak0OpwX/gQjdoRrGP2c7gGkItcLXqam
Odp4PxbJIlglEhrEzb5Fyxk7aDUwEAFBsayqhO2c3sDIh1BUY7/a8EiPYAUgfRu3
ByP06wvoyY+zb7L4dqDrUYqy0Vn5ayt3gR97Q4YByjQW5EG3v93MJmmo8tqOKNv7
ku299GyrVaDp9kFLGZDygiU1mNZpOH6Zhxpsn87E72mLxpNOtbCdE8gu615Iv9iC
jMKqK0OEXxFOOBF1r/sZQ5CrRrkCoVBq1Z/Jm+xMYygWeRVNqTnczdZjFVTRqliQ
5LtMhG45cfDGfkVFVAO2Na9dFkNgmiOixjnLrO48aqzCrGpAAum+DMxir88e4z2Y
Hvc+igCpznTFxSrdbjaq/GFY7FSVtSSX2wgD8Fx9Ne7Ad+QTsgKm8sWNn+hWe1BB
FV+TAIS97ieYRY0pNw5RYXe5iKtBebNpoejB8oJszj4QVsnTywRqEag8E00RSECL
71scu7LoYjO7ZC491ZapTQN5aKepeWm2Q/08Ea1Nzkgd419kgwFokwh+nSFnubmB
+sUxzt6WbD3YdJ7k74trUko0tWX2z7qGpyyVcUFJ3+rzzN8qrW0N8z6QxE5JC0U0
YAo/VwCbBWnm3cud9G+68pUhRI6IRrUbpEioFPecFQkqXI1Srq6bkbD0mKtKpKL/
ah0G0/HB5nSTG2Iw6AQCvfbRLrtUdMm8V+mZ91UMMUdUrLk4YG+7vowWsGbhNFct
htrsalCugTP8SLUkxSqxKQZJWtZJ7pi5hiKsI4x/tVkC4UXRO84sqWf5eyA62KZN
yKB5Quo3cEcVqFNQ/KgaKxgFuZTazRRpQPpsShFxyO5G9Y/KdHAXwxZWEjMoBpku
Uuidb0Z449rZC5U3ZyeXn9rF5ldylUvkbZjqadhdPz48gASv0Cj/wO+zDSjggsIb
se5MXLT0nvxeHBVof5ic9V+ez9bRc0AvZwRYxwO/AJAYX6Yqbp2AOvPw4cGt4mxR
GRNyKBWXISuwnqVT9ulwtkk5R2cXXql+p1k8fPfdQRAnZQ/bSDJKL1H6g56ZWUTQ
ZartJ9dA3PY6G9N9NMKzlZ7KUjrGE1RscYxamX5nECiCY4n2zg+sHkkcZVycWaEO
F6cX+oDb7kXWhy7mvCTVYhRm3GO2Y/z7yooBbH+pAoD4FwJSVVqVMKSjz3In/cyl
bln4Ur1d9FEMxePMYBywFo/jYmKx2vdXjbgWGg/cr32sTtPVKPy2EgA9IabHRlYM
PYXb64ebO+wLlM5KnVPfEVxMfLgh1WdTfOHKwL3lWabUD0Bg101WIvWQRek3HjwM
Gg2ca+C+BU9g2Dh0RPdAG940/gfE4HlailetcoHgV/A0DbSmJHxuL44ZYu7nHKpT
aqgq6Pa8Lo3xeOqaHAajhggTVdQRYuL2yDhre23JcpctaY4aVAdZtqATNtyEzvCY
mKCpZClQW2symdzMmGY0ym2OXbEZR7jLvwm/GzTf6eElX29FvrrJxXC7lnTHOyfq
dDMH4KFpPvdQDp/H/yGDFcSl0q0eUG36ksc5LOwXTv2ccf02LF7gIQWcp+eWBgs4
9RcButgno8zNdUpI1gYpsQbXCiANfZxiofsjf0YjYbsOIX7c48sAAA9MvMsGfqyM
I9whUSEEkIeIss+/n17pJXU4U+WdaExUAds2HmSMfJFeB02F23m0bXTotgmBVyJU
kY4wqbDAbAt28xttKvaHva2d8AIwkf73IoCL/B2SFxk3R0qX6TwENyUHFg/StoNS
98QrwlDRjCTF6YX1BEl6tNnLycZlnH8iBhvpSnybETyrJlZ7ITu2USUeVIWd6JZi
IMyYqohb1p0aNNe+5fU+r/nIR0x9UImabhUcmCuBKHR04dWumRIKvgrHjyzskd/5
VHqvqe1MmEGdLjhCjmcx/PmhqrnRMQSRHeCID8MbVEEBEjLR5EJxWB3vPftnNZ5c
4ffNEwOV/mH7TFPWPpQfhMBINsOHsWMEmV31xGkB4Jwob5Mhfd/UztynU+FPKUNx
DDwHeduwTLULaVx0arqsZpQ1IWjT+jrpysi91QIUa1j6v7rnYkL1FIcXyVXvmYBw
yVF1ja7REWGW76VByVddkwNKExICS9ZQCisjAys6AzqA8KFj+q18qC0v3BuVP5C9
3A+rJPAv719zSNFH+VEtRT8E1MGR1evPAowUyJpbShY1TqeZDFtZcOoJru35YDer
DYxtgSXeJt1R4TuandA/ll3x3YYMNh+zXrzMFVsj5fA/ii+ChFPNFb+ZymUHzVoa
YDrJJxS+L0iV0QEVfWRK1+7j8eNwX1/9tK3h1RVPnGiQ5CaWWy1LHKwM9DrqUvlr
EpXM8ONcGryqA7Ced49rayAeMqdsRofiB8jBazoZkZQIaeXvxc+Aa4BQ5SN3afmw
JYFCpcHYd8cZj+lzr+oTQhC7eD2oTQx8XTQONzy3xNb5BnCJzU9XW0GZxKUeqGL0
vOAgIBxjPX25n9ab/wEJxoy5EzBaqFKvR+aPDR7l0zz21wEydv/GhSqOOwoZdgcE
xbwRHqLBWiJQn+lIZhiSWH+jXdYSmDjVEydt2l9CaLOvTEvhgvElLsIghmD4ZhaS
NHCsJL4pJdsbLxQUgbnPHwHWEa8tfM26Rvl6htXIWqLpgzVqYdrDsnr91JzFR5Cj
BY32R5qc5pSOtedijzMOB3UraqoP4l9Iv8GZL3m+JGDoaAnf0+LFmVyW3neJK1F7
o3efmtL776NHM1L9Itfa99MWG6xKlUAFeJ3gbFjSaXkLIF/UndRdOiuYhQ8xpjhR
Y3rzPerh/YqMQA2xKd9N2gr1+U8YrP5wStimiDHyEicvCo5TSqi6qwz3sukaTHar
jz05082tISb2wujatUCK63c0NknAslbUxEeVkO/7CKuYC3Wc1UNbAhWVRR3Jsusu
Aoe2vO7UCoRdDYwQNSTuGNy9tO/93nglK+lZAILH+2oAsZ8A/cw/Z3ywAxH7j+st
tRCHqoHAeQ8qd9JJMyY7h4MgyISU51fZ/736fqJH9yQlttVS6DINO4CwfGmyDiLc
+ETn17RPGPX5Z9/4Jo58zJ6RGNquOwTebBqxl1CXJS2xWht7IJqfzBaFCr3wDpa5
5nxa3u7gh4zt3eUx9eS31SlI+cfL17InRI2RdJitd0zn3CeiAiSx76DxH929xS68
sf7s1+isL3bupdGqAMO7m0xJWorGVDc3to7Cf/0oZAiKVQJIEZ7tmcCI+urlSxs8
ywM78JY1S3/C1DPoTp/FJx2sPW0xMClgdX0QCFT5A7a2IP77wohsA8NsPjcF8PCr
e+pcTOXEYb4ur7hExpm3yUoyQUZo3c0t6OkoV1kuqcm8pMir8v6IQ0LwPwFjKPud
3uouh2Yb8IdhBF/1tutHQmndtg5pPqByzfvj91oG6JUjuPsmVg/BxY7xn8TxSVkL
BOoFphsyaAupq/ymzu90wOEFK/SKAhrph+8amiD1sn2JQGMmzWhO7QipOhqQxhvw
EO79R/ZyXxWtEpjv+unRjG4Ox3VZR9WWG62tzjLT4JAxstnWebFs4H33gmtxuPlF
FUMqnRx1w1hO6zWazPd63wZPjwMQi7dYlPVc7FPjaH94QrIsq1Ix4LlknYbDYE4O
nxMHHhvVjfYBPb0iKBa5X7IUGxev5OjriTRe5+4ONVtkld0Yhdc9XyosVPCWAku3
4Qx9mIg5hUXFIACn6nW0O9adZmbN89wR/ObTQuHwFezNdt0Dmtyp3pqZV0t+2DRX
Vlpp31r/vmPq9onQbW6ho9/n6OpTLc3e+AdrpfjEdJf+vnQx0sB62/RZtdAzrNqE
FYV0mthTash435xpnaOpshOdrKaRR7612mCLJ8E1I7/hsaNsux0tYMdBRSX9AZLW
M+S5IfXKfMEpYds8dnG3BzbYh4cY7dUPFkgIoeu4+LFSNOEqMNXcFc+nxNyqyAJI
fsLPBmWBY3MDkKyziW0sZEvH2VpaNRnhX3Wl4lJx62HicY0tyLE6Mn6Jqgd3M5Ss
RrpgQYkbhfojTAO4wksS9pE6LFyPt7CfiK3WNU9iN96dNrmOh9t8ya/ugCaNGRsh
GK3fhroCfYqBt0ZUwDsjEIsMxt1p+DgR95DNw0TR0gTlD3ULDJQzbP+X9i4Wi/sI
aKowmxOli4PvVumCS2htk3Xr66xn3385alCIwdIGYn1gqLK+CVSGjsmmadDb3tjA
mWCqvcaNjZGnQ+v5ZKkk8+8gWWcG4TfgHkPAMeAHevBUS0Udi45vUPn7r4RKTqA8
WXwa2hCkdXYdMF/WogRZWoHH+2qwC2F7lkXPlMBfXGt6pxfJxTBlzUJO7gIXDQuX
VspOBDPsvWfQcZZRB0L8MONeIeSZi8YkbdrQqFAkOHMCTwfWWLOcq1MyK+b4Iyr2
bLMRSY+tErT8F0GiPxovYMS4xIBCb48OBMaXTIRK/QkaKwm+kAXDJ+E3xbTrkQev
MCguhNFYHy4KqEjVyWfPZHcar49DGIqUXadE5aYboajai8hIG7h8PbK1iligFAK+
aX8W+ktWDDJJyy0b5DfR8w1BdOIRfMPI9Ges+Jyuw9sskqTZbXaAIYyACnbdzIO5
Gqv8EK94ZlTwrA+fRtDE+OIjrowN85ey4oPQLBfcy0rrY/CIvKKPE6ZbPjxWybO/
TujrWip1q0PW2tffiHPSguFvdKLMIqGeNYjWvMwGYDTm88XBbz5PpPhraThZ/bZ1
y6ezQmnL4YvkpIwlAM2ih15X3zn5gmtaix5yZBGvx7KaLi+qQYMZ+4dSJRlJyHW6
DAgZqOn7Ivv3LKVUuvS1ne5YE5b3iCpHbLduxSsAgGThGbztgAhrmYU/F+BnU1X8
Jcj6GmXYaj+Sk5sXzYf/anWl2xjW9WOWUjjDV6onLvJecg036BpZDn5/X29Ay3EO
VJB8X+BB6Um7R570/1nwKbuRXF2+69qzwJcGIJLf0Nf+962I4fC/uORvhdMZdAjJ
qfPRiCUZbFrh8ghj38fMNGfMKKflHqiB1sHBXy1avYxxyOF0iv1B9nGUK8Ues06L
3szNINx1bfEujKgmlgvz1JUMD75pQBITNc5vwUoVvFlIDV0ZCn/394u7zug1okVR
av8eoE6K0FkAUCDuGaI8QT0nGbEGLE1MbZe0JdTUuFxiD2UBS6qvkiMEXARMcWpY
DBYapTCAHZ4yMQsIuatC1ATcD6EL0lK94JvNVJezl9ohxizkzHP4UdyEDuTMQfNY
FHtmg3JDgJMqUHxUrhlO8O14Q7+oxhmctyfFC4c0kbeSzimqwEdgc/7Ro/enOU8t
QLd4x0jryjH6XR2/tolN5i52Gk62XjjERV2kqor2di1slIHMMsAdkEDEIO1mcX3W
cM5K0rzlbLPWMGFohtqqKNfBefI1qTi464gNbswAijMcRcOk/YPKwbbMxtGZnhQ4
jWP7kSz6Fwj0FsDf8oDwGdA4IF9b8rEWvt0vPjwn0X3Va++hw7QIKzYwGUDb1+Jq
eyDC0mx+DIoIBhMEXsCcAmhxPiVtyRssTbI4RjzkUD0UwM3rRPfr7gfaQ026Hfik
nMpTPpGyS8cUCTIbhmTFb2TF6HwGK6fu2QAEOzri4nWBUEnedO4Pk9CAqtpjt8Rp
kpVPliJsZWdQ/Itc5rFSZFLmDmWuG7DnwRGnMu4463dOu418hDVctS6TfqJRrW4v
I9CFhql3lwsNvzYAQ2TK9Kc9MG6Cw/z0ATwsa7fvR3AJm4KmzvzxeL8av53P/OH/
Dz4qOfYEELyDJr2/hlc8NFwO8CkZ1EgIBj0kG/3y6e43+AVc1ymuSULjICFb5jil
TFpf2Bye3mcUDz6KRC7iX2RjGnOjdSJ4OMW2ZHMwMu2yh6iRrkoFVI4tCKBj/Gkm
p1eQUTni5jZdjXH7vJV59dpmr3SAPgu5WAIhMqbePRZ5BxGXrPhb4aSq+lbLJugl
+0zxocuL6zXIyU+n20NN2GOh4wANd9dJtFpu3q0oaHf/dpRgiwqBTca6o1f+ptx1
AD8sPv6Yx77Hwo5jz7JID1FAo/dBmAKzo82TWVu5pEVcyAzDXXbidMSFOo8E6dno
gxwPlGkDNjMpT1F0t519C6B9QFcZT/r8qvgJwhVx+hkFOHSFcT7LE+Pqw2aqrXu1
3z81gqqkIjk+ID3uKknSNfotzWwqVLSi+j2boXDDT7G36Vs6OoxYWJVao5+Ihj9i
9QiMlSWZ04o+/qGZohvstrcP38Ykv+IWSsg4vlhTJGzo5CGoMdaZXNKl/eIj/TZ0
6PQPvhfEYu9pn+W/SnY7J55iQBPfvIFLWlF1xteSWum5DL0UCCq0vudQ/Lmz3Xdr
ufBZR8iRouIK7VQEUwTEmUc+eJjr629XxNxHLJqzsXmzzdqHmulM+02obi1f7kYI
ntmMShzSagrNRwOJztAkaetPSWOJ5hH6RaaKwUH8tO11kKJXqsyoalq7yUMozKDd
VtnQ8bK5DD3qcnb8Wh0/bbd+pHi3QmPxRGDe3eFPvja7+R7Q4FKIshgggZsayQq7
Q7g917QzFfEEdZE79ptDu+R5R4Q658Wi+U178DOQHV35UmSQHh84VUXh0G9s7jy5
5LivB09oIzj6Z7ztsuGzy4FZcd/u8VPAjM5nxmGcrGYN9Mi+B/941H04rWh9yHHV
7VotPHzgps03Q4YdUAE5k/hY5k1//VcROJEHJBDgZmJ8fILtyBQ+oMpdi1FqqU4d
Q0/tC1AHSL3f7Q+PWux+zWYmbenSjhwkCPrh8R+Df3sd4zqUd+nT2lVHRzpo3X+h
RX0d0ci3T/ONbzJ3Y4MLy16ue4xNeB5ui50yrBn4IDT8Z1k6s+4cbqJ2z0k0qhtF
Wr+7ekZWeDfi0wbFQ9tqlQe0xqAp0aseKDbRjPW4mIPPARERwQH6MsuzIDIEM9tG
+yznk1NIIUV+LFzZvo/3U/sWaCzXWw7GkVgUzjg9dNl7lANQi8Ovt+z1x4B52gzJ
24zO/cKv+PHA9OwSC7yjF76xZk6NxFlUsaomkeqnU2rcd+jXTQ8EYxWaX6rXT5aV
AS97Xt+qEtjUs7t5nvrsQoJz0OkluNKKDli5VbyjaYJPMG7+iOh5XQQ7Uyysk1dj
nxImoGdBnWpfu9w1IdSN5zeFP+Z8ZlH8IpUCm0KtSjvaJP8ooIvDTDliFWKS64YG
SWyBYwWVVNPHvIv0e/H0JP6yQnaTiV9jDxwueVWQWI8v0ow7nyQshT8Hkba/LumJ
k2pVjG0Po+oQfILBVTi/RCMG02cYbT6+FiqgK5xGLF86OGbSNoWdNwnWnYTD3R5+
1dy3HvuXItqCH7gKHDTQoJKiSxbG7K/d7UBQjiuNP3fARRt/D3R0jB6jv9lP/ltT
xokSXL3tHuVttd5fBYo/b570o/HJQpW7snX8QtUDPBlA/9gNZYKkj7KbCHRZrOmf
Qiyh5GRHL3zmw6qrUMTVd1nOvtbxOUBiSlYjk0u7iyvhHyS8I5H0wx8s46hdKDVg
ypuxIdOsWQtO4QIUk9IWA/FmlrX+iUQoMKI5X+dt7FpiDhEo6LPcAKuHjKSNlWd8
+ohVOSn523QZ4DyxxO0WNM7iAdVc9En3LRX5XFaD3yjAhmGWW2S0ioVIyjMWTskI
oRtsTXxsr97DhtDL1qYGPpfdBH5fRdF0KM0mLMywfDN68uLbyvLJPNxdLE03pKr0
tOZ11KOUpMFjLGkBf8updJ63bhu0mqBOdAdfSF92L5ZXjYe+j6G2UjIogMfrLskv
q/Pgy4vVPvNg5PZTTBl77Fbb2u5oNGe59Jh36a2vR/csmPK9SWJjPXUD5EJ7jfsu
pwwoQjcOOzQX0W0fRry34o31uBlJw+lWyiY7dNVn2RfWGDZhx6JzfPqhFvtqcAVt
MypmwPLrAGNG5zcFZloz1nRLcXcSf9VrNMRPTZOc0GJIzUNTnUjPqYN9OA9d6Kw1
JSo10MlkstRfmNHltirOOoqvWo6mPU8dfNgX3ND2zIjFfNmki5VLu7J/9WayFBFw
KffEVOdpsORAx5e9hVAKBJMthHBb33IejLciVFyb4CB8YIolnvPVaMCCqYH9zmO9
4qq9K7bxzT25VTfeOngaNsEkSoIaLPRsN0ElKSeW7uR4AzerPg2YF7Piw5E9P5hi
uQ/LN8TWbqjHQFuq50F3wSAJWyiybZvLAghwhmNAgHWRrJ2T4gd/bswVgLucAGBE
0qyv0Jm69uXzXwn8BQ4eVB24DuIW8OkPrvRiCYrexfykyBi8poJvIfVEfRmb5tcU
BIy+g9vFyTYtMa/IJf2mFLMIBU4tuXlyWP6Iqn2zTWxRsIX/kBhR2rH/LjqCPLU/
tOk6fzsjYP6l+3B39FDUAvNyaCEzKNyHcnFRrpKMz7Z6KJdtE+deOaJeF6zq2kjL
FXAcVFfQIRpAdtnZm0kPuylvM1SzpcifnAvh1dDrLlU4jjnKa2TGLxt+SmD439rA
2cf5ABKIr2vpx7yp0eMS1GckNlDxBzYSQfl38TKbBCWUug/s7x5FtBz3Fnhhvex6
+YFtzawIS7UHlZ1Cv7WiLWQqN8W+DK4MFY1qiVu6C2GqepxOb6wPbRdMkMBMwwSo
anWdFNeF//5h19GIgDjBgTcJqsR1U+R5VqoiNNKkS0hvlNP8iJkKJ58ogkyMV2gd
jkGDPdHr6HaorwPFNRHbk1crsU/lQttPte6DiMCIHMqCXvzJGq0kgIUYjcgUmzWN
HbdQhoiwMW6YSFUTEmrZN/wEVgc6rJHtej/654LIRl2JRakC+tpsVZjajJC0mHyV
mtsYiMk3UspKczrfLEs69JMqyArpXMv+/w62meoJS/xLOJqcXg0p9yU5Oxr/lo6r
uQHfUcUO4g/fqh/KI9ls6lHMKBCKiOGyTAdBNcRVFd/w55zvBrRnKopqkQnOMPYY
AwkJajnVZk79N7qx5kFA8AYxi4UZy8nyGz108KvzXilObZB0rJpLw3735FmqnLb/
o/J2LTnydbxPGQDfvAGu0x7eV7yttVkSmQesdfv8q9U4cGk8XqaEMmSNqXVUJi7L
mCN078rOpMyAR/irORviuxRUSJXHceostJ2zApk4aMfDNHQ0k+NufvJbdCYfmU5H
GQ9COdbcWU8qux0ihNP4IjqBHjDq1ppMc5gQJw8p1iNku7ID+vhe7HrHwKP60UAe
nMRQrTUarhvk6l5RdczxdfHGZK8FBNvupNDN++rbuZZSLw2WsiUZDplZH+ASdy5+
yZ+Rn8Pc8ZnoJwJbwcgWug3nTv+b2IN3vb95U+pEEVoZnG7b/K6IMevuOY1Vwixl
mhGTU6jjtQbp4ihgl9MZhZjwFD+pJzl+Gaj7mMunEHshxwUohcyYeEw3K+3Cu3M5
ZRFnqdu/loGhVSg8sWE07kNGeLEiw1gbuCIMTU+FlXzmL6JsDRk0LsAsn9NwrLkv
NEiST3py+Bfl6xV3MyMYd0ezlVhFhqowC2CGekPgx8S3mJF6Jb9aofkgRxkknzV6
g3n9LZeelmygW+jdhRabZb6xaCaO+giHwB4AQvlat+yG6vc0G0bQxcpPRTakyTI0
SR7bHRXBPld4vMBH7FaCgNP+pHwIjs3SSR7LV/PJeBrsmVIy+3Zyu3R6B04wNqYR
zgUw4iprOQXfu3QUYgGB4UGzmBzhI46FIKjrhKppfvtD3wxar5NXXAGYFbK1BvNb
h4qNUrpxTAbcOTMRZFZ4sDgYs6dyWfT8dtxwlyzF8LpGzsnnp8M2K+nK4dtkJwK1
4/Qggh06FdyOBjwOu0BSBPIL5fAhNAosGP4hXcA23q2IYrtrWsm7x4uxRxkVUNu3
jmRbP91N4JY84o6sqq3UcfrSMhBH1X6USAjCCEgVOpWhsfFALvKn8zsGxowC+l2L
TTx91rBRwpqG0xU1pkRLCNe3tHsLq3fA/q4sXUPnlphIw0bhy++rxiYZQi7pJRqh
HY7Wc0fhCIA1WxbgnumRuMFRi5KqPOU17Lq7wIpDWhzmOlpCE76ueSMjd4DUwjLP
EyUKfsbZtxuyz+4sqCECT+a+qxbQl204SpnxDb9qGQzQqSpj9uyAADELjkx4XyL/
QiJpYwjNDwrDUgyOG8hSYECDi8GLXOOWmJUkMS8eTh7v440kWdRvQG6b7tqgdGFW
A9VilDUuAqK1X9qf57rMUFfYy9L1ag1R+s1w6ylAQuXMYuj993dXinzZ2j7j/wew
4GBK7PlGjqpkwXI5GzNu5k8H3lEjULn8kR6pKyUN7mFcYePHZeCpDrXsg13PSvby
vAwDm/S/M9gjgqsD0+VOAe6ZMGStfyoTg7uaZdK4AVrN5KQ4seYzeUgu5XgxmV3j
o5tcDuIooQV/ISBCMwk3pqekp6r45LofXlsTCQYru+iyKAtvPBBVzyqiPkkeub3y
HiHaCeUt0Xk3D4bGz/swsh8laSsSlOKnpo8MQ653/9nm2eAA5bT6KmUiaqL3gm4Z
0yogbWcOshpayxCPLila/exXRzy1p3ulSdHFuy+SfpnmhVp2F5JA5OfyZbV3nwD8
smv/X9n1w6A/fcWNGUO9Xh5/MlGe/0LXBDD+X/l+uG2GfDShSlE4pAsaimbQymV1
LWLt+ViK9oLwBg4g2+yReR23H20WuoLEHHqU3qufPuanacUtgbi7mqES83Ari2iH
it5VXG/rVmI7U/s9QdsB+AvBFGSuwT2wutXJmPnB2H8+C6OKly1NDYwXIlsd+j/G
X+K78G0h7IhIQtIrg4HnAgCfOsymgPRrBMq+F8bRhb3dmHoX/Vo4KsNn1OdKNU81
0pIvLQZDf23dcdHUjzEoji3u1xyRYcMZVZi9H6vJ+tCtVC4j9JVaI//BdAiPbjW1
PyBOZbc6kseaF72hRil+Mkh/izq8b/2ZjplBHjQ39bYQvNxi1SG7yIVY9XpLr/HD
hyUtA3XN8r0gYDwTXMp13jeOXf4t59+SDYxZvuUCjn/rbnVMNjaklNlSPw1fy+eV
JcSNEBR1b9L7jul4Ythp+UbnTr5oUNdNtygDZauCx9IIq7Vlo5mPtFYiwFxhd4kQ
tE9+3iOsO/23n5RT8cRz2+5bLHAWZ11dWXvb/4CKDCLiZ4DNPrq2psGJCj3GPjsI
fk9Qa2RTP08spzfbwIjcd6MK+6jwyfnsoxB7cYHzu6sM74yJ7UqNqnqeRBAHU1bm
TFXZ8DZ/+0NoPmO6XSop853MCRmCDAGpTFFTnbChvjI0IWpNYIbgHd3bjRea76k6
vne5dCNTsB2NTL4BZ2SLWcjMjqkrZnKvTY4P8aQlTOc8s51YPlh/kZ3xI+G5KgoB
40d44RVVBZF3z5sBYJRjMs40R4nLwRnV8RDQrShi9HiMcmW6NHcfJ5Xzt8LJPN6z
16ppKUhl4BvLhkZwHyTWDyWtIj0hQtIpKWKgcObn5eE+QnAm21A9/zxkpEOu4whJ
qRYJ6V4QaBzM8rLa3Qfiipii9fVTaBk+OvnD2hRmZYYZjSm21BhsvxS3+xtzNtaw
DUghnjXsuCaQzXbcAGY+MqLUGm6vf2lj0z0vt/QhF4mKRrjdd6TdS+3useKWccv5
+dXe6DG3Eqldaegr9X26FsQqP2cPzAqIv4S3YrWJlllsQhShxPT2eqHtWP5uplMp
Y3cae3RSa09No0c4J7gI0tI6K6S1h1JnMhnzynZDtO28Ow6Mj7iWb98D5OLp9/Hn
9xuGryNQSUtt855pKIjpM+Z1rSNY1Afsi1VwqD5/wjyAxIPZd8fZ6qO4J9VJ0hfx
y5crRyOqDnKrVKWmwpHSpiBmD4/mq/seYz3iyrdz5vVoF1+gLu0DLL7ATSclW2B4
k3Pdu/1m0Zh285ZnBlxXuBo7dZwRpu4Saioc4pR3DPvZRkkysBKEdYcE5EwqBAOA
zOdwubHeEfGIO5EfxoeljKE6pxQBHIlu2XrW5BCwWvqPnt5jae2zaBha0mMPiVdK
WCiym0TcLuTAsRJGt8H1mErZMi0ZXH5uMAI1XHrPlA5KCIECpA1S+N2Z0JAwsJuY
lTZQ7P3nvr71i5wukLYnBiSd7m6BnWMnbLgzTTmBs4GjTUim6jHBN9EdTL5qbfZO
rpr9SgjIulmQMId/8QhQrJbaVAD2UTNMsf7m5iZc+L+Efl98MGdK8Hhb4g3QiR/g
+tfP4aZkLuj6og8dOVzDoJhUNcUE7ZKs4Vyfb5l0D5TmGLOYtP7Gxa9Z64bhTxOn
JWt2tUxoZgfJp8Ooq7zHHH9qqTY7a19klC2hLSW8FgqKgB0ArkCQj3rpGe8+t5IE
OG2jM8+Ehkae/pXlcRVZQQI5Ly5ZzLZuYCxZyNJNh4hH5hKUlpeopKByEJv/C1z3
Sygv1wPAI0DqrSDwFbvbEZjKtvvwf+YAcrmdpjhEmMawndpdGlTnpYkrYd8/kOsd
bHbuzl/UFhmvQJrMcs4mAuqc+OMwvShEup21xynTugukKSVy5fpVfB65+mU6vDDs
pHorZ2qFHL1adBU3UVXwYEBS4LEyItdj9GbnRm/CeoSCoaLmdsX2Tu/Oa0HSAteq
XM07n7KwAnfsqQSleIkpS4JxhbUomNkAOcWUXMQsh5zt7a+CangJje/hFMUtuZo9
YDE4uUGkX6paauzr4mpzSt8hxjPRjAD8Jms+mG79PG7RkZpR30V6wvjNcc3hxuTk
yl/cxkBc+EfEbpi038T+N1Enkbj87/kbQxwcKT56QTzuXkMRAR4jLy0FAYaCEdXt
kL4uhC36Tnq85vNgDWsTk8s2A8gQee41GuUbO986d9Tw6gMqlozVYfLTUHZdojWY
ogBIaMeyELX2qDjOOPPIaUbY2GqdpeBy0K9fgIlqNqj8AuKwtQp8nyplJx7/thlO
AFZxgqlgPNP7XdZQBcZ841aHrfCZEEMrl31jSS6e5COc7QeJjYFBTDpu4LMRDBzS
V7OpwiDkAs8xBqedyIzOTYtThp47tQy8M0t9+vva5q0E/UVg7NuehEDOrc1huA6g
ZHJAKDTLcy2aF4EARIeGphbykmAzhJRlcjmhlnDip35kb9QgvqGRgEmCMGI4s66s
6RgKuKTDHYmqrwVcAKqLppBBidK2wQHjEbE+4p8y4S4yhEuKUrU0MAAv1uiWbR7I
8BG3wUs1YGuPGs8ue+IOkZLxuvjC/KbPm8t1PgEt4v6DoHf+MsPkM1P2v+L4JBlu
yW7UIylpaY/L8xfMxazj7inGAgTh3j4U/pH3AN/kXpFiolAFdocfzP0qo/Pq1s/3
sQeeaTnvdNcWb6uURJE61IH/I03AsZPS+rUNpmymVRLK8WMPkz6LddcN/IHHAdH/
k+QhhlJZn5HK70GjKtqV/biwZsKZgfyw59VOhrVOIRhQWfA4rZ07BfWQy9CVSDd/
VcRUJNenprwFSqIfiO3/x9tl6lybxzya4L3JiA/jXR0s2HqWP+CtvV6tRf3PJBeS
TOJrLngujcSbLjpJjmLjuBdoGyLPrZYZ4XM3u/pVktRzSgBj/h1rrgZFk/YiAOAf
RTL+Zlh3Hwp+YjgRr/w3okAGstHX2btpbIhhW68CxWdUTfCWGzKrMrdJ3VOuz8G0
HovsFp4q0zYYtAhZbZHzXEHPMV1L+1GW3ssRZcpEMDJz1JL+nIJP2w6mDi4fWrwj
ClHPt49cKBO1SkZQmgbWkqic0Ui14yYgomSkkZDsxlu25mH9ZYVI1sfhpPVPVKvS
B+qmnn3whwfUkTpKZZ/sZTUJx9P8Ur3YHbS7uACENMO9B/L51sVBrotir2qjp0XJ
xoHvL9A2skGdoqtCCdvlaqn8sR2e2zd1dDnS9xtwEiK8xEtvCdyo3JQm8dh6YKxE
yykeHAs2mug/Mcx0LOzd7jE6NTQ7iLRM4//2CDyx6FpXsjChDQf0OYJr0UfCCk0T
eyyHEOvCmaIaL9XnBLKGAXucWF5eeOMKwzbOELDW6a4xjJIxA1du3bycQWf67gdy
kWovJbRtZkkaAYZ6zipy7ENQMCXqgN97uwu+b35e8bRp5PuS5XE2J5Zi7De+eu/I
VcmWk+qnEq62/xN3wk9bUTvYD+F1ed2xhdGeXccF+QlJOp36qr9Nl291QjBS67xF
kAaTEr5/RQl7k6BCpBiIhSFBbMmME5iDjI5kiYdKXfk7lct9qY0ODA6f7f02rcV0
pkfRYSYB85pub70flhVlJwLBB96sfKldOFoZPcBz9TchFZmfukecycrBSGbRt322
Rh54tNNv5UYKfHWUdMmArDqqS410cpn1ZfD4566VPMY8JuncASlUDxHu5jOB3Bgh
NZkLbPHSmPlj8H1slkaA8DLgzQEAD1YaEXtlTA6kUC174t/ntFTeTQ3adfKnFuWH
lv0HxdJEMcqwwlreN3rPgV5m320FgnZpWLoxWkVwcfhUMnRRrKh70wJmVhXMQdBE
fZhaNUX/LleHsQ5oPz+kxuc2/tVrHfiEiM7CaUz3DntbmZ+EEkWHIbcgXvsXhzIR
H+XpmJ6OuItm5bvJeX+Lbb3PnEaKc9zIgbumcaAYbmkB3SHcYwtjStHrETssF/e5
pAxs62npMJWupIuU7IugUZYJoL3lINnQtjtKTXTsFOkZwF/mqRQc4LGBWpf4fNk8
qKfO23q5pzJZPun/RP2tGIhBcefnjQ7amPoVDH/SP4Eaf4YONljRkiR3NAOpwXFi
7cGwyIgdix54Vjw/X8cJyTkTNLuvEvPRV/Qolb/6uVfN0D6yel4d7jbnpJoEYnTH
IlqkzjSlGehfh1lzvBojeaPgRbFQHyMRGCoVq374Q2xSKOKPigWowdYDpVS5zve5
m+CiwD0InZ/ilCl/2/SEmkO6MjMZf9VtrXJ7Xt3E+qVt3eof3yhkVgpEgVkRyaYI
T5qkNsh57QsNceCAE3qyiM0OhYARysJalQibKnDNddSke0+A9FarY5WJtf9G8oMC
PlgoyJdZMQO081tOsEsSIL9nz8/BzhiRa1WHiMrLZzkzg8j+JUmQaPbQkkzA+aHl
DQFtQg3mtGkwbXMwiV1VcxkVvKP7UR7MGFL6HZyQDPxvEy5W2pWbMWmiioLuPanm
25wtLEmavcbMirpTSfSyAS/e7QJOR5d8e+vYeMAiZEeyseoujXG6tRGoTLy1jKwI
KnCW9P5CgSrSpCtuc5xoNiddAJqfny+wyxqkH0RpLsRfQat1x92u6YD4n/hCk8wm
d2nAZAh91We0PFnLkrsVrQ/bHxhdCjDJAKmXSxML/5T6C5zASTsBfLOy0EpX4sXY
cQUOnrunaMIyHwTj3xTNk5lAcONxIPFNVnbZYjWD9rT5tODj7lfmJiPjUvIpYVU4
NYI5BRtyGz35T+9Mk9ParIHGvHDSdeJF4Xe6LfwVT+lb4D8ZzdKZ/n7juZrfGbnn
4IInz0lgmM8Xx4Olg0KS3tLfUA3FO/bQKQPo0lgLng8BCclWQNd7T260xovu3p15
Qr54DG6Q4RUgm4H0utv6F3iXAU64zEwDGRvdFN24qZ+mG4fsQuJslGTaZpqCY8qF
fOvxCjChMUd4CYiWI6wdheypkDa2+3DNMRmFkJ4LYit2BB2/G50uWbMxYhm6aBSe
h4SOLPUxV8LqI2kyL43ZZpGZFDhIz8qqix1cpATRxUZpSX6DfVe7acI4oTR4R4hj
zHJfiUSWbqemP39TTpX9VFYepRNwyo3FTb7avr/e9izjOMHmq4BpfuXR3pgiNzxe
RWIQsfq7alaqz8rZSXFGSxUtVAktr3lvFEt3g1aOYcoCJefEbP9ZiS7KpOMeK5yn
I+oZgUvu9wD8Rm9867ewKXt56FWTmELgBFKIcwvKjVjJvsPZVseXQQixYA8h0wYm
8U42QAZNY7qJMJQm+jU4fzOKdbjmCvM1dZ2FvnpmY3VjuCPVuVdglwjJbXZB6sDF
K1KmnMVP3GVyLTKvBqSBA+g//l2qRTmUCbADiPtVuLO8q1B2eUKcjXWM8rW/dXlG
phENJuNSuZZdQHrEnpr6hh/JrAS6u+XRPXWeXt4iBEDm/3ktyfPeJTI9E/6399HP
2qKHKgluKiHlaKC1xHQE0gmN24Xuc4s4/W7ndMV2M1d4suYq//0ewUzkGR+54lR0
GS3Aviyfi1E3S1YezUqm7HIMuxrHkAOs7+MQf/CqxNMf0knUMNS62TunwJSBuojB
sXDTnY0DcsP7V686fqjsmPmvwDaJ3j1lS5VQ74mBWkk0Ixt0ybDDp/XKrI0Ow0v5
RjuaYZXdBCljZVjSd/CcjdVwoG7rPt4+pRycM3/9u1Jxvjorn8JDK7kFC1GlMW7A
zDGoU4amY+pNZ1CQNfYiD4YiJJD9mqeV08GP+jy+6qVChFkJNlQ8HYIN0ltEWW7l
q/oVxh//3rhK4eP6UqzzLmt6pVVUdeVshX/v0nwI1oatrd1DUvphJUrIo/TMErqa
hHaHK70hWoyjjCDiTNYyN01AEuHHZARJH7b89DmcC/8ys0XVTT2Xi4FskOsNnUZB
z4D6cZHchK7iVi1lvWGK69xYvtyMiO2jGDnLgvHem7Y+8MpivAgJ8aWkJKZzZyeI
lDrScrmNYAJvqQnMXbunhvKGqQUVWeG/KH0IN8ECAI6cxnm5WkLyU6jKL32tVlUm
lFv57h3xVRpz77SGoIhEWFtL1cfcBnDKVYhP1lw8i8IXsjTKZY/nugyG9h7F4zPh
PMhu/dQCdF1k/EGKi6YG5RA7h+k6YfYuhj9t+fmrBvsPhVM6LB7+OvfuSomzIEM0
H9Oy3IONNaEXX/g66haWiEqzvvXWJ2qyxzCoSV17uUq+d+jJX3NWTW3vT8RhufJ3
9SlHRYo6IugQKekN87S8jIKtq7fp9SuXAqvytUAbypR/8m0bIXMXdMt9l5MivVQk
RF/UEY4LObSzmDusvli89LtFvpRkwGXReX65wY1U6YG3GhFrfQDzpZdtRHXjf4jk
1ZYQizgMmbaeF1+Ce88aan0EjHDnKsvm4hv8WYZY+ovEO03ORyWzpoWUytN4PFcn
h9hnNoeG2ZtCWGvdQ/YhttS9E1asQJFJPUNS7JbEBInKsahVWSVN+g68BKX/CK7U
XYA0Ews5HaMY6qEXtLYuQhbzcg54330U3VxEhR25h1UdhQD+X397mk8Q+L9FhMhQ
MRYYrZHPHTrBJUY+k1KqZBRQhKzpC23E3PHgYjeGMGHBQtnGnvRRiW1EGJJG3g0v
TOU9baldz7LY7X0pW7uMNnTSgfqOw6bFabD3i+e/SFADOe04Xs5wNZWSFYVNSlME
iqW9T0VnpYqjhuoqwSJQlPZBhq3ILnmIUqJ541YdPpsywCvL/aGvCm3JnfQDxV3c
paTjaT/D+HGA+GdMl5WWpM7JH6d6rVmAByf4IlKYP0Okmc6bTg2Oxor31z+uAL+t
vgbeS6Tfq8MLah5bnwqlLTb9xr/dySsLDFX0bCNVOfCjwim52toWfamfOg3qN/vO
nR23UPeHg+khiA5aeJ0n5F5C8HC8wRXCXzZVIagcVz7smotZcQRZR3eqQ7AtWdFr
y8QwADlNHb6VrzUhDVGEd+sZG2amB577L+J8G/ao/spSs8bYYB9p/DmNePQWXKjX
EOjoaSBoAk9pefQHTOxd77NLecTC5m8mkLs63v9lqOSbUGcd1f0GFzPj6m4M6YKH
jkWxxEqHPLIDblGP0B3DGUhtWfv/bLg4YdpkR1kR7zTe4+YcBT4cVe7i7ZXl7FSO
k30DRJt+fGttMEuyJp1Otv1b/aFn17AOUISIEOKqlL/RXaohV9Oivcu7imCBkVQg
gf1I6U/tUCOzF8uQr0B+c8ieHCeAB3DGlcpNTvWDUoh8u3LPi0cBQ+ASXbhe+TbB
gWSQmCmevBCIBOdf26+Mh/1f5w8tvXMPlRuYmpJYzX91+ZDEyBqbf9Op3NyCUWP6
1UBNiSWZDiybOOaAbxr622Xod/qXvE9MbvX3HVFvoDK95C6p9jG+H7dVCVaGWdyF
iegSAtWspzGpPt8Aqi16vYQ4bguI2E5bpBvIdQ5sEA2XbOBf0pp6k8s0duGXG7Md
HC6i01oy/jeE/mkilptdMtaHxo4NlZXTJZj7drVdK3Zem6dOB320nU9jlEeyURUx
0KMZg9GrJkTBsjSkKwQIAafPZ1HXaeeaB42whbFmG/AAv3UoNlFFs2o3gj5pkRf2
7zHe29ewjDeFJFRUtBHPp2L8c8Bdg4H2aeon+MnCu6M0BleXVjJx8L1Do8ZZxb02
4BD3Jv91LlgNpPqqfuIbJz6SOjZi+GBhDCBaY5y6M57wOeFUDU33RYlt2BCx5Ene
rg+uieEakKnoHy8yzG1O/MZqSxg3gJSZCBs7HoDBITACH9UAzGnJ28lCl3evCTJ4
9sLr881P18IfqOOjTvGnpQdxC4ZaF3nvqz3zBnpBJhT7TsJoeM+YPdgjwxCD2qjb
y4kcIx0nqCdyPuJZ+f9TVdseK+92secsId4uAunqPuSESSiBkTznBuPScEEPS+fX
Nbi+91DTpS62aCCjKIY4GYL9hbQxLw4R1qQf99kzoZ/y9lPDBSkb+8iCGpjtbHpF
3Az5KRdh6mpQwJHSxJ4J5xIQKJXfM0hBUMK9YkWc9T7vIEramcYysmm11jBu3IVo
IRjyLLWvrxGbgLT8z55LbZ1r5ws8pe28p/ne49zngAlAsUPFRuv4TBBzNahDFcuD
SdZ7dyVFfFE3CXfLNF2LFcep7qERJ9ZLEueCfMnNoSI8C+OlODr2Nqu/qxwtFyE5
5vdYAUtfqCJEWyCeRC/P4TyiLeXVY/SZzR5bpLTd2JDxWpC04IdDB/olpAFo7wF8
cGy8FAQgyPh7XZLStZaWoH6bGntKxUV1paaYe2ioOWkiblJ0j0r/hxrUuQJwjtvl
hkGI2AcU4J6dJmeZuM3XCQ2BLjlhkpE5uOK3kSESUVDi67aVf240oNVYVPW5dm/i
x/Z/IytHiUyzCIr5Yzx29JFZedmjRaq6H8EJN1g7AJ6nk/oheuaB7/ppKTUh/KGw
bYXzveTqSavq77gCYdcLEo02dhCkKzVNMTQ8HQmBJhHzOLxVvI9yJV0Fv6yexclv
tnw1ALoIMnOC2bUfvI02inTq08PkOiIrorNii15j/jNKj2ouPUwq7WcqmwOijmfP
Sr1E+kLyLi3CqqfdXgimXH8r5uMz4+CaiZQ6vl9KxTwC8knJcogRcSHbN5bQBIPG
wVfPm1+pPW0eZfjsOzqyLfwubYWKNjx5Pf8jhKwqS/3V6eb2rvOViKyKYQg9qeFH
Z5EdwV6/bdBpJxEm0gKSOA/cxosNlmzbZX15H+I9hmTINlNumEgvZ/2XU3kiQwR9
ceMaCP5YHA+XFm96S/IUVkRZDr/s1uEF3kduhiPcJj5Nfb+PHTqTV5eaJ470VqIy
VXm+z2ywUSxpe1JHeDTzh3vjDs2XwE9dJ9ujGBZ3iqB8ivhYHJD0ZI98y9bTBR0K
g7j/9XJo3VeFiIWz5Co8yEBRSzNHIZP+ixxNcM/rr88EkONgI5ojS/pxIXTp36YY
vFPTCBBUlPp6Q2PzJiTdLWwzGrdTF6JUH5j83pnfO8iijLHLUIAAfXnp3PGzJ9Ze
m5uRhs2n3R0o4OroYg0PyMFLpy6x0PBYaogi8CZAbVkcbkzHYyYIdOuLKZMyuU1e
9BNXxsC8ZdO2/c7YE2uGxZLthO+b/0HyPh6Z0uJTfEcHIgIqxap+E9fFPydXhK+t
oTBKkqG2hehWeelliTkZveltKx9kSfJoFiuTWmXOpor3CuhBfi6Av6bDEAC45Mb+
XjLir9ublihho0qKDmWNzS29Xxzhgsg4mc1ktApHiRBZ0Z1CzU3ReEgZfqVkOAy3
MD/h7m2FGRasV3RVgvGTxwpGbfx0vRGJCbHXqrr+ikn7aeBdkpe9s0usXPpWvrNs
zWmdbPTLM3B7FkRVis1mnDYnzMqbLZdHvna+0NeCWEUbdHF+aPKwKLEOCemuQBcF
Yn/h/CfcBjYyptlPhxvWW5JygE1zFaLfxAFpU2aZH6g8XMaKA1eBxqkR+WTcAXFB
k/Ta56zxbnawUN5s4mOh/O7ZtKfxWCVchvUXeWGrhHX0oPGep9qzJKd99UGMsmVH
p0ElUq7qf37rqP4/k1vhvqBMFqzBCmmtafILqvaboj2tFeeGKZcJLIu5I7RFsGq8
tSZt8IDm77VuO7yc8dZqsnoEexU0LRnspTd4Jiy4PXDHp+K+0bXBgbp3ozCoTQfd
g5Fh0yuyfNPumfpiOrpU9ymnAivNQe8stDNRU7qz4+XYhvJUbfpJ/GIFBBxeaVz0
RdoE0d58pCLu+9sISLzI8BxRpUypt3PREtIjFd15lU+7jJF3Yzgpq/lRw8d6fYMD
7o78tmDul2qI4Uf2iB83bIUv36Bxcfk9w8c6+1h5rb+WA+8C005tWaFekOZq7DrD
+mS/D3iFhNpCrHh4NiAgccinhLPrsofYCCLp3URIgUj5KU5RNm4I3PRgX8z6d22D
ghEvbGL5IbhL6Zb5p9ojoc5Eskt+eI31tZJxQ9vPEUYdiOWimXWQrR1VOaCeye+0
akmHeQjn4NuRFPNd5zWoHMi9nPTnRGuNQTebUnSWjIeAY7pWqVKsedd879n89m1w
Zze6u53Obwla5YxWPOSenNwCHwjtmEaS4+vFse7f8BuMDTKiGLQYuSBiTsDu+wba
t+c+XGE0AOXmpZqOPwfUysXxO+F0pV0JT0z0zOaSG81mszf87EZLYnP+Hs62AlYB
61rbn0jCUpJH1xEUDcIFxTk+kAA4C57UpKblgKe3ULLJFaYHdoeUxMn+CiNU0y8J
UIVgWynya5jqcrwmkezdcU+YbqwV5Asr2MzbbKFj4WNe4OFPJ14z6cWVRX3UpKap
W7B6BNzaLduDe65cRvBZyCt2CneclX+bsIYGDJ3hpO/hu1uzt1tzteLLw7TU3baT
iA/Ea+1ywSWh8Ue5MV5ZR8RSHy7LVAHpm4S1xCj7HvQcB1n8PeEm+un/6KjIGKn2
vb0e7CBFO8lncCFOfVgZpedr+BdGRmB8OXVw9ihP4pM/ZzfuIXSJJIbcEAghoboj
licEm8ex/krJrdrHpnyi5JPmO2CX+iKqhT6xJ5fuEoKKy9gipGl/ghL9+YpSarBx
uGv2M2xTZLSJCA8ZKB3wBLLKxlWGsUs57dT/nf4PJ4SnULk9eFx+gnybbcvbC7vV
52hQHtZjOGCE2Ov7qg6kR85DxyDUkYVmCeHs5O0tefCn9VzpUt0NIyHOc0Tu4QZt
IQHMWFQhbSAAkrPmhqmhs1n38Kt4yEQ3pd7zQtZgYp4iOEEBAHwlglHs02P7R36v
7pwpnUGJ5gkTe1Q5kQnHKXlK7xq0+yg5zJ+FIzh8sUaQokxQD2Ihsq+fFIlQcu4F
NdMmJEizI8aXGvCDKO4aIsYDiiV1f31AGUORJb0uYja8tDZxrGPTJZD2VNmXDWG2
PXTC1OZsg39W3ApnpgkkTgOpi4tfwrug5EPZPImxgT1tgJf8VSUX1Qb7/kw9s+eU
vjqjZsDe085G1kNVgddbnc297RfUFcJA2Qb4FmgwdeIsFfmFD030tQVfBMUy30xT
S+/hFHCncee9YmD0BfdiSfL74hrgDgkPf+HUMaYrdSrIf97wnriOmycDKpyBiCo+
Jk1yzNCYutZfsT7qt4J7a5AF028+KnvTmPbF8BE2+Ym6QrDu5cyXuVecQY9ZWgU/
GU4q9YkW+3PvDCLVtftWlF18FOk/cho6K4TqqGsdL8MoZN4xZpjH8OUVaHG9rd8y
wx+fTUNpw+24rswX2CSiOsjr6d2H6HX/DP1i5OSYjGnE+yqheHF+qjoL2UOdcUHf
SUTZNdndk/bScBvl4gWkPqwmq/4DB1LJZc6ZqTuVxi4jKg6Nm+3bj9LizncolYeS
+6bBu+Uff5N6PkKAXKGOPK7Rd+QSu1kfk5bZcpwR587oGrc7nxO7+2uZHH9QvcFG
JVOyMyYuAAuQBiXzJVB6XipN+xLAalKqoA+ZMIupXGDUOsZvxDeXYQjoSyncbcFc
jH1UH58Co0RTvHLTafW1Hya5sbFQi/LRI1M5Cc4QPmXi8Rcn6wzwms6t0U5PH9Wu
OKRP77sxPMwfCRB4kRBkhW+A3n4v7b79P8wBHV1Czsrv1OtcZiogTBULeTXU5MxC
C5hrRQFMqrfmdJVHmCr3cdISuVvm5+eYRqFYmDor3ylxLeJEIYHj5gQ+LFG6/cLq
Wm+yPFRVr4hOLN+9VXqFFM7Brws8hX/WAa7nz3Hv5EzDmlJALa/Qngl6+QBsqT33
tRuNsvaHUTEkILz3WTBXV5kRpEdezpkq7fS95cvQGG+GnfotK8uc+Uev5ap8v9EI
N4BL2lh0GHE87DeKd6Iamo84e+sgt3jrS0uxHqQYAQyx/pRDSnteHfHLYh5U1mWH
L5kTylm5eOpFzCLUXhmzYSE3zoL0Yflid6usbQmSUHHOkXf4lu4Lsxln1mqOyp8p
Eb24MtBdQsp/L72b2Uqr7UjPcwiZguxdCOHb3AZjys3QLYlFeLlBGPfFYDrB+GSH
16HR7GDYJLhc5aKuTrKQLGp9oicbyIk6lJKrdeXDJZEb5a2YEZlvQ08mM6WB2F77
GOSNaw6xjnll4dH7sfRj3+vWF7Cj3ogZUXAVsm/kFKqxnAJNoVLvkc0P19nF69Jc
oz18SVRGxPP/NCGFFLRQptcZuamCwVhFrdOEwC5ceIYPeYLaaKMsq1vwMHOj9toW
O4m3zD0B3rGcflrwxIXP1t0s9XGuH0fj/gNx6/ZVwuhAjM3cObpoYYMRjTtVBInK
nhKEUEZOFLY6uzlkD9mFlKAJtmZqP3035lJ4zLlAsqjcunzJIIwKASEkiG9LVV8v
u0Sdustg/Wwn1sv08tLqww3OvmDEK+4J5UtipTGMbkcCekTzbyKmg2MkSDJABR3f
SPANhm6Z4tex8IHvT/XMdm7vvcPQpxa0ZZjtblYGCodekv4NhacpFw2a159vIkGF
8fv4JLQb4pf5qzYnmWL75cbe0IYQyyK1MuXopf/7mkBJH4vEF20Bh0eNuFZjXu6g
e9tpBjl1/4E0lYwx/zGH19F3H94icYur3ZzZ/SG+DTqTOIqx91IgqenLP0j6tN/b
JYkoNpxeVGh4mXdrFpdIhS3bNA0Ts+T8IhslE0ZNShq1hKWgWEH2Goyy/2fjMkxX
CJBduIwXwAwPiGJ6AyOTumbAYI9+N5qT9NuHVwkZ6MLZ8y3H9TZfwYSfxsZ+BPbM
AZsv1MtNqQIpbvt3xLxkJxDtU8y6gywOTyxcyGPDh8u9jeCjrkdNldPAp9iUY2K8
nuH+swCv7P/+FqjpzlQrqQEu1Nehjd1I//p9gKgpsoET+N+ogxzRltlVtWuTHYj7
VLunu28HRr+WGAiMI7BeWrGOgLFrX4BulUtKSYFo8G2GfVMG3wfmdPHQclEiniUO
iHjjBLnX/AbBZfLJcCKCtCT6npCPBMbFN9+A/1YzSrGkixaGBK8U0devhtD0loiu
bTteewfHk07+GC3b+6o4nOj+DZjFYHZ0/4SozVjJpQlAzZFU5j0qnHhxyVHHT+eW
LKhkhhcDh/p9ovS5E4c9hA/zfuLtMmxZrQVy7zCDePS1kJj7ZBIpppivQ6TQMe+f
eHiMumN7Lzd4wRB52JgHasqSIugiYdFtfyPtTqQjMCAC583ss1geE2PRTsFeriYy
FX90eI3ZKHs/YUqLIDUKCLr84HRdSvuc5TOGEZGGnRxYN9GtWVVZCNSg/7hm5zs7
6HCElPq1Wu0M3xj/bontl0T3npxhnW3DDA2vAFLjpbI5j4uyfDYBU0JZLIvlrTYz
bLZzyWGHiv9+sUPkaSkU2elKne+uwtACU6uIFFWhcgmkwhxE/sPqHtYEZ+RUKBCs
SsNHjvZNhg4x5k+msB7QSiz99Hvd8cBsGemyXgagegEd4s+U9OyF106y2zse0JcF
kMhPjVHte3dxJG21UliWTN0TdhViagJ6cUOrRWt0BG6rTqYSncEiVrXRNYEU+lmF
69RYnADIdgCVIEK+vzlS3icMkHsrZAjOWiyvTsLjiilIRaZxBTkiEenb4VymYohL
YWP4rtuOOYs4nmRsG3ofsXaHazdX8jrY36sMdKY0bmoUbY0Fu/ovyPP/mrtZU/3j
XaYgdxXDe7aqVrCkgxe+6rvMLDNffQJLGY+v03U3pyiMgh6LrpCtgimGkM1sp8Jf
UOQCIoEHp5rUTKzkqFp2r8t1E1zSbfefm+/XfdXNUr0PWi0ddtqcer6bObX99Rtg
Hn/JfA2UwuB0aRvJ5iHRCt5ldeXKwo17O3HA9NSWYkz0ZzEFObqqWFCfAF/ZRqZT
2I8QlUChb/IxumC3/Ju96AZoXD2zavCRQkFMa0hyKnNTah1pSUkKS7uMzl8N/ARE
XkHjs+jrRx+K+Akbu2IAc1TuIjsM8DPU59gP3e/UhnFuBwL+xudpyaM9unQi43kc
biW0YUEyiUmZUmbxfp8rAtHryeIGQaV35b4FBLpLdTUfmhrjUwRS8QgTv9HtbE5m
h/blJLh8BUOtQlKXZYjp3+x/Sn9DDL6Ss4tnjeg2/x1R68Ue257sEIAXrec/5nyJ
8ZUsHtl5FlBwHeClimzrT42C3gSz25BYhcieF0o4akzoiEVJzuPpfkKVzI5VrYUN
r/jd1y5P2/6nwHj0HGnVISAqv1acdZVd+t7IUUBi6jYkLNpAKxR/hpxJcifmwF0g
K8aR4OJncGCnf3hlga6qkII3gz6rA5hLwpZ/g8y0WcEsM5WUQxNtagleMeW2MF/v
ssuYR0NyJYOZ0WnFx8lENnD/63/R1/oHVK8AkmbcVfMSALSXeA+YEYddELc+ZFlg
Ulvos4IYFFSA19pge1FYLXkd11B9hF9EkU/t3gA7YnudXh3RNnI+GK9eWjue1Xqu
z+eaZtW9K1LAW5Sp8PYd7WlHmhr1bNzWmmMnaQ+kAbYHDIrJuT8A8Y7B9TQePgGi
+TcuefbnIb8Vq4/XTe2umMEYUcTOMkMDp/5bVNPEA6JcEkNwkarsdVGzKCePNvNy
ABcOBbZIITFqKV6HzX0BdHEJxa3+ROnXL0xrOj4uzwrb5aRFPBOcZOmdqyX22SWT
3mkYIKuoN25SFWOKi/iICLjUNIUF+wYcVgR+H4xyaMK2Z1GUT9BNfRmEG7515x4h
6bmcsdsKyb7WsKsbsFNjkgHt/PjrmVXq3NbwseIIMVgqrGYylC+TsV2irBd/Moe1
tQXiZs81izwvNwEATdmvLoSYhyDmsWQ3y2y3BC/aa1cMGDm0V1WRb9NnqJO/stoD
O+C9wEwYbfd0Cqkihsqj6McJ8AaDHttDLRnge0yI/pjtF4elyWQ8U27SlMe1hTFQ
BASGEqIvkETNEaArDiGVCskrBwjejP3eK89uAEPSxtAClqmplSi8f1pE42CshKlU
T+T7Usdaje1pFHlIRFY/wRo0PR4RD+IiF5mAYl5ysEAJMnZmegsXkbTIotKE7RUB
v5p9BwLC9w8s6bBwy3xeQwELO8oe5sbDMD3/QDZPtj6BGU5Rsb4enU53s5wrplGs
/CHFR7w8kKRv0dok1VO561v7X319yvTAKkc42Onnh1bNnt0Gxc+J8qdjwZ7d5lzG
DKIoDDAN5nv1kuUEmKQ7PHeoS1r25tdNtwTFFHo7Np5szFVgvvWACzqDNtFOJtqo
xBDE+tnfPBkxYPyOVvsaixrkft017ULn3pYZD//Ppx/6UdBPRxH2G+JBa/4uOg55
UF3CC9EWFH/f41H5G6h7oNNJJ3wWmmcK7BvoJfTAKwDvZWfjB7Uz8AzPuI5it3FP
sMXW+erDAJhsTD+4Mw9fZXhlnNtB8VNI8KVI4q5Fx5g1T/h95rN3S/17Hf4iw/OC
r2BKOzMcNNX6DbIqkfqYtP73+SyRBUDxghza01AbHkLhE2yEWgd+dYPUET4Jy1k5
vvgWz/TnjrYO5Jw5g2NBNrLCqkfO447x4M5vQzu4EzCLe6qn5mhJu2JFmVsRrXid
MbOcA8ckOO/g0ldWiClvymXnbcWjr7OVctsFOg0+Uwy7sJL9UcZBuwJBbZ8mTlmG
YV1eUq7TX5NPUw5KvvPBt/wUJs/A9lkrY0YN9bjV+ptl1IfOJwkFJqrpzYIxT40o
mXxuk/Ujjg6RZADwIwWlMuHOm4k2L16FgeH+kd0i4ps2HLgcruG77tvFsVntvq2T
oSRt5dLgs7nRDAKnfHn2uRavyx2GUIHtoGdP1PE/YjIeQZKO+B9AEPkEciDio6UL
2r0KPvFXsF5ICHE9Hek5+u9bZwB51KhpDMFn0OOOYkK+hbGuTx70FIePA6wu+vVy
qMa+TTMEviEA3w+yHAQishWPHEmC4Rq0IBaFpfq+Tp1N7AHdUnfRtSrgcMY05oxB
kAfHIyFh9RFK/4T6ZjQnTWrL5PDJEB7rNK9b02fnPyss0WwWm9JDHdtRFzBk1uK0
NtnWjPZ8qar0+/+mkXuw8VBYSDKN8simbMvSIABh3oP0GXgkJiJ2gMI7B9nCFeIW
/AsTPXp2p7OQj00biqIm8dpPAENvDCQExyjPPD14n+MoqSYPsIF+aKHiF/NwlHg1
8R369c096WzG2Dbi2LFfheg20nhxoo9Tvf5CxXT+WBS7X6gChQjO8PixBzNteRRo
oPRkeDSUy34Y1Kmk8cyJi19WVgIUAa8Dy8PvS9B2QgCG1cQ0rlPhg3xT/PfEmTAn
MydwtfUA0R3M+ZZ5yWBY5Nlt4jTsB14YxKcQJSc5/Ko1Xs7k47v1sqhccPi7Jj2H
D7i766sqlj6Bac9L1ykbz9YcM/X3Gj+JTNxqAhzxwBdwAeD2T4fF6mbkb3YDoX0S
q5VR02eiu1KCX2kadgg4S9ZpHCL75r7gbU1v4IMc2FXe+W7UEL2kgp8DSslg2o+m
t1GMJxPE5lt9RhZWSuYWFq4STIphGuVBk+EgzyqC5as/J+Ge5qdIx9Soekz/MITL
sM0JmFDgfg/P6yWT2VkOG4jBGHUkf8wbm195ZaRyQGV6DTa0eUwCpaL3zPaEn4ai
I5U0nzcwiFeyj+iy8Mc76F8P6WK2PHV3cZT1Q3+6Lo0czZHyEQDp0GgXu3bty2fW
Sesti44SBfmqrOua0EL0z0EybnuUe2vp8QnB5N+OTJ1zmvJxVsL/H83dapY9Yodh
Lci1NTbFwVsYnNdcP+rnyyH15SMQiwOE/LXAA67ss0Af9E+mF/VD330kZwRjJvoy
yxMhklnr6DK9lVxEXyBGhPhYjQ41iLrer+2dknH4lKOjzQW0cOwdD9p549SM+G4Z
CyYSVd80gQHmohtPkxeWuu85WEplIyd1S0K2IjqJWlyGBygkK3TEqXD1VrhXGC4+
A6IZ1mp4URJ1lWTEDx50jMkA8s485of1h9+Gx0C8E3Mju302Jewarmatom4Wx+2e
rXHxYLg6FCW5VUa4BH3doOghl/2bRv4KaTEgXD+KLOjIwnwmo0QyHP06KPgvhSmA
hKw+2YEWt/UndZut5OvG7ViEOxmrK7H2mZRUay216ID5z3zwlOUN04uYSyhG0/te
eL5b+UykzdATYKAoKYnphcBJ+oA4zOVREr+8+hMPBAcXMLapLd4pDJBnkp++Fqdo
VSB9NSGPAH5cFBjXNoGRfcAwtw6B6+4qFk+s7VcFBLcBDagLEakBPd2HkFCwDLIB
dMwRiDWE/HvI8eq6N0cAERh/hEKkzHp7mmUbt9AKitXTovnHZYr0BDGjKiOVtBQD
YKmgtrG1/O3boeg84G3fA9osmBX/CXUF1wQV+uEyKckHwR8KluMrgAEj4M0+NTir
IxmJuSmeL/vvNXuPFtILlNa/RODu5v91D5ris/7+KzuzLja9FccXyrDWGoh5Rv1D
6M3+hHLxhvbzl3Pg23CoL0KO0cwEjpq05PBR8BrrW/WZ2hoDRR85tOT5xKxTQBIb
W2llKdzgnWViHMNjkw5eTL/3wGIEcWPiR5mgUAXNTkn9V9cNjrmLMf1j/kW1VwOM
Mao01JVw4q/pj9LNS5uxK5le+WWHS907uNaRFG3CwihSlLyAVx5JhSonYQv9RAg1
H2e8meozcIkmuwwjYkQAlmctmUqNVJLrZYW4JtFkLsoXgwKRPnxcvQCLksBWniTV
AxR4ois0ExV4Vr3PggLoLGRhQOlobFfCaERepNse72dcz8OjAoX1b9jk9wZQ6kLn
XA+JX1gzWguTV7pO9IfuCwgrF0AbMrqhjb80PZ4A0WgQNGWRNHiNvzktOpeTqZC1
nU36TLrItz8yqWoW9qVrJb1iNUGrh8cCRkmBGpL+dd7MdIzgSetBNIGWVfEx4O65
HkrpFxSn34+YflF37dEPr9cneEb5lVdEjrGXTeHcpSNt4jMNz5bMQIAeg2o6dYYH
msGxoytm316J+lKwN7E/HLRz+7b+KQeN335LhLCGD4zVd6sKbljlkSfGr5f8sqKI
FtN7qRDt5GQBJeNXBZLb1P2TMpGymJ/4rapNShIYjHq2DWSAEJYPd/30Dte5tS5E
vqzNXsw8i+5xCv4OX5Zksw55VSUl1IoAGp+YhGn9ukfXj1cp7RKYK0Rz7j80DNmF
hAXMZrTJeNu8toE2h/3UdCfm9ix5zuX3amjzlTNb+hsR1cVBHwPks5sSVYm8kqAI
ug0fjK6kpmorK9wEjJCWpL0cBuq/7Lv6oE98MJGyhUvZOnyots/SUOr+aY9OwwyD
2dakmjNTz1UJQQIhCXtiz4A/PA9DdRPnnNxpQmLc8b3t/jAp1Fq+ZyHB7d8unhBS
jO3jlNLY/A7twTMN2Eg6lwdTqTx6ObbiYogfG76m2OijR2A0bHmkGr9uCmOn6/IT
7FzuVwORmsx7KSRZu+uNy/oWxJEDx12nP/tuBiwBd7W2BgBSXIjmeGcQ1i86AcU/
su+PAoyYlOw8VzFKMfhgjqEKISUC2p/IRJEjLzyQCVdkd0AGY3jpARUHh6Xh6RVg
9awBtJmHxoNTSvBj4DXRLtULdjJtwnQmcbA1olCgYzaA2s23+z0HzAs1fEvimkAt
OkAcN0eeJB2CcPWde78vc/0piO/sqgM/IDrfEJzYeO0rTTkMbdvz2EnLmBUdZItF
gAxgZgm8n4FZPtDMizRONkFOk0Qli4YjlKwOKQFTTDBTQV7s4ltQjm5FYWljM7UM
XrbWOw0uIfJdg6BlenXJkqknC5TtHDPENUuAlmQ1IwipMu/QGQrds78hvRQBDmut
WXbvVVz9LBp3sFsTN5JTHpI7WzVxMeBGDmM3y9XqbVud3G/ph3QB9trWfWssWaeM
b3UAQSdu0OedMTd/ANoGME4PTP+H/8PFnst3H/Mcdt2b2rIWZyjYK5odxagtt8/Q
jukSYJCMvX0J76jf/x8wgQbpo7oQfAne4y2Fmw0gLKpyl884x9p7VmwJyb/UP6jp
0kgiTrYjmGpAsm6IDHTodxi5MRwZOkdyv76JeNteORH4ollaUPE33rAVZ5e4aftw
I8DOrTDPXL51Z3Z2ibCCuWNJXV4qLHAlAtpBGuC6Rzw+tHL7WubaqHfume+nol1N
63wyR2qgcyW/3W3UlWkKd7CZbI9g3FFKlcRDJD//ds84/TqOY82ky9oFW98xC0rS
dNLQ6gT40SXhoM6tG0gYvm0oYv/0zGUX7s81BRKAtrtzVvu5uaqK2koajgPW1IwR
VhPrPr/8269Bk67jBAfEMBZdE1tsPRudo6aGTcIgwV3Onnj8VEcg4KszxXHWnbGZ
6lKANco/OpJ0U2vd6P06SuN5+SOyOn+Hug96ZHfpHHiIyVboziayu5jc77u6fkFE
Jncxez2rJWsV1Erbio5JNPX9GQ6E1SbhrzoWVvM5FF+D6tUMk6GlzGAYFn2eEvcf
Hi6KW+wPbRUVnL2UT3WfZsmHdd8/fmyBAe3Llvi21lUKGa/hir79WSFj2X1ZPE6i
YAsXomGTaU7MMmqMDXIy1Bkn6O6Spklp/2pyvMVPhK6nru1fbbMxLtMbIRgpaolR
MYP2k1+aA/gjLmjbcg6hWaNNi1raHJCN9hJAryzo5mHjrx/I2U0yJZZNF3qkCVmk
xzyBd2JrTCgkBJSLI7joOMAAs73GgCjY7JN98yKDy1jbrd0MgHrmbYH92LkLThbF
qoKrY9M3sR6I7w604rD2YudDgkLYiqGN80nZfiltjx+Jpv6RlLR/MzIfg9rIKzLn
9XKjzyAwBpwk/AKtfH5VCXOpmE2j8iJ6DCSbXXBcICUTuJe+qYK6OmGQxaMQyvM5
argwLB+qNn6uiS0s+eRfKAym+FYUNPKt2i748iRw8DPKv07BxGZ+CTo9ePJ6xydj
QyZURjnx3tVsDjk7BJF33tsEZjpf1uKtTPpSp+OjZ/p/m9tLw7ILnpl4VqWMtXzg
E7G2Oi4GNjNXKdFnw+9C44oZYklQvgeGfNBMR7QT51V5MRQJHqJf/OTrXq89Va3y
KmZyWaXtk8J/9b3Etkau/0Mqm/ivjciy+9Ddv+S+4DaGA8fu3+Kj8BafTBhwdyo0
/B4lBdJJzGL3wV8MPzIYdrlYZQNNTiuN/O7HuSsgORBrgXRlMXIYHqX0i2K8CY+6
OzwmVZ/DQpQGXt3s2wp4o0u6YwRW9uTXcKzUfki+Wd4Bop1j5d39R8ADOeSjJhC/
fGFMjYN2YPqbgj9q9pB4SX9vLu5xDo0ojDKmruXzIzmLKESUXrhIijGw63szs03R
Ed0QVYPplyFvG6zMjxF8Bur62xBvTzz0UGf+MYh6rouoWq3fEwG497W+91lTGfK2
lkgZT6VGIJQvU4ODPcJyFu5L+lWn15KrsH8dZLKwK+vR9iOE1zcff9DwtjGlEmst
bo6KBvceIzgaguQ0NBDafR90HKbOXKPYskf7GUB2Nw4q6czKi3dzgTsbx7xOljIE
gSakNqg/93Kf3uODvAybIpgNhSu4PntQbbTpZZoH7ZBsQ6edrmh8g/XQ4xKayxe8
NIAHPQzQodoVnhLBi7Qnr5hQd+PIeLpCWVSXcQ28rLm+22uH4oKWeHiF99Q47k0Z
/awKGjhM7DOnlJeqIB0kbiK+rsBrr2eiYPIM8LiQC3GH59PQw818UPN5IDFlh0DL
owFvqs9fKBxv0RJBEoiNGiS1aJ04F/X+V20GfyGnUmDaKyUyM4rowUtpfM6/6QPf
wpZoNp2puUabhIYWSyvr6hdKJFEKv5XGZnu6B9Wa+I/vYuqKv43TVcykXKdeEYS1
9LwDGcvsYidtHbnRPGm9ROSPI8p4B57+D/qkCh3m8VoR7e+YeNsEDqnoYajpKQsf
baZGrGBSrBtD/rSZs898nR9atVGp1SY0im9/XgUvTlcrNm5h54Gp5sCk4GkC3QHq
gdFVLgRSgJQbFbGRjyjwHeNZAmNzKKIXEokoGmrdyOgmX719mdpAO5bZRe6esgcr
MUNmN8aDaYuWYqMLuoRFAoyM79kOHyqjUB2jdSKQN9ASbam8/dSARNUXr5aumHWm
5N/Oao/0wHSELserwedD7yhzJw6z4P8ofI+CXawzU635Mh6wwmGI/ZpHcVmzaJSb
ky6fxMIlsTylWz2usOf/rirfPepTRN/UPKjJrmJUN2Ojcjr2X/KjrJPE1KpNEoGX
YuSD9Rhv9lWYB/SDMJi6biC7KRBZwl5c9VvQrbj3l8W6b50pBrXA1nOj90MnOF1v
RQ5dZReCfNYkumWY4iFQc2Xz2zdE7xGaoJg1Y8bL3s5pyqS9qs6Vj5k2W6xJBxQe
B42IaB2v9MYoeihwM3bHnVVA4rnUldGBXGDWdOLKLlFUVqw5656gZSCmXoEwzBgf
NkyvL4UBUojzTVlbIt+m6N7gsIHwrizk6apYs3JoNzbMtymGxxv+fxY2O7x8rIcT
+VNSYsuWEJ/BsW3gjb5UTBswp9173TGXdRQ65eKOSe5sjYmIadY2006bnPBcysFy
/LKkybG+PMYNs2x41fbBpXoVVoN3CExL6UbWudo59UZPS3MQp+iTJV2S3s/DIgxj
dVqmBF+g11Da1pLwR2R0EGV+5g8wSQ+s2n3kPQ5RXz9FkMqSXPmrvs9oQbhfyptD
VYHl8pantiTQIZELbl1OuFaK1DOqM4Se42Xzlss4c/2AwADMPRteb+mxOdWud12o
ef0EzRuoI55t4raqrbXNQhIkNdojITVq4D8309rSkhhKPcw6otbZDAKDKRVetW2l
bsrcKVZG/khsPFGl4STDbQrnx6fe6NH7/okke7ChOzPpeakoYcNY4e1ZbV3UuASP
OwvKJIE8EL6kMyqfJ71Z0VKGf2IXyx8YI2/ScihPKiBEiZIzQbPnSjg1iUv/ax4f
l0Q6oH21x6dE2kEqJxfTKqJ3drAMnCwSV7IbAWI7eL96auWzULQ0VbBhpY++c2p1
iUlkevuAebXL64CS4S6sMvCZzi4Jz9Em7bdKMUf/7i8XMMgzzxPmfnj4Ew2sBCaY
nxkmkFE0Oa0fDsw1wO4DINFqxuWP1lNrIsBKDwBWavJIJLELvrRfSosRiXY4eBsa
KNNh1xk9//0rntWqu7QYi1bznCzxHMuMI1AS/TpdkJu8iJk3VbX+f7DZyeYhLCRt
iNtEzWMQHf8HyjxzCwDdcm9OH+Bvoc6BzOX84pQAeigA/V/LNu4KkNSfR0cOt31n
5w9L3dUkz6B6peC01Ri4A57L/MJKPIJxUqkKz4Umrqfdzio2wLAsCJLZw57v5p36
yr13hUJH52IdN1fDhItKO3r6/9kabvADPBuAF8Z/uD4/hSpzgFnJPIin6iNUSzPP
+W0+5zqdeubdIFntWNeXchLb86TndWzqfMUx4n5GdAwbvQ3MeDnyy+SsYkycvgjz
ccfSmCPQwPxkpm6bzjWwbcrwOdcxf8vZGBCv/so09qk/zROj5o9lOGPymrcEcCQQ
ydOLws1CRnnHiZi4J1PC1DTx2hV4+0S+pgNzjXNC2U9rRsHnJk1zen59h9TOawuM
6g2LT77US8+7J7E+oBh6FlJjJdbAXdteHVvWaLSsUZtNphdVISzoOqtKcwQqQ2hu
uVWK4sAP18dxFeAx7JZ6WWcEDSkYFSdq73OX5Vr6Y9LcOuZE9HDd6cV4RAKG2gvu
UeQGwbhqoykgHiMEq4Y6mg3Fwl8hRQQoNd8BOtWvydYfL9rMJuDIU6Wg3FNa3vRp
B4ot6MFXTmYhUdg7/jMDpMxZmO99q5Xhfjs4w72zkJlPA1qg3yCQtK1MUh8UOgdS
BWCY/JvZRi13CDreW1eU7NVDT7Z+tHUMhp8dOCHX2YeHmYTakg+TH/Z45TMuaESp
ByEsbtIxJl8QJHkkMxcg3EWB7uBHeQM2SjVaMQM+3Zb+o2ZGE1Rn0OWyaAt9l/tU
ASYEiPQorCncbKKVlGTqlQpa5nZe0eYP7ZoVO4FXjCCOSFGPyxlFIXvbeDZN1FUJ
ZDKyU38Pp9kNcgX4mrt7vKl1tfcd9fKpsWcCW+PSeOVP1FGOKIUf95BmFd0rkajZ
yzPqtooflvgQskKOCU81+Qwhxo3VXKS/jbS+9L+69X8s+hYf4UGNV+MQ7bDzFZxv
KptLKYvH5NUYRPCPV+iNjly1IbhmeEM0aKFQlPz5mlySIXN7dFi49RHmsBC6qjmi
V6bIFwxydYQkDf9U+margbgz6YEGA04MSM+EOpShU0hqWnT5dwPeF1FfBPMHmXLx
L8e1wBc6YEueu82CTbeCbWpmG8XF5GZW0mfhJ9M41W+KoXdkoEGdf6Syp4VZ+RyU
MqN9p7/LvhN7YwZWpSszIWeCiivWPlNNfNoSFMpgkFlxMIysKv7da//mDHXssm5L
d1YI3vdjW07aVEfK14Wy3X4PtthiTgv74zD/1gJqgGUB7C30E5wcx2V3IbwR7ORy
F9EKLhZuwNhGbJl6aXJ06X5/pa/LeH4at+Ri3hh+WxFzX4ix3O5l9I9lqyjDnHfO
2puetXorjgOjRbe4+SkIBN162mZCwdKekp2/FIzygzKAkX/hZxWHGQSxzTGSqt/s
Mj0x4jyzr7ZMH8yX2Ba0YmpjQ9SfVgKH6YhvlGKkjhKlj0Vb14FMIDqpAqrUoZO5
iCXVQ5yhhSn0Q7rdygwcvWDJdErCtM4SIN4+j83igtC2YCsMtnm8N9/DJr4WMCZc
mZnau5iBcOwx59FoYKORT9yuEYLrC4LfoAz6bF3rG6KYv2EagJjOPhnQQUaNfNjd
twfKLcBfAorCccNLwpUTT19ygMjP1eul7VKcOug2CDVrKn0029rHfoZery6QIQEJ
enxTcrU+hQesAGuNG12dLLKzYkdrv3/GgU/Bg0UiL7uHp6AI0X4upKrgmBlH5cFr
KZ2uaRelmrf0D8MsA23jscJu6KiI10oiFCcy7VqncFbwt3bz5EEqItqID30fa0hu
F3fJmF601EK5lqK+uKglDvmK9BOnoJrrNs189FhkO9YrDX8K2wq6WipNE1ncI+qs
VaBIaWtJwsWUpGkIBdtyn9bbqrukUpcMJWtZamrR/1AXP9zbzs2qdriO/vZ+VCMA
aUJ3ByL+Iv5yrGVMwkQPcvQIUSCqHYnAb2FerC9fIL7jxKYh48CeKXmfPT9pjNKt
2BNIbIw8CUEOwuwF1ZbaeVK9EVKjaFiwuLyjrFf1JN1Roxb58/7796Hju1AAl4uM
lKWS5jaWxCWfJo14f89wuHu0QcBF9XdQ+3BTC0RFdTW9GqSZz8dLdl/mnl/ZXJ7t
vTbiG/bYS5hBbSUleCQWRbs52BVGSrcyV7WA8zcVecccwfp0k322oKxkX9dYh2cw
sG0lxUvseHS1oCCR0x2b2+6JthovuwYZV72z5IP+Y3shxzOw+B4iW9wPGYgQRys3
3TjNR652ag0EpV26th+17H4Rt6SLip4gWsWiZp8eFEX2tuZMCKSwQVHKPwiKGE6+
QKRgGKIfhURpTr8+QyI3+RinFI7Yz0Yhl6ObwvTAEHmVa2GrjK2lKd8u8gR4L1Tx
q0erwbmZn5Q+pBnCOTyK6QIa0jG3WkCuVORiELS7IHOzfNzW0x68PRbU7WdsYA7l
gcppjsRL+me/hXpvXBzE/XUsG995TMBQEnZLdoswQ1okLC9zxXk9tUib0gAb/I/1
BZWHm5g3r+WQcxq0M5Qm0ZoOE1XgXkyFuA+OVqNSzHiOKzwGWME/UfBSNM2wwdMg
Pp45Epl97X4YqMj5MfuWkwKxshvJop/pSJfLckxT1Jqma7Vylcp2b2XKEAuEcC8J
Pjkhu2YLmvzKScpO1cVYaNh6GReR26lFPs7KWllKgcsami0TjQG2uWkI8QlUSP8z
3kEradoFJL3Boe8urlFNqsYxp2ubwKdvLBW+Glu9eWUDDB3vs92DhHVAiZ7uwjjn
IDyy5+DOwT79771ADCEgYREB+/UNjDRpuxyAmwz5RPqcAYM07EoagzG5psqqpkrv
0WEY/pN+L6D/GEwtHYGNYER8NTUC+zhy/FyiN64QRvHJ97V4LnifX4s6acHpMFtM
nWQLGpAdA5i2/QEM6daMBSYcNNceNpQUBI/tuMPt/pHiWdhKPV2ppFzq0nciCXvo
E80HEXOpbh2FAuL7UsrJaH5DxYddOVP6viQRr6Z1LHjtC3mnYF4kvb2M2pxzVUuT
Z+8LSJ5KHs1yUTwWYLqTBw6N/PmTD2BBxKaBjG6EpTP6Cdw3+CzcJIy8rFc6NIsJ
zLDHZjq/TrT9NdBh8euaNiPuzGOCZqOcer6Oaf9bX7rajTCdrIP9SqODsfr4bcnY
PCG+7xY0xFslR4X0jGjhgAx4qiIPLsoV2rZE8YRg646Tli4e929tpN+3cWqZFO7B
3qtDZWvOSdjv9CgbX7hVbOGXvPesM0ojKvnx3HmbsAWHVEoU2HoGAFkfAp0/7CIa
hxWpAbHTFeZWjsDLiL+XBdAhwOLoG3gC+PH1Qu9TxqWeLOUNLlGte1wXhbGaVpkq
RFA2juUHYN7yHyySQ2SvJsEXnjS+R4WvtSDwBtKwf+FyYrWIYKlZylLfIVyZrCrT
3dw/Pxi7ikRILDTSfBiyZyP4PxCDZ4hOpn/+bkfQOweZPYWmpcDyV3ZOg7vw74td
0r46R248Vrb44bZ2uUrWXuuRzKtddWTcXxOmlF1ufpaBNLN0VeYNPgU19kmOQ3qN
2NGVt2HC/ttIk1m+KcxpHQoe/8iOtfwG2tbdFY4QkCT7IC6F5xHQuPazo4rIS/uN
W8lyZh/OCSj+6zfS9BzMyGljkmz2e6eGmCa0Ch4V9X9VfMFojcLQjEKP5xqq3n+m
fL08HTz415HO681fbBv59kRV+Ma8D3CF8+y6u1FH4IUASK+sceSC5vQVBD9neiz4
RsF4PXWG72A+pkJNnbQehNUUzhmuusVM1RRqUoumHBV/V6sa6HrxrzEsuEJs3UJc
aYD7D8sQKkfpCtgohdSe3QJU9r7pBpClImSIc0kkEjEK6zoFwK9pX7l3NSCandSa
9JlwMQXvI7GlWhKIIlIm0lOaMnWk/On9bKgPdywtcnsK07B1sXSLGw+sXKfqVzQk
1WWHFoz/yBTqAouqoZFSmFiDbm2D/4RGIudVBf4FtspYPFfE0QOKefsaVFSCERKs
WegeDR7xUcNPaO/cW+SU/GTko85llyx0OkU3K/L9YZsC657UkAQ+DTs0ki237ZEa
2gdjDICZUFtop6NnqcLV6UTiHlxq8nPTd2DAr4wrB6Rd69//oFJ0gwFM/IkqTZSR
/QfPprZKmi9ahzZsu1OhTUA9gaL9+q+n18uAe4LIzLOMQHdtvWqxSvAqIy/uHqMk
lDTtHBlTi0t8ihHfXD6banJP1CIgjclbL+52Ju8bVFBZxNfyfN82BpOvip3CxSiw
BlwZf2e/fkoqDWDf0ai2sY6b2WkNvAAwper40P0VKQBRgEfJtC8/YDIE77ibf9w8
wRpXX2kR/9ikzddru5vajtjEoJliIY3wLgsUliOpMIoYVXsPzcJKMMOms6k0FWez
LB7Q5yf1/KL1Z6i5mtAZp0jaWa8ARgPtUlTOu290FSXLH+ny7uuCpt+4FlvmDxq/
ESsLaJkBydlk/9Funa6ze52NGHh4+82jx0KpJDa+3ISyr0XdJgOMVoE3evlD0JXR
JRC0vVLLKUhm3U2x3HIRfHhUcfelnikyvSFMDCkubPjNExqK4R1wpKf3P4PqpL6I
dzNe/el8nWf+CYUKhia0tQ3hRDLH9AItYXx28y/iSXFwjweo+Via+Th/BWXN8TyM
whiZ0fy0P6cUhNng/V2Ceq0sLZPkM1eWnaIMCL1dR4xFIM0YrLDL5ME8VEDyk6xA
I9yryMdbbE2+jI0wt0xZV5WXlcWsuDyMrXlRezXQp+PdACvDX+Gr3b43Al4Q9Cps
gzPlRwBVM4/rKqG1tS9hm/Kuk6etEMJrTIMKZBsduEsC8BZqqDUotnA1fJXlkdr6
vH0aySnPH57G9cNIXrMypNdCT/YNn0OuF1+H/fvbnkb2DH85Ytkj4duVomYFaLro
ZSRlRJmf+oAOxgFlZZQwV9+jXOXQIUpa4IN7YMre72tCCtialMj8HGKZFeSVw1Pr
skmplD0E0AnYFRkQXhagTZnnhZcINfMjHCmBDJKzp4irHxd1Esnfj87cuNlDCtZI
ZslJk27UP4tucsDPpa3waOwtDZJ+l+8+K0iN1ucmwjtFpZYZGWs26CUxJUY7N5n3
MuMXUKl7UaCYXCcoKrES8JxLtyCdNxHxhkR+7Db5VXNLzmDsA0b+/DZ4kyr+Pest
m2xkBwbo8Ds0+TigBs+fcJW/RMLao6vlUYB6po2t2Pncb1UdntJOvP999U85Ha9B
3wFepHR+6MCfGqbf3XlUHAIJaBO/Q+n7A9fiHydJ6n0G3CPg3FfSvUNTFIXdRcMN
jp78fWyUhcYik+h2DAY32wgDLhoVgPKze/aIjHDbOSzeiyI3QUUmSlAi3xftN4RQ
Pf22RNEk6yk814zp0TlwCOcj0k+3eEb2nkOvyYL7YzKlWBNnS3YsrZJqSGnxC+06
o73sFHIhwFOF55jFV4lgwxsGgplXLoxMR58N/dI1xcPnx6iAerA8Ky5yjyP6gWyp
pOF6lkd/qWlYJgt/P95QexCEIwVxBTJJ5B//PiFHn/iuvrb3RQp7YXS4JHfuUtIW
nyNkTlGh5UNy3bFNb2GYHGvA1aBVKaLSdlNHWLZQB00Vg9eV0uVT6XwQSqI8klxf
faxI9khTvtPXvtB7GCwAeoih06T5esPm/VC0d2l28X6hObobtHkovSJSYPSqek1n
fIb22vOG1c1J42kWP6ODgd1RIZ8hOK/bI43Cc1Jj411o87bmDxmNCOT3gcr+EujG
amoFetZS3zmJIAOZvAKgYL1YftVU9z6gaAtxd7hpl/6Y1HFUD0nmxVfV9CN8OpT+
sNdwS2mwCyo4cpln4XlY7Kguf710/cj+kGhJobTawJmXmy1qJxxtcbJF2Ey925ZA
RN+sMLpszgxxNyUWw5b6L6R4jaHr0UndoVt6TibcOSaqR93ON5RyM30KUvrbxmdB
3KYIDQpGK0q32O34C+JWW0dA9esZx9pAK0yiPGtAWYrz2oA0GdWGUoU/5a9PAmlv
9pheMV3V0AYj3Ml7LOZnJxrTCjBlF/KSTcIcw36NEuBSjTFgbnVTI/kOxJ+O1V9r
V1SCg7PglgZFqtAD3PpD9Wkb/xGycVUGfZlRgW/hbxtPQIg0X1Ur4FL97LgjjXI7
6QkUSf27xTsANt7OXzbhMoQctw2wpmEztvjaAnofoEOH/kqcyYIow+u2h0ukjmz2
PyT915reqWPafW+aEMuXPIDOzuO1NKCt7cAFUw40boAeXk6SiTOei6NAe+aA2IBH
/s2NYTP/vyrFICLYJMAyzErxJkrUxxvDGcHouATKZ2jYrv8CWpEwYcmwMlrTpICo
WdVGFrUDbQJEKMS7OCtZVtq1VoSpqk1TuH89Sa7Dh16KNkIRCKH57OqWcTjoCJMW
MkD2W5PSgUx0qIcI6mO5y63m+iQZ/HjLA4OocgomcwzY+Yku7vY0k9ZEM/7IgnrO
gRRwP0I9A8ieZ7xRgBG8qhi1YwHBdeglZPEcvLeTlVhfTQIUQahB9B2STIkDcz34
txB54hNUtYmozoDdktzDXW2I5RrNoy3KUDD95KVYID6kb9d2lWoqTicZ6ea/q5Kp
eKOpa2yoneDqy3IYQy5tiSJXAwW4oy0c3v6uWFt6fT23OiT0RSjv7v9KtxMq1a3S
saKFOQIpcQXu96L1yzSevasuV77KeWpTShUoQpgkxCGyd6IN+STYQF4u1alG8g9h
lqdH6LcFiLKYFZ4onxM/YpFiel5EJvs8+r4GU9v3njfdzeSnKtb3wbm+XIewkWPW
bQD4BkztK0Y0ohTbdMusfx1gW3cWN8Q3MCHIPXxNaraOI+Jzz1GmTJ+GzPpu9HuX
b+WZ4/N10h2lOYhh0UUHicEPwXnCbBDHloZ5u9nvsDSwPx3s7CMiRoL+1F00LOOg
fst6xSCXmxlrXes2hxDlghvSW8yZdtRthMPt3Ufa/cVyzeGlawRr5vmJGK7aF7RU
luSJYbdk94Bh+gg13/ZA7RkOUMlKQ1ymvNIiS9egUlA9fVNwi4bY23EXd+Hjf8HR
vkIJIaJhS9F+vjISZY7Bj7eqda8rKhXl5jmE6a2+d/4/vTRHjbH+ImAIQzpTTUk1
ph85VCEvyVGA+eBv+cV3H1U+5ECknjRdv0rsziIogAmGHywRt0D6f8tKY8XGFkJR
7WMMh6Ww+OgHlv5s1o8aTRXmAJUl08Yk723Aeu1A6s8c+1j2sOovm4WiQZR2A+AO
ee546zTSn8Btqwn/C1prbDloEMklGc4IPzrpb+2p9HNsVBjN5lY1uuWTtHhAeG/e
iEEFLgRkcXnahWcM9u/whSkz5zqTOS9zHGtG6qynbjVGjES/hN3Ns/+Z7ERqi0mU
Y0j5LR5quIl88oJ1A+0RPdBGn6iU7xu0LGDpqFxSF+0PQTtJUsEGe0Tt3l7cDvnu
vEuwNh/ZqT593sTWCzPQqRsnD9jWb49katHsV8Dd5Gs9W+A45CTFPdNaijHvMIXy
U1GJUD3qEJ+G5lu5mf69OYoX1jLErsJVpsH8Os59i3Osmj+CtRGO4pyaF/tgOsrO
8Jy8jQ4dYk7Xaa/xLcMZFXjT/O4zwiqQgI4Hg+sZuv7k7yKY1Prb1tQRfe9vhWV+
Bz9zUhsSIW4AKaRyKQjt8QPlxPAKchINMLL66xoM+SztxsnqI3qCo50895vKZ25F
kVEEEIzkkjX0+XdB2dNV3X3DspQttegeR12B9n3T8/Tv0cVAR4KeCtzOm0VScfuu
lQ+TdV/xXSTcyeKjgXKrYZDygklThNY389J6aFbQk4g53+fVIZV3HiGZA/lmBNwZ
wUTAmVWvdBjh0P74fB9jS1NVoeNtxGOOjeGagmpyjaYQmB5sc0kFuMWcQhPazKYj
T8en6AEUeOkLehaqihy9uivL/yHaOBVSiPuXYjbrImAZAvS/ZqDIUQSP1QXtKM2K
eckKK+y1UkIX+cjzwwe4bfgVYfCh+QzsP145vFTla7CFJAm4BXKXu/yCWUL9Hdk+
xIBshwj4xNthhjJ/1Oq0DK71pt461NHsRwwo27yA/DSpWqK3AEeu82Pz70YH1NDT
Df+WXXOPz9geC7NdKZ7RIFxQ9fjZWXjOP+5gOxW9Lh2EH6lD92KOAihKWaxEa5Ry
0QtBJammGBFmUVF5DZp0gUij+DqY1COx5S5JwQJ6zLgeQgHdeMPqwEhI/U9hf8lb
tggjVN7EwabG4c7VAOzPawHrlad10poFs9fUKbpg1UuU3PMLXRU6sCYKUPETscEL
WgcKSZmf4ZSJgh4MGd7U7pyb/RlXkU8O/5fBzhLy5DBEGo9sW+sE3xAI3SjQ6eub
AVVo/dhksAM8Y/RW22NIEON1pTejQFDRrEwJw48hAIj/aIkXDSh5+JJ/IXsuyIZ1
b3nTXX4qIdMqMtDyhQao/LiRHsPriCj7VTN2k2w7KUdfZ4savQmnVtD9YuzfIyNz
bNn4EMIor2FIjhUFt8csHSyPT3kiesxYjkL6z03xd76F2/aoQY4FnJcQ8AjC8QT9
O3pv5AXdyLHjz53giVnfMelBca6N6w7qDAkiNuaC+0vtFYxIaFkPH/aN9XgHkStF
0dYpfukR2ES6pjKC2+YUMBPYdMGPqsdQTTA6FQSNtzFupUPSf6OJHFGzXNGCs1CH
Rw4vryJ1SFYeNSteFiNAXkpDXiboYcTtRtcETguiAwj7zvhJWt4rUZ13+nkkv2Y6
YesHMyTahkrHGO2Y3zw2GNlgleaYNSSN6iKOvJKkUCqa4h50BJmvxZ9wSGrot0DH
rPfxb5jgCTnOFEpgHE8vD2M8W1oi0rw8P5c5RNWSZP+zvIPBj+9j42KR7T1/zhXw
iYO2E8W/Qxdiqr9QKNtL0MHgNN1Le5Iw1Qx38lHoxIfkxdFD0EPx4uHl4dxVEm2S
SHvnP0adv36+WUbr0athDpX49eXbm66yFmhcGbPtGawEt53BqY1CDy/0kTvQDgJ2
mD36ixBCKusXVt89lsRRhHUEdIORUHTeb3TVD3UKDcHpplvZkmr7QmrWgm10z4gY
vUc68DL4QeLGYsZTED4EY2Xxucy/0YCVB/1RBa+uE+e5Wyuhy/4pxqfXSkzo6cNc
jkRwghHhWCGxZwLcrry3ewqDJZ6uGIiKEPlrP7bSeahs5rYWyeC3BgZYQW+Izu5W
4i1woqdHT2rGzCZe/gFMmiis6wA3z2f+8HvltKTjc63cX6ZouemFNGOQ+JTagUUG
tZNED2+cgjE/SpUJED5UsTnTZBIiUJGExMfArvsbRJiOu5ujTM5NaalByd+bcXzA
Y0gUji5opB+26mIQ/66fejJTxc8cQT/ousTrs8luOoKDlc8xxOmUaNJYvXN/Kcte
L394wBVlGYrWDBHnsisQL6Vfs2xsZusVwX0FAPGJwlvtN14mwIO6a7m0pLe9rB5P
rD1PPvELfyFjf4ww48MyknT7gOt6YimpoAsi5fiFwJBkOTODRjo1rhZRUOSelO91
yU3bGB7fua2dCNsA3og2ZXTKOSyDFZOdEuYLtBT80zHnVGEbsNV4hUQmJWYpdXUx
KV4vCWa8+vzNIAL/N9NaDZmRrve/LMPd3OALm+j109pyq+2Lr+dGWHT9I0YifYrJ
O85CcGCcLNbXUsEoQiSXTOAagjAKtPHYTi/vZna0n3zuUSz2TOpt4FQJhIBvZcJr
BbZcegUsXLkgiR6/M2Jc57Toltu0f1SSbtM5rYLlDgcULa0bSYXKyIgDEf7aWsoa
MCBtl7zblZnaOdQiUusV5Th8hAokddPKbAWKWxhR2lLYpTVsIrhyqh0NPRmnV+u0
IIO01+G6Yi0kiqrcjjk4LahTuh8SFVl7pN8pgMYG6U+xtHojIn/WP4jQXw6dK+LC
Uv/mDiPvACBoqBRa9Evzvl0SELRNVZguMFh5mBGuPQEjIfGOBEW4Eqm47bzSOCoB
KgBUo1rKbMhIJDaTQiNYXWqE8hBZUIwRgtiCUnCK+q8xq9Nhy3UUx99Ye5xypkHP
chQxNfJtLP0IpfaDgvITapg6xDE3M3peoebZHZB/gEbMVRRqgxpJmaJRFIvtvyre
QwZz6eIY55mbvKV/PN0bP/V7VadvIVmASl8JmYubfKez0lqcORxA8jOPq+ZqHxkO
hSQHUQYz3oR7VYNRtFJP1q1obcwAUnaMgMBw7QUGl7zpKWOQ0fasflWHQheN1G3n
l4LTnBUPH1FnAMxC7dLQX+PWf4TOwiVk33+xAYtq8ZuDxzWRvR9VHp42Nixad/mr
ubUxQR7IT7UuI6uOj3yjoSfFUHv+5CXmox6lW8f88Z7ysYWRQXDtXhtuYNt0FQPk
lkrKHcIuq46QX/vi5fNt2eT9jjOxEE45CZ0kzQucBEmWPpuMNa7uKDca+TqdYdvk
t5oM56uXyoKLN+2ihDPSTrnIQgS43Ac/aM0a3OZZFTayaJSvJWrIbHXs87ThQT9g
6arv+TBr9BMYspqLoghBfiUTUG+eU0VImMrzC6Z2aZG7g6pm/T3zyTIp6h+FbgkJ
ZVn0yWPg5kYifdh3OLDzcIytRrWLv6vKvgF6g9bEiujzfrQyoOKcl3VH3XRU2aVR
FzuBGQYb8oQ05pETOovToJmRowqlk46pbrckZ6w0DDbFpO0+TDnSwZfbAeMVbs+q
kBsqBSnoNbP/EtYZS2ivWZK3o637dtFUiu1kjW5VBBwNKAlaPgvmT2I7ik4JR0H7
a8xB3/fsG2b6/WRVR7IyRQEpZpfj4twjaNKHZTKcgi2P7rfz22dOu/3pANpSUq/g
CLh0N4JcwQqE6EH4A7oHuaQtx5rD/8X8ydfMA/bnCo8EaYyJm++UQyYat1ZDCmt4
3Btkgx9+YQj2kTnOlf+dDhxbyPMIDgQNsEu+YxW4M7ICY9cUKX+/UaW9IqeDBL7T
LkSMHCsUy335WLduP6qz0RYapgBws41PX9CjK1xW0zbbNJWLwACMHEnzDn4RVD/a
ZU48aLvG/VeQt9Jqy53IUa18k2c2nYnKe/l2x1n4NlDVCF8DEWs5HTK1EEDY82/5
UbKjrMHP0ymiE65KuVFnzEVGmGYEP3Esx3xHk9xicP4qM8fpqxmNW1RDPU4rKEys
BYuGd82cbhijSYPoegmpsGwNQLv/nLLmVq/A0VW7HSaACxsSar3c5lGIfbYbG2gh
r9O31ByCU9eP2Ytrs+6muHSi+dVAzD2blHo4erLnfD11pfjl2kYAF2lK6c0UuFlz
CNS3ni6JdpVH5Ik3qwk8TbVsmA+YAk8J8lZib+ODix4o2JF3xwKoyyfitPQoELkg
OZKS6mLxkhWSeSYvyF50gs+8bTth4UYrr6dDJ4dX6jzRfE2PBDkNRxDL7kzpNhAP
I0qt/TcWAIicxXuQckW4jj/VPWYCHwJ1G8SpVgWE9qFUNxc2fAnOlbLJWLTMZ1Ys
sLZa7hcDewcVoMBUp9VoIzsrfJHf6JghgBi/lK9eZFEZXj702mYWu/QigmY2psa3
yLLEw81PvJDwIc6GWDLSdngMd7ym8/72ukd2m0ZqeE0txzsmHVUWM+xtkhHmMMOf
7yN3JDa+aDOM+92plryCPsKRMjp61eBY5v4quTPlOyZlAr6GmRPTCGfF9nw7wf6n
q1bcQOQCrzZauxrEz/xNbOqtiQIFLuDS66dH8H8COmJLitd7edps0KXkAodSUmAk
NIvwb4GC+YwWWwIZwblaHPWmBetg5igIqBZ6NuwbWA7+8RMPtq7scsM5KgfpiTUs
TewrPWNjP/oMJN1EZoQGaDP/we5lfBg0vqgbvtQ4cia1vR7h/MFbM7W3z5/+Icyl
9Q0YR9HK0Fo2yjotC5WjGSILI/hY5OsyDB8/dXvF9jMrqu6sjnuJQEozzkQAA4zN
huhE4zllJFW1Qog2yi2VZ5InmWpVS81qRbyl/n7wLBy0X/pcrulqZA2IYqo7Ln9S
I9lxe1f7Z/RDMUpPpox6hVP9tYwBGpI95P+pCyYRdV03/4c0htiL4hMmcHlnT3LP
PdF6Ucq6NWRb8EEWQNfKdWItBtBUOacLUszhxl06E2d25uuftGTh1SulwsZiHyDK
PqLYvesDC97KepqtF9vxuuU7oReFH0DeCwUXTXjlEXJX9le62H3WDEGdJ4SG2wdg
LsJiYXRPZzNhRKWl7AQr7ANbmkm6sWdnPc2c3kAgsNc/u5/eaD3Jrea+CZ8f9syA
zuuKL3omWDtvWEogyfpf2Kb4w+lkhLi/eLYiaRMyOd6t9LeGx8ciQQs9p+HxCd9K
Sc5F68N4fBbPYmu8OTggbu+2w5jiLmPGn8tTzmqzOVnQQOx7zrKNYaDzjrpqQQRE
7yGsXGtQzj+RJkBodf7T64jhFGCUAMhGZCZVIHUm3Us4rbmRoiPwHz8B+MwNMidl
xBAuxVbL7BgOyBIaCrbQsobWnibHsDZxv/z6Z1iz5YwOFrYX0gioNn6QfhR66/HB
7PGTefENOS/6TxIMSeX6rkQbSZXnma5FTK7THBaSG5IFfVqa4GatEGwVgSW94SUc
/Lp5B82ft7N/scCHY4Cnxcak+yaQ8UoS8fiKGH5PSYcMISD3dkDgXBMj6SDhYFOi
t2rZrPzNeixbGhCnXM+icie960LiZUjy21oUTKWzP9iSuZeg3N+5/2KOx6O4aTTR
RBC54/bV4eWx6Qypm5RGJqplM/BGrFvdLxSx1WBu2fm3JdW11ZOy1+hgHlHdXh6e
XcyB5U27xOTb7Q9c+uQ2W+WFYNK41qLT5FzYWGzu2q5qagvuGZbYdhrmiD6t3+Zc
IQVyW3in5/PzVBv17aZfy56AV47gsGAClggKU+I0sePZMcvZ6/oLSaE91y2gVgto
TpUWhFDG84szco1Qzf0LyhJ2nJNu8WCPp8/6iAqRUMOQmfsVjx7Kj6AUKjzDSGHd
+pbQ7sTD0VnazuD6Y0l/DYJWypfJ3LlZfxFA0SvCCgnr5q66CTpaiZR61/W3DSwj
w25Yw27pNxVnlTN1Kypl4rJ5rbP3hZJ9Wcis5dg9EhODCb4OlUCn+Sp4NcYF3xoq
8mwZJ1rAEAxlS/KZSy1D98OzNzzmvCtNchMl6BTwGVe1ECLMc7O6CGCyHBPBstt1
WDNjZidEa/e6CARlI0G6EUl6yTjZNupkHkdI5zQUp+erpKVQmSZu7uGshCt/a2a2
4rwp4eeDNZKkzXE5EQxn/fHfwnEuqlhaJFEd/6MrGdX+g3bNv5s0mAaHLvViqHzP
gvKRA1fn89sJ+qv7ZPAiCxJ3Y93rRRBLtEQ7B3YL0k8yC7UmUiZI9y7lCwyqGsxs
8QwWkjsXs7ZmTZDTkDnjejmMU/90on7TYZR0laEprgWRIm5dpeI+eyv5CBr+W3ce
Q+3VQj58O5UgPbv5VaPJeYP3aL+pYZrcoZNoGHskeuFTJkni7cI7DR6dXtcV5vhX
OV+8KKEjEgrZY8e1/sjWg5xMS5VQIAvB5HoIsV/LukKd9Wd+RHEFg3LjgnawLDPV
Qd3q1cjyNZsVJh5jwLJXg1RrawJLKmxugDyqIJrmBvmUGoFk4697mE67xH4gn/d+
OF3Vn6aetxUCurfKFEEcG5W8+NQgJRv+ywWRNeN2ceO0gl/iqX9wrcjWchO84Zju
oeHwu6v4NeO9pGr2Iw7tI5cvR16l1yLl1NpuQzAhPdNlAYav4VwQwOqmgbLCIrAj
elXBowzEJDCF3ir7blOwTenxFPFmnC1q985DGa9akcLPrpt5cpnqII33G8Fnkliu
BYJ2h5sMH6E+tjFSA4syiNQci2Fh0HBrcN8S8qYJznU3qd4sgjZms5frmHDc5i2l
Mm9+W5HPT5kP1awtquFt0BLXCbjyOA5K1j0dn1JaPV2kqWMtrt1QBSMy5nMzCaX6
TAvqs/fNWOGUqfgHeV+Klb0/jnO28oN3qvQP+6BcugbowmTVirKndCX6/Qc5GsMp
iGLIA8IzxvQNZ0sQjAkPbrv19SyXB+Wy17cs4ONpU1O20SK3tP0JJnm4R6a6Fh0G
gVZSJRZ0NiAg7IR2Vn3obpt5ueB5YmjIKd2+/comWWz9fU9ePevluavfIx5KMX0a
85fqoiG5XOpELNKk66tdMm62pNIZ1QTDIVzoNDd1pDHISv2tAmUHoPjsVvzDZnXL
1XYNiwnsEfgDyjw9EozYBJcEuPuSQnlmaAfVufE/PrHxB+SmeavreTjkMi7Gc7d6
2BxR6xRUUdyPV3Rn9lmFt/h3pyTQr6RkBmtrln30sjT7Nx18DLwFDIeQw/Y/1Wtd
nAvM23n26WoAFZHF6MpGkD66nx6P2PoYu8VHRVI2lTekSo8ivLkCHqafTz0yDfIi
pLUGEF1mV+yHFW/Iiwjdj9jGs5qqmTzZ/2rQvUoWowMSG/7bGIw5e8wzNa9d3PAA
EvyXvv4xHs3maJ8wDxtCa87I1VQ84tmZ5ZMbRysLQFGD29eHQygqUFydDv/6TR8R
HDYjfEqPFhY0C9jncD3DloY5yKIBmqolKvVYLzDkMose04+Y6OQ4PXZ7ZRagO++o
UPufhfeNT/f7etMO4UYDjvgTcQL50kDgYhziCEZ5P2tzkL0A8KK36igqxPP+X/7g
FI2jlfP7l0l/lgW0Pk+vIeVbPBHHj9O0fj131975TYuusBTR9SavSLOTLuQidfo+
F9hXGjeKS0n2ZNgifcWRkpfcIVH7lBiOarbik/620TsMMX9ds7mii1+4Qob4VdZ0
oMm7oSXKiApAMYrKow5LOYn2ZUkRo2U9LMeK1diLgHL4x3tYJOSFR2x/S2OHtufu
/qujiK0PqTYjFNCfHLn0zAQ1U5GzouHlmQi9JUd/QHvjNkKsIewbSOozfUVuixwN
MR5YwThKvbxzusaUHZl5Qj3sxjK4ulYR6WF8V3YuIxh0D1y4YR79DiTuYKGJWw4y
SVH8KTW4n/uoHK7WaWSvjeUST2hYLrhz3/kdnCmw/bz1YUFKfxiBkVTWw5+yn/K1
0WmrbhmG7b1lO1H4ZjxgFk8JQU+HC8TE6yIXiPJ5ogeU4Ynq3hYfH+LL8nOelorB
1y5MlRy8C0t5po1ji+rbjOzSq+PuIzqMDeKtC/TX+ql/QjoZ95EVj2HF/qeEQWE1
faYWa6A9zWdVbhkz1EzRgbhOlIswj9MVssx2sfxCZYAuLm30kugGz3tDgEhizJj2
kb3m4lLEf1jKuih8m3TnqIboQ7c0nT+FxGXUqduvP3c=
`protect END_PROTECTED