-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
ZbE4OWcusoUuuagyi3Fb1P4c15RJ3Ma98+w9MoYI/xzcyM10jewaGZjYQSJ+PG4+9KRIsU9EYU6r
SteuoMl1UV9RniVXhk3JfLljKq1flKUstVQrSWyKNHRDJE368tRC/USj/YV405a69V2ibsSOknwo
sZhGYRP8zj1JUPqetKzyTHrmpmmgUIAPyxI0ouK8CgL2zjIdxfjLEZ5HgKh0vle6FunqHqYa9vbA
lhuDIrfBe+W7RcOtTshncyc39Ekb0ZJD/FxQ22d01IVyKbLV51XjVgzndULfmcGNAgywnZhBmzZ5
NuTBL3hk2PhvRTWcSZEn+Yiyi/EEpQowDZCMMw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9872)
`protect data_block
9LxQzgWiu7YWTGuDvMYdNIgGQwP9KVibg5bTabm9jpdhkXPu3YRW0+rYRvsRcmA5lsnVBgQL0eXO
wD9/Rh6swkwBiOikJz7aiWCOborvQL3xEqBS2xcDkhfq4k3yMrbOAnQ8XQ9s7YuUp3AOgUwjVO1I
rl9vfncZZXj5atTAXfBtIwptn7B4SXqbTawxjezPTqbZrOO0r4mva165gVqsmZ84Eb3bY/CRpVSn
jbwzM6nVYj1ufbeWIqwQPbTsZ01rZ9RwIqu/0IBNf5sXab3t2Di+oArUr8t5JF9Y2DxOoi0IiMw7
XCR1aFgrR5kKbZKwuMDoaz9n9N3AyY399ZeWKNHINPVIAXqL4Gv/k3mhyJElId+t5hcFdIoAzxfr
qLybMVQf1o/aFvniUdQG6CDfXqLWa36xEv9I6djQzINge1g5cFnHj+6vX+dox8ds2C8LD5nRBpkK
ggWu01p4ZifQa46KRpEavNkQP4/Ty5OYQtyAnLpXTrdZOw6N33KckQylAE2uhSP6tIv2SnQ0MgwM
kRKkRWApH5YWKneX7I/ldLESd7paWt8LDreni8f5aHPGyM3s7DNWGMf7imkJTU6t5dco2eqg7B8P
2ArBD/ep/xUJW5SsxiFzzaX4HjBOpQp51ectoCGdYSj8MWuscdAkF8A7ev7xQtckGGkn3wr6U0wy
cfsvi4e5mqeAD59tLJwzmnq+e3InE7sRAiarkINygVIl7YQ337+oxbGKgrcsXwd+8KcJyHwBcqSP
NjWnubqWwU3pCef/2FxMHjUae0oIkDuJK08zgJ1abtruSVVet0M81Qc5ioskqDOrCiXsu4fEwD/Y
i5YplMLPq/T/zyQaJ8yge+c8pTa/mrxokZGu0a0YvcbltAEB3sefNBf7ZAFIhGHMNZmtCuBbLGoU
hzTzDfC2XEesNUR3GIQ0zWjyssbGY9cTCLCCWvYCM0XawbAAyq3yUPu+tE9toN36od4XBeQLPRVy
wUt+832sVB93r1Yhx39S9Dxr5V/0szO0KoxgF4HXjf39+lWmrCYkaK3OLWiy88SwuVmDsNa4fQzR
1IAOhFIUprYC9NbhAFbUpIEKOlVFSN2nrKd89x7CvBMxogZwokDwu7ofp10u61N54QFOn+hn0M3q
3BWg4RAixQ0FnI6WcFJchDpG3kGivkq8+ZxixIbfFUh6+t7Tnq5WwD8YYM71HhXn1vlGV8NJYX/P
GpayNYZGbo44QPVSvxSOJSGdqFwMvzRTWyXDzfYAxpNT8iqXnMbMOcJSUhjc72qakGbSf7lm3SE6
W6/qT3uoG/mQTd+u8uOMJoftrxgUMeYtX68oBtRL9xRNDu8CNKWwJXT37RSvh8sG/SsVrM2bUj4I
3zd73UHIV6y3hUyxDabmxRaZINSOL4bMtftEFwkHGZ8hwApPDtLOZXSK0got20MaZ37VScuG1c41
V01IsWDHYjjjILluNF7eYPczj7VrJOL4eIUuYqEkfxOcIzd2f2l4ExzkR0WlC49iA8Fj1Aj+/AYV
ykLMAMEcYO18uEwmGtLe+up8CTxHbfPSluInwvvRoqb60tyuWIeQW86ElowmKNjWfibj4j44gT3q
IKEZFEnVpNNR7ygHkNYsrss+9teSvr27VmbsObXSsBgWHMlNaXgs86PofvLr/+5BorgQe8ftmoYe
jgEApNSnQJf38klNhEcsj8xq4hVgu4TLKetkHi4aKbNxwpY7ignH6a35jUr5vmok5vH01/vIM5Ab
9nIagjgZQzNjFvZOAkxJryiX9NsxWs5uM6yYuFK/ogeQXGE+l58uArHWLLHhwZRtqBAU95sJw5Ci
Nn6JnTS66uGwiTIORXGkS4aQOeORkkQZFJZLfHdlnOH9Wtv9VLkayjEdAxViXWZF5ktigLWoFJyP
+548pJvc2/zCEfFuknZFeL3GsSyYmcdXJXzEpsEpFt2pYQ2b1gsPqrI7b9Ube9zeTE6GAILyxZFL
+94/WH3OF53YyZ4N//JYYKqKMcdbcYxipqZMpsj+QGPT/Rh9p+N+GjV77OXMKstBdzHkWDNK+QNE
yJsxwOmsqBEWfDjp5++jDSXlUn2HNrCvCOoesmwkNpTGpYFBY5K4tc5F/JGmBFU7GzQx1NyfuI3n
0Mzdnv/pb65AJ3kIjrJm42gH8lG4J/ozMYpGDH+CQ/tz097GbSEhDomdYdwjJAj4CcXmULU+LID1
pDsXqmfqe3FlLpxBEYEjNmyLWYF9xcxOWBM6H55Sv7pgzX/8ZOosWgmMU1z01TCnOBgiGx7bvnPj
oXyXWglVcUIu8W/58Gq5h9Jlvj8gLfBldadGWsVYDTYx8XhvkJ3YmKePu0OJNEN66cl5oI/za4zz
u/ZAznRp8lOGNUpjJZqbvWKR9XSE9kBz8kLPrt5D6dqcI/Do1rAnaYxfdfYR2S4czdFf+2slcj+9
El3xfMWNa4HFN+WBaJxTkwwY7P+RPwQ/IOZQpi4UH+6+euUT6UyLQNESUUsZCq2RNObv+R1gVMRp
REVH7LCwHZ+T4PDqZ5oFSpHkG8p8AGiv8qurRE22LsWMed+hqQ4H9N55HtvZZJZIzQYqZzE3uhIN
DwZ+lLvibhjq2+C1QcZNF7sPxEQriaJhMAFOw3J4LLLtWgpu2PfIoYA9/Sbp3z7gI6Y4Wq+7HC7A
2o0o63mDoi/tej/AnVrZ8f4j884YmHHjNCFeSdGjdLm5J92mvxlch9DQXxZ1/Zb3lhxA/bvkw6Yh
mhRpvN+ml/5PhHIygF2LdH2VC5gjuoZD+kvV/NSpzu06+pkFDwV18b/6xwJW77Gxk9BpF+d3Damq
UFTZi7Axf6H6VM2b5n5dVWjLbhrrwWNStfPyFBUNS830hwacn+cLpDwa4FQDh3iS5Ay1bwgh7yv/
g9GN2siW7gMOctIY9aDhb3SHVkRyeeGUAJcd4tTewBy8pPfvjWnuLzm940rGd1obtOWwm5XHyoKJ
MMdSfkZhCAZCOIyd094qggF34oU9bQicStkxOB+xJoIZ1mr/hL4TDeMOhqCjKy4/HR+Sb0535uWD
URCNfDuvdtj0AD7kX8e4kmF0s3xAjKPNmIM9heBWcIXEVfsZEOJU3hpfm31ymVLxMopGqULT4Z6/
LmWASy7uWUxNCHFRE81Wu1WlIXCkawo3dxs7tJamfe2PGDVdcfycMXZVfGbVksMxENdv7hLiyoql
G17NcGbboGOxKdU0hKtEUUKmJluykDQNTm/nqtUkBhGFrc5SGl4bWryg6wlFose4SxsSbCHNlLTj
wZPUdEeL5DEABdpSgc90C9UaNBbRdD+eGzeXm+81cs6UHAGLcvaH3WsOO0yUxM7AbkXpKq3uUWrh
5E8CneR834WSPtXrIWo4XY1xOUVN5+5l2NsQp6gf4En5w0044olCIENUS/VkT5e+cTdhDqwJyX5X
sv0H8oBSw7w6nBjLWByKNi23920+pdY8ffIce4n+JSLunOImdBhWvK3CwDDzrWb8uAQPsCBik85o
JIA7m/O4XS8tAiLTc8gDKbamcMW64Gn5vg2yC0eQHQk0IQk7mYbzZdsv5uLKGi7Ozg0wknIzJ4ns
bT7W4dpLqJz9Gt+ZVlUb/s2nxruRLodXNHDPCiH+4ruri60BDND4PVFDivPhrEgRjYMDS+ojSaD1
a2Glzrtw3FpKdOtpZAj6dWMEdu74twPDblcDCPJfPJzkVkJAplDJvL40SOJ9yI5uyaIxnf9zK0A4
dkJXMlv9CI2B4M9GLytqJu5p222Qcdb5FvqzbKyUvNAfz/U8f57Ulz4IzIFQWCAYSN61BUEmBRR4
+L/tCoiFvDS0L0FjUNEFMNRyNviSKY4eiFNPO7j2cPfHDedCbykUevYT8Szp3XhY18in4fRwgPxs
fO24MMx4xWI2jpxcVkm7/czHXoZVl/M5RzO555hwhW+NU+sNCbJqK3TeLY+K2TDSuyxkLIbOtS6s
qyVzqB2epP+535cQUmizpwWU3lG6JzpTSiMoxlDkscADDmSdGneeg6ELIze93Ten1p9GOWaqvNaQ
SyTysanL5gJ0Q6qdPak+rQzuD2cA8L1q1RXpHFzxNcdHroE8ilNMgqj2Uq8ph1PE+UIXPh9LZC9K
uKsU8q4Fv6P9Ehfwmds9Df9IFfh+hpjbaQrmkBZYH9aqsm2TBlIECYVdPPstfrwgoa8A2Ao8lilW
6FbD9sjFm9SEaVFsjnS76i3+CYDOZvKabnyrprudF5Jf9hANs7UdlN4bxTeMajirrm2cpLe2mr/h
Sd8C7u44Cjd/9mJEbA8v+Q2gts6Ncc3jXmeNSqqGY7D8tcLih3sL7kh3t+hr3FagYeZ9MQi75R2g
QMYFO10Efmig80w+Krql7CqiLGHKupo0E5/QZWs6ckQCg3vWu7QYL3VBMzxQzJHaue8kvL8xE3hG
1Ynre4VlpSdn5KWDKdKEP2iNtEr7xcewf4ccD8BZboqYF4ZTCDADU1DnRmsZSB//Ce9bkX368qBS
TwECewzXU7OXOXkb2NYe0PLP5uB/AQ4nOf6ZPVi0CrXQc9bgfSzBJXygGz6UE2ChYZAvcc7hfD/9
DWjd2kdxoBADimNSwbr+/Z/BeAO3mDDfNc0iHSs01xu99F9Ng0FOG6GR2vEYa2bmAzziaUuEEExv
HBUsdTD14nbQWu7ytobc2p93Q0U2xMCPBf+1DB75vHGWYiUTaXBHOkJXwOb5V3TysP9Jk2t39utF
SQIMkczpXA2fHE09NNqBuT54CunMKC5xY900XWFB+9L2JgduXDvl2J3PfEYRvH80F0/vIN9wSQr/
CC4TR269mVAIySchXGRuRdvIVmcTdJmTWklH/YKhmDuh+kiKPdnlKvKqrS+iZYQ/5rVWQcWjJe44
XRNbccAMTeAz2OTfvuSZ1QftX9E0Tjhp2V94fSL3gAmXCwAOiEk5xmJHMrDdkgOy007PcxFUHl6e
YQV2UepS9GYRp8/d9nGDwzV1Md+FeXjTJu2W6Ag/RgR2IlZ68jvYAx/0lRsxfOwk2T+Fo06FCRjJ
8tRaPUmYjRUpIZxmDXMgg6V4hgZ73d5p3NLb//p5Hb6bC3XA9nfJg9rwCVrmv+K3krXSPCnZwP/x
0yQdUViC/RPHvNNQoMttHgv/WOEBhIxSbruiHu1yymxCy8PWdZvlzu1MHJAu7++BkHaB0t81j0Ar
/vvPgFVzN1KN99iHnqOvBvC1m+PFylkcB8yvj0jSpOQIN83HRmd9odDIrSyq9NWRXA4oFWfGXPzZ
9HuVhkE+EOXseW/I9Is6Ww2iafLPde71Ai6wI5kdKUBI6vMdWrcO8+YaZQ0kNSJGZLZwB0fRtx7z
MdAiHwMYHsrFCXzychz5GzBEyeRQFVHsQ3Au0/kQ5d29eBHGBYH4FuaXUYhQjC/gVCVst9RE9eVD
qWgpYkJhWCun6lT/nYQDk4CvWapGL9lriNmFS5FZZb1RVhZckDWke62DAvJlJJrWvYCzGBRvPOd6
LztYioA0PjbLk+r2NZlCYbJX/RuBK/0mvvXeEo0Fs/OsKhfLbyaAikTlkoFcViEwqzLtjjfwiqFY
1PJdbPHr+lLH4Fqvq2MXFlglCHYhaJ2+e/JaVHgzI6A98+Vwhu/wQx4sSXGWDhMIvF55lp46cj77
YDIsKlz9+RTKnU5g40oQGosL3DnSR7jEU6tHhG4OzGXd60V0Y7Mly0OP/8ToHeNeXyfWJQaXL/iX
j1tvkXytysvBibTS63CsJ5sTlNEA+M1+RBnEF7Xj+7bRVrpgfx7o+Kp71wLIoN73tRUm5w2gXdpH
v4SkHwl0NLMTWffiNgY4XFK8vE2IVaYZz0icYB8ttnh6putb//9dF1SwYU935HWxpfF3D3BzxmBC
QGkp1D6gPq4j6hGVzciViipvZ8bY23UmFZoAwMqjlyHhNKP/y6LVHh/mEkPjMILWk0qKgYreF+5K
8IsFFU9h2Tt78hvnUAkr0C9uMnrEbB79PRZeiv1DucmYk1IUbn4N3t2+uHc4+lFsjXvKV+EadrRI
I37iGa9g1fpzDIELRmHoRVfDwszTZDqYazxqq4Mr/m/kfZiZzFvPWniplJip8b86Q+zQTBud/eEl
X9zd3j5egH+FxWpH1UuegxWMBD4+bQ2HqF8N2BUH4ksPS1NbPLP3+XSWia5mqdth+wQY3NWR24OI
YWXjHLZ24BwgwJ1zpyTrAKmqmn/xXockGBkiLNAgINVR/WjbBqiwHstb9Vf+/l49Se9pmw2fk+qO
Do74SpWTnwwgNlpJVFNZBCJsH8iDPcm/Lg9OnMstUuKCtBcCfxUEIA1oAzV/m+q0M5Ix05wIfITu
NAwhs86eNVgL0s/DOJpgbIuKPd7aiaIdFpHhzZcEApRP5Bk/Rwv41wkbvacjfiqx34JYWVHwLmc4
8gfus6b/BJLR64lURHXITltht00VKMsrXMys8vv/1H/EM6vCwGvj3HuCe3RoNsmcMDffTMt57WnR
g5sZW1g4rQiNdfmW7N6hn/0QcBfU8BK7QqZei8F79zy68g4U2TC8jxUmf2Vwl0GNRpiU7QsPnezp
jzrURz5DCNmPWmfCwVg8DKUESqmDzDDFun4r5MsicyS4GfiDNyDxpG+eIKjbrUv9uf0aP5yhmqgZ
mjL0K0j92K2VfVAVU4Zzyb1xudpo/p+9SiFQI6xbJgkcdqk1TxM8g6kLqGmjEotws5Zp+BT1P7VR
kRxL7ACeZ8WK9ne0B3/faW70FFjvsT6qq9aKpOMlYF3k0Y9naSE2O7IMBkjxgKuE9FzAuu2iM35i
LJOvnI6YP7IRwnueULM+OZvzbQzxoonoqnaxmsoSFcEEsOcg/WKWQRIK7YWsRiezaayt2Ds/zC15
zJ8s8vaWgpNl3YQI+/ddgKWKLyoZc76CPVUAQk4IVyXctX6V1aLVKiFSLQD0NmQURXvsZjejKaPC
sSlBR9LXSUdLvbWczDz1vBbHDM0DGyGWpoClnKqSPBmoSrun4Y9y6aWsT/rbQckAEfF7zqUSdKis
rUyhfeUM6j+Ano24VNlziUggi3pBop55hrYiziGH88+hOIDR8K9LGGyRtM1Az1A3A5XGWyoQbqq2
Wf2YhPZdEcjA3Ciou7dPlfgO01chYw/SHCde12F2fwG1JDd2eSV2xKJkJDZ+Dy8WkD35yFUqVzYQ
vfLyPy/m0u9e8vlEjXl8yAxwmns4Z0AN60h6/fRvGCIipeo9UIbsTZpk3iCjGlGEF/5vmp9L59PS
EKFkZ+HTLdlHxexb4Aj4gxridR+qwRtGBjan764Z5TXe/6772q+7AvMXClrRFb/8E8XLl5Sk2byW
dNNudDw1YUNPJ8orIgj3ZFqvZPsioAKfPdyTnMT7+Ab5bcEpUFHkYNNKW/G1QRPYHHX+RO3ewZZi
It634N6x7RP3Lju2fHVqw+XYU1Byco8xVRBs/DJonuNAMqHh4gGy0Ax/HjdH2zE+I7HM1w5+PB9I
fTy55pWEaxBFFZM2GzwD1+PzcInz5yZaDXgfc5kQsmM5l6uCcS/a1I+DbvUDrPTTjCDLQLplhjgi
YFbjUOxxktVUyAshvRYRf4zKLsBsCC2PZRNyOlC+6+hyXdxBpHRAO92ul6nvSbxAvcTmC8d4TTBj
uab3jyJzr4Hvzs2hQXDnbYUij9/Nw+eJpSZhL7qxLb3Fo1inSjILkIrAGwxXwn7okK6dZ0ZYsa5X
671Sx87zRt9LOWq/BPGHanjZlsAJS2zvIqsaa7oN8SPYNMDmJ14er0Vxsx1D3AoEDVHDbZGIgVxi
34L6eHgw0EiXONVQPDENpRUPkZu8aY8jOc0QqOgra7+It1AKXbsiu6dyaPGgs0yZWq42wkM1eXuK
O7KJetKjTx2wrETMZVTzkKfMiNlIp4SwhK+CFYV70UyTweDtoFG4kanQVS87pcnYM6RlVx6Agaxl
bNn9BBRmOVrKm8rXT5RfIGSBp1ceHM+LWtKksz0/U90aTPXHwqyloXbFAZpwnIq0+f784bX3cECL
tHtcF5uZ69ynrWH+f6dOgLLzV92W1lAyvhNIwL79nC1lkUuRzCkc8uIW0vKPDEv6SvY9jUoT5KQX
sRN09eDmsm2lsR3ouNuXVdtCUf/4CGBfIpQVr8jrsMJwE20ngxTYrd77PNBdSGcI/9wx50cznwSn
grgeX52WbFhHY9gApHDpTvBW7u7+pqUUU14CiTTebSng3ZD7nKbiJS+VHOBdGL7qtHLR9TKUgxrb
6xkLH/XogokFPjBIjKjPy64q4C80i3UaJXPv2V+JiTvMw0wrNhQRyl6b3c3R6T4JcdNWSKzXmGnp
5QRpwtx3itvvK2joirmSD/GdBdjFdDIAiRkMKJnZ6OifQXUbLyOIUmj++672yJcAH8psvowAMsYD
FJ5MjoEM0i3yATqjvX6xFDSjoq8PGf0pX/Af2TRM4kumh2+5o9LJBS0U0AwbKRrQl/anaif9sMTZ
7NRlcyCBo3wUeJvjjWo5lIXxBLypfuCb9zCsYtNFSqE6Bts+yovfOaZlnOshEIJBxNbWUaf0fmo+
kB5lmdbvt9mcRrdLKxDamC6VEe8djukk27Pii71rdjNdZ/LTeh3V7SB6b7eUAnY3aHTNKEPPphKP
faJxraYIlk8Mk0s9Izx8f1llPe50z9Mb/MTkMahV0ILyogj1O2U/YFEj1+N1ikgprZ6Uc6jce8rv
Oph5Q2vRoV55UJE6TB3ZjuRKMriYTqxk4a8I4yb3/HIo+/I0plfcn3q0YdQPkYVXD1at+Iz4wjuY
LY5MW22269Cgp1Ymhc6iM45hxWL4s6h2nddtyleDwpZmeoiD/ZAbSPvgQ7ZfzwzBC0Spl+j5At37
6JJeTVeRrRjafYyCh/i1MgikaI8kUJtLpJqw8M9XRLHJESnfcSmIp6SMEABLn9taqFiBrcUCMlcA
Yqqf2PO3wnLCRVTAsu69hE86cGcq77YFBnSx8FsZP/qkzjnYrv00399KGepya4hTrX/Dt0d3HCAT
FR/9dO4r33WNJdCx+/poeAlDWsRIVCpCph0HnlzOzAuPlV5mx5wfhJKwjEdktoFMZkWL8yivQziL
sa81EKdtwittt1JpYpisUmEaPxa0E7Gvvwbq7ACot3XYUzdvU8we8LFAzdjoqAZQbQ8Ne4fuXBMz
Rc1doAYM/gRIBh+ldWYRUwAhsVd4fx9nX2FWZwCUiJbrWGucIW6bqlwL4nEchrZAm5Vq2crhUMmK
p/PeVN9N+hNHWvY9PWaG0NcD6LFOaiqlVtsS+wZsL5Qrb210KeczY97XD+/Y4RqVza5uXih2a8ZV
aZjP6InoBpWhsYXRpLrWWdjXF355uZ1duTK54OzEHI6yZBoo6qQkuUxJQJ8PEJHKU0p6bLXyiujU
b3t7G3rn5eSOw0HBwJOAFcDZbj8J3XpAaKOfjctXXPDWsc2GNMCTF5tbruOw5A5QzqJqImszqVWn
TmWmgv/bmqsJOAG5q/r3J1wgLqkrN9oNxWGoYUzgEdjKitRuukZNzqG9yFZ/nUoKJSe7V2N9njIN
ekiGxkgNyAvYCeXTFGn+PDYErusJMjToxaDcyOt53yrcLlBTdqPIK8sk0nutjgnkE/busE+Wyvlb
SXIiR0pAPth5bB6abv3jpQIltqf2VuMS/qK/ZN8m39VQ3huVCeSLrlqY0ALi8Y9XJt2uKrvtJ8tz
6ktF1xe1snO0DNOWqtmwN5AMdFZsE/TMOUh/2QvHkXWhpvquEldBVGig1n18+NbbTltg0nqCxBUN
uZGSh1qzlF+HB2gV810D//088IdEVNowYUEiRJFR140IJIuR+tM8oGAqWWX3GqrKSDtJXRAhZ+Qo
SWbM7jp/7egydDAf5b5NHiGW6DEE+YbMR7fZxVV7LpLVhtzQ5d6YbW2RUBORAdq6sXEJQwg2Z9WF
PExh7A6Bxpma/h79UfeAdNLEqq5U2v4dASnMT6XSKs+4X72oD81VKY0T2yf5jcQAEzBIOe2POg51
YGALEiAh2bzsXXNqSGMePWpBsjHnY/9Q0OJsSE5aNwbqFRLkxxla85l/GuQuwrMJuA0z9T/8H40a
TaAxc+HZimwapxlIiWQj94wr916ru20FaSHiSY1PZgQg4YLWkF1tb4W+xliYbbFwAdDz4dkV5j8d
xpuI9X0zPK1GMCxUfBB6ESsETVMi4+dmM9ZCmXwXoIvyqauh/MUTdXvO6+GtzyazThcRHzsPOoDI
bMZGjJFMWIuH4F2uCgct0HJaGmhxDEwZdet790xOupyMQku7AwNNSek2t0lHvKm1jxaTGCYC1JgO
sC3HBkf0lM+b7yikOSIIWIvpENZyi+x6dVJfdzPiTTK0GDWKXq7TAVdyvYmIwdrs7cJKh1E72cfy
kggqSfscl4dU6hA0PH/3ZyjwyOY2wGHOZFR7gkXp4+KNWgrYgrQv9Lor0/xGr/dDwmDrHJhbBSe1
WMtEct+n6q9qVOWahg7mQja/AnJBbKfl4x7mhf81PLoO0NtIzCJPz2NKN8pujGXCVh0wHTqtjqjK
4Iop5nS9x76o5Xm+Olgjitqj8P80ugfU+4DfO3Yqo5VPvG5hj7tRXfs0zQwBWxCOcmIEEh1SGkJ/
F/TKmVUFqCU8kgeXMij/bOGm1j5kQ7b7CldKhRsJKLCt7+Jt8cIe+5IBl0PfaVdFHgAcZAdr8H7F
FKxqcBgJa9xs1yesS/0T+n/4YMqlqcBVALLz4FzP+ZSCHdXH+HAwsbpR9amWmIfE8ERkKU7zsTJ8
rYym+ynYymGznAxmvIEm81oxFdE8jhJXyFVeB7t3o9QHSqPzwb3PHTsjxvePOLiIzN/kbDgB2qT/
qZ/3t6aMzIRoUGfksOzH1N7DncYZR7Gx//qbnMwEzCWAoChrsJeR3MwENxsuwfC6Baj3qm8uGbG+
W0c4KR9dN5/dCijm7lLLWRmyLzo03CTPo0ijJv3ZtNlcebiEuZLPNd4uSNv4EajfTLNqEwqPXTOm
JYgjzBU8QKgCnXSH+lePd/o8XJAutvOiM4RHmHaLUiU+b6lIp6DZMSMbqX3aAn/OPrkHKpo3ABQe
hK172TeYkmYXWIAjWqUoN588gWKbb9Zd/lCkPY+Q6W/ptQjHCa+tY93tgySGTx1puMiN6FGtao/G
/JimuXq6/akPrwYCHhkDo7j2WXWLBtqanJz0PaZ1206KlVqPCnn+zIdJnt3SCnqbdV9Tvez/aJaj
qtMM86zCWTU2DSNRP+LaplUK8ezvq6D9KqROJ8AdN6ffxRD4Eb8S7H6v0gBZetydY3XQ6doFPcia
90Uv3VQrQssvgVb/hhgmX0bAWyalkpqKH/v/KBearywkG+Db3X3ZyjIA+IrVnqrfyt8kft6Wk8dz
KLqkRp9diHXuaE35xaYjLu5VxAtjHXigPpHUWq+LN9QqW8I/cuzs8JIKzdRjp6MQrXVszndY0uXr
GzlOfySM5R1Bv0wqHXaUW/N/gCHeGB0u+05L1nivpvrln+Asunw/NljrnzmIf77RaBOsnfySNEiK
v/OZlQBz3NIhRYwmNzpWmJayHuttivf+E/9cRAoQpQBUYEP0o/cO6kBAB7eSAmRgrmNtJuqiZdYU
5QS64xXeSV579OIt+d/G5aG7Og8PYf6KbJHIWUhNmK7Sw4jmU9RDUlMGXDo646whE0+QitPOtg/K
gwk3fqj5QBwDV77aX+qhEFk1xHVM4DZkhHRPA0wrzqsyqMdTBokOu/LMky8RvMc6oopQkdkNfn0A
SPy4v/6Au7kZVUm1MOW/HxOXJX6qCx7xHWIaFSvf6t4WKlh9MPoGyHcDZ1NK0czAo8kYFQhCZ6j3
i8MjBuG/7TFW1EfWjekGtzkEGw5TtBCLC5kWkKLV/mJnFL0Madk7MB9jzC7PVqZlBWPKtxQ9omIi
WVMVZyMeOIfrJX7JVWFKDvuFp406YvYDNYD/Y4uhCE/+bkyY2kPNbUKCI9X+PUeembxE5h6S6KSl
oYnRnVIKwU2gf+1IyaJGpY/JKinv8tcYPXyvF9xTfZlmzx6X6wwNM+b37Y1lidH0a53Hpr/tlwrK
qLuCpSR6xsBuaqlsZYcybUOYpz0Wgd4+9QTPp3VWQYshsmDDLsethvtCdKb6c0kn0np2gsbnfgfa
jMdu86N/+vxFv0UQKt5T7zoI+yvxH+JY6FhkOU1t5cuJmCh+T1lOiZqP1qT3ZRMLYU4DB5gaTos6
VydO1iN+hFKptTsLTbKXvfachA/+H4n+aQ+CvrHj8Ka7Un3vRqGqPGRvUVdfOUB4gMDVVLYjL/E7
Iln1vo5FPlyfHYQkdgfgIXkdizJgqtxgJMX92Yf7XO3HQwcX4T+B/b9VfTteS3ZHmhWDtAb2T3VU
1DAE0nSEWmZXuJzSYROWYnF/Gz82Pv+j/wUyB4dY2PAtRU5tSn+G4HR3X1QDTkd4t9Yv2zikPmWa
N6rKVvz6yvA2fyB9lUx2sVprKTxnL5KOn8jbfVV2UTQF3ER1MCYQNUSOL6JNss8k9PKSjgm9XYjS
E78n0E0d9yKU1BGr57mzdezkuwLA6WaLjXwPeC9J+Zg719UfR9qBDF2Vm2nk0veiQMRAq2zV3dfI
8BWeaZCV4iPYZU/BdnJKv7ZZbp2/6KlK7RWaUElha8RwA+I32EjznnBvxTXqo4vtLhqdHyoZ7JDh
1bDB/BCRNEH2cLs6pfTHrcSxbi5KIrRJj2yDkuvH3MFTLS368KVdGEJbgCtEL9050q3nT8JlQol6
W0vXSo47SC1McQBonVoPS5EFCwF9udGiLJAKLEmbCwbdd0RzU6TLPVLwa922r9AwIws43YanlBk/
rtf6CYUPo9qX7xqCmruBsbzYa6QYCDr0FklHT8OMmpN5cyb5WflII9SrmrHGJ0Rkw+UjRPC3b2JJ
+az8GPIMKrOg6pcw7PDdeoxGXom0yCzVfgRfHsSPkrFyXyV36uLUlXFpuVIAfNAgd2KQzZMWVPvN
q+g2lw+lGTLuN2NgVY+j4aeAicuyCTeUHRygCgqTWLY+sArBn7JwsRUckaBeoqJu3uGqcWqBTYnt
73nElD1ZAe+zTIc8Mp9oLHY5AoGnUmVzK7usvF5UxYp1hAD0d73J+wiIcOfChrSulZS+mMwSSoQj
j/CvEE0SvZiKyXLmBaGbHI44jTNs5punsnoVcjHjGGjUyaZ5wncuoA1/ayNXmSaXim/6QXROSmk/
bV37llzlFyq9dbk=
`protect end_protected
