-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
HzUedcYhr21k2I7avA96f1O6lpNAVAIqxG5SvzIve6lfHveo6uDwge/QJ6wOOdix
Q7k0SdCeIZdApIeIec6dtTJJ56UB4dsb/ErLL3gd4Tr1PxmWK2HKjS/eqAXYQjOn
QSlnZf8oRv1J9agUogrzrOq85L0IyCmCvToM3AZCFrLNrsoGyMfBNw==
--pragma protect end_key_block
--pragma protect digest_block
A9Loa+0X/m8abGIprv8GUsyG0+s=
--pragma protect end_digest_block
--pragma protect data_block
p7zzPBgQ+Jd1LimVs0cSmhY6uDHqPTz+7pDewzl2FKJvpT9Hv2Hmvs/hVMfrVv41
00tw5SR9YGIcRmd1mipCbb08WfezBjPXpcS2cG2oFaBnAAMQTvo7d9Gfe9bHaZZh
lpCVe3MPSsEAsLOfekuf7gDWsCbq5qn5x4wyjhCqboM+AEs7Q5FS2g9MGOKtWRxs
uGzETMIT5UUWTxz3sABPKTAH4D0z9A6plKCtezTJ2PUzd15E/iZNdrBednvO3fyF
Q81kK7SQnEjvf4xwzw1K/C/IP6eLolvzdA8LrnQVO2zarwzVpFadL40DbUdzfIuL
HjXShaVRh63zhOCzvu9kuGIzcUJLrImG+CW0MLfzf0eUimb3bRPtLVB2fCM7yy/9
kEff1VnIx6fLbahyTCwjwYhjtdMaVzFYrQcjnrOaezTqeimeZafGWCgRTAc61uU3
49UHrsdmZUsL08swp0Knb/MwoRzeUYqcBNpIdqiKWPsx0789nteCPYTem5EXrDTQ
SpGSeIYebVUa2RRMmO02Q4uxKw3qgg/CGEnMuOBREJ9ZVc0S3p8QCuksLGlupHuV
EPNg1g4/O57Bhqzg1UGs42hHYNQG6vf/mnUT+pPQYpA3pwXlV49z5LLDknSPg8y4
txrL6BXw2sSwNA1UdXdBDENEfNqEauwCVUq5aV3h9uEgxAUtaGt1ZHoxbnMdOLK8
3H/9jsgji585KbUNaQTkXlcJBlB1MzTbKqnQr5ujZqAVlazYBwX2eIOLFLPHV02G
Y8ul+zL0HNZ0l/I64n0Q1xJveDQmv97tC/o1khIdZEsgPwYK/fvcoArScoJWw/+a
zg0cthnQ6i1EMwGlWwIMrOWEn7oGP/jKLQj6hqZlLNlVvD3MmGiTL5bSJ3BWCM9g
AFkuZ3Zgz14cNvHZQu2XQ38uYvRLX0iRagLew0ig6I1nxIB5XQ5/OQL5lzjGPM/o
wJBZlFzKPBGuhfBFjU5y4SGAnNl9efgEJxv+ucSR7o9ax6FWEawRArpAEjOQ0BWr
fC0tKBovtCSWKl/ajdZ8zwMJ3LFNTfbM4ZHUwcrr7U0aWoH/CMgphUNYAwbXVAX9
0q5LIoOEz/vNGHuwazvMNBPLVM54LIkQ05PikhjnJxLj7V7hh61KJBih5D2QBaFc
LWJi2K72nmXy5/NPnxbOU35rq9wu9WfHh557j1ruYeHJWoCHNhdnzPjCiM4nzDE4
2L3DALh74mINUTLZYnmIOVQ7dNj8lbH/pj9aYRO5qGqdRgzf/e/MNrZYwN24e29b
PIBB7KCCA4n/tO5XxdvDDG43arp1QzcCiHXyMSeJNxx0DX1XaR/kwPp+/XcF57s8
AVyQmeKsl4CDptQi7aDBxB7dC31x8w1GRmWnVCLwMzy8j3KBIaU3SNC1fOWpkUtA
CleGVTIFRZHR7wEOV8q55uU5QNAfsTYIPGekgBLT8AUP6MSp0kajZrYcq9sHaMjg
HQWHR5hw8FwOHmC8DJ5BYEnptO+rydLDFPxJ+N10qFkiXub0d6KbPcu7mMfiEV2P
JbunfxTdGNaL0bF6c+phVp83BaIvsv6pkLpF3+4zzllod0DqcTE8vffdgJTT9Vik
so7uujOVSsq0JIhLu4yvH1vqx9R1Px0rD1dRu1hYlcWYHatlJPolV1Yd/BqNGdRj
LGH1Vbhn7MCCtN2br/5Ptn1M2vSJbs56U9rJUIVpTlGfwtftPsUMLDJdGqfL3EtO
2t8n2e/K/YgkDArn099q1N5ay1igPHxQGZugku03fUpgIo2zTH6xSf1caX5osdjG
oWjc1ftvIYYUhMgBEZObDOgJ3LYXhwF6HlO3orALEaPt3ehrV0CJhKVJvQKE/6pN
Mg0sn9YDZdTpxCK81XavzSM7pxlV/BEHo4Ap86yZ+RKBT/7yhdzu6iTrG97UCVJ1
M9lgCGub/x8k0Hy9GpPArYns8h5jBhIoFMLWqydfy0KGsfwbrANHt2RYoMkJ8U/g
gPrer3BBvxIgYCyJSe0SDRQNdqF/wDXCmFnhGFKCXimG9G/dKJ+XJGL08zuZPyN3
VpNolKNwDzirf/+kd8bXB7vOPep0BNXxW2k9AKeJJMIKS7Xm5fNsHaObMS/FH0a2
gMasjNOevbmGA7611Qh9eYyVOSIIkBGkasPEvhEdX2F6jnC7zTIGp7ZL9ZwcUSqt
V7izAWqBarWMxre5bSI6HRUIQ6QncWnNc0zcSLTXDl6APS1ct2KNcWyTt5NxD4jF
TWLBpd7MwzK+BCgUwkwI15rp6lyuPfn31bq8/XUPa3zRbUGFYC5QpvSm4V8oOMOJ
wNSm1VQREPuSGmItciLG8T+A7KWmEdY1ygrDDZaMfaV0dYhOwDbp+ImaCOQsL128
aZK7V1rB3qWYLM1wrBgm2boShUpwQIZwa35wLDJvyflV+4IXnIu2CvvACzOOQ5RI
/PDuLDEuHGocQOcCKMXtNlZL/sFlIDHuIjVIm9Ing4TCJMlL8W8WuWehLxpvmaYz
jHpaS7iKyrCfm8pRvzVHfjD3bzxsB/rB3CK0hP/UuButp2LSE1NUgBbxXUsrp1vV
Y9gZ7KT2Wxdw4xUz5P0F2SEFbMCZgBbBG9t2gyLg4bQB8exCglq40nHmW+qmWAh/
cyaTqQjYrGRDgRcuE3nvBIRA74vZDGJkYyLYCnUcoHKz8AptPocOH/7wya7ysVke
P768LtIwxkOAfBqNU9LuzDOyLylP8lS8rc85hCpU0PwfoKAiy7jvk0qCCoxbuzR+
y9p6lYXdVQbp24jWo6w+srmKgo023wvoDMTlU6G2uVDjUhfSxGPT1EyTQVMkZ4NN
yuFNzwCW+jV5Je0d30M1W9n/kcZcY0eGxO4PwXkZOBX5MHP5xhTjuC0zWb4RRM/6
45k8w9xxQeUJcF7pTNP26OdQKtibnvObNxCqYDP9Fqux4iURT2f9KHXEb9tH9zPo
wc4mcC5UKk59GjBceyZ7k0CSHEN669QFLOghsTdYzi8xSMnHJcdaqul2/v/QkCmj
6l2Sme86EA2andEd4Udhxlw4QvPNALwQrIIpYP9C7zSn1PN+vYzVS4iLQl8mTuuK
jwpbD+a7VkarB0Opd2sch5LGyP4/zzKqlW+YT0AEPbt8O8GnCFcA1CQ7UsrnWikq
UPuqzITwoCiFrWX7ihzxnJsmfL4bLeNpeAvYYgUTKH88aXVDvYp7GaVdRF37bMfU
AAXtyRKmIHhLdMW050NPzBOZVicktYW6Angn2pTB6FMqi4BQKkRnFhrAiPwtSccU
svgNi7e2O7CKxm/5jIOf2ngBxZDrXMdOwIn4jc+xqsGqvoT687ES2z/lC2EYV9z6
7a7+PQVwLJGxxiMsb2jvNJOoiBfsfQoC0n+sqaIl4aGzStaVxk1h4hyJANWlJ57Y
i5bAYNiZJF98tKUbW5BYqy4GAxSJ/EaFeReUxE14wAf74Qj/P7Y3TMJXPPqgcIuG
7DQ8eZHN/nC63EaFXjuDj5s2f6eYNtRoKxjHMQF2Yxqy8kjIe5A9QbMDGddvG0UN
woMUSDBNsTMgb/jWancoflk2t+nZ/mHBcd/7Qnv2K8uM8ntT29lfFI2ULXPfC2ev
ZqdIvpfHwov1Dt4FiKIpvuU0mzhJjSglt++eCsdORKciPJvdWclXs3lJBgveb/8r
xyyQ3eLXcdtMJoqrF7F8Rnw8zD+YoPj5TSbPXEwGjsio+HFqtE/hP77p1Qisenfy
oIMmuFI8zaXpx335whnpOvVgdaJtJCxMAOYybh0VBw3eCPWOat5XY6OOeGBD+MAb
vMFnAoTU0+oJ0d1K01MqM71w6P8oZyiCtk0dCGD0+kyjbc87q1gKc5pwY9ST5TzZ
jkpHxGjis4PukJwI9iWWxLkGRxn6+vfIvNB55P9pbl1HcjoNyNcPb2c3AkCTbTYe
WUgk9xHlpWiElY3mK5GD3gJggDoeKkvhC/18RRupr1vaUX35rvMWbmbzOgzniGJJ
BsFF3DZzwmKUsxIvcMSxA/xWLVf0a0vR3bqCHB7I0HIH5iLVMacjhwwWpCv0QiLH
dScsdAIJHxl4NRVyEMNyX1hfT4LIEA9NcKR8SjOeJ4R0bKF1pbrJxWnxi0IlvtqD
HUPixIGAEjnMEXTroyh7dIEc7Gy2PeUoZobn+FqKpVJvSNPevlzH/tzakZs/FrvM
UTcO+x3VDScgGOPQVbK+bcYNdC3hg4EcNLPZMKh+Oofqi3PexrYXabrlv5abn+Wg
Mjat4+9H49cnk41bwIOOksDLZnGct4KEimhLMiCzpsQctv82cQmvEvLhAOVknSHl
IGzZfrv+G7y4ku2fmho8VLwsN9Vl4jeYx0d2ifiq6yKqyBcZTbseElhCeK1m39Y4
9CqnJIMOrbmIX1EvMnvusBtAZu6tFJpeZVNpFxfasJi+nmuNyfa7bbpLm5AEAX6k
kqPbsfslhu9TwoFrddc56gRrSP4vKSFyCg2dlJKeAzNgrepVzTU1WNdQR3uzJSMI
kOBcYU6lO/vW34y5bo3xNKcc5QmfnEdwEadm4JXXKuJc+C+JoEx0ogf2Jt+g5JoU
SQpRZpYrQ6M2tHsloNudkehfpgLAWNJhkXQPIL1YY845ny4oXnWY+HazPucdkHfV
GKAxx0RVpRn2Nvsx9MdBkER426fcpF3TprdcWduILDdU8y3iLdDsRK2wDjs1VH7q
uTXY7n4yYoXHt8K/MKWz38KTGYJl5Yho1QGRr4SJb8Tu+kybk8JrCnNs8/AO3oii
jrYFnPfL+Ouhd54KH9lfP09ltHAchqZKEh4oxru/DHTp43vSnLJYhzVmdycLxck5
Y/r9yLKD+tZ+6TusIv8Vc3LU0WdSSSIRanR/IwtBcnnCjgNrVKDG+HgXA21IOmgX
gCpb6ii5BZQvLxuQDN6YNbIQu29omuvx3hQNU6uXqtfV8AngSPvAmLi1zsYhtM5J
nYWordYXxFHjeMgMsyuXe3xCIEBWN5rf1sr61fG2N9oLLiHatKmFc7ZOvpJRSG2X
uxJhQP2Rx7+WOjvzP+j5iesDqr0dzFe18bTo1UTAoTB40G3R+uzFtlOpHxtWgu0x
ZFrkEcw1Z6ek3sJzxQ/CI953rIMVbFgHvos2k9D9VIN0DzLgzwkx9hMdkQkqg0ev
A+uIMj6SKfySmo6Vv/b/oFZ2Kz2tMRQl56YRblzFLVYWdLyV9Xyd5mKH/UthE/S9
MMlrmq1DwPc0sAGv+PGqZPvLpBxF5lCSOgW72zHsVgpCkowYr6CyC2rnXGpDYyRX
o2jqGWQ/qPoGsUK3dU3189FLAFqOaLcAryndTM25o4TbxVt9rbsd6qK48WX7tlBP
JrVz2/AccnpwHO4KhLtkLEoSlkGREIIdTlpd8Qrqxqp+Jg2shOCZs5HQ66lkHvD9
Nwnu0ue1gJVROcAk78aMvzpnedBl9onK74o/dxPVMfI5TVo/HsxeZlL060Itp421
UGIV+5ggxcVXHPh5FL4tzvh9wScxrVnLvj27nnBXrV2Z6mtgyPGQ6Vk0XRJICk3n
r1sal4eovn+DnqSRrN2VTLb66bCsbdG4Am8e5zMxIcx4alTIt+xJKS/HJuRt2PHg
NBo3ynPQwzsZVLMZLcZ/fxLzn5wltbroarw6QgpU/LJGPTfMoL59aF632fh8x2hY
WY4lxmU41HUaFNYRtezaFORQ2UR+m6XafxacL81jH5CPEDb6VnMPlwC7IheAWyBu
Ra5AdSllhyoomnq4mAD3PmRtWCRP4R/EZ11mPTZvxUehn+J9pln9Qn1HAIljr949
bqB67VQ61s3yCwd1hAwuQE7aSlhWg+rX9tdhwrtuVFZ2dUi0+yH1GkufwOQaZCtH
RgP8uljDV42wBfCIHy4NIzuO5s4DlUqS09hN6SRh2SSzJrrvimvd/TxbymC7ksMh
vNBB0zaqRaBXHEdUCZ1zL6k0BRUhHrHG06+q4nUybi2eUWdAByQ9lGMkVDXzjM5a
6b8N4oNxcaVbkMgod4NIEVyYQp/03YmgfFaE5ZVph+znHojpfj7YmFe0kNL+a7qC
86eW4ajIDq3H1A+w4kd0mRynQexFMS6xb99WpwKPf1PWHvY/eGJW6dF7Ib7uG21b
dzhgiLp7A176q70/KMv4ZN3jl5jyrYR90zyDpSEb3r9UQzSCdwu3mk2y6v58a3Bt
eHNiibDl2CdyAks24D6X0ns6WxbFNorQfkFekl1IGrAgLWMPCJbPi/QRp3nLR0W8
l0HvQOM0x1J7CgooaNzldcGllJ2dk8K3fuFlUSoxbuTu7s7plt+kgzXmfB6C3/yC
eL+GXorw1ACpsZWOiVb5wldxxNWSegnPSp+zHcft5ESNC97ePvYG/rEzksVH1pEC
mhOGjpfvk3UgR1PSx4RK3MHw3X7a9jyuuvJmVtl4zhq2tXVrSDuV+RYXDjPqCH5x
rPQEkkh+7KdWTGop+L6kqhGqBmLfKRCBh0v+bVTRgos3ZEecKI2b0BN/dsqWb7ur
DJx3xHZb3q86LDpx/z7Ieyqwj7fC7SySXc9yS37AeMT3mg2zIyzWH+yWh8Res+oK
w+cSGG9m99IFLtAFmYSDv9Xax8svdXkSENOrZOq5LF6jYkK20b/rTI3pEErHjiOe
yt7nFxu8riceE8MYjSpd7A8jFcjFfPV7eY9cqIHiTZWK3UveYPbW3CGb5UrgVcEd
KIDUXguoaWVNWwmdwGe8tP7yeRfV3KgafNCKokTijHl+iAViTp2iPfYX/YkhCsk5
bL/3pp0eqNnDXvC7e+Wf40kEoG23iKMT1z9C8ZjHwqUB8GCCRZNUqniONXPUlDZo
IspISLjwdTV1RHxUNkV8D3ra1pRneMWPjcaeLpOUbcrQZ8WPgIMdi67GyWSz18qv
Z4mClNOowBDMGBzUQTGiMEMsm7fF1eLUWtP3khNzkfQgnjnjQww7Jv35/yWfMYlR
S796gzXP2UaWGugTQMa2oU+1VOBD+P2rpCvNaCfPEJ0LvHn2aElxOSIu0YB/Yyal
1ATxn8i6raobJvfCRMVDOkVjP3jkmN5dr/BKDW3IPFhPxoYbFBaSyOH30kgHIuMr
zf5Q+ibMYIQuT8sFZfAoQfvv51uo3z8S45STMaMRls8WbPQMVixry7fRifeIYvx5
Iq1oKDa11m+p9nAhBTGPwNKy+UpFm2yuOenAud4NE4Z+zshCnpJAm3XctMYjU1am
jQRWBcI4+9kEDeIhXXbUuayaV8biuJrhuHrRS0vZUZpJbnMeeUFSKDLg1Ky9ZHio
u0oAO4TCxlKvhwTTUpIllGbH4A/NjazRpkNNtpnYkgwhmvqYJNaOA6zf8fHTpTqQ
45ZAvRMBia5W8h/VdO4J7o2kIm/iN7y6sKSw7rYFvwWByqwEldmdqaMs0Gg/q+XK
CGooYMTG1zPoIYmd/LYVZkiS02MRG39w6Sh0iv0EypQwMoBR6EcYMQ7xCxw8pab5
eN7nPLefZDHIvYrz4tUaRhX0jakR4YSkNudWlwc2q/+M5SRwfQljQ7WB/KrrCbEz
8WCgBlanC9IXq0AfC+Ni0fkErikMhgToXpw3vE44JOXhBe6eYhM2QYsWCneKbQZA
V7ggwUOZvlgX6muRrm+QwPyhf9R2qTHFVuj6QIfs8xsIXmVDm/wugXRce5Lb0xTf
JXzDWADx9zrFV5S0IurSpkwknSj8shv+B5JiqR57pt69yArQGl3ek2sFIAwzaZXM
oCvPLyatS7HNhJOiNnKrhGa6/4acPU34Hd3BJnnqTqtEKowvLcv9lxdfljLS+oLP
JwSOzNOtSjv/i9ogEMYdGqojA0LT2oB1XqY/y+c/Fl3YyXKeOmCnaEWmgUQMaazh
n8NJoD8mF9Z8d6wwxFDXqXKFUv1OZdvBLtdXYN4UqGnvTHJwYDr6vjm48jVMzjvv
zFpWbJYRzn2ZoWRNkqFE03rx21s8i4L1ONOWMWVfIr8quoRml+UTa3gAbK2kLK/S
iRFNo8HaBOIMg6dPX4vDqIGSvcrEoc1a6P4hHHiBqISvfZdBPlkfgRl01xHHFNkI
VNdJh+4/qn5LSs8FCILM/30Msd879pONzDeycp8WsMGrl2gmtENxGhKlpT8+t1pz
9R66uhalRtGDX6jx2AeH4vph3yqiVznh4SqgjugDx+ETkWXVYwwvn2kpSSqOBGA3
3YxisOvfUSIx0dIalTb1zV1twcwqgieIKIOR7TQxDHYsgLqblnoViu8WG2WlZbWg
O/nJd/SLOHwfYAZf+s8tH0VUQZysul79RD984mP9Sglw8duKJwvPJXRtUl+avwUx
jIBYO0Hd7fMZ/SgHZo7TY6N3KZMReMvzCeFd9jhP8gMYqLDZn6lTCb26BGnumZvQ
h+bV+qt4WhzcZoUq3suj+t3hFKn24kgFR1z9J/IkxuRNLVTwMtELUmpTOeHEBElG
TJpvriRNeptOPeMZkXx2yy9SGLhB3mkApo9v6W+TFcGzqzStlbDAAgSg5iebO97j
zsn+GYq/3aXpYsol/EApYqGQ7eRN9pcJTWxm0K7m3U3z2F3mdwRE7cB8vCFBSCNp
y5Dnhbxi5DejJH+4NRCr038i5dfZaq3EYjwVu5zbFIsGf72nv8bxbCj3KtkEiH3l
zVe3L+hiE9yTJexFThEBQJvG2+FQXlahQSg4M6pgqdXbB7UrYuoNh6TgzKnKBTxv
kBAtKTjRVm/B50rJpDu+sDT612Juq0jDjhUWnmi/1CfC6Uo9osQKjI0RKq89+9ss
8qBvUk6bfGRtFt2Mu43cc5iGRfzobq6B+BNHVHwssBb5qz4nzonfvwq96muICA7w
JlxH/2N3enRW88zwNw6DWNrPSeq0co2EsdlikEb/NDffhuRU68jPRyXFhfYdr75+
GwUHtTMIPmJa2mm3r6dgRHyHiBU7cL+ASUS2KqGm5Yoeo9Zqc7qe9c0wTYFyKfzW
McxR/KINti7LTrDAVUj1HDGcjAFcOr8Q4R5vjbEbFKNp9kboSwp2BviT41sUCqEw
eciQU59ywXBYWYFbXk1ZobxCxbdPQd42Kk31RGRi0UmvZelVY2ZD09b74RTezjwv
te5iLlNT6jeURBly0Fp2MAqD52KP1bucn2DJVctSKQt9sU/jY1Krr1h7oLU1vFGE
Fd8VF8X5luREPfkR4zaLJzcb0dQMDEk50GaL+P5VjJ77+QCkhMJRTlMBDTiRJq48
e2+yTCkDn/jtCxy+1b6iL2bIMPdTrMlBk7vlxF0Q3AizOjxqU8qEJ0xpvCzyLtr3
r6XU7xP7/LXJUrZaXd7GcwHWXsa6M85GhXJqLdg8FsuuXb3d2QCu17iBrl8H1bsQ
tnTHX9PNI3N+HMjkXtBc14ThD1cnntk1A9yfdFpOBhZaIeAyhBmanKhtJ15cdrML
7rs5y5YCZz6ZaqLyU8lt/lz9poME6djvIMKJpjqU9Dk+vfu9zCTSUuiWl9FaLTDG
VcrLsjWTtnCsG4oq+m+nKOX89nAH/8GoJN3wLwZ1X1EYtAaQvSF+u7aSgKa8fobE
7RtARN/R75UlEkg/3iD2Gp7U8JJD1JuOYFmEMyZbMsrhZpd5VVSB+z2k/6BZprIN
a6IFh/gJxlYg7lCKcNwheWBddFMd6Lf9fyrFXUoiMGWtw/J/F9xy/HtuyxnFXOuu
awLAfBt949LxDnXKKOSCfUE1lQR4mfOWiVu148fk4GwPLtSmND6haDsAV5/e1++o
iXsLlEucI17hL240KYLUPlOwXtkVvpOH/pTu05gW6BBsul7H678XKV/0NmpTUIST
FskX+wyPzxauSSo72qHfWr6rriQkNEyaQjiuy2HUhDGDhcqMeBwvhCvOnqTb92lw
TCnh5rk8nMEPGcU3t8GDhRHn0Yp80J/9+GuLhJqPURf8T2Yx9Rtx0Bq3AFu7FPZA
T8QWUM/91BvvrFMaza43IihIMswrJyydofiXEK/J9vn6TwWmqizFFxgA/Z0aagId
UZDMbmNoEro8jvTqqF6LdWn1AVkDwNr7nR+kM9qQ3OzpHvAZwDJ9hDwTz6lX1oDL
u7cXKAIuOS4KjP3QmMXnqQl13Ixo7ceMv4CjCPybomho4osxa1D72aqH0bqMtZxf
sudz/LMsWYUFti0CPreLdlR/qPJ2WNCD2lv1azs05WSoSAefLsSdl9DV3xAsx4MD
cwb0RVrt4nyG3S9akuhNOOLXkNTQWSZdFA+DsVDfrSxumuB5qH/388RuOVuemQZX
Ka+TVPxK06SJdpkS1dj/et5Rnj1k6A2MMFKunJqLrECo2BNNN0pKsGhUmuOsxT1l
f6mtLmVwcmEJM4TkUFZgOWaj7sfm3MrckGRp96M5sd/BBmToHJAE0eWCmrabUDtE
pW724IlrsoITZScA4omc1lZkafyApk2pjDyXYSWBjM8pD8Lg6mh1yxXHzxOVGDeB
AxKPExKSKfyDtOeoUDWKVK6MNPwyvePBberSFdac7FNL14LhGaaik8ST7fv//CC9
1Q/bIECI2vP8gj8u3ZTRxdNtJPNke/H8eo3SlGm+GOBf5KEMw/XOHPgsELcrgQTk
I/sltWaUOTGLJh+UzLqlYs1OGLK9B8mvqXrGFOlk6U3e/cOcZCyBoUjFH0mNVHB0
OvH4ytAKG9KLAxIQ+wpvNiFHcTVgqtJ1VwDUysjZ+SqTbrQ5ixDMLIsGcMRXpLv4
ngRl1ClkJbrxzuhp6FcSvzI4aBK+zDTTOlav8ojDov4F6sJaVVRv6qZGay9VOr1a
XHh6Y0ONhK78fYpKUn30hLbJvFCyfTBJDq+4uDzds1hF2NupGUEiIfrjppkebr83
QGDXDiLMKFMo3M1odVRzLV/tOXEJ1+gedO5kBcROySLaYtaHPwlqkRUhPMDx2ETk
RhUUvpAPxMYSFDDIfo7P+Hd1JrfSPxXA+2Wke1bFfHNYduFcB3v/NSMc4DdOK7KX
mx1BPmPnFXh2gMqtN0I63zQSNtIC322hNcMTvD+RjTZifM/GnGmYEx842LR4TIII
AMSjfPC9Pceclek/eZGI9mTfTbYCQklhR63ib7meeUJNuBQHK1C1BmwlUx4+Q4HE
/7nlnKKR/BpdH/qZIfbm1Qkiza/+BY+E6QXNAErvMDwN75iGX5W4apt6eFqclPEQ
3k26cxEJ4MRVqGD9cjQM1Gaj1Frgq3+SbQ+TeRcS6pfoLpJh+IX5gSwRbWG5KHHd
24Q8jZJI0uIuHNsRyp5YHWWfrMptA2cyR1attDlhLmeaX+QdtvBqo40M7GNC7W3l
Rh78Oczf3I8UCHcSpMJvTRrLWBdPGYjWk3wDRlKHMmFKfwqur2MXiFhXJd/S3pqQ
q3bbWSn3hDc9W7k8y+79xQmdB/7J6U7MtFgMm6RE9ii9Ipyd+PYyUm/MpVRCWUhi
eQhulAzE7zGih4TyBP+iGtOcYcWoxBhMiOThICyVTmoCkixmCl5Kd5VSqYQQsi8d
8q3xkGMQFl184p0Gqhpa1w1zmta26eGZT2/RGet0CNBaU/hKOOtGynQo2NDkX2S0
cCTQBffaq+uvnzChNH+8ETTaadfXaBa6oR3quTCGODRflEoDqs3PLledU+DYJRq/
oSi6Hqc5ConkX+lIGScHoM4fgezL8IlZwtW7nZyqz6YmMkQsmm5Uwhk1RGTsDYGA
bUAdEY1m3ilyk2yPqLwN76F6a2xB3asmjnHBGJQKG30XToeFKtSpVHW2HYHcjYI+
0IsB8bC10y5swTq9c//5cB62bjEsJtuckv1Q0O2bxM0nYePm/bPgqL5hBNQRnoIZ
q1U81WSLv8N7zbj1znM7jfVOMktQGadQKGMKrcAVdBVzN3u0bjQ8fWDiJ1F0Tk1T
SEM/D9/NwV8thlxSRp2Tb/n/MU1zX9ho1ma9gFDQ6YobUm4IY0bzbGm3MrqWZtn5
i7E5ih4nyt4iUe9WaD0j9VE3rgfjTXGYTKR2/7Ihza3vjTKFr2f9ZHMh/Wvi3yiY
anIeoOgqK/wOZp0d8Vb9gA==
--pragma protect end_data_block
--pragma protect digest_block
BURVjB44qWIcP9V6gj0Ua2cOJOQ=
--pragma protect end_digest_block
--pragma protect end_protected
