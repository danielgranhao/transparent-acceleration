-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PnrxmcpX8B+Xo8UlcvJfUkxO1Xqr51uP0ToP5HsM1lf9tLUj+HyKQK3/4Chpx1k+HOF+8WN9eZ2o
r2ruo+LBb0jaVs8MTVixG0MC/hC3OZS0DXpwui+pH5eI4+QkeZ2wzc5WPwTvbFkKarYoXWGGMU36
mImn6HAh/RjQjm0U2WODWr/FmIhUwfgowAAFlRGozbK2PeYQ3GTMu+3aGSxJf2PBjt4gnuxJDg2U
aZTGDkfgINyDPiSVBmdy+DoOpof91Wj2mARjOp06cd/2Za7cJ975rYVE0TWkHSnCMQ8EOSF2rELM
9DCQviUeEz9Vn/xvl+FbN9fSKHL4BJgMfQUImg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 13056)
`protect data_block
9yBjH5BtqnYnjLZudNACzLf51MtkopgwTCW2yD4nDBfC5IOc1vcFTeS62puEoSddTT2N7soKoxMe
wC1Q5AUEEwBWOIPVOO14ZDUBbOmGBHvnKf+gmjF870VEB4cXd5yCOIAcEsZri5ICAeQYZiD1y7mD
QO0UQSRPqe+LoJXMTih24CkutI7/joW3MjY7Qa5vrZsOoXOeJM2HoKCXz7TauFcLCqpkVnXF0wJW
w3jKAbQRcA7UhZHV2dKLSVNYI772LBVkzsa2kYdNp+fjceX6jH0uXoqsjQpAMsO1MRAvoWKq7E9K
GLOnbOLUgL0pBcUKUwMVbba7oEEYoLy3x1pv0D1ZIRMplcA9uoNTyl/0P4SlWj7jdekR6GQvt5OH
oYh/ej7pknzvSQ4/qIFu3zquO6h075jIn0rcUBqOFFkArSwegjRVPfEVw2xH+aAWk6p90cwvq0Ev
W9YdNNbxJVVEZsbvkBvoH3AAY9tkG9dsxWL4s3BS2ny2ySunb1HRglZbjT4mOJpEfJO3gVsNHPIW
E1AYcEBYFyEdbKOKfp4SGjGkJyIZMsZMikGR1Ilutq69IFqUMgQKNvt36dWUB5zC3GF0f7am9Z2p
u4f7biRan3sCrBKHrNmdNcxlnjO4WVgcG7z8YeDairwR/BBuOxn/NSftOJrloXvN/av4qndaodET
HFirHpZIhOdonoCtJf9erJjL1VVRvCgME8sMiq1VRQNj0VqN4R4e5t4GiGzNV1LFBX1KXNk4Hr3o
7/EMKZncOSAzavg+Dz9o3FUzUJiZsikJmulkXYHhlXKYxRfjT+s0Mjo1XtXl6lYL7qxJNnqefG6o
CoFHRvOe0xnkraVGCM/As89girFvEq4iUehTYue66VeDQriMLzOi5gVsUZ9HXIzAzri93JpQ1gOW
5BQOqT3L4dESHq5nC7iE6jsah/K3/mciaKmN0XGgVr0EmFskjdeuBYjHxJ6TK/jZPb8eUBlfe9Dv
Ye2W3G2xZ/DIWx3onHjwmS6X2hgUVAnN4tEWHwN8GEx4Awu1Pp/ZDVJf/ZrFpBdeTgTeqMZQtwoV
O11jzq+Hq30RAEYHtYI7enSHQYQMRZrQTkrdF4cYM2yoDjfOlW/XhpWZreKN7tYBHriU7xMtk+OK
xjT5dMONur+gY7aR+lkvpXFUwtqm3a3GWEcjTsYOMhLYu6wXcvy40gSpaTN+sveBQhpP+GMfVZn8
CdWztiqkMNYtOlOORemfRF8OTC1RSZcBqA1fu7B1GGTHCbhefgX+gq/6mt+qqtF+0bn8PZIoxdfm
Xxja0rBRUgDh7HAuW+P25gYIVuiAF5OhTddTwkd343OCRP0+iojNEopf+24Ib2uiJ+RwB0/MfgPe
0LXCuc6JwjH8IbrtWgwDxOGeyMOYjSbdCNpRyCXim9jWjnuk4ZFrazH9AoO2gYatT9UsgqEV0Gef
QLNBg0d1CbqUU+PQ41NiGj1NS+4TwGs+CMhOoFQb8SFBoKAo/n3xDcihNWUO4sCPi1w2kHCFY+Zh
qJTsxWKsCJj5ZVRL91PtaXRgV/hlPpcCqAxOVfQPNXD+sInmcmhTZZV+0lqavboJh8kEdBdn7/EU
q6+XXsnzT7fY3nf0JNIc8NjL11JpijYdzTQjGWjwb3AyGlkEK8yXekS+o/E/v6uqB4zP2bGA97Vx
D10ZKYRGak9k5zwswNLJL3LVZE885JlgHqCVQvCzrQ9lR3JjCWck4fFvXL+sOohCUuXyAXefXvA8
RmuVAjgTMnL1MtXfuaEnBf/7T22xPRp35Bi790KIOb+lxEzmX5dDJ87+A6aaG7AKnOdQh3F9JMpn
WMxQantYyjXlB0b5CpNBgEwOJPi2nyU5cqFkSSpORos2SEVMLw6NfhQ8Rt4l9IXJfHTcDmagGfnh
E8fELxJrQhEDdtsHXl7nACBAXhTWNi5ALpVXvohhOYw/MsvL30U4uWOroIswrnlGdUC3Fz3xKP+g
v9NzUxgH6RFaRwET/CXtiBmCUPjyGTC4jLWb8CcvxJzNhFL2+2zbeNsdud1vAYymMvu+Lu0pPLEC
Zr7/NCb4LXIFh1hSVs7IH2h4JF5yD+o5RGpEdFhPSKHATH/s2S/Qpa6ERIdTzgPA7SbdzMg6JFOT
iDKh68+eU5dN0Atv1wFJ06inw7eLN/tl+8gDOgwhXBULQVk34903g7jmGe4w2ce+VGsQvn6Wu9ph
1xd8iOCInJijxsxsWHwhvi2v/iIuuRYIcDdMK+KMES2+pVGF7z7Wi0AnU1rfkYcs07ZXBwXoI0Ap
jjLsnni/KyoZmA8rW8++oqzYXSSIa0Dm8D5KMBuFgo3ZmoiEz+yREuTgTIqLudqg4Gptn74yTvng
hiJ9t89weGuZGsWDUpFXUfbBKU4nZWYpAmxjoOb/t5abedcpTWkYo27f7ruwkyu8+YuMmpB4/X8y
EOvCBmJ+T9+0SkWHFdO9QRju57XTAo0TIm0jNGgMqH7vUI7t584kSIAp7OyW7KCOQJ88t+7f+JYw
MiKhbqNKwn13JIo8wQgfm9WgBu8TlaFn2srydsf+tWG3tA+UXlBuN8wMs8LyfXzKhFDZXDBEC5Ls
c3Z0V9AB/3Eyu+kbGgeu2XAKqGs8CKC8wvkPmM2Ou3efhFIs/j3+FzklyEDwiiNWLXlxnCOiC6WK
KNZ0t6qazo8P2FhpSBtLpgZtvqbUyl3RqIZQuAE+RC6OZWEfuVUdVZTjETLE/jubC/OrPnr4Xo59
U1o2esjy1CnsLPU4YXuG2CXpApqaeKixcmYJgMmzlI8bVkxaSbxasSeRCmx2WfrngehQ/o6sFY6G
0LLDzfUBsHG/D/MPWZ7y6pWllmOiKBehkxN0ts5qryv17KZdBKugPRajhj5VP3lG424Drt1DGMkE
H8O5pH18m+heqvMfS7d+yZYyu65Nv8QG5W/4jY5dliNJJAzOAt3wfUY3ROThkOFTI3CjRsaZhfJx
2yNbUvK8GNNVK33mo5KIg1l+IeC4Q785HEE3wLePJqwCis+0BOyWAO4z+jm6rXvVeQfAFRFZDqrO
w7dyUi4tTEWPk6WbZ+6LVg/rln/vLf/enpB1McB2D+LxlQ+cZjinq66nbzAf9ONQDUcRR8vB8SXO
/+LgSgjH/G0bfBACFyuUntHqU5PPC2mx4TgapcTLtJpJ/UMMnF1NN2nMrPF7dOpM9hT6ir4VVg1E
ODZMpOzgT/XhLIC5BTBvVJ//WpYDM+DIFy21B11YzVryzQfhH4nHVlkt01Ppn0vGWto98+TX3FVV
9DzsoDezBRrxF7ocJMU176B1LsLS7CnML9EFoz5eBiJuZwOSC2W0ZSnoYB+UeXiYFAbOdptNMjRu
Bii3TEEJZsU0cI1KnVfUDmB5dIYBmmokt6xg9smvjp4m2eeWtCrtTzDFdLXXDzwOc0BFTMlonj5t
mJpp09ajBQzR+5+uJq8H0Y5FZ2gHGJVgOSy8xYO7ZP7ReHL412qDglC7oMA6PIJ8+y/d8p8BDZwU
QfWoYEu0fsbfrNfPQ6TxC2zaGAq60my0zvsqMtBT+/RJmV2oHf+9UG6LI4oz+G9hTEwdr2HNFBG5
Y5p2klGJ8BSHFcEvyl4s4zEmBSISp1GBis5wRre+JLXCkuoDKhBtCiF+pvsJhYLzy3SSuW4scfEA
pcDb4/GX2gxrxlionDLOmesXV9sg3q09HIlrYRGrzzapr/WEgKof8Fl/SPG79JshleoiU0g/nI3/
6xud+U6Bj354R/0ovmtM2AKzQLQhIozLvzgLoFVXaItRCPP22UH+eLZLCYNCgkgnVmH0bMgqBukt
MOGzZ7AJcSC7PVsqeNrV/f6DcHCI1CN1kW/TfftTEoQfyXa34ZOM5h/a4FSG2GAt7giv3nR8Yq0Q
voQsQTu5YvZEm7Bs/wVuMlUgU9I9lliuHS5XScjSemZbcE18P/la5Gw6gdtgPbw8TOhNJNW0ebnk
sjVMl6sKVDcFmLoPlL5DH4JXVJBa5sXeDVd3jH+GcbC46fkA2wZkhr1L5c9yqlQ+GAhBpIGSXgaX
qhf+ljn2EuopluQUC53lBv6NaLLdmGSoax8Oj1gJulppGxM/QvFvIftDgKCopPgNkKcWvkDyz0CO
opJMNuXDniW+xCYW0e4p9yDbpK3034kA6oIgBbXtYjITjyv1/nbFJEUmZ2xQVtrBI7pYrlJIpHt2
Z0VVbMC8aKbuZgFIJFnqZCeq9l6xStvQEoZz5g+sAE3RbOO47wjAPJrDaI2BEtuNj0qe6ySfUZHb
uopr/GHn2NqbILaxb5tSlFG8Kqqlhcsv/00BPy82YF+UwoR5WK3AgNuvSELv05XxYF5p6z/4z1Ra
mQ0R3NIQsXlKN5Gk6WiZcip9EUamrRmifDEN8Tqt802MjCIr4To9+JJzn0rYJgUJtqrPjynkH4nf
yZdRn4w/qYimJiB++Nt+6hF81PiqfuLIi+js8QGZBGlHQSiX6UwPxgUNZLmC7/OrYJup0PFlXGBT
/m3soY1ptOHSMrteQBvPmDc2vOxTnkOvHydCAx9uBTcFYsxc8qOGsqL6drfD4C7wggFSbGiUfSXL
kKC8njybDjgCtn9YwdQcxN9CEyuecl1VUV5wV4Rv4vpfDkkPMnZYqKvlKuL6HQLj7siHanuID2Q8
kF31KqsaoYU6iEyyZkdT5RbamQX5f6CuzXDmAlzRHdQX9AhlvK7MLx7mTrWIgzCtoDfqI80Tmxxf
jr5J4QSDRoJk5648UqmpSWY8yTT+OhjitGYc+k92baS2MKbCnkUKtMDMbbr6GYUmbKB9j2U95PYV
os+pSiEMkr05YWJAkZqSboMvmohLna9HleeUTsRlAtUffA5NYlXyCBj76V+GL5M4LnwoVvN+7Usk
1zF48t5LT/yqW3ncjN8EAcOisplV8SLzaI6cUw/d+RyrAcgXvx5uFVMWjMViSz77yS8wbw+sbMMd
plhQHgSowe6cDLwTiLCmesEHZyM6v2V8XyPVvQ/W/2+LmPH13sQPeaLg4LMPaysjpzSH1uGkuTbo
+SrY/2SrABWgueJMCH/HgW2Y7D3ddftmy6j6iRieA8+/I9mJEQ7YOdVqQUavFkxhD0g0vx4V0yCw
JfTvMesxK9usBNZbSelmc+iLtOdA8J7jJCAlHo8gN0UJHSTQZ7f51uegLWPc6zN4HoxrTDxdTO1m
SEg5sHxshS9xrpkO7iQuV+3Hz1WwepIWlYWrdXJ7ZwK+P30ElYbCiB20rYMywwhLxiJiRv9LHW7E
gV0X8NxPelz9dJV3zOPAHWaJXmDx/u7aalA8NfBko1C1h9Fxu8EKDilFxSP7wySzU3XHMsmOj1YM
4h04863Ll3Bfde2JU45KAjgy0lhfxX36F7g3sr/arua7711l0fr+Np5pf0VjmzMrBujRUb6xuv4X
FBPfUyhU2kJkZUudhy+YxOuPJWEXZYvFXT4TDBVOFHv+myIHnflE86NEA4wQNQzzoGhlbs8xbBHX
bGPneDwYWlnUWhYbWgpJ7q8s/X061VHlCbvnjH9mAJ4Qg5t++JQiGCZgsv53aZrGHgJfYtqIQ/2q
kiTg3MVtLZXC9RM+3ygjGJciSjmd30lHwHptneoWaLBW4RWVmcIoTfF8Kz4+FKf06f8IJjumo9Ud
hyrhpAL1yq7zeGeemC2C+C2KE/mON14Qnz+c+reUWK7hIiwtkO6iGOJjo/T2dEu81GPDKzqXQpnZ
I/YCcuLdF7LIolVw4G5RiGdYF6kiP248CFGwe8TBL5YOJCXRBnVsKyU2gFYyMH/Hze0Amy7u0xle
t3OChCr4LR33sqIQ5TezIPSC3cgzPa4p+SqmHFsXXmhBQQ7b9xba+TjRMuubgQiRGxnscGm6Gk6W
BvzUBEq8chq3mZWGbrvQJLHF86p85zgETGXymmYUDUWnhOhf5DOv3t4S1+8Sa+pYyhOT5kp2b+Yz
GZBJko887gvfkUitn+w0sR4V8jL+RzCjxy16ZqTJZqzuGYOyFxuiFioyz07kz9JjyWvVfwQgOL1U
qQS73XfN9PQlvS8pcQ5mpw/jBDZqWnFhOmVrD6bL26nNKBl57XsWBWpFS8zu7DLkQqHKA3ik3R6A
ZDalYLeLlVIqvTC8hdZzBdsuS1DZcDIkgU8W6nkg0GahCAH9ALNt17do7hzgLRCD9gT2i3Sew9NC
6vbZuOz/GI8haWPTTHPxku7wq4cdVJ2tpvcNu506YzBvcGfK7rB4AXLa5vl1aOLPcAxPlzrbVkTt
d0h6kiT3ran1ymobIz+fA6LGvuVt/dv3Kv+GaiFXPVQr1iHidPDkpfw7cwF1LWyMjB7DZUMOLkfT
Tk0+tAQE7vt+feGj/MF9j2XpLig90nXf3mScUo4Re3vpGxfR7VeVJPD6SwEhoJfmLUs4LNyMiDHa
SmDNLyDofDLNUqwBNGTXz9wNsH6k1QV/VcNkJAITIpulAqQt4vOJL6qmprhoCHatbgN+qo1EmuGJ
SGhM/DlM4oTNNSaMqq0JM3wsuubmSXExYHDKpAHLmnxpHV/W9UEfbL/UFzBfj4q8b3KkM8evoUYH
kGJlV6vsGDiGtQaYWDIXTMnRzqDZjdAdylJuVmKe3oVy79sSy9ZHGSezfPT9jbS/CSFMSwLJ70N+
mAoHCros6XytmnFfiatzkS6URE+tt17fPUP96tulhcb4635Ax0DRBsAGwx2YS1hTL/j1N1qwZXTo
D/JPL656kckeSqNIYs5mmarldcW0XQWqyV/Af7hJJixGnTmcEz1R0h5WOw+HLr8KoqdwaabVQCw/
Knll61TXmWQ6tEEmlcb+7GOPIBqu0nPYR0BSAWH9wWpJA/UxZZXwbwfDWowu861KzZ75QFF9ayis
hyzgIvvU8aZI9cYBBLSoH/HwfJKPuVdJ0QUzRZFl4Mt4XPb+OBVxURe3I0jvp7zQ/VNtK/uYWi+Y
YvQFqrclnSXv95wTKim0u78QehZ9+Dh1qfwIzRatKzcZXC58Q518lnfJzBKE5VhR8qx9T55ebk2k
Yc+8rtdgmcinflTOqoipXoygVPIE65P0rTWYMKB2C9EhpqZAsjBdyoXEpYgM/3/e48786OJmlDb+
H9CRgjHYwt/2ZqieF+/9G2Gce0t5z0xT+2p0SewTZlbLkWPh8j6b+PolVuehbESgOWdwJxxCpiEr
BIM06XHgOx7aJe9jTUB2az93X5pyI+coorepufKuuy66pHjGma3ZuBuNVTNHTN7CRRtZM65CLDqn
sO4866pF8QeFes5P2vl7F/qSSzoby8Xr+KfVR6GqWnWNk0c9MkBJxQ/fyO3eUoTUNPBCC/LoU48i
S3pNxI2L+iomug/PW2YJkhm4Q16FsvGTVtxDJfchU7Hvqsxu36qEdnCedh9RDcrsBpFWzyWJSTX9
oMpGgKe83B2VWCgLzCE6BetrC7coMrL0M0+fM+aOKszo+M5BtsL7YwAHChWsfwEgxJgYJeZha3Z0
ZtS1M2ADGEUg44Ceup2nY81u6CVelRgfSMFQr4haLtwcatfZ2+6D51Z+7DAvE8HciWHc5o+A9Ty+
3coOa7yKFE2NRrf3vStugLdtObjUZJTcXl8EGumgOTRF7FPUcx2ZsOXeikW7fMcdXER03F+XpmsY
fouQE7TbxLWm5go9YcoiU8eig+iJJfxOEsd3n+hSHEGTbf2qrVMnPAKGxSWYzzTlsp1ODzcl4BXF
/Clt3srQ1YoERAlxqCHBPzM8hfChz5qVxWnUw4Z/4V2AUfb2mg6MMW4hNqb4mBYAYiKpjWEyepWM
UUEHQH2iAnEd9HFq0+GHGr9k6LBbWnpko/Yd8QTyxcbRrns04RVSsOB7Ib4a4V9FK/WvkaW16T/W
UPFDoCfhTvk8COqJbi9CeaFUmIBXaU9HDmZQIA+Aw5fi8jrufnxbORQLGqI0Xz0U273wjKhHVaSN
AOYKBmxBXjzLg3kBZ/JCj6KNRQNeZL1Wg2QFZLYr4dCCOrb1YgmU8FaXlFzRUnB7tHG1ZRm3gSMI
B/zfldfVRLKVWNrxIobLR0KMr/dLZy6M2mmsFq0D4JmOEcAdcMJTTKqExsXiUejz8vSwF5omm26L
WUXgWsSc/b45CuZwBNkGVUQ+iHBA+1S1W9DTlNdmRvdYKD08SgFXVMHKlHmt/fUDmUVeGHUQRVZ9
kCJRGr/eGgcpmnPezzvdz+Se1WjZv8xm6d/skWFDsu9ZK7brUvsXvoj+eF/NMrveOGBOgHPjEgn4
TPywI4FgzoSMK1ZzzFjS2ihTqsK5L2h3dcsWZeRO8psze1JHG9lslJF4ns5EGz/CZBQFnUxEKftQ
0XZTzZ1gaiYzxcLlOdpI4x02AGWUiJy0taIDkQdU1wpTEQXmxYl3Gz6bIgVBnl14W7kBL9H+QqcW
ekNKMYRUEjqPXmGMcz7QI7bSpIRN5OE8CdNDHG6Yx65ruaNQD6Br6k687sfUeZoif1xe1dkGU+Ea
vHAzJ/S+oYVwg9HScACpCc8s/AM9eQf/gx1nyP4AwmZJpeHALGdmfBVwr9BocljdRjAbrO3jgkcz
jv7/Z8PKEMVkxTKgCopXHiFUY8v6lAgukizHJZ6C/vj8ugVs/ibyjCQcgnw43pZVD/virWoJ4Jxr
hnhEQt+el13g5TRRR0icHtl1hrR9E8ZrIe3VzNosfcto4IXYaxv2d9imGQYWFmeVYJqspWoBocLL
5DnMG9eEJKIe357PKeANVPAoL5tfQ73uNj5iZF4RxxOU/NB7FViucoLFsVGgN5fwynRR290e158g
eqslLdGcdoAgATUr3p3VDiObROzwTfkv8i93ZZTt+HItls2jqrQAv/SW6PVR36f1Bsb055L+fnTb
xJIYPyYcjp0LzSVkXvAzIFVLm57xnwQGm4YwtGnqf0w0UNyDC4uzkMt8oTrxBRl/DFWLgum5Pad6
ULh7fKl/BoiqdfuPRvsCbVFzeBnGBOVPbi1MIu44qtP/PyhuXwBJusMtQ4q4RhkviIGLkGd/fvy4
v1Md5IM7RNz3Unxi1Hh11ggHESzu4ZIfNrh3KtDzmy8wA0ooNzAISGtNG4AaNKsGz6iMlhVaGocy
S8R9T2ZLGys9/9ifJ7/YRm17sbNKlVm6vUGhI1z9/NOoHc8fVJOyrKjMRyMj8VSq9t9XGWFjNyPT
oVVcrd0ZSsTeke2N/IAAssxZaxTW6Ylh4IuELn6mVwxZiytUlwGd7bHWs9SErrAyaN+Lwtod47be
tjjrZ1R7AN36dgwB+vZdHpKy39Cvml4asvOcml6uNUj7mEZcqirOOqLUDxsEOIzPpWOiR9Arp2kt
5D6AyxpaVfmb7FemlZM2vnLbgFPmtIVJTYUL3bgRQ690NZArizlG4cjMpHhK0XezTmNl9XCt4iaL
wSx5fi3a05ELMEioZluD5cMRXNYK4uAMljbyctgsYFxCWT7ZAm6QA658NnRncTg3prb0Iw3XCk4K
tVV2bsDo4x1t8Xw7GCsGTghhHxRt/L5lP/7Tqhis8p0fTarUwZ2h1v7rBLCGXHP2sUx60pU6b8zo
albuqbs/84M60SHcWzf7wsJQCbrZSd8Sc6bKRJPxPVhwCFctzONfp/HpcxlsHXswbzA+SX2UBYmy
cO0ocyLGWqIUePxsKo8l/IpZM4kbiadPlQfp/heHhqr1XgkpNUxvW6XQwfd2DlVqZkFkse3Al+a9
TcN+Prd6ZYnwDn/vMQNN8RWSUA4XFZnoQcf+fp8FcTK1fkn+pyX4DSjwgS5nQv7YrLJUOfpwWkP+
haKYeQaMpIWJ3wHWs32+y4V3xdoDZWsVcYmdgSXln64GJJFHNlcVilXLQ4yZ4tO4G2jS6U3DYrQk
DIdElQRpKN5oaBpoG6rB9xv057/S7BS/TrpZLQMwt0S7LU2Y40olbNQqpyzCTJ/s1DvNRrHVObQd
X2ZPSo0px3Ubw9W6UN/dy954ueoq6JGvgip23EwI6jWSG+XMj3sWN5oyhNZGxisLSzkQK6NdG5h7
ZUdSexCVZTXo678SUjZfAeWQhhO+KRXsQDr0a4iZ9tjXYkPAJH0WDlo3GyHIVKD0Q2RgDT6CGMxA
hqrbU4uTaoaoYaDW6VT1KfznP6Tu2UylWAqmU46yDB+UxcbIsuVK9LIwrJX7hmTFfjnAj1Pox8+P
kL37/9ygb0hDF+PB3l6eLnLqYtf1ydloT4w6fDMj+PTUxpplC/0K0NSK/A2smGyHJT9a6K7+3XZQ
+LIyE9iJSXNp/oGNKtxkD5HmCJbLBVrHIk5babQ3DrMMH6z2DApFBrX8OR7YwVnz7cwss652aFMB
Yhh6xKJejNtqfHv+z8ZC9TNBiN+uZ7H8AO3tdHAfIkxDzq9VEetSmqGmv69e92KJpzb8Vebblsxm
QBoBqeHwS5MsLd8ka3GlU0Ne3dRZ2LiVqYNMo725Qvk51kkaB9hOxtfbJHl6paZsz5+0xS8M5VJT
Xpv8vtZjDPtGTSV58sZLieZIvn+lk+4P1e5vNwJ7MClgxYmoxhLQKDg9WYctOhC5iVfiBnk1Mgw5
km+71cC8aHoFvK73hMvmnZyrlz7UHQyy/of9ZJw8HGgURJkGcALq1DG7vzds1KyHz7u8ZnhhoazC
fAFKPnQTdpncPscbLKzchVtyQMD8tEN4sF8hoMHhtexORzJ7ur1AemVUHZY5WxMTgKoSBaDOXzl4
BL69uMN6oMRnvSSnlA+UboChhCTT2txmUre6v1VUgUYHjjtD80GTW8uvREXtaYxUL05l7KwY/cW/
zGFfnOeaMSsju9nufD5EmJ30+dcnfZLs/CVPQjBN44L2N2EZ047TkeNiatyS+uMid+00CX/SkDnj
HD23A88b3gkyMoYkKvtTLwhyfRrGI66j3IHNfZTXLYngumEOZQbcPn1WE7g+jSY4N0u6QtMiUCTp
ApdFo3lw1OVMHFkkh5SIuJePZE6LAHQaTbxDESqrCOsucVSEpvjB8vl2u7Lr3f+Ycw1GUK6dwtvV
3CI5H/05vZKEYd696ia6rha+6WuerdpgmbCcgPh2tjMeBfzxbTdEGDu4ZcorIObWgQrJPJaQVzL2
Ybw4SJDEvsQn8UJPXthMl0y90/SqGbMxgnXW/LUgwWfIBTgvTk0NXpAFwiiiPlQQSEh31dgrFkeT
MKOupxUkO/UKMBJg+du0MQGibEK01rMkDcKO2yaOlHlQJygZr5Y8rO/u4/52jlZ7Wx9ZnqnrEQSM
1ssaAfOKgGEi9ojrT6Yl9Eg/4HC1DxvFJzE9szJ9LqBbpvm9s/FK7EYDFBvL7O09pbc6Ane5q/vT
D5dKmuSVYBmw0MS3vYXg3CSZyxznofI56tPm9Xndxw9tgtvqbm50F9wImMtnWVer19HoomZ1RHPp
xdwLWkULullcrZLboIzGjNgmX/C3i12TznjwBjUsjHvBvBdjxfk41mHpupuoFVnKLCPip+cq9ZhO
D7y9tYXn9mNLq9L8Fw6NC6Bca+H/1GooZEk4T0OQua631Rr5R31RC7UHVOwxvCrOT+eoVb5UAK7A
zV2nWaMYbI6LNenwe8RUOain2TU3LhSQ/cZAtC0Hv6XUG8AxQ9/o2NP7nDnpc+3gujP8BdGz1/+6
zKhRyy0+HqFjE3EcSFghrHmXtxIDIhIvGGy3/fTnoGx9uLHu9SDNfZPpcBy2AD4R0khdo7MOseck
/g4Bpk1QBeguGlwbC1kt3JFivtI6BI8qjUME8AOvMZfQ6WQvYo6CgzI+zEOohiMRNo/tt1p2gFOI
ZODLhAhfC/qigaTnZS9RV9ZEHFwYwQbpz7zcb2hQRl3s5DPDqZWOjcv7C33AfpIu4Hanrh7AYhOV
6Qb1m1ISEM/pxbXJoGY6Uglmqlz3OHkE5Yc6vqBwvBKabFxKb44hypgDWyZQuZfvT9SZcJ2sNOoj
Z0maRl80n5oOdI7D7BaIbwwuo8od8oz6tgOZGpNX++8T4i1cU4vHxsRxyrUDVH7neOmlI5kXCfwP
rXtEUaV3TDFdraP/c9HhDcYPIexwve9zOU7CnQYd+ztwNJeH9z917MhYEZHris8ckvKSqFNcYEp8
NDkktipNyVjw0HBInBe3M9ybut8QDB7m2u3o3vIA8C8cV7D28QUOZt7nVWDuQ2gFEyZP2Pc0e47i
m7NWu55OGyI8ZqYu6ki/3bfBOT1n3H9uUG/uUCVoaCJxRv8GdovI+kOjNPpPF6YHcfwYKj9wuWqe
Y5JZPnKPS1IbsxkJOUR/wvbHf6S3Ul/amZsiOvvADygG2VB0fHYFIroRvQgM/xrnprd79ymgVZ1r
WmzG8KV0NgFnXaTcwE4/0xkv1IwkbGboMHizUPD+TWit3C6mky7Qfls3ue2DYoA+24P8ZkVeros4
jLv1nXtmsZrJldA827e8Ek0GIa1xN1ql8j+Hy4xnI1Ku49zvJdMRMW6lMZh6eS0zhUQx9385uNCE
oSsQTDSvRBhTljKVkMLo069fx4hU5HHWlvGICAnrrlyXFwc4ZblK0VOh+0/+Acw4nSLKWfrtH/WB
q0K1KFMC08LX4tqEwkLIbbhsklsYGOVioGE7h+9Z29jXEcU+AmURqw1aZe8GjE5kPOJkzBlks7d9
ycieiS4vA/X0DPptcDwvoM5E3pycj/6r+ICDoq68Mi1zbYsTYy/+nqtu2Cm3b+5dntz9GG6FvdRm
uYNGkmzu4nl8LQGRsvLhpliAvNW5itsCy1x8vWK9bJIW09kY6I7hb3NQ41DIG9eb8k+XXedPvZC3
2sRJr4axkBpnNlyshEaI3OJkqX+N5tl55jkl6yogdihLvQ7Tm8uERdtD2WUGWC1Ihz3rJsWnQpja
PYd5tHZQvws0T4iNbvS9zlLC34VRGe3u8yVJJkdPegjszqidPNXjz6HfzwhhDztNhrEdTaMo9fhV
hoyspSPGHmG5DagUCfDQ837HV1MC1w1seCLSYWMY1DF+ULeGLHa/No/lZb2WbhLfel7Ugk8/6cZJ
S23+RBRcQY9/xDM/8lpbQkmgxxDofBDUfJQE6uWoZXOwGjSwc+r0cRVgM0/MHJtHK8eKIUu22JNh
MHeffXWoRezJZGuaC1rHxA/XJ4MEcURc8NjrQqnw6VuaRtGB7GiguFivwcV5qTa/n/G6uXh4Desi
2nEulRiR5rchdp2lk8U3aXTt2LeEWdpmEZ6oka8ZGfNNbXJxQ0kCMTcyL1bpn0rjaQAYwme2ETGN
GjG0FISRCsPTe0SoEAilFdAnzkCy5RaKbVDgUIfZZbYPSUeCs4C+ST7qFWiAWnFYBNUWyj991Gwc
nbuDfwXtfFDftqtQloez8orl5mFt3nZSsy5DtRoZ86B0YM3RwfojIIMHs3i1GUt97SE8WcsV1CCl
5S5VzdxMUd3f0+FlO3j5blyrLldmTE5SLuhGbfVEtx7IFcbitfNA6/ndnFfp9TFKB89NvpJnX4fB
wKWn6rvIRxB1igyUmpDLTPP9/ONNpHRnH+qypbYbwvluZ3YQbpKOLkR8VOkBe2elKhmj/OJecSeY
5HnPJJ5NR6ofqd62smfUqNu3066HLuKlMJRYEgxllnXjaJDih8lRhPQ5DyCUnqa02k57wy1+nwP7
IP+qaZo9FRzqt/7OV5mm7NHsIbFnEBJdZP/ZK8mNg2l9BcLRlYDxTh+/7nN822zRM2rQP42FtWR+
X1az6eenGKky8isLbTOjvszJu5tfozq1fBUCn+hJ2JVwzvoAkDNnT5auui3tFjveqCdAER8kP+mB
rGr8YZ2JYEgZAhQcpurCzwNxl5f6KjUVcEtkz8RBG3FbtBKzLcV5QrM0271TUUXkUiduonM0teOw
JQ0sJDafbb3AQScIDbRPseBtIQMAW8AfiVXMnEWfjHebpYSUP5cVoD7F6D72lgqK9wvFpMexDIKr
xxAyExYf5CBtajwliIfSHQwT7ZGwgwQ9dyqyrOgA3bwJmpnBcQBA5AaxnROzDLwPLzsogn27B49M
TjGIaYakmAADhCAfK2ZgHDNUe0R2MadCU8wzmodmdKodz+OyB+Kc5fKNjYpGRUAFtaLj4sPKbYhS
gsTgxACNUATr8jpdeTiygau8kk7X/6thSSv9KEboG+8LSdHYrJOnmsAsz9WuMsznP0841M4731gm
b5EUFbkOBW7Zh3STKNcs9j4C7sUm09Xqc0ydQSCu6DAXTGpLIVwSOv+tK81CDMNX64lR2jshId04
pVgf/qibRT9iHLqTaVwWKXU00sbiBRZR3Qsi2wdaDpmnp6A+GPMWkgJKG8iQk1rHkblUREdjoFpv
LU6w0GsMk7nL3PNossDvp3eeejSyAbTz4ruJe5OQHQ/2P+dQ6P6gk/hMmboGUeNLHLZZRoPdlosd
CzKjaOUwxBto2xN+x5SNJuba2pB46RcqgJMu8y8A79Zlqy1Tcs4o8Irb0GP/WrxpwQ+bXjqlWagp
+yvNnIMhtQOCy3s7IsJvWcKLiNU/HhUXAFeS3mmWtlEbxalaKIUmbwt1PZ+3kJ4aVDtkZdAoq9Gy
+KoL7GhxKNwG31pf+0lpWxFKUTbm25Mq65q+G7CPGlkY5uctngcVtHTpBdxZOIO80nvfYWaqmg9U
C4dDX0J8za4U+lyrQuA5+0VKT+OA7xIgnkNG2hWAPxH13jn1boDvW12LBK8ps6qnX3BZjehvp4KZ
b2qYnJ0aDIPFBUVjRefOrIzKK0TKUAhZ2rP1x3YWS4BvTW9lB/Y/ICo99M4w2UbrxS0zbSip3g5s
Y6AawwuM2UJ2HgirKqUcyyPTey4036Nfk5VOFrH+OiuBtlhFCYxT3H0q64C+WO5k6AmFGHLEyTGb
c0eDzk+SytdnMP67CkiSWmK53IitHELf2MUmK+iE2F4jgkMow7W7ECA3x1McSmWY100Fmhc+3r2Q
wwDTaXSQY+ew5OvoWQKyjE/lrY2KY7nrA9AThU4mDWW5ib63A06T9AA7ZuheRyXcg8QajFpXCKIw
b0B6dujrrKHAA2hOOigJZSgksGkge5B/MbpSeqclh5hQTtAyOn1s/d5mvQtL77Zu7EFLBByKwiLF
f1jeofLu3By0bznZqVXzV5n2ZykVNMa+ZUCfM4OG/8khfSuxRtkMBAtzjo53n06tyBh0zyQvG0+e
917M16ZiZ4UO1NSGXIA9UQ7kGKLrTkkviakB1vMMPNjgcBnNTchqXVNulnlYuctmp0rq9CruqF5q
wG4uazlbDrWnZmldApr6uI1IrzWBWAQ/5k6BkhUFDvgOXO4bIqcl6rONFM8bSscN5rhOsoB3+7eN
XvUXkxjNZ5gXNzPDKKYk/EpqthXIwLw4lRjACjBQ2JgDjVNZd+BdxQlXvvhLe8XiGy313ysI39Ev
t5V86zrn1C1FXCa4YrzrWhAw6A9G6gnZARupfHCQKsOamLrR7C0UZuodEoKYaG2Qmw+/ygHUWdPq
g+kaxUHg8PJ1phe1u1izbwNi2W723y/TdK1rtyCAHmICdDCOBfvyG01EW1PCJFBB9cIaYtkzDgFN
txU7hd+Lj0lqbuf+kNy0k3EVMnWJL741th+VqWa6qss1sQIvswSGSKieP4cf3wlPJSb+DwWFtYDU
sdO/DREaYSruGC1LluU7Uso/tRTsfq4in0E7Y0/BleIxOBQ+J+Urk/S6zkK0hi9JdZ4c4wKYOLSK
DkaS5oTIQZfssTleHNKE+SQUGCqla67Mz6MAki17+PaCes1ZUY6K4ExzvPgf1OBQdt+jcvKRkyDM
AyKOT4vyYs/t/7P0x6wgeqo3ZcK0E3j7MTV36RgSXVzpy0J9XaSJDbLGBpY2AYEy6a9H3lVbwSL1
hJG+6QP70eIFfMkDJCTGdu1p61wejWQhs6fbyiE3OIcAE3aRFff3cocEoxi453XVzNLSKcn38jmB
cO4YsPno7hhuGpp+LT8XPUKYBowJ94sZtmEeW+BuUu2WTnNrDi2QyBR3nyMKnq41xd1rN3He57Wr
JvyUW9kE0px9CL1DDzp+sR97p3dDd4SYbCe+lNaMD4IbRawBnwT6EjIyXN6Fl1V6jhbgQyVROrRI
PqQuKPf1xiiNRb69Tm20rVA4/J/+24A0Ok6HkUAeb366fg96DG5Io+FWvVpyYdCmlEJnkY8GfANY
SvRjHr+yo4WNJC4bs/TALJ8WuEuuB6MFZiMITBjBk6UOcbXP8fS9a8FJH92dggy4QaSf/+S8bWSk
xWnD+cQliN4yapi4yrSUTozzrpceX+d2pXF5SS/PJoEZdADfJU53FdTx7ztxnS7EQDh3P+0XC1qz
Q1NIO6f7zPMX2GD4Aq+DGJy/GCZP9JTy3LWorm80lPTBAKEMH3cRH+z9m6x5uHMUS1TOK86/wa1U
O4qEEXolCd9/US7fFZgvJVrJGtkMwEdmWd6/k6xbkgKAk/vXXbBxqfW/Am7TLo3EUi8a+qMPgACz
df52l0meMRDywEBW6hAWupzSvYL8AzjwB/k93Mu2IONtFpFk2LgC3iWLEhXpkwn91lhjZlqOEGqd
5/aGXzJiVjUI8XGCthIrAfqpYwofTg+alqxCdMdg9RuQtPoX8c+/QVYKaaHnHRpdkpUdVUIT3Ejh
YWLozEYJbgcrs7bRu+WCzzRV58wWLlWBQjOi4VvSq1IyfcNyGTHwuqC74VGAIRrTB/MxzTsH5DRB
vntkc89D9gLqrjOyXpD1Ihlq3DyfQFkFCr/VVvVecvBqaqA3HOpIZwn0mw9/FqgGtgyzLlPSNVt4
qBB3oJxX1Ov+sf/MexnWOEX3juyt9deAN7gFsjz5tPnMX74DH88Kard4zzUa76rwvknqIWJAkpfn
geziKWDaGqvWmhLMlSF1JOv5YZPiQpj/cPAF/N8kJKzF5WPQ56b7Z4k//A2ZzL30xTV6b09NHE83
m4KA3dEnw8vPDELBYj7MbkGZ9MG2kMuzL9DoKfVPxrBJ6qBQaSaMAh3gik/pTiNPuHASpOIqIJaw
p/ayTzOqV0NoPn9EcdfsMdu66CA9t3fSsV9Jh+J7JSu+zy/ANiX67o7ToPGzpRuogILakU2xCkKI
tfw71ALUN3rrit2U0055G9iwsafs+aj4hzxIYSyNzp9+ZtqaecXb7j21i/F53ZkRkQzqfk2GnZHe
tefjCTk5U6nfW5jp4SGt4Nj9wC+jVmhXnCXq5iC+keMkQUNOlNZC52VMqy2I8XlWgewgzk6xaP2G
8HIsOoqZPw18g1fFJIF4wfLDFxe7NhCpj+ptTzb8B2v+Ti8y2wgjDZFzqYizf8rFBxRM+M7Bnhfj
hoWEP2AM3H85R6Msk5OpioSWYXDgXB8J7iTxhI7brbsAn2NgV1C3k8ZKnfMe8of5+PgOUYo6Kv6X
a4XfsMJUMnkcg7e5UkYdOcWkbARFZPP9+10xxf4DSPDETiMikz8G1pkTcWzX+0yTwH3Z35OSNHB3
PVbxiNTnoml7Jz+7rW/KEeVkCtzArCHPbikHvqJzs8PQSayP+UGWyazCeGMIReGANFVNI5ZlVsQu
ebvJ
`protect end_protected
