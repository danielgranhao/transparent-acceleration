-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
gFHYoB8g1U5gmHFRhqCcTwub5DxcFdtlTgf8pPHeVTAtGD0ANvGD+95mNhyFqf7y
CQjCU/Sb+0xokKDsr05HkS4bxolDgd/xlAHKT55CVcJLdxS/9262OS5A4iaEf7A9
F7XiYSiNSKEEElHABwxD1RrdgGR0jRvSLOhq/0pBw0Jm8wGecNuuNw==
--pragma protect end_key_block
--pragma protect digest_block
WJ6npObncJbPp5lxFD5WPTvf/hA=
--pragma protect end_digest_block
--pragma protect data_block
pjCtyAqSpOJciso7prjbNruuYuJSeMeCK/XQy5820/pqTqe0/2ydxSEH3G1rJTNg
hWqjezTQ3zw5QdG11sJn3A2BbSBC9Q9hk5rmGaV2BEQILlWmnAszt+mT7TYqf9Lo
g1ORV3QMGGASxD6tC7yoSe77Kz7PQNgV0oIuu6BFzPnv7R/5YTrDqKberFFeElfC
v/zxGtYfXVNQWbCyEqJ+LXa4WV8hWRt1VtC5opvlB/vEz47gHTso6ZngTmdq3vHl
FU+qtDNp0LOC8jWEN4IalHGrRiw6tm5yqZqi14xcg/dVjmU5H2bG3TcupYerwAT1
zMWuUMQbuZ1GFl84fdHuhMmcwMkGQlPnuBKw6iXkCEBUyNQuZxmhrPJjrN/cP4LL
cp6DX+BOARnWeCei8i09N3VAVFqFo3lDexxWUTJEbj4tCAnraKd5wCJf+2g7UsKL
ndf1rg5AgK95GYk2m3gFtLBap0p29TNYslJiDBuYUXHRq5hAENKwZSVv/OHaNaQy
5dJtUthSAw33eSG5pgYoVxuLLGdmhHijPoIxtYvuzdefrc79T92mARGW2UdaCsUB
md0mG39A+IG0TiZBJ9/jQVpwpTcV7tJvYme/buEEdJt6di7VqHSqouBxi381Nqqm
+rm5ZFpTHFbpP9d7URurkmvZHPr5U8Xh5ypgt7w0lpVnyxzQV17Qb6qCHW7idSey
I7Bc0vpt6ti4fIvXnq2qEnTu2NHCfL6SZ/89wlaAVNgdysF1MjXI7fZE/+atKEzZ
VBGcJFWsIfUaRwTE8xZcNL+E5WdDY4c/7FT9YWTn8eS5OctEXhJZdNUJ/sJBdxgs
+qvrsbP7VSAk22RFvJdG/Cega4pi2PxT0eTt5YKfau7C05JC205n7e6zi3nAk+7K
xwHjyIFFVMwzkiTy8siWNlGGnZ6zQvF5B0NoI7AjYAyvfjtsxThYh/bHAyMHGbU7
G+V/4UhVThst8A5CWgn5f/wiFlN0D8yp3ApdZgPn10xYCmH5D+mk8S8hvRsHb13w
e7kjTuF1PkRdW5hEycnuYwaKYGxlglqcAkQndsBmGh+nmPo5dpNNrq49zv9J7cpM
tV+lW1QsGysv5Ngm/2DxkwAs8r3tFDGmqshizgbi6EP0igPRbZ9XCGnBkou2Acrk
F6cItAP5oEFB1BDslNZal4bg5dKp0liEmwvTR+B0RVKwhbVYobYrJsU6ZD/opolq
Nkuk92sHb8fxX4kEOzoQTMA/e7hFriDcssj0XiqbNRSgYrUQQAyrz9EdTRXn2jb4
ar+YOsOWYY5k9dTfEqZK1gXsyFO3ibNQjRZg1HrtHycLG+gdFASCrDPD50Np6g7b
qunqGzycyygSfSvUoQZb1unXNZtPWqh+xGgq9ubxN8d+rOO4mi4YzDFn9cOIzs1H
oYDglKxAbRjSMctR8TMfaUaYXexIlhqEhA18elmXO8FFO2N4+IncbdaLsh/Vg3kn
S3ghI5bkP9/QxK3inN63foCryo7O4EhZAjuUI81MScXPlDYsyi7TpUBNze6XG2Dx
AtHu/bV63fZJ17fArFTPb5y1O4GWDd5zcddD3mmFh71JJPHNHYl/Ja9uEosXzcRx
kIrHZcpm2k+4H7AoQAKVypuH55mjU4RfC5mrRf6pFHZIL3D1Fv1hCWof3hOT21V9
pePF5zijx/sRCIX7AnLOOWVo5dfy0rpxZVvED4pZdZt9Wv/h81FDCkFmJafwK5UY
7cAB0jjb8O+tJt6CAJf1dAhmIqRkQDQJBghaV4I8usdvzTHDQCU66eiivmUFJ/Mc
s8/rifwEEDn94rkBlG9pdXqqtH5Diek72iDFVQsFw/EpShV/h6qsFmwVQsZeHGkT
GIYGO+bb9wYDZatyR2MnXUgfleNxTm1gc1Z0b6J3ui5Vn89r4sXfyeOJ6mKhY4p3
awoxkBBL/eKTig+q3C6sHw3CJXDobyrPfE9nE05jYgTmshFPPqzHOkS12VBK5B9q
whQYEoKu8j9KwQCxQqMuhMSZU2A0twGv9O5rXuJIgJ5+6fYwkTHMXQSqUtSqX8ZN
EErML8PcjqLp50IRFNxAb7Io87xEu6vaEC00FmY8noa1+xa+PEJtg4WViOQVZcWo
wR6+GhDGrlMxmNIz3SdDGVBAJRzPUYsdkUzLXHNAbeVBS4MT5elpAqQagCliyObR
It6a0/l4SKahztO6ycpANwtHfpyHxgwQV9YY/guUZmX05VMcuDM1uwevvdoSJBgy
2u1q/AxQjverTvwLN7zHErE9+fy/XmN7wzfybhwJbfGzO/gVAZySifyTL+nYC1NX
I6p5fCkQIz4fNGJ9ocfu3cFyVMvr2BAKIpSOQBdTfYCtZBfVtC4KL6G82BmK40Tu
DuWnCqyyVthYPr5rK/BEWOfOkfPGMKiyMamEeAwxXVWEYdrpwl/zwHRF+z2cHlp4
AUKRDQ92gyJ0GccWqKeNKOC/SeDAcECx4li1SglQl51ixEsRihfe33hQMXpX4YyP
qtawW9Xp6C9gQjTulQ6p2+gAmZENvl8PmVyXq4bYHajl+djNT5mAhPhWQKfmCP1L
cYrzjlGrSjqXvxBhwx97Q0ZxQFgXsIRnnWxTpHtOAwDW1FCmjD9wdXkv9NcFiHZT
tFQnMgpVI7Qg+jdJ4Pte6Vfl/jvTFhJlnqwjMpjxLRRWkhSajQ7ZTSNN38gNEFGm
Y0mSIN4mpdbElOwLAUqvPFSrC57gVpSxhr70hgU161J2apGf3IwoNEfoJzpAQC+N
GogOeWF98Mkkj2ErDT+M/52BTERHnkJgEaB3bCerD/VPGg9z+Lf6kEXjKWWyLH78
UnMckJ2Ilk10ucqPNXtNbvw8Jk7gpAnEp9TW0WVpCtTi/TZxVIcCQ6jX7Qf/GPCZ
X7pAuyRTafAuBXDNVNMd35hHslA3GeBMkmlMJ+KNcptoUbqmegnqv69nlHhETVMJ
7AjcT6Uh31a7grzfYrzfqVned8SKjtsAO86lJu7iImeZD3fN8Xrgv7cU3+p4BvpE
LEYAJuES1CvcOGbOLQiOCjggVWuCvivQ4lS6Bhl7DuhuN6hHguSUHRx/Npa0kjCv
T9t1lgVrgnY6b4/tRmZWjbbNDNBcpwf7Bi6WZc4vvymTdwRFAev5Z+aua0dlogbr
l47l+a8ygFA8rqPzB1Puezs3taKmYwsem0GClGfR2hbb2QsFP4MXAyMcmEavSi7T
F/Bq1cysJ8fdx/XXhhyki9Ulha8lYvM9fyIeOu+o20PvohNA1JktaQu6Jiiogh6f
OagpXNmFs2z4wTD17U4O+yhbcZdlruVT5K3B76KufCPCT4dlUgoFJ653ruU86xHB
hQGT/K/o8m6FGPEogq/Bse0bU+aFVe+OE+M33kXvvh6GE2jDVz4AU33wnEZtRs7t
kgwnnSWNiFhWb6Bu/Zpm21WriVHAIZeoEkrMGyPapF8wtZiePRXQ6ioIOLmCKbdk
cFpvlKAf+aTJ7hhWb7QVyAS63AqsZ6YdEbrDWJQ4wrUnHA5Q98RTXYcNjf+3mwJm
AuzDnYpDjnvQyuVdOoojYmYyC1k4WYZ2vaOpK8qRPdanMcBVlYo5dqp0R3lv8Xoj
CxX1ohyEWAahkkeJpU1fQDv1IqzGXMRhwUnXdBLdznVvLfBDoIB06b6J8/iju8hQ
dgnNVqJTLMrrHCopYYhwUjyRCvI5Iy3kHNnnv81N52clAWM/NvwzZrrQXuy5AI0t
eNKwD9FJ63CxWcOm3QxBp1PEQwcV3UPCJ1N479wEk6C9bj8IjIMMyhFGDLZmRdiw
0VJvKBswVYrcyoSeL7uKd0vFbUXMYpq0/yccqXsKOTCYqu3JBmsqc9kAYUEPu2UC
TqI5qY/dfRKYma+1Zj7kICHgDOqpD/aNymeMbBdbzwzJqUyFkXk0tEKAoLvbGK+q
gRDpyK2aresxDovik2XgnHHzSX4ezNkd4NscjTNQV+WxwFKRPzDkhtUXJnWvLCI5
/dxbF7B8/pZAhiFqqd6yvjxUtLXqPUObnJPGX6S2lMnnHpdbaRBq8BXPF8iX/9pU
rq2yghBz+yxzHY2BbKk+xrRh0vQ9LPZVYzu3EM55omgaTIpmQdQK4kOjgLhaPn2Q
2EKRRLKj0EHVbnGuwBKIBFCsYbA4IRLP7rcPRONSdMIrPLgSPWZrvewyqB0xsZjl
jy/+xKoxlwPcTdn9q9mENQXA0rX6TvIqDHVsea4jbNHlSbbyqfvNLAschEzZWlAE
nLFVaodnxah8pTesc8HlLRfYyVMYTODUz31qjSI14Y6RRvr7bWBelX/g6hUtqyiP
U6MrDLwGpwjJdH661HvZ45mjayy00WdWQngmu8ETGycONsMupDvCcAP7QBTdo2mO
b/oWnj2C9mWLXnCLcKdaal7KF1UxtTGgOsdVte1SSg5+AtUd14gJih7g//0h21El
fp1SYz5IcRFwoTo8rbakLsA/jEK1DFJIRWKUKnc12Z1drM0bz6teA2FEeVYG0cYx
XPhGelZNBeZLur8jQFN3/cHbxZm1+N4zKbNuXo1feH2Xn1jl0Gnvb7qkWyQzuB87
5//S917OW+DLDN13QujMmf1J5ZYf9bS+yusdiRfGPWI+5F3/qeG8vuiGN0TM+lef
1eAU0ErIxDjd5141waRZX4zAo6yesT0DiqHZbZKxk3hc2qqi5t6275GfdnjTs0Gm
gvcY21YaU35xFcBEB/g9bUItURbfHrwWtw5F/OPFzuz6kCMDJ7qzLpF+c29DaCIf
LD6rKcwxRt/vqSMVvtGMxqVq61ZvPpyKbmgjveTSpZ9zstA2GmIsC242CDGBMCtb
xpd54hlV16bnM/0iQRV8ZNfutfNDSwtz0nsXSWnC8lLp1oAoZJsAkvwOL0ThW0CL
FKcqYdo0cGrBTct2e+XcWLFxmOGZqUXBDMCWS+plzKnNzp3ONSt18zrKeW6nGLKD
hzNSwR7RLFL2Kn6vl1NBIJColsuOI3pPWBHscCJwE333UqJIDDMQS7GW3CmS6UWa
/mpbZReD1PBia0Vsnxw+S5jHrOf2JocncrYN45aqXUNJhzs70yyKHGi4V7MaVF9p
i2tsPafnIVyjQ7e8qGOynyg2cbjwy32g6J2GEWxfXN1eAIX9+4BRxsqpKVnSNHIU
TN3KhExTbwVX5TRbJ8P3K7KGqOlaoeed5DOzuTtbkV0XFLjGWjlysJTV9LY6WXhq
zXM8scU2kwK6196YwHzsuASxVgIzuU2dsiSPsxpoCpB73cvJMCP5nh8GSceFPeV1
JgOfHPnQ0fmAct5TNzj8MvImjowNWyq7fA9Im0munc2mXDQGh/qPQW2znNRe4DcY
8eS6jo50mcrVEjeBzA092omaEsVKvvmHNP74T/FEZHY3JNXs4HxmddivqRBfPHKo
iQdgjsvD5L32jA6jeBqQnswCLfTZA2N4NO4I5WvJXPqJ1m9c1lvTuD6nvI1iajY4
OqLkrcncHPv/6BcMIx0PRwEu2+fFUE43zIQGXhoPHlDVw7Ii2nshqH/rXRL6owJC
fyABBP9Pe+7LQdvFcY7noO2XedGV5ZkywmkcVGww7yfn3aBNPI5aBXZ+X28Zie/9
szi/ptFquNF7IvRzkjSYvxsb1WMcLAYJR4B4RraieDq9vuZvw6nd0DUOTf7XfYEd
TRxFZL6vQ92lrhTVL7tgTbTNDPU0hTKKnZ/Vyhgb3avajTdJ5ANoG/64TxH1VWYQ
KkAIkdrWD1iXRAlx6da1yqJh7KRlSbgKHpuMW9AOwNWSXJmbh9ldyPp2ijEMa6B5
ptvbm74PkqxtWsMmq/Ac1bvvc9k++iZfS4h0+QnnyCiVimqNCrUB4+SuIFRXASIh
Z9X3NPHBlUIS30P33muLQv3rSIV3F4ySAeQO71Fcjrn0z4ZkupgBDRqJf5MmnbRM
rB1NNyeJx+Ep4xPmapvJcMOJHbXneAzkdtXDYY5eahhAVwNeQKTzKd4scDX42nfL
+W/sZK2XUuhj1P1iYY1Vz/ql2P9s5dqRou+JjaJqAPLgmek5iqh04fytUGYnnnj6
3VLVZrUsVgVQt542RQy2nqL2jQkwohm/4RIyIFK6wuYafcuCOKxvaDET9sk9wBgH
q5JQT49lSiwmmzIcz7kJCOxB8m0K8zoCR0YPbnfFuCHi8n0Q41pviI4u89IzNfex
N+C0uUI2gy8//7S4w4zpouCnTIn2gkd5SsmsWsjRubyzo+9dNFuRNr89BvUPuQXp
YqRsUBr1IUXiXS/H23dapGjvVnEOCuvEXXhkStEPwes4GPtKrzWFRc2yq3zWIu2p
GgOHYchRF/XW6ZSfzgQ8kxJYopwY/BUPEndX9sAv3rCCNeNb+PRPQUHlHY12qFqj
3LM2Sk4+HJaeoseUv+sxgPMJXt8tKhTQpQZ30BXVlFfQlNjaEs/Is6md7ZYXrpg6
fVoiZT+5IvsG33AU6GoTOgT337FLR577RRSdH9S5NJpIMG/4Mqv6r4pAE7N2wBmi
xfqD0yy5j1Z9pHoVGoPN3baCMIT5R69uzzIUsIyzkFvNep8vUmTnZJgc+KwmqiBd
aQ6C2BK8ZASj+LIImR0PUDQHcHx5J588Wh3oCPQaphQC/yobuE3gLS0a6vNPSux6
73JojUNBkXE0d3CunpxQgJNHi2gB2wZmatrnElgAvXAnXPh2tTNN+fDlNHCAE368
kP+K0pdJsQ91kJBxpYa5R3W0UoTmeZyFKGe43z5R7YnKhUkGGdB4Vzgk3oK1lll4
2UVHc4hDGgIkLpe/c5A9EZwg5aw5kom8rF+jn/oaBxIIlkSrvDzD86n6SnZG93qD
hjIfgrznCL83Rt9lUNaJzGYv7qdGEUJmwnBvGtXfVdjEwzQ+d770xKHPi3SfxXT7
Hf99oxqd/y+wOLVsiw6IkkxndXII61kx7ByzN3BADxuyvfjkiBDz8dtRKLrj1fiw
wRNEn5n6jYyC0YICa5Uqni7hOFtbFW3ywcHv+h0GnJMT90zM/iIyx2M036WVVFw8
grxZAYZIW88ZFUNX3WxuTu9fJ74Qk4if7Ho6xnU3y1xr8h0YuYMwAmLnDL/zc8pT
gnd+NTsmq1mr5cpwvp1F8JFDCZtgz3NyKns1fGxTYLjU4wVkmAgpgCgMtpOdCrre
Y2fti8q4gdj4Jhg0E8wRtvcZyAIagG1bH6X8c4aKh9xe4NZZoDaEOMpnpOzxwPfH
H9Dm5PcBx73bFt/KWRHJUENVKNZPtmOdzPqm/UCrXJc4COq1YOgguatFchi8StNR
aDmisUzbpZzUPIhWdTndGC74wBQB8FJkNhcD/CtpXmahrrly9wr8r9ECQiBYgqEw
Ecf34BxGL6S9OnS4XJ26ZWfMXEKkZbOmIxNjkDa+jlPzMFLjmfsB90JJ5hwEo784
6jA1lc+NFxBheEPcjZGnAblfkkJFGyRVHOSm3FwZl0G1EmsYhEppe0HF0Njoe5pm
UzCFtKn5ArYqzHC7YdBDR501tbVuh4QwTt8yuqaqMFiO/hqHxjvmhd6Y+O6e0PF5
kuoqLhN3WoAuSwXfrvLT1T92qpcopqvtyDQqUBzs3eUyiXXbZ6ItFMq+F0fWsYus
NnHDnKUMXg1xitRGNLgmjatO6TX3QGraArbcBPmIchLXbhVZpDXW0B7/4GDp1Hyf
vsdgh3zsDlu78VOm+hxwDEN7aTdTkBzzOkz5OSsyJEpbFSIZ6X+JW5r5XN1mTm+B
SsqhMlnaGGQ9/3m1BlHLoQO4fzjE9KVJ4F+6jSm+/9eeKZIbIS+y3ooRYY+Udug8
n/WVEqtk9RVL/3F9j2q/7wNCgjpG1ammcAl5jTKsSdsmgrlxK6QMmr9unFogu+Xl
0DTQEJYYBLR7Xw8HOyP0GHUDri7AoHRG5MLho5ZqMz0=
--pragma protect end_data_block
--pragma protect digest_block
0h1JF69L2Jjc9XwhQpo4IzJXyJU=
--pragma protect end_digest_block
--pragma protect end_protected
