-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
PKTUXkJwECeZ4TieuAhLKHsZit+G9wHxrRa3zZGPG8YgS2t4x8E+QzhvcW2TLBjAyJBdWnJfePsa
H69yIOcGmt5z+WeZwT8YXpTZbR8vP1zN8nuHeKi/HOQNNoRnWJLvpj3YtNFkJn900H4fBLCoqe5e
B5fh+ihxJ/l/Qa/pPUyTZhPxe/Fzw9LOH422lu7fFNgHk3NZ9hD0Q+vpSef1tQtZVA2iTJX8CSrb
qrHupb8bi0526n4ZiKLF30UeOjOz4xnzPIH01xPyRjkZBUNsBVdPYUCiZD254HhC5SnWxdcJWXDO
qYFj/UIo1ozRzI4bWuiQyStKdZ0zPVaSqS4PQQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5664)
`protect data_block
rNtav2NfT2malbuyGg/Lj4vW83Ztn4KqoJsxydN+UogDQIR0ejf0xL6WFar4WFyqFk1pMqRCIFI2
At417ONikDzxDXws1l1vJO65rk2a1VZ/DADXGGvHzbgqfvNPtO5Oxs+KlCnimktC/fAwWVd1nKwl
wZcxDypBq8Pau9RZHGswI1TLMvL1nTVrPrCfydDowkzbLtrbeqJGc+52UCUqtGv0pGbiz8/XwEKh
URXrXw7Y9nx5GdNpHeIbRdL+yosn2R1v9AAYudPzt5kM7NvDRWiEAVUZjrwIJjoq764NxL5AqztY
VXmLZS3XzJif9hF3xauStcPzB0JaueZPy/E1iAAqFTTxfSUOl/VtJImoFxCc46a/MdWllS64qrRy
xAxx4ROKolZJw/MJjpRbjR+0eDmYWtIT4PCX8rvVg9/j/eyFUEMybQFrur0tLdo6X8yGtwRefm0Q
PiEWws9dfKmDV7oi07UkGzY1QbTZpyEJtLTAIrRJrgNf9WmOwNfbaavLkuLq7UTdra/hBiutLPPf
9LHZ3SoQw/OVEl1CFgvwprM43C2ljUfqzP6gw69R4sG+1pnHN3GMvMG/3lW5RbPgc23mpTNv40X9
1Z/UH9V1YispOZc/tY0ojnq7qzem1OZnb2Vzuhs33iO2pxdBgB4dB7yd4nnirzDWzJCM+OfNvimO
iAkSmuinxRpSwj51dgBYrh/InXSe1ldfufdwpc87KDEdmpaR4XPChfLdUIDV2UcNmVYVt6f1pfZT
i/C8ahJoZdcS0tUWnqNrEHYKy9U57irFaAI6nDQdZ/fZh80S7QcOKksl2rYbedEp6gadNbv25g//
KMfNbLHC4tDipRNs7AsNaIEMOmuMuteYiv4sIPsyQtPug6553lR2SDxuEIP7C2tNcjMRh+fym7Po
Q8CpTOdpG5AyxTUyiOxC7Nq++z6K6PDFjYh6UEV6HbFQAL9V+c5C0LNasdR5mSN9oz/Kf5128uNH
zNcEI5I2VSLMmmboffSYkqbWfGnycD87z2KuV81s1Mnr7ZwiV+eBq2chHTDpRMBmVBnX5qMQsech
+IudPnEPayXldzOg5EKEktRaWDtlhXJ71TexhIdyB86L9E8p6wX08w14okHaSb6Q+tHcpg66QpjS
Khbj+8qh4qpcnjmr7fzWSYHCLjlC/I7CMBsp876R/8bzvssYOXQcqSlHL01eYEUdEbkk+UvaNEdj
fWakOg+RPjys4oYMx66dhmgUl6wkbKKgF2iVhn1lllBn5Zi25CTqKdiqTRiybpbeynMIeliYF6IO
uuSOJHC4W3+Z5HB19/CBFfKROtsF50WdJ7/xl9/euxlpApqHiH4Sepm+NTaQ5hgekYDIi2bpwBRr
C2+E4c9vfA2Je51as8B5Mt8k5eft0qgcNmJ1tbiPBUkyOBmY0xKyRlE08al2FTqluokj9MK/7Pbz
ntthg8P0etbQFB3amV1R8zaA8gkeAO6kucJKMew4jr+NKTbhqJFZ2HsRC6Zm1zjK+O/k9bCvZOBf
eoFjKctyNsfrSXYiH/3g7lJgCOzDoDvRb6oFQZXgDHa+2X8spxncmanGj0EI0LDuc6o+CBQSqxmN
2U9acMs3mFnWyIu7HDzLvVQKBhPVA+Xui3+ajGJgFoa796ccZ1oz6m0xnv3GKA4WjX/HShkMVZzq
IC4mIKPiCk5vYLkwXfF9Jy/JNH2+3LwjRHMkNhBTyUbUjjKN/2nzDIVAvin0SelUBVt9ZmgBXh30
HcK4PpKBJr6lqMbLsOXDNGmmyT0C97Z2H8oxDgZr9rvfi+tiNIBfEISP/OI0MnvyFQfFHwmTafbL
9HXnATN6pmx5dVMcQuUxp+MJaaWFobdYO3YkZQMGlSxx0CexVgjVPWDN9Lb/4JvnJHL6ypNxRq+y
kR7hee5SDILPARgtbQVQyGwKamV2Cu/BmTCjCmzstXLubw4hLmyHOrQ0nTGszEGh9QR5UDILctPL
2TrjOA0q6tw1wmFjnCgTrcjw3MIqcKRqYCuzc+o9n84ziziSOCuwEmPocmHYZJ9lgAX3sB9JNk6K
lg477ypfdib07SdaSn2gHhVJTZbjJZQsISUAMTNatJJ8X1hUDgQJX/9dGcFQVXT9PdvavHN93LQe
mPK04kLXKsdVOaNFcoEfZah0OxcMY5K068vC0bKBFW5uuRDPKZddWY6AO/RINmO4prdw8dHjMNkQ
rXw+WqL5kb6+1+kQsWL7NsBTJGEfzdM+UTQEb0+0lwXblWn6UzB/5Q+2UE0xDzCYNdOe2jEN1dj7
eHTwDWRLYmgG2biwl8zUr17RhD3AGj1bnXOCbU6Vno3tUudkSF92aYsAPvTCCdxoPvNvBORqQVEL
xO9mwrCL81FhQB1SB9hkGUxywu/v1T7vtZFr1CYyj7YyPkUJYUEIyNf/7U300ZAfwk+QVmYZ/3oB
oeWkQpzyKt9jI3hKJbQZDoUGheYhdcx3Q6IOfF/RSqqXPdpzb/zSspDrxHiumHW8FgHVj13ap779
J6r4bt2mEYfPl2BbAoOPF7Qe2UtIbgX3r/TNI9QFiSdJ1ggTG9YR5q25NQfWna7m4WNi12qD7Sm9
FJu0QAbmNgHR5R/EbIWDQiGZE4vAQfpjfaF3RQax6KVXLvGggVcoBSAaHTmIX9xYvzFDmmOjVvyH
ZFdnxZJ/AoMFFmkO5/112sbN0ev7Kgny6e1MKTrqibGXubxmPtOZ8xh+y3XwCn8utMBaV2+JpQWO
tjdzQHe6dYLd9x3EOIODzQwlzbdgi21EaHq/TDLuoPqb2IDc7u/rHm3cDpFKj9/1HLfneAGCOodM
VGjqqgCygI8nt53nBbDvoQMGOogKR3Mg2lP51tjxFXcYch9QXvv5P1b3uXNZmAPWfsqmHS1CJXaX
96Z0ksVLG2qs84PhOVj+wP5fn1pCGBxWuFzYqZTgEJ12O8CX4EQEL/bvFBJomHA/I6bVpV6nANWG
f7QckbWpHsOSiFPG8YpLI69m1s/s8JCsfHD/O8w3ycD8GoMpkRaCk6XX/V0k0U2CFSitntnEAF+U
AU8Z9zi3TiXQbCjN1/7jlIXXicAZm5IImdfpn93PuYWHuTFDCVf2S8hdhDx5Tbk/DlJzWCO339Nj
AYkUN3ATHtdrHJSiKRBchmZK77Kc8C5TDYmJd2SMuED2auqGuQBbjx3Bnhuhr+e3vnt88wCZWDzg
e/Ci7aX+4+CGpgAjG30if/YA58w9EUeItS4tMROetqZCaphJ7aiCUHIdj4GCyHiuoDUMCZJkDkex
+TPww7J0Xihzgwx1zQucIDTUNQkJaZlb3AgoLij/EgHsPmtMnjgvwV1bjPHQNJylhYghKm+JYqpU
/vMnKCJ3yz6QNKO6hlf924iqeKLl/rTTsxWHWqGplY39C0XW3gsVQKapK+08DfQDggG9h/yuUDQN
tA8jrzjRNe28oQNSb7VVO4JucALf2n1urGKHJEKqv9rfI18e+2qAmrymMyly8dz1MPABl2XwA6BE
3GLXg+iddtiUXk5T4VAu0ImY3soExNx5O3IQvhFbh+8e0rszmh4Rm+RG0rhNUkRkYGyzu2e42PHY
3MwhysuerRj1YgT7LWwwANScv92Jd9QqsoVJI+WP/VN2YJ23ZFZFKW3unFthwO7tILP4HoZ59/QA
vH8FkfbTf/xBV52vIREfo1o4L4auvA6HDgW5zZVFlipl0Z8OUZFSmFO+cUs34a9od+I3LrdCJ+ZN
qyUZbq+4qK8J/+He2FeuVvj1tTet8ToVe8QqNTkVdFc9UZUz/mLJneFFJ/yZXqqHS6M/hxppjy7N
lFRtVMD+++a65En/7M005J/9fiJCgq/zxpL6biEe0MPzQFTfxw0qNQSllD49HoxjLTq31JOr8SF9
uW3LrQQWr6FPGCOV/TyLKcP6GduVAhaqqteyN73OTtF5206fDRcDuD1GuNRuMb4EBVcQ0uCHGEH/
JgptMgvUefjt++zXJ9YylRM0nFWQc4rYEmV+Axd1RnyVpM6vwE04QnJY7bHj42r73cpRSZX5hCkt
cQnnxjzCvtfeReXl3lqsHrEIAyCBuVMzNd/1vHMbZPoOLzMsxhtH372FUtYvYEymtbH5XYLcQ8wo
/2zgK9U/IX3PuwLtbtW0WYxbbaHNuVj+2LxqnQRtNJDU8J+tmJimJkkDpreLtY2ra0lJ53SaWMBc
rKRqNCY1X3kLlRFLSQvD0mREvnmuW+culMOK4DrvLo0H0e1jVbL9mfnFd051qjELRRKbAHW/VERc
QFiKEzKEz1tH5jhID3pjt3xcW16EzyYv8Ami2whjmvYidQLN9YOkA9PSym+wbrmATNCntR7fumEP
m9DlFSBSDaABfwExEuS5VheKKODJAmH+LE2a+iI4LD1IKrBmkd+RchS1LnZ78zCtxVWvExPGqRPY
0kElP7ZinfjAoE5YdtD/XkyjOTljvWcyvsO+tQNC6vj5S9eyW3q+3YHw8euevy3SxbnN/xBnTw/4
KngcjFF1h53g9Io+Ln1QQavR8cmwxzRVDUaVwTMddOJ7jgZ2wuto4i1m9wsHoFLCb3/rB5d3OxIN
JUyfyQnkvTilwRVOEodRKTTZRoUDIi9VnviFSI5/ccDGxbkZYcFOXIqf/LTvCuTPQwMRDMWfINlv
fol4/pUAuAU2GwUPbW7fkov7WireOa37qknXIfC/e4fEVAf0bMgNFUFUkisQ68MP8/56bhKOPgez
AB8EqDNvIwZeYFFUT9QDrovbGYx4N12vClJ/tgEzEj6oxAxGfOW4U6rIpAjJB3dQYa2VE32fcS+Z
vL2j7W69LBTuYppSUtc23nVJZ+yR4GkerA5LGsJVpvkReVTsoz8Yk0IrM9OeEbCMclnjobx23XA+
DY4K+O1kPTq7kukDc2Vh+EOhzZEbQjFRhuyS62gfHuOzxTeCV1BoY4ntWT+wrucz6gpfQJleNpH5
pFp11jhxsDdXDd++ozC7fO0y9v4wgQ1eDuxGNVkrMDAdkLS1hIDKrGPcQg69HuLjwsE64dQ3S5f1
OLBUpTzDmMv9BmkyaoDdWPIg1XrFnwPudZqj/eH+g+ZPuk5hWduHGENT0eva9d/OdTFV73XqvZ8S
nWVMUgxIYAME6B1w8Ogfdqw1oJtZypVC9gWT1Bb+gFxtVR3xY+2YcjzBaqcjDOcne2EKczwz+uZ6
Pr1RsQWW+d6BM83DOhRHIAPIGs6V1QAbDLr/QqKF+EzQLhPPgRrQSHjBGS/F7l6Qzwj4n3+SMssR
BKmj/CutQRBci4ZWYWVswalyPF/lCC5MEv6y+UnAOoMkcu26woohfS7lL26LmgaPAzhk/LLyVM+C
VeOCRZx+eiSrazyub25cqNZHC1lfhY5OO5kv/D7nj3Zswfh0HxFUj5+sP67Uhc9kG6V8z+p4OAj4
NClJpkX4i5DWqOyp/3RNr5aTLmouKqVzVWMBh6LJDvoFU13Zhv4stalY8+H/0yI733lYUDdDHH92
IXKjGtyxsHFQz4OhKtjdv9Qoju6nihGkXF9jAdqjVfPX7v96QHIsV6Vpt85ys4ejXP4VUJhyThBo
Egk0Xnn4pBX+amHHec0bl7UVz1/m4myKXC/CUEV67IHeMnG4Ok9XYrQHvkiZEClRgwPTJTDunPUY
zVZN+ddMi8q/btxiUISx7H/dFxs12BkWFV0iEKUInB0Tq/jP3Ij5rPCWBnqCl5oQQX0Nr/UaaFy0
zhaQ4M7KSL7mRlk1OMWh4zxTN7YuV08O7YXNyvvy3SM99g0GOs10hEsyUy44JaIyowwxr1n6qF4d
JW34fXCdQ58P62Ue3tcL6zCpHtVRRCO9HRz8k7ZZ1lFVKtUIExsIgQt3/nKLcdE6o3cZJxCbbWr+
NIpn2ec0etW9CZd3EBRJXrVTa579gGThWQMcPB6vdKSWYSbT1nXxdm+oo6Ofqz98BIXX4gUjDwN3
m2q3MHYh55Zds+lnksEk/PiTBXeqzCvQmGXuUBSp9LjYCwsyO5mNLcEbatr8LK7yrjDH78RkITq6
3j9/+8FrnVZGwFhOUp3L593IbfIWFqil6r5YaugQcmjkcKK4C1fJRcAv0aGbj0AzDYf3uhis2Ocb
JCbOLDJN/uBu5U9HUG42jJyLUJ4xHIfi447mpTz0oQ18+K3/tAXIztHvml7Gt406zVAoTsxzLolh
NGg4dYlq2NOeU+4NO8gBQw0HQ0UsoUPM6pM36IHD+ETmHVO1Y5RBeJRgZIv5wCwA6Y3qgXRcgA+M
KSxTSJACqkLdtzvP45R9vuTWS0I39NrH/uFr0DBP4upEm+JTkcQPCfoqWGFoM9mUY3DuZ+3ts2K5
D5wPhRkme7MFAQK03ORfWo32mtg28eAR2gGXmZTsf/qh+SEJINsYtOoxbn1+v2kd1XTK+v1if5n6
+TyMTBuf+l3FZdXGswFKRVXRO7HYLutRE0qDBija8cxKIzN1fYMQSSUhW4m0fAc0x994uNdfIcyV
2l1J6NFd5JHecVTZwJjxeYxmZCF9huo3fyMVtXfRiIJEeiLeNryA3nXY5Gc1/r0ALoQxMKXVRG4n
YrZjeGmfDEGLQwC7PjLwZJbncNcwdICoOW318dhOWF3ApW4tm68SD6q4cKtlt5GALNOC8OAj9rUg
oK4csFvspaAo/7TOwZ+0WkBnpNUiS4Wpki3IA4Aabf8cnsuAD+4IPx+V9buerzMiIwyRanWoS2IT
yfwL8N2pZs80DM8IO/u2vdinW8Wm69qwdys0oSQm4tMKZ2jr2cVthwhHlPhEogKties2rjpiOKw+
W2rh9Q3QNXCiz+u8XDqXVHLCXgy1rBLOe5rEnh9VqbU0FKQn57S05KO2jI6y/iZEHhYzP9ppkWXR
aS8labMAI10yvx8qk9x+ao/4kmtrT/hXacntnOXw0RRPN8Vu1EM13Sw51XEu9/v1wH+dk4ZUv5Ox
4lRwSFXMC7x2TbLxraxiy2KK3h2WfzA2fx45Dp39HMewFNlcXr+B1h1GmmdIcNulkh+vJ/KoP9LF
81WBv4v650cvXeAfq93Un5lw9JIcvZ4AUZYfOna2Iy+hjbznImOPLyd30af0w5uEfGerq/mD1ybK
FRQE2k6+MhU3p5jVLnL0k7JJFPKXb6yvZypCPcqez9nuWSfjed+VnDgd+OXutOcFTap8qw3ePqKA
aAu2jFoWWzCh79eXhIE9as4biviZ5pgtVvaBR0tjYh345qwfAq2+ik/T0D7s8omdM/QEw74sX7RH
1N7UgK9mb3UFH7WrbdcrO4+u3luBNfpGU0B2vMBOnu3+mLbcMs1D7Ze45PHXEzpnDv4Ti3GguEPw
9ml5FkJxeUmXiauPA4uTi+6SCr3DR080bBMK9c7cA2+5v+100hEJ7llA/NJizqvB8Xvt6EtM66XB
7iTNSXmcNy+ps9Lwh55TmdGXtDbHuAGRU8IaGWEudtp5RTJYnoKzSoGnwRqdFe82917FT07d/r//
GiFfrNd9ty4+R4G5BcHRIouhVQI0uBi1+bff3BwTr6I4scu1D2Hj08STXqI7cTYFblZme1Xd/bdz
Ia9fGRCRdQbeZsxthKl3xsCJpORC
`protect end_protected
