-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
JNJcvL6OS4R89OmSqlsbRWSmqjQ79iwYWnzrbjDcuyp4csIECeK2DL6alsT0+bVt
8Y2oJG0DqPMXvZBv/pamn9lhbuP71dJz4LkvcZnqAwaACd7B3waqEFQ+E8iWyK5r
63AnrYAmLSn42NMwnhjSyHr66PijzlChnpGtWv/q790=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 81689)

`protect DATA_BLOCK
8A+lZ07UvpTkMzeDYSf9Z5ZM5OPE0e85FwlDHC48Jp6JzqDkR0T5d3rrpxKBiV1D
Ze4qy67mEmFa4rnn4xY0mYnn3aJAiT5qRQJBANVW7HwL1OG0c6y2z7kPy+Y1YsRP
7eLJBed8/SPTRvzNSgTSIxgmfftuW0Xcts6tl3ErQ2P3exrW+DtY2f8JKb8AUgN/
Mwm51SuIKQmexTgM+p7FRkpp3vUOc1qjItfaBhaz/mfuCXmjOSrizQXan/OVdvOl
lg6S06frif3AX+91lANkXIXgUfJulQVvROPNlz2HLo8PT2sJpyAH54/5ehsgs1PC
6OE0VgBm+V1f3VjLj1Dfk/aP64OGtM8PCmtz9GNZs4Bt7uiWXY3zhlf0Ji9Ko8Tf
tnnOK6rtx35+/pPL8/QRuX2xtsl/SYPZUZJni3BDCru48G1n/pjoQ+YhF2mR7h6e
Q0lYMwnkitsAwdQPxx0rdT0j6YcDX5mLyq3vuDnzJ3zaJc8Zdbpk9moja6E6xKlu
+XjB8YSlr4FLW5hVSZqAdkU7OwIBoQRx60VJLwKYWRcQCztTwLOTt8Dv2vMn7WiO
SW2DqKlzXrnSzZd1tn+w9aIKiVWaNLK+4YuE0wXtAWd3y3I79Z6P6Sy+7wggbJ6K
PT7vf80OxrvweDozyrkK94lNNuBiRoi/tI2EoX7KgG/O+VTvAkwkhcoNaGarKUBR
RdwnHHekDUtbYyRzl0605NTSNUgt5bxyYE7VxcLioozc8RlEip+62P6t35tSSvN6
RjrhpCyeuTRzgzUncm9oTvb2wMTV4skqmkoR5zicjuylFo9MMiZvFW3Kii9LiVxv
uUxu9wupFZnxyVJYxVGZ0hKkf6e4u+ch20BoMrKJQLe72l9+b388LtxH9bYYqEg/
asWV6GcDnldbonis+JAZ9UTo5LyaEhAOlvHPnxF1w7m0ZF+Fjj8cIqv2F5k/UTEq
5PVXFxmxnPMWCyvDWhXA78jixRtu1/3cIUNMYx/zC7Iz5NO2S/Z+ukn56X95JWcS
KWrd1QAkbQpbZittICQ756rtM0W8HyJzgjHZc0tnCfOeNDnc0U9C4I50oa4iP6Np
K9pJuJ+I+IOzDI7Sp+mb3ylvd3Z68nXCQw+gQNVjlYIha3gLvUPJSxvZ+2zjGYsD
bw8FWQlyGBIffXwCdQxkgnhZWla2LI0W10zVnHd4DWDqfPGesxhAy0h3mPDG4cyU
9bsN7akvPIs97BkK3dRmvJkyMhhqXMRvCCgI5e6jDm85afNm4eEGCq2kEWeOqHXo
UknsHpGZCNK9ww7SOfV9S1se7atTDr1lkmDgFNzkJVWSvRDgNp5/dvVFSyRA2o6R
a101OFOYCnNuJCszQFOEeC8uUkonz28XJ6EGAkveN0Snr68e76+rdCBkDbIgZLkL
A3PQXW3hulkPhAgU7DoHHmw9cBAix/FzFjYGqELpWERDUp8bzvHnZH1aKmnZDagv
/iszOK/yDh5gumOLReO6A3qY/9/VTaKHKGCF991i9Rn6ZCB86H90u2MntwL7LX9D
c/SSxcGXRDfy8ycboR/FlR41/n93RQvrjhrVq4E8Asqp1P2JNqQ6W7Y7knK3Oqlr
ZR1pv13mbU8e2kt8seWa+zj8P+0N/uS4xap2UeLemjTUdiKgdFczBzDsuchTD3kU
A4Uci44BUq9E+XB4gH8jyYg/bRxR5u4pK7oMn1emCkIacJ51n24w908hJ9WLZCnH
4YfRzupqsJ600agXbPX/M+rTq6t6VmbfKYWzjK+CvGAbdjVc/ql/1+0GrcZh44Fi
niLwhjIWcHH5r1tsYGevb1FQGf2FhAk/VViYQDVjsMG5jtHsKsysXyDqmi0OfOhQ
7nYDcd7Ii1z7DW1Wo34t8/O8HJ4en/crYXX1O5N5+FESy/0i0NjEFqg3gVHyWGOx
0OAMO7aNsNxJt2l+DeTlMDMd+rxUC5ea3ZZkromcYbXONjdH49+LoL+MCtdHGrIb
UthFDErtvAaRil5ij09vNanoGQbvWLf/e6k87h/6fha7it621bhGCoF9QICDwB4M
Ij9d7hB0X8eLn/WMQQLLPWMpSOGut0OhJ73rM9q1cgjAmK3frA5aNxMHFN/SW0Zk
Kn1l1SDQsAqqVyUUx2VuXZwpblsusCCRYvUJBv40g9czOMup3fWQTofVEaPIBiHv
ObMpPyLBXa+dbJ8cEt0tL29poIFqPWfMlkpltHZoHFF5SVn7VnZOi1aZUnBPP96+
X86XRjfpv64YuZW/4NXtBdOU0/Te9bpoHzWdngvV8ZFq3ZCktcwoFWyYD6jj/7O+
qHta7Js0lbiiPaqaBt3RtXaDGPzwcxoXNchD3DfJYj/AEqtR3ecfWg+u1DX+QhW7
2LMsHrKCnOrBkzO9YUtm/5SYSI1dBgDm/iRIsMmlrgCQqBhLreMMTxmPXechz7+z
BGg4XIodSiw0NfSulnz4NGnc9bCJRzNidGRH1Pfd0MAbqKMNtgP9vux1gqpDVur9
IYy/2AETKdukVACV6FO6Aychiq0aQIwV+xtF+Zo54EcBenTN8NKLafXu22m8fz1w
zOsjVlyxpT76VwvUfaEZVna5DILFKWvqXxB9TtPWGZd7Bd+3ojnY3VIa8J5uBNZl
6XQ96837yzFnAuf4WoojttWbp2zDowJIh6zMIA3hPNCvP2YxCTZjff3H9lam96OU
v732TX9ztZ06AR/+fLhT6oD6mu7wrYRnjvAbTakbzmTsSeH0wD5XV9adU/xHj1+d
xoXe9gJ8e7yUcWTjvUvTpMz7givbgj3uGMF3xRF1n3KsIwADUkXTGnaNRgCOTO+9
5wxG/rNenaZT27I8QEBiBDPItcv4Qwg95oOeKjzg/NJZMlLdJyTpNgMm2bHUmIdP
YT/aPmBDebrsh46v13z/jfDCBFORuvP4G/hL3lH0KGm5T7a2MMIV+1l2RpuZic1x
U355lSZA6BpnZnL8KkSR0FM3oI1RdcH69CMzSXjJPL76xEpB/ssS3bpRMyxPj8tR
Kvdezwp/082f948mCGyPvD1o8Xil0cTBr8bZxwfsSBB7dBhY2TKNPLcrzSsBT+WX
JZJkh3dSrnMK4OTxL9XxtxEgmhjjesyNl0vPP92keBVnGD9ggxthgaq/ZX8yvTC3
6Sjs5BN2ePc0WFjKQWFbMEXRuQHc15EDDXcVN1xMkNFCq2sV4YYgHqsPpobILzaJ
EinkuO5zrp0BtzdmH1d9npi/cpoFhTjedFb6hwjAHg83lVhxf9oNR1x/royx6z/V
v2tBv2BxHcyyxdBUQjGmTf2bKvVoVk1uxPnyjoQvDB9N4H3mv1YfdCBLFXiDg3ks
V6YZqXVEYSWvU1LpafB4iaDE3jow5zFqu7lAjUt84mwDE5dC3Rl+eacnFmHytFTm
kPgxwh6ADsURNfGNs6CB1RiB+rA+P+loorgHHSkUym72sRWN3RvA7yRrG//SJghp
L4YP2nwuhstiUB0XmXd0J1wp6D/T6PIPhPpqgf30G6CKg7cxrN5dMczMpuKctQR/
3X/b9mUCyOZXoCOkWbHhQh5BMKEgxhO6QRbSo2au4VdhzOqX76XCEXaHlPMp4Uxc
JEOsBVwdKjnh4MamrtQTkJSv6wftxPb9jPpHFBeztePkiKB2/wmFoiW+qmGrxFRM
ILp81VmShiiYdtYPLYuuIIfUTpMQLtesz6eTFnWsKEFjjH+gt5QjfXx9PQf5vs79
oV+D7GNtQ5Njl+sJXO3YPOYFCMapb1SY26y4D6Q+Q9MIRQ9knvaX0uL1xmBga5LU
XGoZcErggX7ViXMpASe/DTsuA6L70wtJoEoqQjB+W7jy8OFUoWf5dZAo8Xx1Zw4n
sd9NWXijnrrtQmcQrBgdN1K7DEytHO/0eq7kxsDB2hTVM7g8omWXRFXmBWQEDIKC
RpJoNPv6LeihYXPYRRB4ZSgZB6JOSBPwTTygeAMBB93dNXNV0rNCzmFzNCEMw13i
L3klRG62sOD+GXRFADQiJ4u2BE5jobpxsxMmAkN3RPkGu0OKCayc/G9nqkPI07B2
KRzxKbsbTrB5jnUvaQiU4q5VFUoFOdVv+FPT6dGNpN/uRez9LA6fXurGa8ey/6YN
uQk3hlPW6NsctH6t8HrhsCUA0TpNKlvX/7m9yao5GV3vBvTvxsijbq/O1GkCQ+P2
lFRVGeObrqWZCPtULDFRnoNUTYV68AOjQrmC2tDUb1lvGM7pi0Q+AlCR4S+zjGgR
8BAe9aOdSfzYw7tzw/yZ19Vul0b+WxyvmkCHtwzH04YMn8+9r4fHF5bXr/j3JWVc
NSq/MlEmwuiE3KM4LGUOY/PCu0xpxhH8Qbg/N0HMEEonbxIhx6E6CUkmRK3RX97a
ZW7jTHO1PHm/VTI9PIRqZWTQXjB2hLWarH8Rvv/YGVDY40eVPJzfe9sp1MLGaJAN
FjTnwbzjM9kYiRQKQyQG8CXojeAlrNOaGg5BjcUhdX8962MYkVfQXFqH0Ww6Wm1U
UmERXAQjl1Ho7EGpYGJWYTVOGrdyDS2ydTPyd0k6dS+rgeYof6uXGQ+9fwGIRdwk
dT4PI0HrcISy9hhQsysE2hbJfMb1uTj8SGvOhhyiAS6g58v6TJ/CGYuy9kB2uLzs
sqbJWdk4KiN02Sn8JWYwv6bSH7ZrY+wyG6CtRhbpSN5MF0SY/FP1kM3z3W2JEi6J
c2tQ42ToC7yVsx2LlJ9v8XCcYZwgeo+w1TLzR6xLvQVFzd6g9AzyQv5gLjnh3rVi
cEll5DrGbVDCb8qYjz2EuLAbGAzCr6uQLtNEMXwvuQyW6u0o6/JAzkRHcj0o/ARE
4Qp4HDBIat2+nBN8qqcWSSRXLmDLeRn2lfWZ4Ap0kmVkvx76RQy0+jL/m0Gi4iCI
Tj+Bqd43ST+nINCNb/Kh8rhQP/PtxaA0fObj4fp8U/dvaM6R2GSeHekFBELbFL37
5UMjCc0jFUiyf7rE86xLYQrHnTjPlAuocWqZbM0YHZInO4kriDPWLbTIePRJj/NO
WGuNlUbF1i6ISEA45+PIO6AvF+VLixrJZDETabG8VUSZa7xHO9w7O6SeXy6deNxF
29jIiiBz6IMMYO3ujrulzmG1xDRrAI6b/+M8GyCHXFR0YnUvnwiRGc40geUw5y5h
5ySkJbiCYrj3oGvKzitpbuQhECTntGNmkn3dHHB8gTO9BMsx2XY/TjMHcsBwzcQK
lUTc4yc35zjmjH0yR7LS2CZE2XkHo2hTDCcIGC50Y5DJHH3j/qjfBSlZGaIKBCky
1aGt6/x5XycpB4F5aHEcyiUNt2VubvT3DtLEfEGVGhShhmclmeaNcxQHfmcBlBaB
/zO0nqlh7gWO57Pa1l3bBaGSS+A7jXrEIV0Fsx7LgXJ+KrhUDneWHl+8FDpv/PXB
67hFLOyLT4kCRAjnwHKSqmUcY5fFReG5YqJ4OJkQVMAmaQOs1HBcGoUagALRuHE2
fTt212JxQ4xafdYPxEbSTagWRQmRMXry7g0x1pQHjphMBI8nHtv/cGWGqQCu/5mk
p3oBRXxsaJO1ZcAOeB6Mr9b1NeuZqfMlU38Pa0hCSzGxxZ08okB4L6OS/ZXAPvRB
tIDecElxIhTMa8UgV/hN7mjizpx+3kkxuxQ6kfQI+IfuNtyc6O648gYN/esMEZUK
iEY/oWzlZoU8l/wYWRLzZQXvxpn8PYBenaplGVuLLDTKMmSgZ9GHi3gsB8Oi2vzA
Z6q1/zziuy2FlFrx4AN/Sih1b0dmB2xDBsiROSQEhNKHRo5d08ER42JKeZ5IK0Fb
XzV02a11xydJ/Iplz1s0uf2u2qozrfUCJ6Wq/m8PGgH6VIgDqMDtkA0wG2FVS0oj
B8SVHpbV45gmUrHmovna5dtvKHNU5Mq0G2/M0jXGeLGui95XqgLKCj8XqGnJ6kP8
n+jlOdwE04qzbEhVYJ0hcBoASevAPOJL4ampIOlBq6seM4xi4XaDt+Mnj5ETtsnu
V/Rn1BoTbRN0RI8yGw64KjyPlPGziq5MoOVEILkoasJs/HuD/PMfmV1Xf7TGeh7O
TjgyMy24AvaOaWgWX/pzraVLkC2NCya+zs9ff3Am5vuQHhvODEYjVBUAgKrH7cLb
ymfRLE9tiqBbWZp0Kj84KfToyxQCiVBNkoTheHVKG3uakQ7bh9EOjRnKxLkqwL8P
rFVHmpBTe0GKFpXstCAAKkHq0AdN8CsaDYIG3k6HpGnjNUSsgSU1vBVLA/hQjjMU
kOJ391/6rwOvLVNiVOveXPHF97V0CNjhHuk4wVyCW7rx3pDQ2jn0IDP77dPVopfe
rfIfBeyeLmKcGvzdZG3300tRjrOgJshyYvpqi79+ZcuhFqVVqhmzYKv7pWE3HX45
IwwqzjEL1zlkh2biK0qHfY4Oao6aaoFCdE4hCdVAp9Mc0OiFHaUdioGScYnk6DRI
8cjepjixHcgTC1yJKASMFUppGmDIz9XyrkTVLosq0z56wAoU48RkHItESZq0C+EO
nLMKpKTxu5hFgZ2BDnmYgfWdwl9J8c0N8FWCbhwRchTDmz16yOAwGlinTNyMobEu
NOzW0GCC0pTvd4QCPkOz/OjUTyxeh3loLRLXNggvaHEBTy0z5i5ZrdizVEMZOi+P
1nSayLU2vY1p8zyDSZwYxdQjeRpYYpi8iQ8KTIgVUsdzVnz5lSEVp4uKrXoBg4qr
oLNoP9naN+j0gef+nzJGmSyQXSbi8Df4R31GM/6NbxwlqbPIQYYJdHdlTEEeTShf
c/ep1y2Ndl1IppS28+Ukml720NhY8Eld8W+Cn0EL+6RprrF4CtSjvGQ1+t1bs6eK
waZ0oSoEvEMET5GCRvMKzVkEqaYvdZ/Itqa8X1XJYO1MW03anHcdeEoF/FyZ+nM2
3ogEVeMdG98oOQaHy4Jv0HCTDRxkX11Z3dCLR+7dDpC9jMetToRbXOkI+nAOAlyy
+bcZemmeTRgftbdG7/PQezNBeFeKoZx5uLcoTzac5zxTl5mVErRXYVxPdHfNFKvx
bk56VwNwzUv0dgUTN9EBb6nyKr+egJcNGOIbtoAFOZU1rnR0qsCZ1r24m37kRPLx
AfyxUBBd0KNfNIGfCPe3t+BC6KETrnzmFmxc4HXU9+7wSa5GAG5lAwuqQadOU122
RujGbql84W9gikVtm9boIKDxeLE4pP7Z04fBn0H7CTrGsN8YBLKuQr/uVbz6vhmw
gl73hvMKH88/q8wCaiZnhUIqjpgqgRzZ9dfZRiz+Ew8DytdHaBSRpljjXmx1oVF8
DtufJCUCAa3SuV6+YQZ3vDtLCt7K6zkqgL4qN9catvZvqHWX35DVceZtraOuQOK+
mJW2xTYLDT8QLQcsmnBRjz3wr8J2qRSOGbOEW07yYeinh3k5oUmpALurPT8a0H+5
+deilJ99G72r0loorGTPpnES1kGzRxSEf88XWZ1hHqCNEnffnbcsbtnQSzWfPNi6
tDjr8Jg857zkMn31uUr6OZxgOsJTB/rOINUk4UvTrI6dyjID77LJvCv+2/xvfFpa
gJD1Pm5396YyBRuavmB3WRzNIctZ0ViwB5DZOB/vOu3QfcWtytpcV75bi0i/Ixbc
dN9WiIzS5767mq87fG7Qy18neyARibzQePsvl+FV9W5adyb3B756WFqxxd71j3jA
YlrJHQiOExbFXfjtGvzOxQRgM7jmnUH2sVfStBTLo1ZWx0ohcP/4PJJlEmvoYhUz
z/t2gDYhsdAtbIfTByAgnokGqMDY9fPf7Dpx4vJmgA57uah6gn8NBHKcTZPrW3xW
t9uBccOYmx4Yj42iAz74k2sjy0SkvUPypQUjOZBDD1gK2Lb2ay5OZCanCPuC9F6t
L6ibDpVKlkVEIH4M/UXFiEzJcF68dGCjTRYSUzBFKVAUj3jHP189LYSsshIq7bGV
X/iTSCXa2iQQiqlgC5SU1r1gdvEyzBeAAoH6lYtFChd0kX/oYe/CSlBtrm5cDFrj
NlylLizIsf3rCwQQfEVD8mFRIDI8tru5sQcbDbf3O1Ts4tiRNk9m2D7M+MaCtvUP
v24u6s8mfC82C/dhz0E/Xtbuu+Z/5TW0mKyqGMOEPYr/NzCSnCvKcKARttdkoh26
F2ZJTpI/KDlImFoCRsx24aEtzpKVxlxysu7RU1gRBRT9xF10Ahwbw/7GAFscqNN+
hg1UUP+BaKufr95dWnBx+YEcHSjb6/XCE7NSukDidx6JbGGsOhJYI2MHqMyJ0hgh
xdNaM1RdlVqEFMIvMrYSFoNM1SUgg62xYdhqiv/L6H5uspuOuveq0VHClqOPTHFS
sBfOHs6jkTeBJlPEfG9dTZUCV3hvh69rDhvaLG/vGbxxWerGHrgj0XF2hiioIYdr
xOgH9pNneRDVOXEfxnPzSu+v8vVbn6tITAZJl3cib+snwOzT2FTsJTS0JTGOyEov
kKavZdkJZQf9dURLVsr0wpEN4hrU25D2Z8XOmaEcK2zUkENrj38DtiRSk4eKiCyb
UBeazxh5dqt/cDwA/rTaS5YXuP8ffWNdUXJlqMt86WxKBRaJJpKqd3MxGHaujqvj
kX0JNNPMxLjhh4gMB6DPB/w5RKQ2MWQGZpQ805FQwaVl9gn0FHUCz/KidxbhQcwD
wjnszGaWvyWr12t1ikJ+DdmokgMaOtMZuNVP4Dt4SDaoAxtK2zUoPHObKGi/qvGY
DhGjj0qjkQL/J3QSis4XPvrq46KmGQOVZp8PGSWV/kVZVo71alERdjiCYqlCuiH0
H5yXQwBGLoZBerZ5L+KuvpPRoSATHYriCYV/7Nu93ODroQejp/rhn0ungBh/Eob3
dLVKfXGIO0whZH9vC9iuHTlL2eRUIoi1PFcLLfrMuHpsb3wAkXhzg6FO6Vwb2ZMd
rMNpOxvV335Gkkg9mh3L93K9yUaV5FakuNbspZLpMSSnIMSk63smFTlSUlrzvpi3
AKbWcKnBfzWJYRiADwxw0rpvGJgDT/HLRLUOgR833iUK09vO7ZF6a6QADM4e/bmp
UoC20unP5edDcgZjJnPsxVnkJP8Lrv8BY+rpSYHEuD+NuJn3cEBm2Z10lvBK6rGl
VwyIYdyqtgA5IcrGFzKyHea4RsYX1rhbQlJ6/ridbskjP+jCaIOuDcqShJ+hYw0s
Mpbm2u82Q4DBRnykNjzyH3Q9mgf3feyYGqVrsQHkQ1MNVIcEnnEmxHQlSMESylfa
xYGfWI4Dh/y7maH2+f/CFz2P4AvZiGkkgmfoT6PmraGaLT6jBfplrLdybkbNk7Rq
Es6bjfziOlfFRJOr57v4chfmYJloEbQ/d2DrK01Hs1X7krcVHkF2KCPTT8jy2krs
8hul3yl6qJ+lA73kcACxVkXTB5lVT6XIV+FQk+HZHrkOUNmvdgq3LMn2N/VJmPqQ
4qauSenSPW4k40H/wUHB+zvadMRzRESSFPbpicxTzMUB5bUY/Acm89rKHXe6Ky/J
LadQhxuzsmKu9y5KjPWFduh48RDEy8ZO/eLCjsbn3NPJvVll6PLihEIug20Y718W
mIJdu8jy5kTlHyhg292ZPmpc+kya6oS/w2l2a++GjKyQrvOxgXROCHzh6sSsMDVD
uGSfwzWJORQg1luY/svenbucLfLjpI22qTTlk5RcxeyW58A00VUXs9g1B6YfSVCC
OyWXxBykppOgXHwb/Y/AtVfP1pSXjcftJ3aF4vfyEMOKKKWKpN13KSF/UBNgTf5N
NXJDrJ2OyhXHbplIs7f/G+gYqr2yklky59i/c0WF6+2Qa/ig+zk0LvPkzguePf6V
GlIA5Wx+zZUr9vnhBzvAhm0p5VxOsykYqc3wCItjcaVA1rtI5ACMVl2F+iX1M2/q
kdrmn5XIW/hNxulnIXaLCvBiNkuwElWuky+rN7qLAtMx8o0rtTwOiU4we+uzU1eX
s5+/IWOEbU9Pfqc7A0EG3urAxheIHGzhFPC1bm7dEQHD+kfUqNrw17q5k6hgnyxA
gKRzmPAYFFBBbdphKN7DDZNHQP406mzed8jRKzH22D66HRcEEDSll7HL0/TFi2bU
PQ74v8pV0Iwl88WNEC3Z5uVsgp/XkGc8o8nAxFRceEL/dDXfiGDn6dwDhD2pbV0O
aOKZpEcG68DHb5uzLlU/K5VVulvhklOzVF9/05/8ok2F4XHL1NeTxEWhvSZcIJXF
Cm781Wvd4wUkHHMtHwJLp7y6tOgjUmWlxv+HVCbbR9MfVkSsu/vKc9yoaG+SxN6V
dp2Ua7/I+G2Zt7p3lHIvS0gfU45Bkm4p4tpxCby4bza21rYzDkvTMBZ4ovq1QZdP
dm48OLOwaICeTHeh92YoBKx94gkoOMvOODm9n6c2j4ISC+Ntdfz4YJ79oc/PYJf1
Eii1eFry5DXJZg8O+tNikl8/U6pQT9Q89K7RjANlb5Y7bAOT5L8Y0FFP8JU8NNwQ
iyeiqK1KLagGlF+dqsa8EJ016x7WuhTDOHN4LYkdfaCrePW189jw+yc6tWGDj6gq
h9k+bVBKw4+b0AvDTsZ3vHnKQTttYQH7UIRuYoLBFlmq0BIO9qxM+5iY0J+pQZCH
yZ1/PQefsI+kRZv581lbzZebl/03UWZAagf2xZaHjMT/WiN3e8YYJcCKRtTSu5TE
h34fEy4ydkKDa84st7Hfh5+Q9Vc/P9cDq1uuqXp4PTzUNxt4Tp9V1iIKuRYbPUTi
8jct8La8XGchx+t6L6QYAiqUhb5Z9fl8K5IrkgqkS0gwhVibJ8Wxzc1q2tfv2/V/
lw/II19mfWo70tDMW9MoLOhJ3cR1evy3xxXmQ63KQV9AVANXhl7n6nkSLFqDF/Bq
wj5PLvz5jjPQtc6Oag93Gl9wjfS7ZtJTZ720RVjijmrFfTZsFfw/ttglWYkR3MrJ
bX3kqFdNNkSeoOQ0JU/AxkNTa/IpZ7zvgVwuECiLYabI9mHCKuP3JtsI12JU01wQ
3fwZSZHHPyTCeABuSVtVZywEoK6ffdOAk6T2+c/qnePItcd3P0ZCjD4Ak5AwCfIS
0SL1JMAwuwefu7p3fpyAVzTjoj1n/lOGbqCaFMiotWty8iaecKP3+sY0EsScaeuw
0oUbOIV34JQ8ewDI+xXQkjkpxsxBAkGP32MM21UR7tsPoh7XwX6XNNbTwNQG711D
hXTNHi/yknQKRtdi5CEWhS7HVhvGra6Lwsympb4hsk3UohLkiriZjs9mdSy1PO4J
+byWpia1HD7ghkVcklbgwwcm/ru5xyJbjDhcaVajjxcz6f6aiG9PbnxSPRKKeKA3
+xeEK47dLn5chLixNhmKxhfs/AfE84F/XwTtm9ETdTBy4qgJSIEhy87AW2H0mPKG
Q6NJoVK1d8Dqneu9g8EeOKUbi7uMIJZAUEe5Gnt/+SJ0jMv8K4I6iRQVSwA57wsb
LxR55d5b7ZQ9nxgvJNkYOPTFGp/BXCaxbFZBWbdxf8NXgGEF5xhfjCELARgmPXqC
80Q+CtOYOFsLE14E28Prr7PftdZIbImcCE85ThfVdZzwir/zW2q0v4sd+rBG0qcU
N0/8wHtwLowkXAh/rh5MGppyQdrSKI6Yz4cYxqQYafsTSK8OsQ5MviEr7+Tto+Ku
HHDzv9wChojyGvRGxo7Bwz3bWOU6798efhpxw+6L/+UqzI9lFEnAb2Xs6Dg0LxaT
DVuBqsHlkj7Uxru7i05yuLa7C3uUrKTkalok0odeKq5osQVi74EcXEbEgFzyADPC
DqC4WLqpBvr/wzoizCFG0QiXHOkHRZZxTZv3FYuAKAeeIuH0c7XU0mbZJSQ50ChT
NrWt7ZOxwz4aaAfCyt3yHjjcDU47vNYVPBYfoa8DGVjlob3EyN3X5x9uGF5grsHY
3SBhGVQ4v91UnY6WScuzkJNoWLkxMZp7jUsv3xQgivCrAO5CMcVenPwuC91A6Kqe
gRa1UjGlEtzyxqzhxs83HERQIKHyLJ46jzwAc62PkLX8mC3aLgZmYJha/UYQ0+25
Ei9roHtBFslHmdPsTeW3oobpaoSxDNNa5y0dLjcf4//8zuOHHidzKM6Xdcf3NUE+
AjZlubUqAdSyWU6mjJkV5q6v1qZ9A4+evkRc+Nj59dhDOKj8FpXlMjxcb2+4ojKc
NIKEmBPiyYbbuwYz44SxILmVf5RuUYeHKHiu4NI8oCMffTFvE9sU0PDCjSIFHFYQ
MNYZTa7dr/O39BOuLbgQcWZQIvpAAoW+hRNttR96XhO0ZcpVKJj5Z/8WXmZv6KlX
CYEGffPhovFRTDsHicHrUX+jen9cjTDkL/zBpLedITH2fpi8DTO1Z6rZiNJL6LSJ
o9Iaz2py76sWQ4LGZth7Bgx0Q7Izg7PsJ2AGG98yANUlruhVN3kNVSbPBdf11x5D
3GMt6pttCanJpilyaSbPJds+jVC9+jqq/Ngb7TEPxMNsK6aI4dDTWc8cdWLB4WFv
p5I8pAJ7O+3wnLo3bVLXpXMYp2ILDak2odBJGUYDFUGweYtwjwZMl9z02GTi/cvG
c/LBHq1/HO7VewVtYkBwC4Bq+9VqSieIdr+YfKC5ws9NqQ8KilOOyMJJg6CyUahk
loGLn3k7L3ATPJHCDvLKYvUStXoHiZ8Z5M/mdW2pVa76ub5EHulfaCQhvJ8Uiwmx
zilRIOf14tN5waItcNpKz4xGMDMkdcg8xadEp4IxXT52muz807F2YmP5IIPaKR/C
AWQ+sEx0z2g465jc5wNlvX9PLHQ2rGBu/mmzLSsvKEaF/W46asg/ChQcL6KWfLd9
NF87+rUr6N9y7cwNltkGFn5FqHU+K35D2VONClj/rEghh0MT9bRxZDEPglRkGLmY
xe10qBN/l0ZLj8/QLBjpNAx07Kyuv39J052l8fb7Pif6jgZ7Lgxf43SqVsLIrr+G
84UvIhE9yPg+hDOYGIGof5ZE0aq2m8SOVKapVgXVcpanmDwT7FRXYUol9A7jxite
HpOF9naFn7Z+juLOR/xtmp+0438+FU7KLTXLh0ckc7MiDdsREud/JHSkfWMPtqJb
L9/SyJ61R4fD6f5y7cLZrO8LYAJfYDDAgXq13o27ezslANHJGZXt+uWNqtF2uy5c
UDoxIG5WdjMuywnX6DFiX/fFX1IJ4RSKD7f4qkJj/7AYbe7Don20Thso4ahdilUM
24OX9v0oeejVMeGu36u9sAgApk9wvStYro8xL2bebf2I0zqMW9fhvebwGJIR/nGI
yCD9qYprcTiMvGP3eOYxbQjDWK1IrscI+j16l+NDbiettyqOgnUGiaACgw/VRJ7j
6eKO9+sDnavbKu9r4equo+tSZIAdv+kWfvYpSKL8g25CayKZYORYpEHlsvmDCCMx
1CEZrhgaYMqNDI3cuLtEBOe/KLeEQc98A1KZZ0HDuO0Osi7CaMo0MmnBkGpJBQoq
DhQ1cB80k0jHffkMiTVTS9y/aJmH5Q5e0RSVibdRCC0EF2DE3UkxchKkwvVCwgb4
6FzKSYO49z7tkBOClpZRmoRy/4Ck8WcIUlCuePkgkhElOy2LvH0Rmza0ZWw1EHOi
ybOEUxRu+A3VB7pSzmh82Gh9t3LWf/s/ehmRentkr4fQDB5etiEW7wYa0J7ZyWov
/iI3xIrBZD+TJLAkPhbg9Rv7UdnVsymSRTl7kDVxVYJuK30WXd69W36Lw4Q6mcVV
Un7CgDxPKUbWDUiqhsHAauK4uAWj/giEKc9Kcx1PWp0UD61rPO2azDMHVDozNPHB
4+fnkC36CcEAxBRmHXHn5YMjpSwPEVT4C1FjQFAFAHe0k4dDP+iu8XoKNPaGNjf9
EW6wVZrftZk6+mFzMei1c/KHsjCYzTM5pQ4BAMFqfPQLbtJKi75KgbQBUIyUQBc7
SHR6yf3YPy73tB4J/UsVmDxaaTTIFOPoN3rFxDcX2JhBtBS9jcdwSXj3rt+nDe58
XN8WZflJK/ZcU9vDQBcU3gkpI949zvQK90cMVAMCqDihus7Ki+GVGV+6obG3mCRO
lJ8IJXRyUrANhb1tECwnPwRULDqPR92B8eGB6HKBiFwjzLzBhj+3Y6/weNHjxcFZ
qC+KjjTigBETr7gGP85tOvpNcTjmb99Vb+7uwFtGD4MxR8SZul66dsftfqhKXi7S
1e8BZcg9Mvz00V1gOzHrFjlF9Y2bdgKNYbjYneLW1yevWkHUWM5nEW0L0bS935jV
RrqsGXbKPb7aC7Bsk9tA7/H0AxZw68AFisTzswxl/R18NmLZyudH/bdkswXhMfHT
DMZxMWx/PFt7JcxNtIDD173WOZcUPsy9xL8A1jfHhyCxgb0rIGk/jGlz45BssDOz
514w7HOboz9AaVvLU9kVZmNyqglQWIf2eqVt9H7TKcunlF5WxQ7/SKF9MGNAzkfh
YETl69Vjv+48Hzp3HPX0p1V+HQHVsQueM5w/mHehMYgE5OduoYnYKEGGjUgMrAKt
iROwjcC5zeZlX2TU8x9j32kGs/xpPXK13HMeZCg9E9+9fCxpPk6mRxEfnx/Xhtjz
kG7SyAkhCckurc2RtlZU7zl9lZPz6QxNBe84WjsyCBRRS0xzN3I0qXVOCl2+KqS1
/pzssx/RrqMLvx2GcBTDurIeVznJVAPqXZHK+bjdH4sAyPBBdO1qxJfU6+3IvYT8
64DTbl1Za/dqScYF4drlMgmKWth/2rf2Hee+hyFtm+GB/0VYRzf74KOQal19PNKA
cHxx1nTnGcZqW7+N/9xU5yjMHAVOdMyVobp6QbKvmoJm++lgmVnSFuoJ4UOzK+xJ
fER6O8moJTcNUlI0xxTSih1QrV33ymyceWPszgtBry/wNTrgaBts17ifdM2rjvR7
3YjPfw6sQbmv9TgllN0XPxDHG6LKJ+iYfNOnmVj28Ajab4Y4E5dwZnsvBEALVece
URDVeSrjFSlxcNCq5hTmn13rT5jmb/wp1meB6gPcFbcudU0Lr+Avwe7lHpLYg/Kx
+eKT2ZXt1qzPE+Mq3fm0pQufQCCGINKLC6Ba8FiZ3aur7TdMfFhfQNrAfwVJvdFS
f7NDy21quBUAsBRB6QcKTL0NGaKqUQEet+RQbJi2GtztTk16ZJWYOSwuyg6P4WYL
5Ja1yVPJfHK/zkUWguf0p0o+aIDPh5k69hFnJp8M70cDhDxWxutybICFvpFNZETc
pUVY3GsJsG46Sm7w1Cx8xUP5Y9HLe6fh31Bp70wtdJbu1Cjud4+PX/QiUqauQDfg
e2/v+v23DGX7EHabpLhFbrxnLkYBkzwE7YTTQ2YCIdEX0AZJaKVSZNu2ctmgjBAJ
lqU3H6q/6LjEqkw7o369tzW8JcwJIvHfLQifEMD565loFciKFaidEV5j8ZuI/laV
ZJKNg+kTLByhPCUPoaEkXWUzAfMq9mffWv7eJVSJk6SXN3KpZKvnBKNuJAabsBLs
twdJ5Z+vx9UtvAnkCp/qyPkFEiYGsPR5XnQn3T1mEop2M8Nc5O+ihJ/3P9fcuSGf
oIUL+0o58RMk1I0/rHX0wh6mUyKRgjTpZigF72qFeZuGHGOX1JPAGm/mIP7DokZl
Pty5lr3Z0HexmuGVOtqYCFf54ByppHI7Gz568jj8BYR4s9UIF5X+Mz0Utlb8tM2V
KYQANxNw9+LlTBwlv4A3er5JO3iBF/cQ8s1Fd42tJbQshUbugfxqWPEwqbgz+4y3
LMgsSOqos+tWakgcQyY6dXGhqjhVePyhvMrLAqO1S9rMH7sv+atpmHupeczEk3/r
Xx0RPjC9tHqZIrDyeqiBc3SGNufXf4zFsv+FjtQ7O1itXOnVuDI9JPsvjZQQfUyW
1LkG4qs0FNw5x/u97siUscaRrWIKU39Ic3M6DBS/HwfwiJZAXXTl23mzcgd4iO9o
To58rN4tygyFqQKyetV+0zB6gf7UB+XM/bVyK4gVM0E1wWnKnkVatnbMqNMzAhAP
rhz11RTC9PAo5BGFzlecxLRWjCRM0aoi6LjLO14PSGMfWJ4ynMr2nFeXyMeTgB7G
CcZ/j0+3tCFHM/+VNpiHdBtVied3DnPG6NrXmlj4VpaSjEfJZyLFUqLgHuri8Gh2
j8U/qVKdmSg0sHB5n85HUWaHQ2VQqTB1S1/GPkTD8VRY9nnD+9WEscwlhiXYiEnL
b/z8ceZ5E2SPmGIv+hY+K6cE4YU6hWcVcK460//PkhNmKYhNw91Hetxte/VZEvzL
vpYE3yYAJk5UE5coONHyYLZfzksMH5oZ0Llu7b/Sk7VrS9lDryAs2cgFKiK+yOnH
StLHkcCTdnk2KL7o8nZPes9lsp4vbbIqjXj0tH7m+nS5CQxgt3Qbmhml4LfjbOBX
yPQ8Y2mQW5GTkV69M/3xW+ez1tjkUOar92Zi/sRMv0mAWCJHplxsJxRD7CiKiPbm
+R3ovaDfv6Izq/gL9QiKVcghCV0le2pMFy5m+z1J9QGljA8F7G1CMwKaby6h6HG9
L6hK3Hiu7Sw3BUZypBV9XKo5/qDRp0YvKu+UaUl8MDNokgPyiOXen0mpNRWGFVZ7
yVwk8f/jAXMlD3o9AFHTsj2PwXf9DKJCyZTNsmtrN99qX4ag1BEehzoFrv7LgKXc
8sth4ioerz/wKwRSF8mVudpTsKtUe2Okat6c0Yq3hBoHcJw2VeIKHqS+G1rsIV90
U/jukqwmFD3r61a8KQrRwzT8jMZhRuN9lbcyVtVhTqCqWwHC83kZmGwT1l5GPvuk
dsLXO5Kd5iuTTmGcYf8UBB2L+lPUDXx+3vKdxHz41CxI+w4zuNdFhhEn/ftC6TNL
gRPk4/duV3rEc/ePgfcC4kkrtWFfMzmeoHOZEdAI/12JfvCPuJFWdku4ML4WIvbQ
iHXRwjuuLbHeL1D39JrJ6MrpfB4bwd/nMz//BrEgOEG7d4NPcu8StkN0qPbLuIbQ
lr0nZU/Rg8EqkOPZVJG4zQrxXrWcjJP9Ik9yaHyKSHGR8A2J5f2apIVdGQ6CpheF
bk65z73knKQd3SPugwgwBDt/k+gP5cdsYwXpJ1lorUkm/FbDt3fZoqT9rBhTqZW0
VDoMxR6OcMo5cWpmrcb7LfobzSyV5Wk/iyhgxLAyTvL8x9pmxYvWOWvKprcOX/07
KwcQC6CGOc76x/WHGIbqJCNXbQSBc7oNAio4Hy1JNhwHMiIT8SqYgMkZQ76B3OoX
ghlpAxlKLmvRacwJ1JzHYWF8dMQfWy/wvH2db/5mmH1+/ieTnObMconIhRoLc3Z9
whtFmjhUE+w59N3c7EjTrXB/EmLCJpuIIq6o7ZJ4zuuRy3cLLfSPh4mtke3nC9m9
3Lqh5haRArCKKWijCg1INEe1s5R41xibBWobwSmg8P/z2m4fZr3n7zMkKB5tcrmq
bnxEuWZ7XFAseYSI2gEWqZabMeG1N1vdx4gXrEPX19C/WrLgTHFNbUF9jd5q6tjR
p727hEk6SvkuIBebB4G3WHj11q8gJtRFsAjdRi7ZnI9lN9V6MRn7o2APwxcVuqth
v7zyj8sYUBhBsRi0dYCTT8cbLYr7n6sMp2xGqBtQlGlmGj6oguC19/jLIdoyeumT
sWo0KO6vVxSaCS9roC/O+he8zbOml5Ec32nWJXoExklVFxXyrdUhY0v9RnL/a7Ur
yz2UMhjGIx9liibNgBaPBs30G5RTWEr3HTrGaJGRXeughB1wG6GzHF6/g+81jce5
+CB28Jaw8FtkKQGmBw6LnLuh3HRMyR6jIcATwsXfqLwm/4W/sDpQ6tXZMOIOpsyo
vQyK9do6CrBTKIATLuad3sJdg3Wc0PJLS1MxekOnc/36/0l6MoA/cXN8RTjg6b59
wBeKD5qtkFO8Xweuzxl/m/6P5qkABKIbz8O/ahPXIYUKfNJ/ITS8+tJj4RxpQRtX
izy85ZjP/c/zV8skWgaYSHuZMqFi4Kj1kH6HjZryNrPsLAtoO9uu0fK0s+YbtbiK
HcEnf5L8uQV9C/b+QG3GKkXcSUORZ3hEgq5ZmDGKZa6lX61Wk4GVi9yECPvq2v1K
7bK3t1CFpW4NCrE4H/EqbT1iiviPFv3Mfte6ceQ6J8Q4ZQosXjksrJDIOP7DKWel
UCXR8AdpMQgSFHxgR73/ikNJzFOUSuiWQz6Ob4h0kzg2PkO6ppkRFdVw+guhUUkt
6fjl1/cyhXy6m2Y8USgqDGUAzknuRy8SgyGkE4jdqTW7pIQzsCdkH5QcCAsAzHv1
rHFp1ctpQ3MyfhurXS6QCuGA2W/geMky1glzfp/xlzHcQdOUObrKpvJNcaPjSJro
imtC31YbNW4cG4FhbAInjjFbhQxKwudWt4svc45r5dYi6iZr1ZenphegGsJjX9z3
ZGxgjJjNsYi++UCeTIom84kzOK2ZnZpr80WJwDR/2581IHUKkmxUbdTPtoVGV9wA
7bPgs6QpLK8U5WYYWvnxkp6pbmOgjTVeejO/WZHC2sw+UDnyIqE/gSotogtjsTp6
q+tdCynAyU2smTh45cTDWuq14ZStMP1ycpPZL2viDvTgLhCkv6E8WX+SythC0ewn
/LF6BhIG6bwuRiLnaOLCgs8A29ZYKfF4v+id6lEa/oNa2lvR0GiNrBmpmLyCTSRm
Gg/nhAo7tuTeA3kUpSEbNtXJXKRUTpE7dSeauzxgQG85aAcVKfLZQeXhcczWxkUS
GkcI755Tni6gqdSweVRSOTeeIuJm2MtLjgsmuRHfON5Z0W2S3thN1xq3pYFVik4P
U6kZBx9ZWbBKCTZHQ649GisuBmD6YJgw3h2Ge6KXLQ49yDBwRq4D1fFSKOczRkpk
g56rm+fZpae/Atol2X2WrlPjKvE9kxRedZpp//0Er2OfARNpyUGC3NQCa0lGz9oA
3ytnOwzKsMTiAiyRz6GVjnAPNMGHbNhSajvZFzSECN2vkZCiHmeE7ajDa1GDVAwO
YV7b7AVt7raKgJGx7vbNiIRoRGHlZGJJdRCshWvjaXlNpLerJw3ESWk+p3X7Usd7
Ha5mkiLkv1hUUjuJSo5iMplyFYWRhg02N3b0EOslboavE6Smg050slcX7cVpt+U+
1zRMAdj3DI54UvFKOmgGTA6+VUNBoA/oLAdLqIlx/rSsmdZhbZfNWaCaJ4MK9Zqy
/8cD2d9NNEJy6y+lCkKVpLHR9w7WNTudyV1FBMSWXSGTp/IQ5+N5/Ry83/Ofu7wr
hjjBQXpFT59XSX8Oq4/0ECCzpHSDWpXSsdO1C0mGfLZIDN3VJK9DzMe9ObXTTSu4
/H9/d4r27moGp6KAaMV0Z/RyLUp+RKE4taRH8smEvLOXDXshasxrJXC6Wd1tF4Ze
cZOumA8ZdGKJpNx9lLhTHkxrzeAGEuhNeBLJyoD7OG+kibTqwmOQorjxoq+rD4s/
YfaJ3sLyTYeCUC8KxhFDqEunM47T1szDJOsNlWEbyb42nHYdk48pCE/mNY0VS/6Y
QZYkwvPBXGRhOvDmF6Y4NbUVt7ZFcRdyzEAcajOaIZmoXNCKpPKEnaArCNDNQX9q
9VaiTqgwOXI5BTqJYSrivCrMF1h1khbBbF9ybnx8Wzz1xQdhBUGXLml6kEtPdDt2
SSupnlNNnwKdM7S2jTe3NCNpL6uvOGXxlA0LyReg3bsbcBnUz2bozLCSY9a+FdP/
tBIWR6AMifq5mHAuJGGZJ0vtHTvFnIyq0Rc/X3YThx050fS9vCuZFnR8QMwiBeD/
BHT74WYx9rp8ZX8vCUChFgUoIl8iuWUNHeIV5nWRL4Cvww+QjCBlQV0bbxIakviB
VKo7ITOdTLWENtwPqX0PF6BCDHp2g8xqHDm190aLxqVraBgrqVzX2oCGoQo7LDbi
1VADTidEaDG36uPqAtJeiK+icaigPexjOCXaa0NYeEZrirpF0xsWcor1E4mU3JNd
kt3CMIKZEmg+EL0XN3daE0wWjCMMHL4nBkVM8szoVyxC4WjtsR7dlwP6s4/Wv2ye
qPpS8LIJLCIbHDM3hNZgZt9JF8f1ZWi6AEXovtKxMEfGlKKx80dokJxM5LXr5heu
A1Kpzjarq5HNRUfkI/ghZJPRL8vDziOlzHcVnjkWDXxG1ykIbqgT3vKcgDSoBxmg
odayLLX8ZAjxC5hUtPr3eBjt+oFh6PQ/5EDzdhhvR2XfJrufV79DmRalhfL/9QQB
k0dElpJ5Jxn++WPWh/Gxdek1jlxkT41axMjJT9Pjk2b+AO767OYIHSluCV7fpsw+
6CkH8RAvGJ/qfOEXmQKkHuoW0cm6cYoxhyZLFqVz9md11GKu6XyflIxSuwPSBMXe
tRgUOV2b4GWI4FHJz8YbO7tNgOVb2XS3UDqkvDXdszp8Xm9frFaUq1kSt/cxlObs
33zUY/h/0KWveXYC4M1RmSq75+l0E3ZXGdar705lcmBQPK7D6mAZk1HY/67oNnfC
CoIdupuq7K0wjGbEtpI8qwEk1QoK8MEcgTH7qiH3fbSqHebxzMShjbTxMW5rcDeh
K+KQOnwog9UMLl2SZjX9HSVpqZHqoYdgx8jHldpyjBBjMSnOEvYpgf44Z0XR4Ilo
eBZr06JLfUcocI7lG8dVnptWQFu8hLMffSyV2gHbVpvK+uU71r3G6FoMclZrSXSN
XzY44Lwv3OZ/S/bGpEzTN1DNANvG1sqYZoTYKSb+uUZBQsGsaUg9a7MngvkMIhuy
Tz9hPEYMd19kLbrSZhvltLkwoqiBEoVzUppvzLVzni8aRdtv6PQyfh1OtJN5o2E5
AT0IR0wEDALdE9B3Gqcsl+njx149ZJZCwtrw6TzbU9dbRdznf1PppwrBefXEj/0l
QPgdoPaRXAZnxI4PKVK8reuiOKhi4YzvLtnCXOlH3nFOV08iqJTAvUNix47ai6vx
0UhgUdkaHzRjDFaeIjmsFtLI0hFAUAC5Ij5p0aQ1sTWTd99KSV/5h/d7JZO3jiK1
DUtzuTOrZ7KzxyKP/KTHAO95fw1XmY7jNGiPBhsuU5gTOKSI33ad+pZ1yGtX1S3o
R+J02b865skOoZNLBICKEZXPPVClqeZcxm4e79WjWQYi3b4NIAH3MkKogvhHAL71
afx/USqN5blyZVkEzx+mAmFc4AjFTSUfwGW1liocOi9l55bz8+Csa9XnHL0YpJ7e
VeG04NIqfBEl3FslTnDGgEzJSEroBNo4RGl3cmnt0YeSIu17RKebfCfJ9LGTusqZ
0+fJdhpK79qn1DaFU2tXe6T9/9hoDVMmgSb+Urg7v7ivdEGBnDHc4PZl6tSLq7ZH
MvAG8qgw8n4DActk0rOINQ4vEuYIzBVhIGiOabPmAMOlvsP5x+1pImFObebcfqGN
ZUOnfYiZMQGa0itSfBIIwrYqDVV+KB1bnrSEl6G3TyzAWYvVfU4oDlJqwlg8AQQJ
UXl1wPckr9ErkPNqkKX31wBxCTk0zYcvm73tyJUt8AztbuUGFUuP/JpysMhPU2L3
shEjwy3U2AK6X/g6ZDDARm57+NO6PQdKUnVd/HVkVDahSr5bnBi9pVQPPjOHbAYv
ypWkbJTHnQkQ08GqMnH/0qBRob48BHUvVJNsHEldtmj21YLOHFok9IE9AuKGqXoF
5N5tGjoVOobPFGpkc5NJr0B/50RKuHAtF/gISdEGqmHKYFoIXBqAy/qTXisFxVx1
LgHCb5AAJpnAhoS1I6gx8ojRPZ8SpupYNz8CcGYA0dzunllpMnzEHbRnh3vF8zJu
2m4PkJjT7LfOkd/90tPPduljwYkmOYDDTgNE5tr5jgvVz+Kp+O0HSmKRnYIE4JIO
aFjJfLp/y9oFJhYkL5QoeMXfZVFVGqR111qkT4U9rHg/R7muT4JxfhKCpuzO+tQg
UiqQRpeMXQ9ORflhcwk60d5RF1oc4R2FS4XrLXQChPe1GyNF9+Y4KIDFpyIv9yW4
wwQsTW9Fbzw6kocwKeoY878eImi6RErdCo/NyzHLVzYrgJwM7hR6Drys6W9jycnA
oGtnrcGJlbksUeSG4kUbrDUXlTx88l62zlGB6HYGAGQPYM157FdlVd+N+fIXd/MB
3AHAKsIjwlYf+C2J/6K5Xkjs9Xqh8uIfJHZWQ8tku09BYm0wSxjZENvkY6+BxsvD
tFd4BUuALoZv4H4QM5WEPS8YKSCw1Q1foJdcNUxmKgoad3egxyPqhH85hrFqnW6N
IILx8i+ZAL9qZ+cRCHXDfpK3DHkAlLaHiveNHsUtqTYdxSX17PoEmAmglCqZ0/gm
p2UZy+8dnsRSSad7j6cCsnVXLW3voE727eb3X9Pe4iXPxgzAaiTtKZUtEyzHY5v6
uhG4mZOs53iRmG3WSoCPmWe68KgAHSGEsS5LA8qtklU/zbHYbnHt4H7mtUnmvNBp
2GghDRhm/fgpLY0S6+9sLgeQSTiqzKSEbPMRN3Jj24YQHpAP+exNgV3MUVZLUOJI
1sBaavYi4YpYB7LzGUoZ+Gabba7REVq8Ihner2MCWZLtGvdgU0yVRalv73KJ/5BD
FQhrbTJboJJR8Qs4jvGRvAEDUQv91EWElaupcQFPRBaIQtHFqKixjFGpqFGtCRVE
DrKf5hQUmVtHeTEVBcY6d+OE17app7xVuYPNTkYBWaUHmYWnpbzrQlu3yddLiCo5
i+wv7MxRHyKidhmU2vCeXi5VsB+PPk1qwpIWIiEjI71+MwdysYHTzeXQMng48JOF
zgDA6xWhbL0TF6ZvQGAl0PIAduEMZQf+BgzHEpeDSvveuSfJRbdDH7NiaJTUG+1v
Kj5ByKi/AQj60vXZW3UgHJtdcYzgPDMHZlNzzHYDS7DsHPZwj0iwz0Iy8O6Sph8V
a7xo55JoFK4KtmzaQjn1h3VYvIQc/hGlZS4ABnZzzP0fHVR2renLhspbYZV98hNK
/PFxRv6c3z0pFZJh7n8Sg+5lKEvxE2Au1G2NJdM7ffS53K+OdHGkH1xsQksiAvkz
QZt8zueF2rbCpS+6sCmneX10s8tYRSWfmrkliG24v9NMCd0mcPWAmBIOXDZC7IiP
qfG1ByXugDy8D9jnIz5zX1sX8YCTw96kirdE7bwIhDlDIiXlZpVmhEak4IkbuwiU
YGqPcy84xQdPAmdNiHnsZO0g+9CgGGUDGG9aDr47tGUL3URCImlUMUB0P4V9W6xE
6UhONkJ/fno1y0AUw5iUzxXbzgWGVmKn78bbiwy4KL9QYR/ORDqWx7UhmaiD6dPH
MSd0JHPfAIzdBIFV8CNIVf7lEPSrJCA85GyO/RMy+Nt8LnQQRJbO96jCsegtL94E
s2Sl5JXnIXwPqmWRMJd5ZbNx4uuSQhUgfWLpmLLN7Zu9z5jyisW8okLoGqj5y9tK
3Ln7PEovfFaJUintMnAVOCKKHxgGmwQEc0t7xBvoTG70h0RM/u+zK7EJiLOVEjFw
yzfcCux4R4RY/fOn0E/oQRPVU9Ot0YuofNYnZpmUAIEkqUqk+8/E14vuvNIXym4S
vvcvHMvBffqKa7BsECM3wR0ALjeEVHqWrDvOZt63KEwAA/KVHp3K84fzhYA6UIZv
WqTBoQzrQfd4k0GCmX67oSF2HO6m9r9/DYMbbgkjvhoGI8pGHGMw0r84SHZHURYm
tVuBZhs60it1vGON2/hKKsFBYsWkOkLhccGp9Mm5AU4MhqEFYn8TU3zm1+FXdFX6
zohm82nyo9xYXiSQMI3qCRXmu4nzwDo9hUtNpqEbiklD0RMk6dPAKsSH8hysahKU
yyfLN2QY4fH7cRkULDbkTvJRypSu2FwiWZcsadOup2Yeasua2aQ2xyoHFnYrsV3f
yMg2C4iFCdJUt6K2QNVGzy6tpDs7tILR5TFIR6tolSF98+GtwlpnrYSPCRW/1nyh
7VjjlUw54rFCXuxlsvAPnsObyGDIygyI/zj3FekmeAkmgvIzalYyHxxSBjUlmUFa
sR1HUmWvam0z2ssgodkYWo68wpFG6KWsvUjcJqfGtXGDWv999diTo7FHMLIcNbDO
mvT9yDKGlmDUyE5nTSN8aOJlnAdDWoE5Zwb1nAP9CItS4/cem8h8MTkqYjjbV/vY
n8tjDYHy6YAe2lmR2zCxWNwAeAsZpTfZsPb47LDyzIG/y/LXCwzK4FX/oExsEAx4
88NBWdRYAE/IlFwGYvMcMZ4ISPOTP1nLcHkB7kbvez/8Yp1fRpkflkntgSOhDem0
xvA2IdU5u7ehWtrkoGr+3PRUTzQW/WGHM5NkQqfThOU5mrVRlAO+b2l1gy2/CorW
nYb/+7tEHAEWPwd0s7a/mLFs+QDnvqxSuliKCoidw9E+ZR7HoXU6oWmfq4kGJjf2
b6Ken9mycR5gkME9zYcmZT5r0f+pmIM1FQn0MtedEXi3jJq/GnbtGjpxbRmc3zti
37f0MzFpnV35yt8tHO47qhveTosQoQ8Oa8CmZ/gxV3ssf0CB5XOJzopPh9+KXTEk
/+Lbr/XgoiiXlRn75gHPsCLwplA1VsWbGyBbuK2FmOGpJQfmRnSHa0s1WGCdQ8bW
x6DDmwbtLRNwWRzyAZIgjvqapGOoxs0rAixCyFfuCWUeYSlQWwvsLJgO2QI23/GC
x1Og3wkPFe47Gb3NoCEEkqtIVcC9xV8h4v7+575on+eJ9ZhBhxp1YEOT+kYd99Sd
ZBeFTbwBD0onARrQIxiHGxbPogirCl3y3+IOgReBjDr6k7cxVAJPpPgfdq4l1IGe
jQTlMMQu6TmACPmGSrwS54ptJlQJLwey4SfH01KF/8S5gnBL8o20Rxq0Aj8Ems89
H3T9EBOP8O0UonpuQCBFH8FHBqCGUQa8OW959LzrpJgTEGzSsnSxsYXO89SKVNU7
d4iKVlhfjQ5Kg5FVyOYJPA32ZQ5mMGRGhfVlMI1PJdw9v1z+PPu/r6uGstNnC6NC
tkX9JPquKsXFPvfcwT2Gb5RBQgflMvSmW2zyMkSbY4y4k2X56ZHth65u2le9yIvu
JbWzjJ8JaJgIHnLv/TQC+m7q1U9MaBgSWZsR6Hn1YcxMyAyODq52JPyS62aO3+ll
sjub4R25E2obeknlaxxIXpkPd7zVXpw5QVkQLdKYgF1qt1Zvpx/cc5w68W/S+v/w
1KmGTZBstO9Ngr05Q9mI3fAsSc5Nv3241AGrrWwE2VXlMOB/HbkWswGpkuiule/R
8btmcrhyEqi5Qcbu9K1H4eB5b+3QFK9ioloVC5tWO+CXlYE7ZTYW+qknfToYnJ4s
gNBNFoSJwugrCL2vI9jJ/4IAbkcyr9trQHDr9LTCURomFh5uCY618p8g2t+RtSAj
28SrQ+43GtqjKEd64oFfVdfYeBd0JsozES6JNK+/J+6TVYqdyIR+UkIcNaWQcdqo
WnpzzS1mkKl/RybGG4CRcDQj+ZoWalTxf85r2MzFzeiR7hdiCERlpdZlkmsTCSR8
B7Vr2Vt5zSV5NxmKsmEcoApQBREdF5j8q3R1MMu6zkdZNO4pHHJ0cwasPZNW1cc2
1qTW7WjiwAPa7cD1qOw4bLuhNFzdiGYMy6cVNvHeXyGyhmZvND/az4QXkhbXIGkv
5qvR2wGuSwxjFV/UXVf4DjJr3MTfTOwF+7QZ2pTFke32PbrrhUmvW1J6zTwUY9GT
Se5ngn+8M1a4ZtFCGj5TZl0Kk85qXy2cdsXph2LZdoHds41z9MnVrM2ZYwkhM0rw
3WMgVqLENOsNV6RdEy0wfdSm/6m8gt1rpPo7UQytnU2g3QM80Gfb9L4W4o/F1g/x
I5+nVbBqPkw20yGmxpSENszRqle+Ge0sg4JKBWKbDfMnXBUC1xNNqY5JIr/OxihP
EoNFl9mXMx/kC9gvZOw3oYvhRUaHjjglq0BH6wfeqWTLsaILp0pZbehxv8qxBxTv
DWAlwio3g+bIH/8Z2p6JKt7AmRM3NtTWNvTIkMx0BY6VfxOcpcdd0l45mrkYZtxz
vf/huVgQxWcnGM6XLDZkmqwApQfWdXgxm8ZqA+walaWaRRD2fFr2GxQN8g+46I7K
vB0dxNSyM46golShOYBew8MhVropNNCTgpZzDK2ohCTJpKT5kvhkeLQjyWOGVq+V
w+lN0a+q+GfhJqH5PRjOaOdlpsaxkITv5XwCBzlq08/uG2BHFIAdDYGeXXjNZ9vQ
H141PMEkUeKqdjSHK8BwQm/vmYt5R2sGiVq5zSiVjJuvyD+duO5gNE0RaaFJy4D5
tz3kZN61OECP8NSPSsZekiCesgTkvTaD5bCb3vlax5tE+nOpI20zzmQh7Qphsbnk
j7SZHRW7EWlTekDLhLCdxD3ky4AL7bpdbDbxmigyrv2yUR4+QEQQdUFTBxRhecuk
XJDAOThrsHkddif+x3Et1rseT/89g1TzvyS8IK1Rigv0a4UYh43ipReEThZ6CpHH
s5GwIPavBkyz0T43YFZcIMxK39mKauKwD27FnPzT/DZrQG/CaM3E018uUhlLNQtw
SkBdA+Dr7EnosuljMGeHH1r0QOMFlIWEQrph9fxCiFFBPpd/yZE6WrkAkPV9SJoB
Q6RLOASGJjReZyuucoADwiX48Ln3taRdZi55qPNM8qOdt4bOMBUYB77m4SiZ1DrR
4O1UsMVUPyL8cOEIGWHaQIkXV1MAZpbez7zJ7I+qmca/bxzF+3D7i6Rpjscn6A36
fUjD15j2Akvsal7ncAjI+oB1zN3H3JhjDRMYCNIE2APosDMt2qAph5RANgFtX9Z+
lGIASWLTQJWjYaI1WAKYbVu8Y8IrsYCAXdWi8/olWtw1vg4DVTAR+6rtgTh/qt+/
qNcYD94uw+l75W2fVQV1LKzPhmFZA3x1fxxjKge8vJdskJE3bf+mRT7hzVyt6JQt
SqjKcnsTeiQyh2y+znFkEKefuDRBJY2G6DC5w3AQ6Gs6momVwQrkzmVVwkkFf+RH
dBDIHMnIDSb2MVxXy0GHfj7Mm831SArdVT3Hkfkm0P7l8JqRM0t9V1WMCwRISuJP
06GIeJs7z0KACzW3x5s6zczkrFfYUgsARmxqPB7eRth/IvCaTDY4iW8E94fMkYZW
zWWqJDwOCSf4Gs9/ib/1yzc3hXBmwVYU+yuN/nDRaD/jrxGHlL5X3FIU4J1gm5GS
6aEixE9sVGF1hm9NbdKfMoTqBViFfZoIynCDp5ZRkDdhVumxfHmMPqvA/J+QbwXP
V0kNj1dL1WESq24W9CjRpjImiX3o7lv/FqVQCFB5AfNsrCbtP6aRkKcT5CYhosNn
CWysMVZtsOznGT1cOFsP+6Ctlbfkn8cE0ZWLYujReOTea/MqwR5Bv0him58WZJRN
Uow3hkj7gYvrKQWxtJJ5DT1l6X2gQgpZLFYj4fhJZakDMHqPQ7pW30Qq5w0CdN8A
5iypbayjDBWs+O3QTRHSh9VozKCOrfs+hBmzw85mF7j7pBfDx4nh3VY/ICi7at/b
887GoxtfvqCiLKRIGTQX6hCjYOCB3T8jF1LGcNbf0+BpaXHd1h1s01f/VmcjV7RK
7kr3+l73gsuvVQtzsGCd1wOpvj5i5uqBELucjbIrrQ4vzY4yDb0XB9lMIcAp4N+B
SpTRR1W+UxdJjXh1MS20+0qmAYa28zWFvSlxGPDhbwTqm0etrQp6yWbsR8HWWWcr
TQaWWCcgRu/HI4dRZT0PbIZehmUVu83wHYk1lsf5MQrMm0umSanBFsa/JdMQVgfQ
17+e2bM6ImoztPS/xj9iKomldd8AWvlt+1glEfxvM/TRaZI0Q47bY5AmW6spLWeC
eQ0d9i5I0DkhO8671jTpzETGzMX1Mqgo8iocR4Iqh3peBjKdNRwU0Dy8XubXgqB+
a21H/wbr0yOBNtjoHMHEUbBf4h5MwW03oVhyuKNaZqNYrOPf2mgbb4QbZwzgGS4c
wRiLaUreMVSjWAGgln34xFzQ9vWCqoouQC9OaVBWCZb1y36Kl6w9lJuZuZ0MJtvC
NZJz/2ymZwrBosuuxiY4CxShuPO+5TIPRG+EWVyYSEf1iPIm+n+uxjUrhv20n7Vf
ixN1uhN6+4FDk9skp08URWBykOoFblSYvoXkog+hWKWDlkF6oZV2cXCUP+LuxBoe
K3SCOenGTNAIbui4WQkJu4brNiyEsohkYt1adOyMD3qER4rNEC/Gi7k+VpOfjfhI
ig3rqW89AKWHvKB24dyKH1jpl8oP42WgjqhGzA30UyfYJrCIyDloe1jNTLKXxenc
MFR6ULCJWzjIjLN76lt+QnM2fh5Q3h00nXV+g/hJO6ol4eZU1RUH9/anPGrgTycF
E005+dyjTB0WAmjz6SBmhVQ41g1GswJj8kKFDlEm1FnYHrSNsPaabAC2nr2wm4+a
XKqsrvOQ7BwoPAkYKxwvI80zZdsYj+fSNuFHRYZPOCBFeddFuzEEtbPj0+aszvHL
fL7PmkhRG36KCRc64nboJxbZ0JmYWiT6VWO5CqSgrnB1T/NNffblajfAtrtp7ee5
Bb1XYEhOStnwQbcHt3pbKuN7OydmsOS/9ALVPn29THSIT9YLeTBCH3U3uKByXmPE
nf4Pyk0TZx9CtqChMUYRmbSuthtA16SK0ffklv0raXJOgXAfz7/OGqvkC3OIxblI
1bdk6lO1tNiBfCqARtFZn2SEBOWQ+aLeUUuurhTbs9kjqEP4jCKetdoIQhW68v8m
ovyekJRk5NIJtEzCGg71c5+OmaIkH4FlygdQWJPMKPuii60FNdU9lsDvGYN9UAe5
6YgWo805pdv1mu0Jq76pPtD20vhXMqTUn7tnEBFpu4A6Gp2WBVMza8rcF1tkqHZK
Z2iaQfNGmCAXtDu9dIAzqBMTDxys9FsLm2dyDnYfRLfYgENuzK4Ww2dbJFdnsXKA
WH2JAfQjkA4bDKdgSQX4R+5v+VsIC/EO/FVa5rjRt0sn0dSVm3lDG7C9tAEyB4Bb
Ri7cveYbAjYlrfzDOLGDS1giQqgiNBXXWxWTI6FMqQGUbrpsPs+A8UccnRSgt5LI
usQZwnotWi2jP7jBYBN6PEKtqB4UlXi0R/d8f7oEtOO2uFLmVgJWshyYLb5kcpVW
ywc1zrj4VBk9oMXujdraUBqeIkKGZqbZgb/u1z15X48LVx3eoj07GCxsLLdClX0A
YG0xAPW0YUQzgzE3oeTw1RqSR5pk0UO8CJTdvfNE7FpVzZfsGVtrEzP4l/HMLe3b
3wqlvpaK65moDPbKhlgUWUbc+hjq8fVviVu25obWR/iWi6KqaHl5mA0xh8xJC7af
3EiE7JLvVCDHJwl5E+duUMSXc3mDgbmHpKVAYdJOaZWscd5nvFls48ccfymUclUY
FbBPzKCZ25LbQv/ly0RQDdbY6yV0g/HBAQBP2MShpzZvJYdoiQmhHG/Volnm9dm+
gOumD8dp1FvS/Y6CvQ7cTVwjT2cKVNrQv97CUKoZO1E5INKxuJydANGrDmLUU0Uv
IF4d/mqmH8Z/cM2XPmfOfyf0ari4tj4jcJwhnAQWW9N0GvfuLQgqtabTkq7qOIwO
icSfpgYJZ8p06V7BbyYMjSMGwXk7x7tOLqo77RxxOILu+/WgwDy45/cmxAz0DogG
4DCoEW2apdMF7HV2XgM1NlA6ZTDiVN1sBtPN0MlgCIKVMylkWrtHTacU0+gh3vKe
+I/iDvTnQdm497edF38l7mq5BVQU+2Qz6d21pogD82c7i6EvM7miHE9tTeQvMGXN
Yb4UpdFjuanzNAbi+ZeCxmfHqqN3vfoJ5hJoDvforCDxsH4hLwvTXgZwHRc28Ta0
cwJjuCliWnBm67rZUjrCYhtBYt2nRR5urTkDarddsFPYeZQ7VhPI2mekUJDPs4U2
6i6qcw+Nxs1X+Hkn28wCQEz26+nHt3JRcXZx9iQueGpst5jbz8sX9gd3T1qBYFoG
X7NSal0UhRwT00yRFZjEie9+KnL42pS4FiDPtQbVbVINU61ghuL5QHNfqgGFuISb
n6fr2i05wz3oE6QgG9GHvajdIqy1tC4ue1cuq3fhCeF/02bh8owDy0HuQ38b7o7c
uiocMZpNQt8ZXIMBtO8hqlqcz15lAiiDdndkOUzc687HomkjwjsuoSipqJ+NRZId
wlUM6ce9pYf6ow3JZEFcMQnnUsJFPSeL4cIT3jHN28np8bkGEFytKUWUIeLO2ROF
+UIZ1FoTGk06uDMOYNLBZhVRLrj2WdHeixtAda8Lb6jNY+UAZwxQYTRztxjeVRVd
MOhn46xKb4fJURnX6DJr0CKcIqlA1Gr43j7k7HG9NNxrrvEh8ezchuioKJXoUIgT
JW22wefxChYAdLGoeNrVKj644F2nfnANTIMfIKdicL/n1EIso/JgOYJZprF6CaDe
Xm6EMFyDGmGJA6Qv755vLc2QzD6zBBWnzHxPTeCU7ILMcKgBQR2vbBYkR0JVRDBD
XmyzesxV1eJ5ZfJ4XfmaVWfsefUs3GEG0zecKb0ujNtOVHDtZfg1+qHZEaUV35sH
/jeG9j6by032b3KrqwiTHkAtX/i5HpemtrbmGrUFJ3lpwScifqz3ej5CitVYMffE
X8JkXDvAkkdrkKWwJQkMiP8x6xYzMbHuBiJUuHU0HVVr2PlFf7sVzN+bpzPQULUm
Hql2dnkl4kAbcIQIyXgZpyAgTtieeRuA6HHgFRNLoA5mQnB9VgNNZX6sbe7phHOj
qzwqtIZHGaLv9ICl5EbHoW+pMpMjQwI+ZoPISofwR8f+7y9EhSi7Ssbf/GEK1GSX
PAsl1ErzWVajYjJILbIDlWBp4rhJZflzcPXQhEejlf2VbVHi5ytqT44zhhRN/0g+
L4t6WU2tyaNI74r/rumG27rwVuRzH8N75OYcgseDvOS0lbRA9m2xsj+2a2QqjpQh
Zzi7Ome9tum2UVG8JZQ9eRjbFLdlgYtjJL4+GyZZGR1/muDdCeh2+mIArnF0E3oZ
ljAwAtCFX7dVbJ436FWzDm9/ShPMloYzGjpbvi2EPod0wvlTacWkXFuJowz1zsob
e4eOORvv51kTR7D0KLalZNAbKhuPaLRoeCqCVN1e+DMzqFQnGe3Og1w7yFHt/Xcd
6EFjHuqnZLIAp/AzI7Xu8MS9rVINcg3EKoP5/MUnUdUEfSUBP5HznkNNybRh37BU
VLz7a3JaITKeCFfU2L55KVWZIkeq4+R2HsaRq7GShj8I9KgBLqnd75iKtJx6PH8u
PD++3MRnzpmblDCPfutx4Q4nKFGJ17sl3XUf8Ht47jD0UBKQgqlT7eI5o5GDfGqr
K+t7iE2UHB8FSB+BaDtbWCUIDwhQ3WVQJ6QZmHrQKW0X5xO4bbqtx3abXcKhuonk
F0EKSJzr+caqJFiZMmi4zhHM27PvYyMlt+nllW+/F0bEU25BYEv9I7ezHORs8jtK
2aqI3L1mt6b/H9WCl96APCk7AVHZBDCoVYNcvi98bFb4NmnhpSK4Dy0kfe/0oHVy
fZ7X7SXM7uJmxzBPxuS5k5hcQZm2Q7dQYXhcmOW1fReyOPlatz5tBFC4FcNfxEzl
IqKyK7hIdFQQXErDdmhZ9YtF1cnYCOvOjpvrsVmq5WYeWbRSq8NMXSIoFrAKtR40
Z6VlKs/mi53pvPET9JX81E+aMBH1iPrPniXQWsZiZielKl79St2xbs10HhX2HTxB
nUHCIS1vK+UYOTLOUTKVplbxTEFyoUv0JvCxONCSba4oQiRSosbJxbJ5YKF3oMyB
iSje/xk/6W3tfohvD1qv2uVWfjE/vbldM24Oyf8JxZ9fbacktvftYuFMOJX6VBK/
8x7oCDjderYKiJu2k3mTKxtce99dpf8OZHGaBrnYTD89R8EzSVDzW1NCq/9JW9pj
+c7XOH/we1rWmuispHTw1E/IoAGtaADcOPl7cs0q41e3cdegDwcMOI/H5egXq/Ji
r3lVyiLQhb1949NdzBII2CBi9MYmYWKHTauurngUsSSQaipXMJhDLDbFUx3A1n9E
5ff8PdLfrjmQKnsT4VLujg+L8l+DbWw4NJXyFp7m+Difw4pcl9mnywCeLBdFVWzs
svhrlI6sCZh1wimJVgPkT686EGHCrFRSelJ1nmYNvfIHANsl62T+o+8y9kpmbqfP
og9WcxMWMe4IONN3wmf6syI+2seMAtgcnhm7kCR6HQHFvSEQE/jPgA2+6VXZrEPM
pyCV6zWtbgo5c4rI1U4MMTUYbu1PwkXz/roI004AMKAsNTFeXp8P+lDVOaGp8rDQ
naf/+oXU+9jPZ5tdbxXYzBC1hOuiEAE+7ideKbhlT8ZG1PCLsrP2oFKS6sWHiyDT
v4vE+7mVWKjdQNK7w+6K0u1E3Cd+49MQK9iUq0IWS4eaZvVhirJPfZXO0dL9lqNX
nfvKWF3R9oHv22p4vtqrokhySDCE27ua50HcWeicPWQEjv+YTyYvSud0CGgeuuVF
11nj1agAjiF+wR5e2lOqEQnQkfGJsOoUZnzE6GWHfyiFmu59DyCqXjV163RPZIJV
mog3Jnt4WpAuwoUiK3sTwvSrHdVsqtx333znPaAi4ej7k84ccRQDVC5kw/HzRUBZ
H/vREXYkxgWL7ghwYSNNXV87rx1+PrDa6w+eTzNvQK6wo0JM85BzNrjjvr+pEsRZ
khfrLhuvSZd0UKmMueK5LL5I/pQSKXuSPvRs8oKRFsqBKua7NLHZSpQ8RUXvb+5O
uFVtoGd8/S03gi4lqPKOtTbB1mXD60emvqwnxxEH1zLS6xgeB9yKXIgHFyONNT2G
HTnqAiDYzgUDZd+RFpTqR27pcu/SI7lEtBU+pFVsliuh6jaRooG+LHkTyPWFscW9
S5DIs8DMYhFtAvgr4ep+Iad4uYGQBNUi7v5BcoykCTL7ewE2PeY3JM1mz5aNkZOk
SuMPK0TkFpBL4tW6nHSz00SC9gi+0jqrvh4l4GmJ2hydJI5u/RVijPK4zmfhsEqt
OLraoNEKZzSpt79NLAH5NWzZ3pqy8tYBUoLfpRx8X1FXAuLmaaFl9KDsgn8bseFs
07wxzaYUCakAxk9K4brEkTvTwV8nKDOugNZdeauLBxHg65eRjqaJNroqdXM9N2L/
8e/cFZdDjyPruT2e5j4f/RzzXAaUaVdlGjp/M7VvaYVcGWJfyh0PNtfB7l30WzaE
9NV4686nmVlXqWE6RLFKimlUbNA9N9lH40GnWx9ucxSbBrD4J48BIAeHY6WCigzz
LaV4w1k05hoiCPTNLPnJiy5yFlc9IsnTdiTxulqe8LNM70sImzZuMcBHW9Q7Cd5u
iG4R/ukBF7T6+tui+vrSV1zOTiQwI890410kPkXnVAm2oUOm9dqMKDITo9IvPaGc
uRfk/RDZv2HOuLKt3rQ9B9+wWFVTPW1jEw38KIEadgtNnmitDpbIXcT/f7qSmnAb
8Z1+9uc38rhucwHrLl2ujVEcoUc+3ODYLNg8fVTOI7fXSaRcX2LMqqjVTSu44HZf
tXkLgmfgIBhYy0ek+jPQIltSyOQznLWgvxlIjthCvQ/y/9zWW1GvU1sgOEjL8D9r
0AQ0vNPGAkiKxspEh6Y77uExuwe0FckK+ePnqw8Djaxg6yJbKOQU8+ayotm1W+M5
XFJJZzxD/9sbJ7zM1gEN0TeWjj089eolSzwTPjPD3UMGLgYgZC6O1ACnAB1xTCyl
4vMqkyMWDWDeLzNnhypBqjN8g+T5D0iCDPi9FjbFax0ZiRzy1s1BfVLFNMUI8ETU
4p8nd1mlBJ6VVzDij9LScVE2M5vGRRM66yqpLpJqLlexeg6yApO34BTnF0x+fzXr
GOSq/Rmwgavzxl3r82TtBskPWxGpa8nqsLyMXMkonmqNrdtaXdlkrxWgYDWwxzBQ
Ic1HPXayqIxqZ7r0uNDxFuDZPpr+eKmpxInOK25gDhhZGcyHuG1QsY93aIWKZzFa
hPUM188iE5zJz34nvjcoJlFOEGLJ2QeGjhWvedSh9od5P+ibNERN5nHyjT1O+36F
IXx/9IKeafBrIubhqd5Wl4l8+6obnvUdCi1MSx5vUAzp90W/P80BhGMSf28gC5yT
TeWZlTSqcEk485bQHLy7lRYEOGkoaNqK/TLG6g5z4tInJaJRUkHurW2l9zaRktt9
/cbLtHzgBTiKAmXi13GEMZlf3VHhWHiHge/tuv008jsClldBLIgJ60/TFt/h/mxi
7xhwK4DVpopogAxI8/tisV7lLptj5XfKdTuif3m2skMFVgf2CVJDmqFtRyDuh8oI
M6pGwLATvIoTTBTwJ9FiIRFsmRj7v7muq1YAlMSlX8Idze5W1vmz2tn3kexFy0Jy
tDHzmQyXVBaLPLGXTMeWe6/7ISR9QVRWZx5VQ9Lkzk2R3/uK0RB9WAXrLIELSXyG
T9jkHjksgwLAeEs8s5sAOd4x5BKJm/sAINn6H/tB9aoCKUBZ71E1n4wCPkzvXLG2
iV9CUp/KY/k4RRwVn1NTXbrFWaWw0RhcZfwXhS+5vnn8RcLjnCh3Qy1MjVxTlIrW
QZ+9+sT6xh47UrAsnQG5vgdbsIBoR0hEkau+Dikq6yRiI6TnsbKb0/7QBwxcJWCw
OFZFuBOlXzC+4/SMZoH3LzlsisJB15+kw9/kn6ghWdBsoQ+rfrqeqHoP6rrFEwGz
KnmPrDuDT7aQaK+NF7tH5bstikaGrlUvON8swPQJcEling0BQxtMvOXeW1BHusyb
dMdrD55/aGn6I5NWeNcfoVOHyYcHBzXDFoZnUeH7xFDqRUmvlhyCtRFWTDgq2Kt7
p4bja+rhzwkaA1XNTwvNFklPs7BP4J5cvv33EbWgzDi9s7/MCxEo3riJeXoc5w/B
FiAXe1AI6Nq/ZWPJgDWCKfCTR/1QdC1YGGN4X92uXmw4AjfpCWukAdinchu20f2R
QRDHdia4yVy2/v/YMyX3jFYm2KsJbB7nskJWCpYsheJkZ3sePDDathTWH1E+CjBe
YbDSrC8rgx5zZYpWb3H3Z5/4W4tMxESWhb9l7xkTE34N7lL+uOuVh+80odZtxhYO
Zv7nA+rV17vCJFjs2IdwOzxpGBiQc5k1S95ApRsFJCpw/tq0kgO4y4Ba56v5k853
0cz7PGxVVuK48oGnx2Q2sr9LyiDUzrPwu8/PCx8Wa9/eILDdtEv15lZv+9VZB8Fs
vaUDP3dZL3QbwL+hGnkeWyr9CpTlvRH3XQLIqmAI4YFB2FfwnFcnrdPt4o4cyU5E
SK1Ob+xRp/wQKGMBtYhud9CqYNfvFglri1/BqSfKwNT2nrEcSAY2Yg3NQOGU8Jgr
KgkTKq3xho9Sx0d/UvAoYJeHtY1PtvEu+hjRlUMktHHvu3H4thE5E2moG+/fG9GE
j1jtAFQ9IOB0wH42PQCNymuVcZKm3AQmRyum/0ubSbUEZUZS87Hp5lB9c7u4cnyP
6sB0t1dqB1iPtczRrBgBs5qPqpEmyqRwbeBm1ReXqigdtImgLaYbgT3l+l1r6ql3
3W7y77vGDuuSEci6BLQCxS6AH16jTh63NIEWm3q90Lo6X9e3W4OH0hZdB6M/57uH
8vmBBR7jhyl6folqZUwPqjvPJiKkHyCOZSkb6740lVEmWnNzunBFtpDAZgP6TDVP
20ITjc20VjYRVBUkFi0E59orUBdi9tMwn9WmrkCc7PjnNipd39uTGtQ+LLuI7iyR
Aj3mgKheqdB5H0vKuVmEc9gxNfhqex5ZMj9W9b5nvLNwlipyaMCVOOh3ptSEFRpV
0mxj7YPxnCxrVcAkIKXR0L2aQAigQO6+lCxpJ4Xj9IUNzSRJmdtY2XwoTogu8JTj
TX64xTn/naLINP/opQqV1vCj7CajarI5Fv1GKzA/nOK81ConZi1D9xRi4NsIjN3/
4E5InsobdNKucUDjPDXTS05Ds7O/haX/2P6OmVp49/Pa9V9IBs+934azWysMhNKh
O0z+NT2SYq7g9wEHVbrPKSWMYFoPNehPBb7+wl/4bpB2DTmWfzJiqE2zqMK+CcLz
+v0yQrvBucHVWkHK6ATTulDriKQ3Lkk65KQmA8nkh+ntJ+1Oug1FdIljEAn+SQuP
K02k8Ec08XZDPqYzCkNG51kS+Gbg4oE+FEXwP778k5VzN1VvXBmetToqub6G5z3o
OrCU1xZR/jEyRVrkPxgXnOVaynpLmxb3XYbzepeK37WfC8bQkeQoVPjo29cwSujx
9i//SfZS8HYkkGlXyWUKO1GRyk5alUNUT+qN4aPvQE+Qmu8lVwvKhhG9FSMjwpqI
HmFnpqwBhl4SlE4YwJTjX0O0oFcbKV5tsPmjbkB6yMnAtQ7q5AeZqxjlLjrAby6r
9KN+3hGyzttW0ipTMT9yo8WSae6okrK5/NsuknHfr9COjevQWHiMfbsNkf0Ib29f
LZYYBmdwte17ngiCmuZyw2repolAGREIECy2mjrIrCP3mVahCSEKO8WDanCYx4nh
LdiMzFHF1QduR7EMHDxwQhTm2EWrnxv83CrB8OR3r8Xs8+3zMhxczlBroFEvVY0j
ygU4uoh0G2OTmgS8xFDf2Xc4zt0VGt8LJOoIRepKIwLghUKYoNZDlEPUaVeLmcIm
QVJ3phP3D6Cu1pUyHmhDH1fCMz9Fx4Y8na7vfOXQc43hfk+iRUxOWkuDbpjiMEpG
bBTUUixk4Xp7IExxKiRUlUk5CaKnGzc43CJxQxDvFn9A8oJmKVm/g9/FPZnm+Rtn
mIK2RyxMgFtTp4XpXIiJsTrbpEy8fONPwHxm2/dXRuVhnOgqEHpbYeqBlnghSDGI
GZNNfPzi+Fw01GpDoTIlxlFWvOpRBY1PKh1usjvpw3OYXuTmhJnskvdHgKqali28
G6NNUT3WnmDt5X2M8WiMKGZFGDmU7L7km8RcKkE67UWpCq9Yq/xabY4O/uw92fw/
G4SyWueodbMKUiNm+s67A6W+G30jCxyhQwOecs0av3NYk+tG3f5jpbnqrKHPSds7
1UYm/8l/TmV7hqnv7Z9lqMv2Y2NYZfUEiQfNFnqryqVdsR8Yl+IERQ14YZZeTB5Y
DDzqb4Wn88theByI7iARRdKSP1hRXd52AkcpMPLY3XqMqpUK63XV9tLrxpiRDV7W
NkTRuod9ML14MuvWs7ckd3MGanI3/XnMPo90+ChD7unJ7AU7HQcZI3ai8VCb8erb
InaI6sKTkLt4yQR4wS6u3hg+68L5p8ENOWfLcRcU/mSTq0BFFgMPOnomoPkatcH5
qw7DRK3hHtacdYx5hH8d7+oyzVKb14151cwLvoMvZtIUtUE19224pnqwFMML5xKw
FhQqe38H4PU/0lTkwz7+4DR4y40zE6cWv46O2WnxY8HoBtvTiZ5+cDggQM1UAuv/
V3JC7OFGmyX37aW61I0ExZXczTXEowoSBlgmb5HxbPpDuPtwUljdDSUT1oacA7ZK
XkPnxiR2XPvrsiB5SkKATyG/04g5BDh3FHg/xv0NCpj1MHXU8FIjCWaPbCclEeYi
nBgABA6xmb9f0Najl5L2dGSQWrnXvTj9VJqtwhbOd51O5FxIABB0YGQw714C41XQ
ayxm8jxJziA+PJRhhaV05xs9KUhQqkb/b9Ksy8LRCgJVmeq+Ot/NsY/9wZjuNjVh
VNlRjEOTw9SObLNEgyWZtHoulxymBxcEZGSzQw0lW9eh01PhIzcki2D06l20kuhH
GOCO519/haylsaw3qcPRI4CHNlQBSEE+0Kzd9k2eV138z99NE78/IV+NSQTyMnH0
JwNS4M05xoM5mSoqqM/ifCOYVrYqBXb1ryjn0gHYuZLW6uoqnP8cZ7suNzy6G7Z5
waSKPN26RUZS2C6DZ74NyPYc5EceuEPnYK6CFH3IaUrv+X1/frN7KytYI9NoACOX
3iEDj2HAGJc/DwZna2ThyphGbB127/LpS4lCqZhoFrbgpzGBlfpPrzjGW7MgZEjZ
etr2kfo2fS+GeK2LmJNb7aP4cXcbACktlX9bRgXNryC9Uz4zy7lE/Y8/+BHLaJJ1
my8vfDA7vakjBKp23Lrn8uoo91uWR+2STR2BZ4GWYpEB/GvOYJb8WuBkB7TLq5Y3
fQvZTSkxiG8HM2ErOP4DnaX+LQkfuQDrmAhGhQEDfqVeYFbpGNzkzqSvNBg/DpGk
0BELjPUE36v4g9Ffq4FD8VkrQKLvh4A3MtwOiXKNsZ4QLcJsFEp3d/5Rv8KGYhoC
ivaCXUvcxsH9ZHbHF8ozzeRC8UuafmaNf6aJHLnUnzAzaYAmRZMOkn6yTBKi9ArM
2qS0LHYmn/Bq3ObmGSvqTDu6QKUndT7C7mX4gevDscCL0QDY6gAPzRuORPn8X4Iu
vovCYLdx+zClGxbueoM0ZC3Mc5gUbXPD1K9DAQ09ueWT4mFHNB8hpAHg2jscHFOU
t1+AMYTFJJBAvDgtL6Pi2wSmpGewyMkdmcuvktzjNoDSr2F7hbY44E4w4HLu+YVg
GxwqNufaxbRbb7huouEre41NFvuEP6YgBJBdwgi80g1/+f5BVuDTwCXnwlUCy7Wg
LL5C8LmegKFbvFCpqojPpfRkQjDik40BEtLzzMcJ4UZz2cwDmCFTqJz3WHpF0i7C
Yf82lQGrPXWvs1U/tW2rp4OtUNTwbn6QSj3tttpXNvrIu3ZdByXoj6s7qozHHMpa
jp7hYVUlI1NIGR+FsxtPt1Q+9ST85vUhXq/rBseEuSrtjxDQAf/ORRkburKKYe6a
HxN40lQdQ69ObjLVy+XIey5my03EXS654K2XcMVSG9+65K1cXb4/abEjV/3Fercz
yw2rVVqjVUQEccmTFTon71Ka6ofboz0Y6AkVlivYntKBPbywSa3nVfthcLHI6rBp
tEPoc+RcOihQZvDc8sxb4/TjAWOJO8Bwm4+itV+b5g3X06WUD4m656DH0Kcu7X7x
SymLpdFvKOIYErsaak+LDS+trPI54kRUBZYObehmQE3pKOgevBi8CoenzEK+Rvrl
5YgFi/iHD8SRNmapnM8MyFXXUS9xCsY2J+cfqhjztEAYbZBZksMRZWA8AgnqeXUa
vPDjgWHqPOVrQ4ydVrG8DJg771iP5cie6lUKkm0A8AijQgHFr9PbVAxIFM5f6cqr
KmMAEoHviQ1SLg0I9IHQmQruPJJv+DZEm5VAYBcTrCsS6DdfFtSQvxNFgjDrSGos
ROfaRy4jOOjbhBp5gt9syQjtdfGjeaGV6PdKNkAfXaJBjRksdXZViYh1PhMkeYNp
Mm11jDyo16aH9U41zvicDlcP34pbBk6Q+S1tVsFUI0B4WXDlewzk93evtEF7TSaR
kt5133xiw2D99y/E1vqtJXSJN9wtDspARLR4uQgGQ+lANGPLyiJlTAYNdozYoPpb
yr6Qri4N40rTYqinrLVVpqAU1Mrl7T4uKoAiXGQQeg8ee5VxvaiVr8W/VA20HJiM
hXD3LeLSvk9O+piSUGaEp2QuuD8nPiPfIV1Jcz0EbKTzOcQcWY7Zd4PmMZJ8p9SE
skVQ+bdoQcQGLIff1FAU2OO8+xLwh1Z5ns50E2Gi9XZItd+jqux7ZxtNRcArhdEq
gJDMlnL/d27WT+e3fRxsmE5lubjZvK+0LPL+QNumv9KMy4IuDK6ujyKrsZ/ON7af
qn8TD2EiFNrdJOeNvnYxH+g893zrD+MGwsyXRlDfxFHGQuXf9ImLFtU5+kRY/nA4
6xvkhRy7nJ5eTP61SRe2ZONu2h+xjo99PKzZ6y/Rq9zGPNXRCc8Xwc5JV5uqBWIY
/XHlbGV01DS6f0cVrue8MbYfjvslNdOcueisLxKETJ+Yw1DngSWDDLRWJlDV23r8
4vYnJaBa+zKoq5UeSu5clH5M4tLeOXJCvCLx/MBUX9Y0qgD0PqHkHwIMSGdU3OUS
4xTbZgu3k2zz20bjPRV9UPpShR2MCER7S/AhDwy1XhalPGXxPCHjCezoXOatGyAw
UX/kqFW2L/+Yk1HadPAEsvCvQHgVuVJL423mXJ6RBLrS3GoVmEpndrJApXN+QKgO
n7V5FKUkuSiyrmq3lI6lEJTrFXcdG60r9DP9djjoqMfSKL6rG4UIkmLfpuSGraxG
pZt8Y9I8x0nJ1vWg5fovWjq/XPII1+RLNYM01o16LCpMDcPjQx/jZQrZwOTzX8H9
SyvoFMaONmtB1JIiQ2VcXr8vjBkkz59h+Vt5e3tzDLugnHAbk6Jo3zKxcZ019512
FXLnPw551dlxpJuWEZQAzWrqbN7XoALnhbVeiU7P7VAtoFqS7t0tiz0fGKm+4yZi
SWev9vLLike7zTF/1sjnNhitf0s8SIA4Dtu26BGerscGyO/G+S7OFKSUYNefIaJ9
C4xad8GjS14uu8KJLEDN/QOagV3b4QZ6wqaNP5/WwfKR2Y6K7zGtxvR0u/RC42MP
5K2DK6V5UYkor9d12rqWzupaE+oIuKdzNLlT1q9RVUEUUd1Pumvzw83oJSCXmzkO
9bNjM6H4uLCcs817+JJTG/HoRPkNc62mw+dbcNXloUr3sCPKmhZ5D5CygmH9zTNw
dbZC4Y/NmZYOtT8I7RdnKoipGLItMu1n4e+2Ph4dfqzsnY13WrO9XW6BbE4C7Vv4
uxoZwJt5Mtf8MEe08XQaF4udG52oD5fRJjnWxsP/cUGKEKIZlhyIa2PfsY/EbAff
6Q9LQ1WH61X69DlOp3vqurU2w7r7ULnT2cQm5+GUVDCe0u8/xk3w86pY6Uh7Qmrx
X9IsJAY2LbjuMSBBIf8HTSoVdsQ4AWQw4cR2meEJAx1cI7+BT2WdYHfVCCK1fIer
DF5IVZZokDy4ALVgEiUJiNnEYm3hKEzQ0KxGpcJm8NyMIiy1/vaGmypsB32bJgMD
wTqJ25pB/CEmLfjPtkeQEZCu5W4ZnCTbFol0wyJl5CWTUMoi9z/NykimgYUaeaZP
zrKsufWb9SXlWpxvxhLq/C2AQ6vDgNSnTsg7smw3X2D8uXa6VPwZeHy7c21YhaH1
rh/vyrkTyqJ/xhKWXZ6mHXjBMTcS2gmOkypYWitkEWGXzE7H3O/WDxAcsRX+uLXG
fFcA8qc/z7P9gBX3H01HqUnWRNVyFSvqUpPwolEoNHX5EdIyJ0P5oBi/NgLGkkGQ
S+QK9reA3vDTaL8Vgk2kcy1Co5HD9j59gQUCBtsjnuM7A8g9i0u3neuOSx9xSw+r
5ubWAtsuiQvz4R0x0NpbnX7tYvSkQwkk8oOhI3zgPn24BQ80Fsm5Argm6woZXYBm
daJ96YKHm6fegNzJYSxnEqK+oLGlN2u34Ptd3JcyajJHB7MlMPMDdkJdlxEsI/79
G5WI/7AF47WYKKIsd8sMifNFYAJ/uf3r9bN8b68ZL+6RirOahFzeWIHn/RKXeuio
MUMwNtuP1Y8Gps01RMFUBh2s6TqAwEDEiz7AR1taKWQJ5rPSUXQubXeN/k05A+TG
DvE8XdXRSSBNoj5G7a8JouN8ydRxz0hXu+7FQY8Njt/shi+b4+34kctq4F0bprHH
2F1RIDky0Fmi/JfebRmR2QLESvoNCViRo7DRnxBiA3EdrD2OlOshw3fqfT5poAPo
q67ZYiCmpAdenFN7UfsLQrM0fXSSXWBjWnwTEm+S+uLIbedm7A/xV48xxvNPv0E4
8I4clxz1KSeyuoq/YwLyvoQIQnsaOBYgJlBXh3fOLEL1eetd03bZKRrg2nS0LD9+
P4QXaLH99HmhEbIyPVEI6M3KaLVTCf6Kt6pfYSR+iNFjUy9BYe2pMp9BF0J7CILX
MInmEiRMnQXou59AYcpJAXprFpqmBTDwt7DGUMZ7XeN7WHkBUASYHKODalQ3ievb
/DLexbkUyOdoeyg11YHOkBM3IudT/lCk8KN947AxF15NJtQdoQF61lnNCZFkr218
ishrHCArurU714hQ78vm7KXYE/Fhgd4xX7fB/JaYr7AJqFPo5ZAdYJajMVGytSsI
cpsp7u4OmUTyPMaqmIQBi1KMw2vOuVjFDXEP61ZL0iHZjnngD5ozh7hEJLongUUC
1dt/lHKFXLIbip1dtY6+xEqs3QXJQC4sgCTsLteqW7NK8SKIdQBiJBpMYxWWabQM
SpnNQtXgtiNm2meirEfzRZI1bprwP/mpPBZuM9yQU/dKLbLXETDGatKJDx6nIgu0
2BBrwJmJzYs0mJx2M2qNLg9MT3PzRsAGngTgPMeuIZcRQ6y+Y1hUDPd0RnM885WP
xfRWeczjTM54+WpqXXZfUBY48hgRYWvmiYwPdXpD/VrtO0c2WMk9k5vjuyyp1lYv
lJZpa3sE4O/Mhj6R7zjkhfW++MBq6CnNGquNoYdF7crPfWPp+oWi5luzfJySofge
1tg8MLFnw26NjIjSStcK0G/JE8DvfJvPSmN5o0UndWCSL20EuuFpAGT5+PaEkxNz
KCG58u65Uq5+zJ8du3scfjaSXj4tijVVJJ9nI++lNmj2myWVOK8rX2q9gxNk0jHg
HGJck1tP8zUxKSRT7vzD6X1oRqSszIIAbV89WRY782af5WLa4SuF/pk1Azcih14u
0YUrhCOdFTKzLpg4qTjVURbyNZMRQsp/3a7v3Xh5OIefwUVqFpCw/3W5nwoNttek
llfA2ZciGKtoncDX7wPZ5/dHUxnQV653UYFRehCLFndjnTALki96RP/22ZU0e9n8
PYiSFsI+h6jCT9h0aGYDIomQ9rcxoVKh+0NRSU2Vh03SpTYgZxe7RVA+kvYk9rm9
TRGqF4KiUUr22gBNNwV5z0ypzMV+aVr2/FipklMtmboxPapvW0s8xIPbvv3UKghl
wD7iGH3zf29Y4InEMDx6/k02cQ6FbPGPRTk79PukoNhtAw0vMTx54CTfZOJzcNra
Ho58o/AekrCGDxY0Oh8Wt5Rf+AaUZt/W9ZJVtcP8cW8qMM+PFaVsv8slt5G09Vfl
83Jlcoc1C6p1h/HhxeHFYfxoSBN/1y1q1jCYN5Rprl4xt+u/A6odWmsifMEJv7Wr
jvyN93OQAkWHo94GmPJ3HnVNkFSr/XzDnU2SAYW/n+kDUCM0IWo7qhMJtx8gA7xs
P9myfungNdB1NzflhodM75FMd73sXh1BJqv4yZotM44QT6l8nnFm7+5rW8BNFqDD
oNTyoAfyyMlU7PX0Z30iNrAoLpZIqdhvtpHWDX5aQO636D69YcXO9luAWNA4K/qH
lv4hnpelfX8Ng62GM5MEPn3r/0cGneZfpDM8e5XtQDP9Z5Bb8t68dwQnbDUrIVYo
WoNpg15Dn7Y+QYPsUqeX+dS89NPDp7bHHVlUeYBYzJ65aodQS27maaaadHJq9R50
XICvmXjoT+Fy6wniirJJsoFXxdMJHMScqT1seiYjx4uEDj4ENr/b1j/fxm0kc7R5
Q6U2i6hWboYWKAVHVQwB9QiRR5RGp2AyQiBSH5xSMbvX4QyN9xPcUcLJ8BWIPqAC
BJ/+0r2MjGd3RNJ4qx+U3MjGSHf/0c4qolpaEV1GR6yThSwOMVp+OSXNmRN9W/cL
US4/SG+85nV0iptJDHPdCpnLqvYp+aiJd/UoAuWvUhkq8h4YOm3TN8yoWa/Ny2ym
YshRgCf8Zv4+IqJh2BPrV+zTZkzk7MrgZmA+N5nKSAB+wOwk1mSI8LCd+iSCnbiC
P0YncwVTSAynDHx0B4Wa1KWVNVfun9RwlnxmFF7p/ObTJZxOVtZ5BE8uRfz2ZdvL
Z+UZLMmfXxDLTxE/zpEg/rz6GEC1QEQlmxUt/HrFIR/hG1NT4xKqwCUPimo7g1EM
7YzJcZXv2sUtgNLjKzdxk47eEoRdzMBzDG2DeJaTDbCOsfLBC8rXuOy5nwAzcu+a
CVnS0Fh/fOPs5Kl96mjiiudYTlycZ9gCHDbb9/mG2i7ENlb/QV9fyv7QnxTCZ7eE
1Z054v9SGuHsabaOpmhMcgToRaHiosaKFv6kQVrZSKicnotveNx8x5mpnoGxm9ij
xOEP6IsH1Us9Pot8FQvWJygoZLUd3EzsxIJxhzp+HbKa6IEvvpnuCLXYTZVmITol
JO6A03Ua8GDtumVNAl9W25LpS3XnDfR+DlT3la739hnzre+DHXC84I+d8UdiiOJs
cfsCFB2Hw84soJFlPv8zXvcFn+O47J2LsI4SBaDTeT9Y5nO04Ge2XkgTaE0wExAs
0tf5NpA6h/OoV0fndS1oK2whenz3I1LilLMJAGERmW9zCo7GY48N6Svl2EwNHjc4
hmD1YolGms708o0U8vO2J5WEPRa6RP8haqMCjbQxrcR4s3gGbiyg1GpyTQu7wzH/
yerp7N38hJFvyIAyh4/O/ZmtDEd/agUgug2nZFvygu1Fi8WN0s2mnZx+U3EGmvau
XY0sMEbQ+9Zk9lnhdPSjr1XLX13ZulbmzHzD7Y99jOEsPO39JlpM+qccCJHX4O8T
gM/txzujwLhMVJqdyTBuS2bDmzgNyPX58IRBukTOmxZM86vltkz7A51xTabFUZfG
GMbw/hbCmqP8GmN72U0ZdIz27zgO3wDWW5qlvorWOVgaJvAuF7VAh2EYKT4aybAC
gIDhwfSAx4ZwGSlAuFNixJ1GVKn0rHXVQvCrl5Z7ofnDoz1pInkkmY3nWcuZA3i1
WPmRtrL8cvWb+/TQX1xf+Yy78BU3bytg4sIJ92K/u5OMXjCdElXY5ZfIsx6T05Es
nJcsbF3yYdf307mzcd2ipgkRK1wY5NSBlOmDVF8qNRNUoJ4ned/OGMctSJ+ZnRWS
CAMR4a9x7RdF4ZWqS9BhVRx8ZQdFOmFRaG7qVYge6LCu/ptdMIgomPqgc1apJesk
mwtECbOs7hubF5bOWRXDr7mQE0iwSHSAAgmU1DuliN/e0NmjqhxeKPHJXW5Vj2P9
6jIoj5z6dDMierHPjpGZBBVu39Q2qeyorVUdc0P0PfYm2kA5WJiEaSFobFoEhHVD
/BCj324ut+UUQW4aUGR4zg1iMd54qiURbZIpGUQUV7baV/ixck5S+FU7tkcNCDKv
jswf2on7pafkUYzDBQdZU9RYLG1nCKXqt3WqHTzKEtL6ysjq1rTVU8BdloTVop/P
00upJm2KISd3kE6NUVKCPaLF1QG2kSf/0Y3TPjX1fV6ATxUkvMv+Ps5GjVZnmYNd
Q0AONMWy5Z6ykJS8NgrCPm6q1657WZdvKj4TWQhpa6kMBrM0TxjxwxEHsDPqG8en
DDgconyZt7yINviZbqRBXuFjdbuF9okolsQTHn2EqCgsYZOYMKCPMUusyfvsQwZT
fV6rIoyi0rPijX12Qe1/Y0IcqHVwkbZN+K9jIVE1dJuN0VzVKmfU+C2xPPUlLTyR
m6LLIpYGE2HRoeyxJidTZfzuQAeLzX0lBPaxe7LNAQ5/lIHB2BfJWUKsNJGBr41C
q4M57nr0MukojSccZcoa2FmdBj4akAilX7ks5w8crIVY9/0QKDj0bmPBxi0OAQys
cdIet9h3bPgQ/CV1NUlH7BnLCnYPNH54iAWXi9gxmz1Apmh09fHi5Pb0UOQ13NVU
Q1XhTxEpKVrXlCjpDyjDFO74O7FLcUgHkli1jynhNZ8rx0Lc35POUFWDgN/rHebd
5ZHBDqR5SGjmvGCmy6vw1uhd8yYOditRR0RT0ClG9bxVAN3ykFgvYdFpfks2L5Mq
/jGWxJ82Jr0rHDuzDzdAarPUhOZNfWwjaqa/0l06BMP396XvEdujWQuwpd3X5oBR
m4O71QW/xfWVJF2H901FJrAC0qmDpaZ3+UU7TbDYb7RfQIowhtv5qBv9gFbH/U9q
I1qYHKO05st6ce2+1JNmur7OhDRuAaq8bcYCi6IlQ1Wtyrrh6SeVxL6CQ6jCrFCB
hc9dSdO+ZFoNoG2LURqQU2IUQHn3+esxFjCpBUpgL4W9hL90oojQBIiy2ke0j5GU
zpU5oT+al7jaX33kTpum8+af4Iof4dH0hIUWpr/oF0XpXrAGGEgR4JhY4R7j+anz
ulOzmZlxPXGKULaKtw8N3qYJV54CkOaLaxhW1LQFJA9Uedjdk7ewWp+1GAhyU2w+
5lrwCjnBmY6MD3O2ru5wTv86q//z40vhdaxWOq6h8U++491yNPPQFq2jLnYXhY30
9jdNaYU728BYetawc/3x2ANMC/5p47KtG8RgMq8sW4IkVctia2zddhSoADAPndGG
EjUMM4mhd+FfGHFl4E02viGzzjjjt60191osRNy73ti0JrIdx+HN6wei/vMc7OR5
mwKAsJFTvZV+jUrkQ1cfQ4fNgw1BuPZzdbiRvLotBp7t4q+OChOSRB0eXSVNLV/C
8UTIWP3l6/GZK6anhC1CQrisdmvPHlA+7Hej1AdR+aEzdpSqd8+rEOv4ZIvAiI2y
qv7uJKBne4+1BlgEG19AS6ihySFt/c0KFOhJejnmlS5tJWgQvZmP9oTHcr8io640
tO2BNn/bqBPP6Fhy1nClsLfQURzdNvUtXsCIwWsMkKJg12kP92ND+CNykzePGTfN
UMI1f6B+2IMrV6yzTNrjtarffxbKK9DPuvayva6tPg3Pkz1gL30DNW0IPZu/9+fu
Tuw8DFu+/RamhORXZ5p3wxXLIs4r9q/i57ZXQa1FQ3bwMNg/7Gkq7mqLHlZNBcxO
s1KeTk71eoj0oS//fMmsw644wBIfpbA1PUaZQuX1gGDOR5lMAV9hSeQVY70crsYH
IIpPX+RSzFr5CqjCAnLXqXeDcRixDkEyaUZrhr2T+yyFvCr+ieIjoxwKRfawOEEv
pY3+3dgdNGJDRa8HSkXodvjMeWICba5WqE8sMKmdfMaR6QmPbWxQPNV8uf7hYbeQ
/wiqLgITy6oU7E1K83OBuV8uMTukHBxWfToYpXcCY7HQiqW2UNnnVLqBLHdVpQwK
8Di2F1lbPw/CfwyYUDxR7dLnyra09YlHzFxHU/SE6MyTlDsRDRFFJ2jkgMug2KdD
SJGRhfRxStNMssOce7A1mhFK+8tMeEoB57XJas6cMY6+MuRq4WHzCAMkDWbOCSNY
BYpf7MP/BZ6BQjgKkkl5ni4nRvtFxIKr0q1qIy9oR8ThzYwi3Rw0o93/hUktx1/L
WE1sipNvm0ev6K++AV+MGXrYMRDmlkDWwFjmK0SYldHzn4vjVkDkiNE/6w2Z1Gzu
LGYq7pVWGt+qVYBRCSMts9Bw5Cc/lPZ6MtaUIdkCmkMRfEJ1IrLU9sPlLecoGm6r
BDKlZDqpycXB2KOYESqqWl9+hQFDvRZ44/f09GhfcbWC2AMj4x93RWzW7lE/fXCF
SZF799NxyqYgxbKZMk+eEmMw+CM9sq9j4pb9cs4tyfQByaWmbq1owAiyN32zKhEa
rgp11qguSaBk6/0Ci6wGQk0P6GEcPMZHwgweAG0n0+jVuchUVOjzIBVXWt+pBUai
owuGnDP5iybX91WIZ1qSH23Ayb7OUH6X/fKDTKlN75xaZ+k6/ykI5banBKLjUaJF
u8f3uZIDr0CihDdVP/UIUoR5/blcqosmh79DQKTe3FOLcFnHfRRmlRETVlOj1Jc8
OkFah2O3RDPvDHxgy2A9R4r9WmEb0ZcRBWu3Sft0rO0RI4IPUjHhUw6IKhzusIyB
ZbsRRuJgtcKv5P5vXCTDdf6dufDQR8Hwh1TDvusddip4vfOyotTzqcUIeSWHxjOy
ZBNpv31N3Hf60nXCR8LwAKXSy2WhtrbH7VoB509ppBlRaPLF5qezkkMOg7xRJmza
LzanVz5+zkXxzyX3VHsj1pQONASKRac0u1ZmQX9lSYDxeodh12DV/jJYmWp/a/IO
CJGH6r3w+g4RtybRzv2pHCGfe48n7NKWVL6xlJEAxDEMwGZ0wT/Y/SwxNo6NKIVB
GcK/nbq9b3xzFqOnjAZG3UcCmtNaSQ0B6DeqbbUpAStinDQJLHtY84NxXgs5ZDw8
WeMgZwzt5vMfZJinR1EfyAVrY/3tH/2jM6c6qvFi31WadCT4XZ+xJsCgDv6rsKvV
HXxtULV3oR+78sgy3B0/YawLAQ510i+z2OKfmxOkdolKCLBhjanB9vpSl8ox3omp
Uhsv7tMihXTiUbWzBO+SddO/UozIcbqjWLrf4ndNrnuATpKPzu+o+f2VbVh8SHOY
oVpnFTvzFxSy0oFPUgGMqWVtpiY8g1fMTx8LNos9texX/AHJKp0KfmQcqmiKdCDC
uNJa5mnaVcvppb0c6+KIoPPoBn9R7wNilpTpWV3cR3XaB2gqyrw0MENKwr1b3ktP
SDgz0VefMrMHfLc82EJnGJoWVxHqiw3CSumWQBzJ6+ai63bK++ZI/8agRaltZM5m
26bjgLysUEejN2uLCDEZ+mJuc6LyUS2CQuFa4/f3GbaRPH+wrIruuP9rX5Vqdc3i
td3X3AqaP/d+RrhhpLTiDzS1/QqnOSlxvgf0faijf/Tr9HsS5n5gyJw8Rt1p7ZYb
2CMUo5x7VTmX8gTkrrJ5MKosy7dQHNEI2Djg5fMvEYGXy6jApXFp4LMPVkEBAq2G
6UyypMJUpzJ/X9Sht66M055uxPinU54fnUzq1+70hXw6ESFiZ81MIwCekVoAdMn9
gmyLvNuZkRu0Oq/at4+kaYjfRCmeo9Ysrxvdph6I6sSaSneI/ClpzzTX48TzeXDG
7S+eRb5TR+240m4J0jywJpTi57puCdefHzBOce9aGVDCPyxjESrFNwkMgDibcOM+
8mBnDudLfg5R8nfEXh2WACxXr/5hpTjZAjg1cWepx1DSjn6glbvMS/QVc5vUUSV9
tZ59ax2MahmKw5ldFD4J0SEVdrAVfBRNJN+vaVJK32u+2uFN1Mn8Qf8s+8EdRMjM
1p5Y6qhVXnRcZ1s1t65rmk2V74pI+O4nX6yR22FAw4XYEw3TohHU7hdP1+7m93HK
kWbR01bqXQnf0Ur9Ox3ikcTHcv72z15bkyNUUr6zhwCLC1nnrQZ3HZzP+NOaLgb+
5Rw594eh/3U6VQPv2DIhpZAa/n76ePtwomEH0/vEE3NGjntjCoDnGIlwu9uXcxp+
IiPTDi9xpXFxszs3UR0F9P5qsGaidqUzgsGHWoyR1WHqyROkxVVdZ1c03dSzUOMu
dqPMSLDuYaEJC3P+qHRrZiA3IUEV1ULyBzBgbR/PY6fiSxQT/m4hLfcJ4RwD3cR1
XdNqV3xsMEbMMxdvKqpSeVAJTAnXYa8yuactSZY33zABsTPnis9wGGAixCY+XBio
jYnVBl+sgQ9AHdr7zWqusUIajBHgNV7sXjsivC2GXFdLaG5s8Ht9rkCnvATtGj2l
0GJwJji8/9SsxM/8Ef2Rh75MF2XL/JszbWbgVykOVoBOfkLYB9UHSJyOkaS5R+VR
9HMhMcnsNQ2z/d9d/dadZaN8Ct4Sq29zdbOzPNIzG1hJRGvg2/oE8SlM+oZYrCEA
OZwKDCf7qr0elyJH490Mk1l077HGUYyNqW7reAncC4Vr9U+v5TVIhs+R+btVo5Um
dKCpPKEt8jHD16pdvkAOO4AxRXiyGNQHabBqQGXaUDe1sUax97RMc6SbVo3v5ZCD
0XIcbhPvIcNqB6n1AIoRLJJ1vnyAOIMdUdpqOyQeheBd2NlLP6oyO72wx0CXe4+E
hTGgzjLtaWSY22EumYaYVWEon7xvNKGs2xstAeZChVLUafhLuXsOq3t17oXiLUYE
jrRKdlITd8I1nVNubDu6G6uZpp1TpMawK+qM6EIfVeFp7oXHB3A7f/5kVnIxnG2F
JtpBr4jwxE1KSM/0oS2rGjzcEhaolFFjLpBXWX/Wv+zw8/lVEDqwSazL3wG9q9iw
HaN+huuCPf+dOX28lA06uLyAo6lZenM87oP0kr4SmzSsGAiPPI1Qk+thRsFXhbUZ
qYTNsxHeRJ7MhWDY1o5PvsK8rCVgN4TTUgiLoTcB0vG5qokev377qt2yPXBg5i1W
+uAA0WR2ddQmNHmjAkAEvvp+qQ2pAikbEiZJCt8m3kux66JJIgzmOnzBhfIC+SZW
qvJCpm1XLn+teIx+UYkxnQgMfGE1T1GUoGa4bqkoB1+2InZLEzRSqDDN/y56K978
H86REJw24gr8w8UdtJvbOI6mtiqus2bOcjJK083dqzDQlGn+uZwEh2edyDANGbEs
7G4RdCnqbbVCWc/mOh+hoOgziJxOHum3mED4SfOCxB1s5THx6gbXTKeEpO2rDpHS
6Ds7bsaYefFd3Pz9xV4WAnwTmTTHm7w167p2AIRTtjxzUKSn7vzqGcHeNM1vXGI6
G0v+AANkueHId3NELbzQzeZifCGJwWh6Ws6nEDv2bzLdg8Rzo38IqcEXwMBcgxDC
9OmKM9BwbBAebA8Pcc4zcYcVCW2Di3gb6kTUo6Arjbj/Pf/5KyPd+UMoMQEtyKl/
wNgz+842Dm0ftzC3WGutJxfgaaD0u85C8zvffzHI30n8IAUl+LAGWZwkISDXF6bM
A+XZGGFxPStquTG52LqqKcysuKY6Y1uJtfjYYZItbYRZ+c2ONnND6ELIX/zw9p/3
/aLRTn7HRkGIjg0+sGVVeAr8s6+/huAoj77rHEMXy7Qmi38rAZ3u28IqhEmuv2aA
PzIqydMi1cKG6r4vXdkhtm/oD25fO/bNENHg4DAQWaiwRIfNVFy5N3x9mW/LPlZ+
rGzugpOltCdOBssrN2hjCP3g/4D7Dhc5T20mfkbe5yTNluVHtUigNr1TkXGVW34/
Cfu/rLK2WfqMvHaylpC5s2sgdGxZIFVYHWErhnGNyk3ISpZIrEP48p5YVUE5X05z
hU+GSVZzGa+LFMep2nGZzt5xsytRpvPQNRbFSW6sRXOFlqgJwlP/n7d5DVrW1g/W
N5nxGULmbEwEbEq04QoVlZtNVoqePYvTzd2RC00IQUhUeoIL+TmJSA5pCrRWED11
WkncFyZIZiY4tldVOqjWmVa7ndWsKb0abRQ/i7Aj97Hgg0fDCvUP770P2vX1OEGc
VJ67cVCXkxq735I0lNsN//YGDF8ZyIoO4si1GSI1gRAVecCk5cjLvL6cW++IZDjR
ILtYG3P/WdQ/zm9Co63bx0mFBDhfXS6DOVWMbmhKo7Xciax2DvZbUFoCvcbRbUro
CyZhAsqzhtwRI+7m48g7sE+ExPUgoY/8tFGmx140TY+VX11o8seOlfebiVeZsSC2
F7+zqiJWG1Bf4601pE6iCOHOB6uqLBcOjymssUmg41sPH1vPVyvsL3Aa8zFfZ703
K2BLl7CI7MCAD4nvkzJGoyM0P5ltXExxA127kcQmpaMjr1x8f6MUnpABDQiGnZI9
qBwNz6SS8QUkqZlJ2CiDa47wSpgv6gaFOdRivxBuDOrovCuwmrcrqfM9ojYB23dm
VjnJ5cuhD1TBlarU3apWN44O4usBxyaHqFVV+y3cH6Mc9+VbZ7jDAujGW0nMLxGi
CeBzz2BJRWemN2/u5vX+pMExvbenecL6dALl/LCjuAMNZEnWP6MCEvFWJfmsnxKX
E8A+BlbYWBz4BrIBQrOWKSgvQ5ZS08xXCnr/Qm3yDoOQL2UonX2zt2QLMl4HkYUX
kuuw+DyPaRndlqlD30oaw4PQvgDyIbADTomZ+XCVtHHavzuHzDH7DOwtHEE4Hupw
Z14JmH86/PsD9v1r5HNv5COxlMoK30xRVhB47vJLu7fTS5IperljEBLVH1MfxEVR
wQCOZ7zSAhnd45pEXCle5kT4ul3f++TKwEXdkd9rU4Y3Nyso654fOOI+OmbC858Z
1pilaPgOw+Zg40BWQ3Tv+cEM/S4MpCrGBFlZqM1ABEu3wkxyMfH//wu3BFzKNaEW
GdHwfcWn3I48ZyWX4R77e8rAZxn4aispfE4XyMY5xtXSYF26SwYizkWzLndVsesX
y0eayWphA4+FodS5uzLVFQRD6XWyYsiX/7OGRFNA8cD0mF+xP/vhGt9dr50PJFhJ
0kpKNz72zNjn6jJzi4OFrMgH4rye+pjTEg731qnynf/9Upa4VuVejbmr2wokTjkg
qaFb/XTYsnwlKJPjwnUGVXdAtL7/3asUbZ4xQoSo1U88fouFLrMNWMHsQpHbuub+
DRrA0l6y1FbK9FRL231BQTIzi6QNZzS4Zd7l3jTsgACgYEbRrqb7DsYSP4IUiWoW
8REATm811MeY+Pru1JgOO3hk3q1822seEJZKlBoVgZwAlNh+049ORsZFIHkzZ8D9
LqETjf17qA9Zklb8pkb9RcYWsisZFOmO/mqyoTenagjWL7WNi6zBZbxA7Dl2X8eX
YNK1zhQ9ZvJGUyzODUGH4LPPi3H6q28HIik/Xq+ZU6UQWJ808ozF+e8t08fbxp1G
G7mnldXVa630mKz1ANxY1t54OZ/Q+54Og694Fbc3zBXGzRzIrWDuRH5s2+d0KDva
y4TKz46RRXvX8lBh2cBE1Ngz0DaoDF6LLpH7bGuPpbGc4eKOQnXMBYMZVmnpyEZC
V1AkoLwSB6TJPOL40M9rLRPSUVGwd0ZcAf4AAMv1seE1Beb7vmulImRwBLZsUeCw
y0A8C3BXApF7OwVNhy2QzNzcLmqD0TfDUvepnyjGttcZuFThyuHuJI6+ZLjnjGiR
juh/3tUvudaTbYeI1kd2JuQAB6sLMcaKNo17mYRcsIfKSGSz6RN1UvyjwUtZFhfd
UccUC5ik6OXnSJY8sBKeB/ncHqKoKH0mGgFR/vmN+ZN+VoC+zdUBhtf7OkzTQqtV
jON6sxpCAmAl0jBsjl8F060Fa7rlpoYJKxQZ5S9U/2PRu8L++5UXslob8jk5aIU4
e1lnGPeugJVNzoijPTRL6w+mmz3RhHxCXhBboKkhcwsorV0kWqGWYRQ1mMBlRt6h
BnmsoT32gXb53p1PrG9+RAJLhyBISyCqQV/hyvlTLxRyk01sn+oNG22d3PG8ydiW
ZDwOCTYb0SYDwZw9jwoAPveuR1t49nrZoDZATkHKIGL8kcrVDqllpNRGnYo/xUW2
GIyky+9ss26EiircW5TpGcTrMNIdbQpnKg03B9bGlE64fH0DDvdylcE0PYbdUFx3
71JIpgS7PBVseBLTOxPElgoH4RpptwwtRVFVjf38hCkD95olFV8ddI1k1kESfnRx
Fq2xZU4cKMhePFUngfsXBuR+So+uL970cpKDCSDNRSW65OgsQdgM+a88Ft+WaSRQ
QhnO3503WUtK3AV2rxfgx1NAP62h3y9iWlqJclgesM7fN12CxLzAbG7RB8hOzV/4
WuP8m7mcqaAFWBu94RwmglE9RHWwiq9KRWwWtFwMy3G6CXf8uBdh+ft+yh9bUOv2
FBunwuzU2mNZSR3CVgYFlT2rBdMFvrJWc3llxV4v1Eg8OEhg1+0cO82cyp80fLZ2
dEOAIDwHtaN34/YaxBUMVLWgHCTtO6BcDGpPnefCwif+ASLw31FSjwn60qMxG2dO
mgJc82W9j5ZIQTrRcj4p512VTyeDCOvcAE2SBg5pwO+vF58aEJYrgTiue59Bb3Hn
AMWdiwcSldo7VFUVnrP41spvBV6IuyjK+0TIb1Fb1ehEhjuHImpiXlItDiLLkZuw
4RLBs6kXTECr6JU6TSrSluqv7Hd8RDzvj2Wof5OeBCBAhtac5GjKckjDzgkPJn+u
nx4YY7t35muPq4xpxL8CT01uuBludljC93yVdsJUxeFwpXEm1NJEyYOObIBQB9Ut
t2udkV8TPkUHBf4QSLpBhGOwy8uX0YDv/MZrZY7GVaGQdV7aj3N3SbMYiOmuopXU
a1thlKJVeMKHaOWgTR+3+H+JpBQsmfoi8bNmR6Qhfm5+088VrQiezauXw1ZLmvOv
9Ja/Hd/3+OFEYGqSxdnSNRSrfu9SONmv0PcaMu+DpA82ZBbx19uD8SBRLviJFOAO
BAXeRKLt2seOGYCWPGBgT4afwNR87FWWu+nn8Fd3b187NWJPcgtGEkKVUUdQjlPM
c5hW/g/59d5BLPUDy8bR8Sq0ZEellb9IFLmWenKI/FZFI4Ez0V65gs7w2JVQF1FJ
eXRB4vcplIBNOnk6xULDHPPwAyAvC+q1tJWbOJQHk5rME69nkk4RVhKOD5fHwEPT
dw78AcxD4XLUVRZok3EFP733UvUIl98/0w3J2cIshBaGtlSSgaLrB2YLVoa7S+Kj
LNUACU176xAYBy76kLMMcl1mzmx7fPZ8UC4TfVGrzSi2Px/bJPE/4Gxn7ma7MBIx
O975sXYsZMqP7+hRTUXUQn38nkaOFHYZoz9wkuXGdHWxpeCOSnyx8pWphuAGutJc
RCp7jWc0VRX26rUp0sLAgGXaLagIpJEfiRSB+pN9oIlhy6bSW+Aumh6ejt/lxb5j
YPhKbcEP3dfzUB+0cZ7ap15jrv6cDawwp9haWk0jrq+Q9rkmYDSJ2RTRispuJ1UA
6VHTnEE4L48KYEN1rtUHcn+mhArdV9yChl/T9YppQpXny3QNt94ccxGcu0tyNiSV
egcQNR1VN7KgQYl00yz8DDTYI9i1JkLkbWbZUnDAVrycNUXXxzDz6r5Gi6fkVgFE
uHFHYLLVCwWA5n7IQaqX317Gsyh80Empv2KDmTaE0+fpiJjiRE/kXN9u/+rvM2h5
UO99/kTDo0DwfVJXoke1fCRtjwzj1injqYdmKv6/23d7hHz5+p3+gHcE2u56jGAe
RMPfBZfy8bXLztvs7MBM7HsZImcyuhZG1mkRzqzHI3cAPNQTnmxmpPtFKGcZsXXX
vUlNv1PZqYqbKkByCLMr209qIC1erRKXozFGJ5grnhbn8P+gJKJ8HKaSDeolirTB
8weToxSDqKB3eTq6sx0LecUC1CCZfPDXP0+dGjo+MtdHDqmvcEIyf3ktswC1m8Hx
EUJ7SBFY68j4lGQASrr9KN20bS6FuaQt3eKgv+8u+tL3/dcCKEVyXsNptK7shhhN
fM573/hNbW/aehVctj+wATvde9yg3FSShMN0f1s6zTNgVtY7PhBltGrLkfqA/05j
HQdbDUgWCaqYBDoeRh4yJ7Whr1MmMUrX0gfZ3oHrxmT3ffdDd1k26Nc4fX6jib30
OC1Bu1QMN6dW5iRR3rhI8tQSNqi1+w/w2GytG11KplucvDa/N6mg6JqdqgUhs1b8
LEe5iuy/eJHE7sq/UQRwYbk9P/Q6DzLICpHb85cjmweN+amaCSR0+c9dvuqbYQbF
WUK4hBny6n1OQvJIhEf4Vtr3pJRIjbKjCv+XlKB51PIJpjzOJxtKd/bzqfaDYZw2
bj9fm2jtHwHmW3g3yxy2zWF/Wu7CCdTC8Usk/8C6PZyDtILDvEij458UlYsTk5He
AFNCqhjnxPzF7ho17AHVuABfxI4hdv7xiRalaeIylKxW63dAGtVQ5ILaeES4uWLM
cm5uKcOh5UdkloZ5uDBbG55e41wwNtg+I73ww1jaHfncfyWsQdfnjL/ICiRBsVKc
GRZNqVlJzlHskneZeqHNR6jnktgNiC6EwU/y7MBQqdj8Lmd14laxGJ16QWDv9Aq+
OlHZ8IjfFLnwlLd5cexHOsAPaLqPWNPvIhGwGemwzZ1BTUCEkVz7aBGUT0s19a3l
jL1rVrD36kTd22rXzGuQXQ6/t/X/nMDkiv2LeVgjGwoX4TSF7GOwpiwetDqMMb/y
mYcgL7jqDpk0zWuQbIRQq8wxizMVk32eI3htWPScRAfaLT0oKztNIYPBLGl/DhGc
jeYuneuJ+WbV36qukvR04t3no+uo8g21bwpXvYprqQ5G9L9xrUt1lIFVWXkBK+Z9
58LKJ0NBhaHP8FEB0PMb3bOWYL94s/Vr9YbnvGTPmwcytQViU/Ebxc7JKHrNg1pL
r3rXKWD65x2zUOOJ/w40Y5JSLryTzOLCem/Yj0aRvnU+GY2unt3A5rDT5NYBDxWD
Vg0KTmFeOy1np1Uv/8sfcjCbsDJOSz98WbbeJ0tFsaAKveXsWuX/2eH64tOsVC0U
RZiFxNyYsrxfb0BoZQR/AVBrFDcHwpJTF24uUqTmfp4Nt69HkTCpwUz71AFSTeUK
ltWarfsDzc0CotRdtBaGdiB8/kI3qX8OW5tGpwkJC8bdnQfB90HWES8VKhvK2Hym
ymNYxTDbBu2cpV9ymq2i8fzuzHU7L62dxklyO5qxbVBY5amvoQbQk3C0UHfsw4WD
AWUMJnNYFIUd1eCftTPWGgSLF2HR2nSwg0D3J2KtmR/nMoHFaenkElMerCGwEQ6W
/9bY7npE/w/viuDWvkQuHUFTlx/OU7Qi0WbUXle7E+TeThIZUu16mOwR36PHerFD
0h6Zn9w15VorYBKCVyLlreROEkONgZVKR8m91/Oo5yY5oMTQVQO0HdtmPim7fFou
ZJBBlC6VRef37UH+rl5dobYfsxapx5n9kyhV4WfjoIXas10ccMmGFi6HYH4U9EPV
Okl6w7hRxfSU0ifnpNcwR6Lo0ruMXTplLxFAUkI00r3P+wlaVn88+r3gacqppC8g
ITMxKaAGe7KGM3HADUGq5W9yvJzMoRk6dQ6SsBeM16KdVVh8bi1fx6obU4yw80tF
zhggwFz1imCokKSe3gmUozlAJyg0ruXM6p6EClbRlS9Y2GzzTQTRRB4kAVIxf1X8
lzozkCBcxAY1vEzAeHxu4uphkwD1C3d+622LGSqDkYtMoCMuyZnd98bMN7hq7kuE
gzHom1TDwVCTC/ob8/xg0uxfkrMwW6dmg6bNt9SyoW3J8TyVcN38H159LHHNTuhe
LgRW419AfbQTAhTR3pmO0k+gmiB0wIUapZ9wUpTzA3m6WLDeHgMastTEhVysaa3z
XjqMWZsZRUil8ABbrteuVOadAEFZ3nkvzG6fC3ZaUe9z6gXMGvJ9mhj2S2efU0r3
A1YkQi0gXMupnyUCbfo0aC3cw4vKjQmSjDH7rKF/toZoUkHdSpVJ+Gk9CWavVuhp
3osRpDK8U5EmhIbWIHvKdvDDH2ffEzplMc/Y5kviqy+10Ixpd8wE59POQXmY5cXC
nGYIW4tnE25XeC2BAhBe6An/bZHLv/Cf9Vv2DE83p2qUd+IOzZEGWMTUMrfNY5OM
Fhl4m/VX4OsnAZsv1Kef4bVfw8ID7/CWojyb+pp1YkJd0Wx4BM4Z8M+EhvmAN0uP
0zk55qRJMML6k/iEnx9vwvAsuFCFFyiwXKHHOP3JpspKq07SP+8nGxlyK8fmTR3C
PDHg/UVVFjd9zl3PDGVS4V2bd4wnntCKXRab2FyziPUOIRx9r8ObQ1FFq1ADJ2nF
bJyv/25iASnsmIg8c+z9jioO83YO32yC+R2qeQTiWvnkKOnAavu3pDZEvXhLM76y
glcTgKDxclc0ena3pq0SK822otTqp59P/+txFATVsgoDchh5NL8D7nX95JBhv8Kh
DsHM7B4qeNG/+o0Eppom7EC0ph+Pm4Owl5V4pr87uK8X/CNc5FlAXW/sUH6Podyg
l4J2SJS8ZmnsTrQ9U/vELp9zaT4f8lb1N1FwB9ql7OTYFPhmNmDc2aLIeINa6FKq
8bNFh0BYuuZCC9MRNrvn5rcw+FnMzypjeU5zsOtbixK/YqOs+4L+b9d3VyymgPzL
wlIWQxvAe2HcJeU+Dai8dU6PZ32b1lG3WLF6Tr076cHSGwolJ8FfWq4qF4Ssy99i
+Ks+vIpBzXyOVqW6So4+VXZStRzBQTmKD3l7UOT7dnhB/J11Bql7jQe3XcOKLVNZ
jax+kU0VwjlrwWDVZQvxddxRdvtQbtovDZRnuTvAL3fzyvPZsZR6ludiQL2FKwkD
CGsuK2v5iiRyk38dulQyxwQzqT48VTQiILTs4acbtZich4JqCiY9CwZ8iIHgJqBp
QGZWK+7eAsYNYIIdcQ4qBqqxUVNLfX2Eo3+nzyZ69/opD9nNfeRY3OiqHoLTD8PP
AS3ZSRjmxyo17nK/BFCBIzz/RLxpZNdrFesNWh0wYEsCjjo7v70+3D3puZS/knl/
zSL/sRkLBqPVyLJfwUZuezaq55bqAzhHlNAGmJ0LUQmG0TkppR3/k6HGufLHdym0
y8FCWaxLcQYqiuqugLvsNiOA12IEYw6vwro8HnJL/M5wcPtVZQ9G+wSofsA44SsZ
LgpQntfCtT3PlO95mHFeoR9CfUo6VvTIUNLXTmFtSu6tO59Q1wL+M9z0oxQd7Sxy
GcJSM26e6ISyJJxsSe218v6bCC4qVEKKfcjBvrZt0t6i1gpQihn3QheTUHOrnUJs
vIGhhkJvEjLO7fBf9mhP5Sut8NS7Sv1jutDP8iy+mvhE3NR9YflH7s9R5cgtfRju
oRgdkAFDRhmtT8RcaZNLz4pCWZ6IW1URWP3VNE/5zo0ZLqh+ysBG1w7ufjLweX6V
SE81EaPxRIRnA20fiI5EqIZqdxW53YWSF5qrlFX41a8VWdo9/IbsPUB96esb9Wyw
B7AhKrUOgwq+lxveUtsGeOoD88cH6G/IRoPAiZDV/dfcOCu6SgJ9H1Szf5f447BC
B0apjQmlDgHvU03fwNIyH6NcLKztjjWNSbiH9uu4Wru4/GBCNp3Env14lTfp10b4
XPpD0nmOVZsGmVK0daF7YxM0lMDBVnd9+kewUFq2WgdTNjYe6sUiLizts8DMbnl+
DBxeDgaQXwjhafkmaD0DjCyqtBvPisiIXX3eUKoo32cMvb/S+QJC/kSfkzXNx+jc
I7zzGiiOdS4SKbIcI6mdL5/GnpFQZEFuMxGcH2SPHFvzZ8TF5B7loiYXwmIVAkbL
/N0OV4LUkARKXgoIhbFbszIr3myp6EhJUHC8egQlwkL91bCT6LrN4owAtv0GCiyG
Gmt0VNP1B8mdsysfzcIHQ7aFw/0jXQGJ6eoMa6N/RcZxBvddm+GXnCicDD0+q52v
9f84Q2MluvWBxzdph38J4etflvjaHKT7JoqaHbCs3OOrGHFU9E2iLsacTsSQj2e9
YXzvPKvoBMqgJnVAPDn8FfS/qGODBE9n2/LbG2YEF4AShyQ5OmBdWML4dBCFSA1h
sNyw+T6Pe9zdT4Kn9jUZeWotXGfcxwtKIWpgaiFeiYg4HCrxvotTPyvcbiVWplRX
9kuJVGvbRN5UyV/lN5bIHZPezMz+YLfHaws2l2Iv/Gl4fjy2Vw3pe3s9nKyhunXQ
FUijpBWOkiQ9SxTNrowQC3S7euxzDIQMbAwhFylebgwEnaknzrAds3W33MfsubEv
qCqaRDRQ0BOaO/W4f1dGKkAaw+O2X51E9tpp2WOEZN3nwUGBjH1y8O9ytqjtbNdB
R0A1Vgwob8SRcTsP0XsNpQyis+2zu3ZJFA8AtXo5tMZ0OvYsY3TjGWaUfTgbogxp
tKIaahOUSiLD7N4RhTZ9f6MBYbolBfGBYM9YCMqJUVR/IhKr+k1cAOwjKfAtqM/6
iSI9O76SGUfr0JQA6q1bY2luD8pM0il+92Ry5tYYaCw5qkVDzRWVVIJfuiDlNbIo
6kiCdvtyfZ+lQpC8XdEgASMQTw/GVn7xk3m3j/zgrjGgpUwkyTbjFLxGGQibInJp
+t5+lTHBObLliWd0VqLzRpz1AGXqb/DDTE8YUn9VqEp0zPsmsKGguCeU6xTvCuZU
EyQJYCpbJpcFpN3w70Vy054TQn8u39MNk3e+bJ9HGdOpQkSC9ZMbmYW61cBDUJ25
KeZgizpJ3YPDNg4537CiHn3LwcylSm2zBgBED05zEGvSzwfuXKW5iHKqzWTqpERQ
1JVlFhLy//RbeYCPouLaZQtIg7X+pLm1Ykjp780MowDLpc4bSX7VOyLcRdiDahA7
Fs5kakx6TQCn/cut5LoeHiIPdql79GYMuK0oustjt1VzKrxDBKdqfFEZrx3sIaop
5POTjGXO1Vzq0fNDQ3IpBi18a+hEZkJ0Ig+TzwrpOAEcgC9ED7ebmXKKXFhNGzG/
BpS/Jm/NLTytQ17TKgBjk7fbhhNEGGplqoNZR7VAPp+frg67K0mCiEN+p2CUxoAS
DKOO0qLhngLyvSZbPWy4HvT8PLRFyiGlIwuxd+HU2oMCZwe6b4E19K2gAZJVmzlR
ap3MmEIjVGNTfVcY2bQYPqs2wRfh4lBNREG+FdgJtD5Z60iecWvwKRwma3adAHUD
HqgsPuapzuOqFcKeKDq1IJtSkk2Y1vzN/spRUA+0aYNSqrMQ6SopRkggGGRFSoO1
F1UowG6pSd/YTMUfL4bqY76rHQY04KS9qXInrgpQdoSQOohlLXqF/1B6ziLlSL4L
fKjzXaxONEO21OTMsKfzBQ4GrEjIj/1w/f4XtK0WECnNtM3X5rFla4FD3bn8Jz93
fWYWdewl0EQSYSfgFA15NmnlGLtW1syqdctsL/G9B7T2y4wbYe5UFM+Emo4RoMRJ
KgGcr+Mv4aQQjHoApV1dxctbZHjiF+JXjZYt9RcVFrED9g3xITBp7W3Afo4JXmXf
eO8ALEq8pTJjGYbjTcll282X8CqHO/GL1ZLuaJVGihBEn2So9EBEDZZQA07yjLD2
0keT8Pq4hZBGZde6Xxe+8FP8V4ryO2HGo7PpXfrdBgF8Z0AInAYqp3VoBR+YUldc
Fdd4+KlRQzhreRp6Av7gsbQLW0gHsjBair8u/ysQxSVpT1K78g4SsZwNLVCGUbVp
2DKaGQ18HkUluL6TAT/SC9IQ+2Ck2VGg+W7pfI62NS5wk9tqmmNc88XREO0+XMYJ
3JTgypj6FNOr96SUIOBkj8c4p4SGefB+5f3ErxF/wKhUVo07wMOZzS80ZBuepkpT
GxRt/EeceTE2XxmrKBhI2E6wO50As0bmNn++nSE3SSw73pVWS6I2igFEbVFaDDBm
wIp7rkF2ETCppRRjxPafTzbyG5HjbhNd7qFvvX1sR2qj5B9TjwFI0gp3fsc5uKyx
hT2OrsX+6hvQFfBEnJsv4PuQJhyzcIKaaF5RBjJP5mOHhLgSrdjPpib9z47lJvBN
UQ4V79zUpWwAsdz6mJJCrAaRFTb/g1we/vw02rNWlKQJYWj0xMXJO49Kd21kj5Us
szzz3gjKGXZIiC8KOtj/03MvH0tpsWyWHBlT/jC6+PbNhOVGGzCInqdczwX+Ch9j
q52L/GX6ZCT0g2I1zcIjRlA7gCkrZM4GxXRQyCNsALSYAEf//7UgDG43Tozc+qea
q9AQOEQ0X0MBWRONqJ0UzhyoqcvXUc727U4TyWSjhugKdmjUF6AtMSphsVG1zNil
Tm8WC131COzmVmp53XU2Nkph12Osi+J1hz8+YKCauc8EwO2ZUgjwRiofSoufXIv0
bob84c3FpwSyVMB8wS+hqymJd35Jh9zUrijqQblNaJ+yRZI9YPZzPpcX4CoQtzQj
irmPhjMuybE66RcJrBGF9u+dKg8GOKPF578xu2vmH6oGmuq+T86+o2mKj7gsVejI
Arlm6p//gfsFS90PPb+3JK45Qr1kh7wRa9mEKJIGg1bxN49yadcVzvhmLDiKw7+5
/2zQGMbX+4eF0v2dNm4NehnKmT1dvwYN/spTFGQwU/QohuPQQJQMl7q4ByEqMQwh
bFKIJVMUC24yjpxA5q0uGbSRbzWbQI0MWiNUtmFISIgHWk+bDl5nVDdczQVCc9ke
hwvGwVp89DfVj5S1Dx4Vc9DKE7kIIQLYJCJbE8gGhYZYT5jo9U5eWkxSQuB5iuQQ
q/sl245JHmnMOp13XZEj0g3NHa8qhtpLSpS2mhf1FckNsqpjilBQUCuZ7Kp+I8CB
oXqdBN5SRmKTWJv9HmTaWw5qb1mVKZI7L1ducdLKtt20E1Gob00quwzHTWuq6xOM
mMrkqWQalgklsurrbiDSFHgWoqz7AsCcsYkZbU4vqZv0bSnhqoosLgrR2FywkMY+
ueqFF/HlbzV1ceQOFVx1yXEAq1GtCfVv1I1QhbC1hXaa/YFxmaoRHwnveQROeBRO
QgaVrVAya/Kbs3M6OxDR8M6WcCRYU7e/YFs6yh3kKllpMLSdgYp2AFZ2mc60XEDH
RdqLkdhOvthXrNGRTRi/Z8HbhINgD6/rSD6/qXV2bR9qMdA7SS1jshbQfFva59rr
6rnsb3UZHp4Ek1fdseguIHaK0azLqGOG7D55243OJyumjE1yVQc5m2FpveYfw6NO
FMp7kYtUSFhBC3m3J1Kie7wTuJKVbZ/0LuF4SZi15sHqzhUnFOn5UJrIVYVQHTn9
bf+FoOAPg1qeqKNBf68Z2siUBi9TIyWeAZHAoWK3LT+cHFGVQbzaKL9vaLba2iSI
03Jp8cHcLKupawUFhSnyGHO/cF4Kc/0lGugBDUyDJkz966HVarXymDoJrlvP0TyV
Escaij8yjitSAQFH2Z3LanArq4mqcohlzOJkDImFrOj5sJmEWxV+XjHBeAaG9GtU
AjS3X/V9KT9WVfQqJ72XNiRVUEtv9a1yBWqkTGlhuAPJhedA+Cos6olyf35cQr3z
9cHQJ6kDbX4gnGbpgSLwUQhinRQh5R4Sx3RmQaf0onGZaam462lZt3CJSGTKLZec
iPoLUbCnQ5Lqug+REPpCtdbJueJr3rJoGwUxdb0nCN1xTTpuubzjFRvekVqFitHM
PCu40ayxVW+QTTjQ7yCq4LYEwy0jz4Te4gEZ4nfJkgvg/9G72UivpD5qi4F9gtdH
QnD2G6tl5eJkSA3KdLevloQEOEGUG1aVdYRGrPMSnGFi3zjG5ECeJmSDD5K/VQDX
mMHyS4kwCS88UxbrWEzUVvPZuFmevitZIA4Uv8u7FhuMKuHN3H1anXbERtBESWbW
6Bpvqc9kyxYCQIBOqCDnO8mcqjlsiPhEAgmot34jegWobUvV7R1bL4inO/Tq9L0A
y1zH+PEvvlu6acxcBLpoxZiBrdGfjnYayLUJ2e9crGU4YDYPuDhEH7iTVOJ8CsVV
dfGYbN0GInOkJHPthq6VVw4vL1641y3L69J8MtDQFtaed4z5AhNAsqY1HU2Pyaj+
xn7VFCWQhEFYb61xWvsqJ3KrPjw9mUZK5PrZ43ljqjH7MQGbAHe791007GiGitBc
rT85DC23Ppgwusc0LRHCY089IEE4RlEioo1MvSOozVXzAh6rAlj41OPVvXBXYnef
kEbbTgYDRiTZkCSiFWFa9+AnBTg8gWe6VJi8iIEAAuD/HPwzvp2GyjoAE/Mmlj3d
rKd5chYaiHZKa2LGnLFt/HZ35kZdkZGzYF9bhWtqDtxJzAqsmriLneUE5odG8BXV
MlGkPt/RCfFbWa3BITwZ9tnP5GUHUSURgT7fjyPSwH9n27EVZT4KjcBKMHGo0sGl
ZI8WZyWZ4PdMPEb+06tpwYv23cxASsh427gvGTxexyLTfIzDA3dS8qGed7H7qU9k
LLeW/fHEFHlPS0shwmE9T7QDsa9cEcVMf1qDc5z6PS0MxoK6WG32G81AmckIvS6r
8aQdtIovBAvtTmlo7j3b1GsRWpQCwJggiDClsDuubYZL4vN52iDsed9R/raDc7e9
1gNdKbz5dlbyDQ+/WPVEQuPBXThZ9XwX/JH6cU94lFSkJAMYS4odoKMGyZvhLJPh
QDmDlueGU72CS+0ohahdNCRVkNk8jvfN9oiO+KHn7BsBfIi9pvO1wW+aPYmDCShZ
UhYFEPfyc1GaJDtv1uApT4MNshRJJVf4OcIY5MscOSIR//ovCDiihGPyW3QZJ//9
tCM5aXMqjdD0vzIWoRZxUBpZdQBXD5DgdN2cCbgAlIsfdYddISdyZrD+78MXPCqk
gOqnqh9y72ZVYXOidObrMosYqeX2Mab65zT/eE5fK9Aaj5Y2AFyBStuZnz8KEudZ
BPyyaO6hamN9Q6LrfEq5MbbdmBHil3I5Xrr58DN5nV2YINpiJUoM6LAgIv5B96DN
Hlt6YGc8GMPXzG73QBjznvS1OcyPjj/gFRi8VMwolK2Zla00V54s1FzRWU0U2hs5
QXnki7sWtMHt+mQW84nmnO5zXxMhUIHFN3xObgK1F3VAkUqg5awisNEtRY85T5j+
GLeqwrvxSX/g28HGzY5j3vZfTD8pogywbsOfpkR9Bw5lc26twAceX4f3tBCyu+T7
9d7sRE1on2mHWQFI8ybV5QrmyXU8B6AHR1NbEuPSEder0ADLYMA+JnXw2ormmcT2
e3XTyvx/OzT9RiFzA9KoRhM8XHsG82pGIzkoRB7tvQxxVQyUdXD+XrvlDM0q7+BM
nTOloEMX7h19xZBtX5veaoqnPRT7IncQz4XvTDqh3TrPfOZQb+lY67vjkViIHIt9
XGXnerwyBP7vEtNjm/794w5r6V3Vei2XKkKwaSLvS1+/mE7sFjlDegW2L63KAmPv
xel9lD1+T1KXl4A6C7YsI4dkk1Ybr8a+EJGb07eUT0yZVkoAmVH8K+Ap2m3z0r+Q
th+joyOwZ65plFDVkfct1SSV+51loR/a4dLSgWZ5y2agzesI7Cb3H3QV7p9Yf1EO
aICmtnFV6S+hwXGDy+wJ0Ct9juYDeJAmvd9F0+YSW2AKkG2H8GfM8/vA8OjtK9Qo
7YLN+hwLAX2U866RA8DCTo2pG1WxdyzlXaDb65mds7vXPX/TYmC6G3zY0XUe72ZS
+/tQ5dLjz+c9wrEPZjQkW0WUXdYbN+KTTaDNU/sqJKVViddnNcxRXYQ8CpmN/l6n
ra96CPT0hwUk0hHB2sVy2haNxVMVwe2o3HMzprRAMzfibMKAO7HZaM10xuVanjNP
JXsYZG8rnVTvUEn0t2uceAdLyFKKVrLbZcxGWuuEIFeWRYi+W5/6k/LZORcb8GqK
z0r+oFQPmE26KnujshsMnYwXpVBwKNoaYmwrHmmOGks3pOeGf655+DGocuAZ8NLK
Yum+5G2o1ijkIKbs5s9S7gKIqWaKuxWXjbBQExdrt+Fyop29OY0tCMQc4Eerdyk1
yIrO3RX0/smvblAjEmnqdScJboz9XUflvRbDxgHxfBYJgH3rgPgizvcGiTX1g6HU
EQAe8QgCuotw62SpXh3p1Ha0Ug+zVv86ULf4Zo2S5hY2p69qe6pJrKboU64aedl7
KGGFl+2rcVabju/no3tSqOw5bswjpUCRhD4tCjh4KCxt6XV6G6PyDkYl6zB/8Vg3
0QZwdlep3RRXIDEbHRYGqNvsbApk9zgnFyc0GDjj2Ft0cnQJ8t9Y7Q/s0ZWakhc/
6oUaGwDajDLVtzteuZUgUxJe6T9lKtbG6HLTD8ZYoF5MA1HNIy0MCspmKOe4OCd+
cMVSheooZQUESCDohEIWcnIWx+Sc3CWRA/HRuDkuwAlLuBY0Nsqq1httVkJuvJny
z4ZOnrMQPsmKnopUwSqkLhNfoMAqSRfbgOGE60/pM+yZFNsARLUJVheioRUou/eB
88Sn2DjhQbzgfJS4Bhv+39EhZfet2wK41HMN2Rt2rm26d1bhRJbs97qOu6aP0IFo
5ExxuGFhO3/x/IRKtsUf0q8MA7/ktiNogotWS2+JKZDiJsiUs46oppMpU9gBowHE
emgAyc3UnhcgEj1cTYRGkQWx/PrHHLvs3jCZsnQX85CGlExLDIoLQP+lSF1C/y8E
uwdIylpIfwwdBrZBnDxvcQg84Mb1Kf8PIQbPCH7uIbvd/Hsrq0RihDatbAwq2K4Z
Rln+hvxWrAd4PQe4lYzGubiQehmHwVufveu/F1dAaq80uIKsaHnneJHHlYEolOGD
Po8LBLL5NexbXiKsgeHZBTIeH/8/IJJFwzarzLgoHHvyHtdHaJuWYuEUBV2c6Rqx
saZ4XSwgp28TH/02SzfLfb8KCEDJ0O8tvUfqRIfNc3wdqK90QTr9DqTgMww9y+G+
gsPBz+ASsDxu2nrQ1i3jVbVs8/sUs9x8jTNaanqthhZ7WYOvXpOwBUoQ3SvIU5eA
hh9ihEvyYt8IfO6Jr4oq07OppImJ2756JQygXcEl5i6pO1UCFkxzW2MN6Tlrc1Jd
BCq3Po0yYV0CDIiMhJKYTQgABKNXCFnXaz3aZdAsqu2urbMH0k6KVF2FRJpsyo7g
IfLEjtKMLlQk1HLTG68B097xLAHOu5JykqiSE3TJTJAoaK3Oi7DiLm039bm0v+s3
P/RNK6sywnGF9DrXRmyVG+SuQqNVEjwogwsxXrxVA5LxJxD4hiX6Beg/x7FjU9yG
YlF32zjkbUjZl0KfUQKg3iiyPo2mD0BgrtL+YGDQypj3+Ncxjq2G4BKNZFRSuBe0
vU1N2TtlLKVP6508WqN77PeWhiNq7OuAVp1J5Q4SGLD+uJr0GSKVE2L3Hjl6hxKo
/PcbAG4BW8k2qbKX96DBWpdnDewAPZwu0QwQXTzZuR0HTjHed52nVp+sr+HU3pIP
ZTLBiXe5gEqcKe+mYgEQwxhJzkd8AmOaI+Efn6jRSBfOh/LiukmE8tAXHX5FS0kr
+KowLP/nUTzXSHZFQ3zJySErNwd92WPRigA01uT/2TsPcicUfxFCPkvS3X9ndKOZ
XFoP61xua9CshUEVSyOA18khFPkO6ta8/Dr5VdBLgT+e3TZ+TuJQg60C35NOw3wn
uGWM4Fjyqrh+Ydq1TW3IzlTYFSow+a30a0P6vjNrws2FCBDzpZrtkPXBGhRpRAFw
VZXT94k1PWRvRsooAuVDMpQRw+FjATggN+epaUL7cjNUJ4RxrRCUdQAZOyCLKGt1
yaNN7b926whFWrDGzXZi9mbbe+Tcl8odxdM85ozX4NTKQLbRgVw5K6WOob+WOKht
YlJWwh4lB1+RbwioJvnoy8xFFIAC0md4J87DprXwPZnTGVPRo5eto9dlTl/uDFMv
PTugnhOoFEDS2/zbMBbZecG/OKQ9T54gvLpJOGjCVL9k8kJM/sP8JCHTRwh7q2gm
Hv9KaiWsMloF7d33DhxozrXyenOsAUbMVN9p1xZAgXWyPHHWHvJSmhhVdjs+evBs
5g1qL+2czN2AOOa96zT+lD5SDkxzoNUjxwYgQj85xsl+FFo/UvLsrfWdthVgNKnN
TJBVRjDsP1zcgtkcR6w31RAaV4gG4XVsbJ4zbMEH0WEriBqLQOdHCoTwvkG8XxNo
vxpUFwOcGDNA7K63c5zfo8iHsOvVqASHvnV/L4CljNbw2Yh8tkXIESNmIr2ofKw6
1nyNGVrA6P8y3WgrbQX9ZbHMS/4+ttvDsguj/zk1Y6MTzz8m/qCggc/cRjjEG+ZE
elhfxemKjy3zthv3ELFchkbw/mWruyKDzua0BBAhfnTGB1Ladcigr4pMtDCFyAEK
BPo91yIOAcIgyIqQFd1OjWDJThFS2wnFiIXmI1aUku6B3w9CyYyHPx7/z2pdJcKK
MiFqOlxP8VwoAxqKiuIsw4jo17j1fVgqhAHxa+bBwj87bMnQEaOL/qT2WmU3f2wU
jZdD6HXJY8JbRVQy+V+M7wr4q1yJy9fX3SOiNGVPO1qJwERZc75k9syeqfpEmOZD
JJKP7AiQdCJDJvDhFt6kU8Q48aNtsQMr8ixZdJvJ/5nO7Q7B5V//hH8twCfxia31
AnRDO+VF649RpuZZn8kKevKZPcwgizo+pfpq2e+4Pi0iby15HXUY/Bt96RUBnEQi
j3S9YdOx2nLyKvuU+41PUvx19Do0vqnQM3T35flmZeW+NM0leHS3Suvh90brJqLK
qzjAB0xWOPbALcK+Mp8nHZ/dklFsJ55Nd7snhyLp2/Qa4L0JuS++q8TFeoxeZ4ei
l6kG5dLVWWh0j8qcKwBIIxByJl1HkXWA8S8eCZPpxEl9wDM8md7dPx6nfmnKCfHh
HhVeqLJ7KAiyjqcSrRt+qHYl7Nvu+8qjm4tldvxxCyGvnqOInQf3ZuXDAlY3icr+
IMtcBNyOqGm8LKLJwYfznAMcPp/HaoZU64oEKXsQWYJfypX+kMFuBYj53g8BNVUw
FwxV7xWilz/hqlUZd84NFbJzBFoP5/D/You8L+cN2K1elUbI6/meRtY9disQGEzg
rBOtnGIyYGZBfPuaSGyS8+bE4MaU17AmNKUK+Eq/NNp4UiXYF92VsynXuo+h5c9b
HGtKUTVdZFQjOWK2YDKz21EjbKz/tXQNmPqEmvEg5396Hflm4iNxQCIhUp1JTEb1
p8LDDNZtVtwcu8K4nMCTZe4mhh0vAcYZwa/C0KBhmM/v8PufVEMnSPli9VawnGco
M3AskJGF2wPFf/x+AhPAp2sWzJGgfZI2QizWB5cuNp3AdcrK/0Coh0qPtPh/O+0q
bKXS2R3hZGwiIkhuaYeTcz8rtPy5Jmt795B678X6IAQpK1Mi180BBONo4hnhivz8
THGuwZBsVCviC3j0fNNpqhljXQZbysOhrxGhHjEXEmqbcCydkRf9ksH4My8MngPn
XgcdMg2oxp3SvpThuLiVGOsgKGOTSiZ9n1KxsslI1U+2JR6dGuooQsJE79JzJybm
lCeeFJTjJZbx046eO9iUVgZGT5pZFModKZN4Kva5Kauvlb6YU2LIWOP4pwWvOZ65
sYKkisWS509yvHAwmOnX9BjRKqD1MQcV3MwvtVYwmWw2X2r38XbFVXLbEHBlF5h0
Yz+ZbDEgw8jgUUlJVYwwRTLcKnXmNqn7KaANA/sORBohF4mkYxX9JivXc/IBCPYr
rexX7nxWJyFHmo3TBQJbEuKV7xIim1NWgp/XxJSGwFgdkiKcO9TCxdrsqpfKY7KU
atLzWb68S5hO9u2JFQZvMQMO4B4yZguG4DNjBmGhNFUbKzeOWyTZYjg5bcrksoIm
fhRnrYmk5i8Eu3AGcVHuvIiNEj5BUvG2c4JMIefP9MPZLYj8p3+vVvPgK8xj3+IM
A7Gcdhzn90ib+DPxt18XVyqIBlA6FNQVTQm32IVrTrRA1iwNQcK1aHU0WHGdcKLd
+MPJKamtJEIOQMGzhXIb+DuIsP9q75hK4VCMBOd2/Ip0FYjcmyb38Bje4w8MS6mp
mpFsKYPtEcGLg7IA+ZyyMHiyMSC33Q66L9yhpTV07QhIvfzeuJGuBYlX7adFhJae
sbiBiq0+KWitn8DsGvqTUb/0DWSyZQsNP8/iVAZtDLUqzXwmTU4x80SHv0nY4VtW
5BsBVcnj54YxRFrseTi1I/Q4COAO+WGcy/EF5QGtaIjMu0GamV3Cp5buq+bKl0mS
c7EzobY+EN+DZacOWxQupb45NstWXpg9LSUykxYeq0GN3MeB63xbWuc6N/+cBhy+
/4foH96J0CMHpUJ2kkz6P1yhNHJ+1MIutcShKlLCPT2AleVuvLGjPquiPuG1X60v
+aU4Gl5OUpSG3wRNOCiZUu7NlkiKk8frOkzDjktaC/hKsAfyefMwUPWKCLbYWgWq
47PoWpeQvNzm9lkLOFyrKWgDi1yFPXSi5GOMucIvXE5dJRG93ewYaPlDYv4KAI/0
OmrYlZDwt2vKYanEpL6S9Q1W6NzbqsmMfehrp2hWu2clw3L2JRJ3DuPZkwwrr+Sa
mVznFoOGF9XSJwBh+ka2NCJWHgx5Fbb/8fw96c3AQP3mov63jaJ6t6Agn35uzR5y
GvIUn2CgjCtm8CJG6uMtjyKGcrktsE17MLitrWsUOZAmcvHgj+hjrljHJR72AvAj
00cvKET/Ssd4MBHCNFkphUbM4+aw0WSGPpOcKTKFk78P7ra4LUPCQgnV1VvjV2ka
6gNAGLOIVyif05LZHPtK4jHC0vtDKE50wICDO5h5js7M2IoLNkbwH1NMvrf6YFRw
CZOZMTuiHdut6errfsacHdL9K8VVXC4qYlOKQyBS4HadhhT16UDA8yyGz4f9tFa7
7VBK4cgV9oYDQ/dQjkPMayouZv5u5QC0mvuIEkFkhsGiz9ZhhN2NvYzKW/RX5k0I
vOBD1SnaxfQKf84B5lwsiWKiXfxLYRQK31U+7/Vja4h1MRTqReJ8n4B9vZkvG40F
accFUlpUHMlDg0JFXIrJdycEvacH/ENoVflola1+0CWGeCGz1H/ZTNSRkFKaG/Q+
+bRXsoQwdgEff6PJWKcBxgNrADYi7jd+3tJsjzhlIEv8NoRiverr0uGDzXMptLLU
54/NluosiSDFBI4iaW128d1EPO+8jVkICT15wgxCqOV2EYRBh11i1bsF1ZATO81l
Q9oDKXn0sbMZfRZmJVPONpMiY9+5bSz/S+RyzCpRYSjmeUOl0XKU3yxgf/HntokI
fPNPpDpLeHy4YOJQM221qHbhlcfygtnf69B7oA6OGukQ3nud2PN+wUX4vbcJedWh
UIODXki7fhWGwbR6T54j3+UHeaWQBsV43ES+ry+j8ayazeieA8382QvFpKPhz/yb
yXqztuBGQdIvr2L5FkKu1oTqZo4duG0tsI6xR20JJ9im1vbBnWA/yokHlhSbegpR
tFUUoeMdTslRrSgVOI/vXkrBILqSu7Lbfd8CxpJVWDTmj5X636flkabWfouxPYe+
KXksicmznZhyuqksKF9AdLlnkfCV+PUcFHdRoNbnApuyKUeEZgS6+1N+fCqMmbaA
CicuYlrsMIWvN7u+5BSAawJ+YVfI/ke7UVipuJ3PgPQivXIEEl5yun2s1E9HmALC
Is77+1Ja3zzhg7RT6zzRZRAOlFU967D+A6OhxtQx/sCVouZLvx4SL9JK3q9opcqz
krsniK/bvFEdIOpMufR/lWtkMHsJnpOHSEFu4NdfJX3S6+e6cYrBP49uXAavqz7D
tDHY8HmfUECHTIuuU02bJ2bvfVoQkeshff+04XQiTDdugguz6T+WeXhVfeEnXyn4
NbmQ3i0iJTiPukOrEXoMikW+BOwPaUegY0GVqhF3lAZq9phE1/Dx0ixxxTwLtf8I
DVM6BqnLsbp9vdeeqCeFEACPbMwMQ/d9On39YQJ5n2wYNjbUaFAC8HidCfW8mjJV
fR9DFI/jlu3lLSDE1jU1TGRkXKsNgQ4+XJwhD+vDgk1ugPbdjk/uia8rKRuihlWK
ekIXGsC9XrlqPrDbLZ+cP035l8XAWnpUPyjuOPz9GUx8s8O8Fpo5tIfDLByabPbh
Qhn1ciqdoZumK6/YW7T3UxHhDaAj4zblb8Oh8cvMgoFcZcg1cBmGEkBWeXUso6HV
zk6nJRpysPFAlitvxTM7Er90002Wv/eyO6I2SKa95BLMi6dtb2Y+oDAas+wKmKy/
kyBzj1YVje8fXAjEJ3O9FuGwIIw6/MfpE1lFx94jBOw6FQ/nVs7uflD+Lue4o35b
BpQ2C29kR6/sqY8QgBBAP5DX10l2xhRHvzHeo9M8S/Y7+fJMkZtDxT6NE8OhOu7l
MgGZm1gMIE6HRx9wH1ksBCbYQ9gHf7wS5Yuv1IUmMX/ZWD8v5kvyPfUMTwp8epjR
E3Dl/b+3Ecv+asbPtLQCs74+/kh3FJtlQeM1chtBM2bT2TBUTnedUXbDhAaT55xS
Kp5A+0UHfIVe2Csci4+5WAFQvMj5rz9ddQWqqLQJRrsH4Phe8/rJzVFhYzJcOSxN
Syo2ZHhPq9G1hCMBhAdYMmVwXJc3nvQsZx0gVFmEaP3l/JucB1+2laabrilCFa1Q
5tBXZHWBqtuUdOokSY76JRyhFOfTa8O3qAX4C4H0OI223+hYmrb9KjeJqyCSEyHn
szVQa0VUkd8hVCd9E1AEMZG33+DNI2AWQQHq88bxweRA6pCu3Tijr800qZ8CJ3Hr
/vlXK3J1j4JkT+bpw+8CRbvCr1lqzZMveQz2trfCXD74phhGgdlQQCsreeZn892/
VcXCl8UTG21Mn3eL2oiI4qRZ6P9udi7A3DV6ppJe9mmYOiosfmQq/FiV09YWFR98
5oAyLuhl3kK5Gxm3FXSuGCQtef4Bd5ZODRFJzEBe+DlHW8WNupzS47zb9bGqJWqf
P3a5xEgTXgtmNJABLkZVR+H5X1KSAgmuM4vY+mJ69uFHCdSp5RzQHMDea8e+GKK4
ta7EA2N/sX5OIgE0IYa09cJ+2GrDogzY5F0N9dgAKcLjK5iJdxu8143GTIhRn6yy
FTE5fInI6JlVnjy1fOin+0QEBmUJQ2GQ9+GZNUocWrjBNG1OuNwAaB9db5y/5emh
+oBnfiQluPslTAg/pGA1tAY+jVS4OCW7Z1XxsBGrIvBMLhSNmf1vw6jpwIPzj8Tm
LwhCpRCiLjh/naZ7UpWvoM4E+7IW0ri288l7q4g7hbn4xdrLInORZhfFDsFDC6ef
HxCXZq+J/UkuYC1s4SNhoe0B2HFiKPULN7Drezpz6EvKEKKcZzPTgSBTq2sJQrQ+
UzLfEiJqC45aMZhUFIhIL8GZjXZdLNuLlTsEeVPE6UyuQWAE/xTBPK9AJ9y1fKO8
/my8usImbfXwnuPbsLino1JFIeCMaFbCAz+Qv+mpwpTZpvzywbL/4wizjjcwC3uZ
uFgHJrlW/Mora+4apezs0y4wz3hPu133/iVol++tCqI36Aqi/CyF9MKkGmGG1/6g
xYz+nsYWxbA/PSzq/z92xzAAwutyxF9PBUK5rzdKo988MRaUl+5K+OAM0luI+5WH
yyvZJR1YotjmtBP0tr0RXY0vap0JUwGUt8yxqMdW7nBt0fZiJ63lHBqSFAYU6Lli
IFJhFMC7o314IuobFG4UAXhuA6x2hvP/3vIDH+N9tOTOUnGaqLSydkN9RunMcnKU
qUoric2ncijqUB8I+nNt5ZMBliNVpt8CRvGUwZde1xuYJ8VcDupSPpjcZeIDLbUt
31a3p/Mlyfp2+hD2CtHQxTiiaV5TJXh6xNL+18eL4XbQBCmjzkO9iaZ/JnI2sTgh
xpXr0eaHRoorS98IrKo/qBZ1Zo5sZT0t+vcXjj7xwK8jOvZuXuGNftzt9BOkXY1t
wETBQk2P6ILh8GEHqi9UMOqC6nLGbTj6w0WtBOB2yd5fgwIxTQxgVdcb+k/qdhU8
a+PhijUzErwaxdpor5CSvWiFX09YvWzpiC/jHjsaRm48t/q7nKSgaVNxSnt0/18d
MxdUYtxM0TD+tV54rvwAsyT6gQp9ZkcvjJoltIM5W9KhLnNUK5nLdo788tC5ZiD5
IODgOOUZSTewhsdc1R1UWpvhNRPHOpahEW25EpedxlPZQTinkiuEpKOp2Nej3XfK
BRt3gn8dt+SK4VAz1mUSw65hcLqEdQrgcwERdf2gqtgwYgbZHMUVnNJH+m2RJAQg
8cda3IVsfavT0+sCi3J7vxmYc2Ox2BeHR+W9aTTrPmEXFDz9+D50BkCI3kfhhz9x
Tp4b/ZD8f11LJ7J24kKXNxG7+dG/T6+SBfnNUu2XEGLa16QbvYV8SgZLsF0J1Tui
8lcVo5GUslYbtYD4IDnC/SBjd2TEBToGBKotsd/Z3JMsSqd4uTR2aOm55/v2vrWK
JGUyNVLgTE2YzzQtOaiqMXxj3CU2o3CAqwgum8HnKNs1Vrgbz6lfWr8ov9EZa+CJ
r2mGKGoL+1y/UaHX2fv99XIHnzVEGnHPgai35w3aMhhvY8DwfHwC9HMtaf08wqmN
lWk67u4RbCI1IG5kcQ4eNKD8zi4/8G+F7LAoj6qLPBC9rkxVR4fkM8KqSV8v6lGe
XaxiPX/uy1rWwj7OtDmrgXvlU+seIj+dUsBUR+NGpjAbparlyM1cUUig/QndKEAO
1ubZ9AmXgGiNBv1WTG6FWqdegbOYQ+YBaVebn3EKZWQ8te6F49xERZRXtMUlXPm6
0z04/t9DZ2tqG4qDBDure3Gz/8KlYzK9gjeorzJ0yvayyTOuwgqMflutVm3au+Ba
qrsWBRiuR0pv8ogUrG3PMwLVXCwg/wzIgLu5VQjjo/yb1Ph04AgJ1xQ997jNlsjy
Es6HD2z8ygJM6NuAc1oGwciACmCVXp6zJCdJj9qvScE3uqvBgnUxZplymBYk1TcU
HartNOu02ZT05taAd6se9b5/t20KyFIa+0aIS9h2LJf77Fx2q2NtCIhgI5aAsKSY
kcf5GIgnCw/ZMCldFAqhNAUhoij69dY9l7Vv3Wm+gn9l/hr2tFHZczd4Y2/ond8I
wVshq0Kv33EeP7PazCDxuUmd7HeCvsvO65l7WseUoy/Nv5PNK5R8omcpunDm1r+i
C6dHbjYb14jSgWdg0UV8i5scJiiTtYklgNeWjo7/iZY0OGcKNrKstpX3yr73GvAH
1wpquFCf2J3NmCdzRryOjeNgRIqhsRoBde0kpJ8gjA10RO49WRCsJfg8BSnDR9lF
6O0yqdxTiHMrgi53+xAhuta8hCUk+BedY+HUOe8Xozal6w8/MYFNQvw2FoXRdRV/
Cxwy1Vynm7Ix2VvYrcKZWehOg8X1J579+tDUp8t7DtQfuqURsLrrsy30vsanLzxV
zUbAaZ3lZptYTXwSUx+Cq1OK+MU8VGsQ/k6szY9CN1P0ZVM2D/3axovkv7Cr/a0z
SAvuOarTp3wbFdiQ624nPNGbX948OQvbxsXVyPwBoBwqKge7OTax8IvlNHUUIuVt
pAFTOp9eiq+Rn7eQ9oBnvPcNMc8wPO96JDgLUr3P47zKB8t7hhHvhdeXNuMTUiKB
S3br0hcvnD9aedXCFGtz2vM4SuxCjSd4Bb3gNCDudHPEPPMjkTpokm0qg35wQn1B
nwpw4BRoBFmZfhPgto5mJllaNDMBtSSNOWuitVrSZ6pIlRZ1gwTwz8zhLP8ZsRLK
L9CTUvYbwvhp0NpL8JcLpdneDjzLCYIjsKW+BEzksH6pdU3bpe+sCTfh4NTOhW0U
ilNKR1hsTL+NwgiRoRScchMtC8egJ89uP+8uW5wiMLi+jn+I1hD9IPejZmRmuiyw
vBnKQtJ8MALdyO89tsyNr9Z1LDwxMyOc0D/8jpQ2zjiaVxciUenbpHnaZhcx+3YD
g+wyk+fTlaLFrkzPDODbJv+5NoU4BtNCtt8VNKZYWUJ4Ohyi7BWslvuSNPPJPcG4
j0rawtHoB30xHySkhhduyUfjUB7ISrixXAoCs7EBA4igfsqua0+ZDUo5qlK8ysoa
WdBUcnNvC7hdwA9hQTIsmcLMleOFfafR5JGwAEDlQWJZvL7QVoR08l2r8WhIVzKN
qteCyiAJ31D+rvpX3LUP0pnQxkkNwXS3GJ1dBeFmJPZmvLblr28vAuOSrjzxgqFP
japSQnvdltDQQjwIwiH0HQQLAc1MH+MYGOsrfY0uGES0Lz3+cwy8YSuoPfvOjyx1
aXTH8NDJC025iLhOOrpLcFVAXMvW3ei6UVbGC0CDD6EDsbU/HHF3KaIF0kyQq6Wa
uGOVwu6+0gEw+h6oLc2BOYptymxHWUYSEwztoKheoU8zRHkannPu0pHxllCa0+Z8
GZnqFbWoC+huOL4TCwiJD6DghkcmGbrHqZRfYoHZxQNOxKTBEQQowcOWRyQmdTVg
b660PAfR+1LfMQXOhXnK2AWXJEWdpHXv5JeiEzABrkWjA0wDdLGyyF3rEZ0PuZIK
+X1gMROAh2+jwBkl1f9oddFdVJ8AYG/8RgXbp/Bb8YIwg3mpSsTrY/WKVVHFgLVc
tHIAV1PF6GRElZUbaN+bofiDyf+Q10AJlxWr90QYHLAsIMJbcmv4EojtIK40/FG+
C5860x43wCSXXMJ7U/DLWXeeYsAb7iYk5c5UEdQN7ZGyjBy66cKiyc+MvFwfQKB8
75tDuioKAGEKMS8ebdAiaWtG8SyQ97IMYQTtmM3Vqr47DVDxA2W+zCw/A8afQDOm
9y73FJNBktjes3zQdgdHXgyti+d+WIi3rTFHFDOhi79P2GPRLZMnaYerwxRORndd
O2pLEFxo8Cn351pXf9FzvCMgQMNjpfSTPiRwTaq6MiVJRH+xkes3V84WqIGd6P0v
QiWH7jQ6sU3EA9i3as+aJsxhKkPdPdleGP1ziRO/jIzyovvKPH//uutQbl6vex4K
sZcoP9oQypdOl4tWuiZsGsPRQpF1a+VedHed+4QkuF+92xn1fQwTLb8nSPJHjeVH
eJvQ0YC3akmR0Fj3BtOc1wGZp20cZHEtw/BDLUCNUH75a5g+1B5PQBXQvt3E1AwM
HrAxkwQQeWxG0PSJSJrzSwRb5wrkL5UtxWHHZomsi2afwk0AjVZl4l+2V9+Dxa4o
AqrHfi52cZi7vHycm1Y8awK+GVbeoMZ7BazB4TNMLbn7FK8uKyEa7T4xeL3z5YTt
dPIafA40/a2xwsbxhfqCF3vaKrYvQzpsRpmR34uTafh8GLv9m9VfP9lS58ax2kR5
ThlWvSF1MtMnx1BLZoddhvvQUaQpF0rGFKWHDM/8tfO4MO90I/vjQK6UZutHbg5m
ggPdvEGFsRimqn5tOX2k4QPc4sSFGKqB3PSCQIqMzOopWSnLgZkcAAEB7IOueo4P
NQy7EeIcCAthT/F4DYjGxtT/i3DpIXptIeY4Ger+TeGQK4a5a6V0uxcrF6jbIoHC
4KQiFTdQ+xdyewBto2rLEEi2LD9xcz0U11yeI2BJwcIs6GYfV988PzPbOcetgaE1
Ecl2oW1+SB7zTKJctBvzzS+dIr0Q4XSK17Hhj/lyZzg2Ohf7/6juS9m6GC0vy+2b
tqHh19II0qVFVWSVFDT5r8vuNz0WfF0pVPoO2JZC4yS/TNiPKvfzgQPmzgSxD0+U
ppley4yIliTVuOYcsBCXP6XwbgRd3sG1XLduDAwa6q4bRfGlup+Mw9/2woW0UEpv
Pymz4uDoMne+vmIaA6XvG7UySZD8o0d+XXuU5k3Y0xlAsTQJpfpFvE8tsdCBq7rf
AnnqtFoRh293ACDqAyt8HM1PAzKHy3R9THuuMkFtXcHeYHG+y+QwLvhX+gI9EjV2
BiGSFXgegNWNQxQlVbI7/wjAtWTUg+GVcdY3FI/mg2aDTCiJvsKqLMgxWNp/l4Px
e1mGpDZ0wns9M7KqTEs1vVz5fIp/8oAdjIEVn3+uaQZBQoBOPHy2zwakARsY4+/N
7X3bXF0ei5TL579u/3sO5MgyXCClMBKEXJJaHSjGzD2n9GeSXsOaR4cIjk5CkEV6
890mZwq7phiPpKDdsHWzpCBjJJSilQCcwuVFH8K0NjRQ8VCxsGZRvsi1BZZ88Iyt
QgcKxgjxSIXIfiF0eI+5t11eFEW2TvL9+zF2bTol8tt5WMzUjbTgthFh99qCfD9h
5L+WXn4iJP+O31tEf3Tv5/j1+h9BIbK2yuBTzd8vteH7tLiusifayo7ciQKn4egx
DjwHv+1zk2MWu3FHBEUmBZy2C+9Jw3Ml/j6YKB3gMAu6MGiDl7ks3pXXxoqa+h+G
BOxqZ8Jm64pLe+uXSpk2ARqHZGw5jy6e7i47F+UYcNN6eN0GSw2QElIgQQ3lay3S
qwSX/5Z+kG0S0zSEWpZHPYiypHPQFn8rHKu82U4p5aF4EIx0ZB7aaurMlepvBHpG
lLW/P5d891QzRTEO9tnc8t2wYaNyx3/Wh45o3JepmrQDp/07vY0a9i7oBnoBLn4l
lWNAffsGonJWYPkYTPmNfucNGAUyuz/3G9ugVHWwlcnDH9ueCMJCw06WvEdhiQiF
MVhNJ1+H93Tah6NJOGFHzGaerD3pTSm5Q/Vq1T3CKHgE1Mpv790fbYz0TVvBYSZj
ohfpMAxbTb6XiJdhCuf/h01xSUod5cbJ7dmJmoKDWZG8Cbee9Dlw68wkINsvJPjK
M9Yx7uzeaSGxooicy/uqXlfJ3tJfK41bGHjYWfaei22pZX9lm1jz4u5uZnd09AZa
xF6dt/8JdYNwb+NfSpMS53DYu0z72ELdUK7cYN/t8Gxv7T14hD+L7VXFbqzjFdb0
M3fXktVWnc+JeddzJg5Hv1WG5yMv5BXwqDvJkGIlsAMhjgjCtYHlZQ/XohTtEEMP
jHOuC4h7zacbfPQxABmeidg9P3UEc4Jbbjt0AO5kq4GkDLWXNgnhEOIxNAx+k/Kd
6yHNk4iTc8NFQI2xi0MurHtmLkMFlxv4+JqdjZnBcKEs8QWK8TT2+iLKZGhN9rnY
DzLjZYOk5CmKbvIeXciwq0Ivsaf0xxct7qXIObVcfO3lPh7LxPyXNDXwiV1mo0Xw
YEt2Oyh/yWDFVzE3mxGBIqmZXUkxsM3wH8ujvUL/6slPuxlEeAue1Z0EwNWWmwwF
qWUZPshhBB/55hYB059eh2MJAHzWXEuUWYYbM/Mxb0DhEqgvoqc79eb/uLG/DPbf
F7duP/b1J+8QV1Xl4k1a8VsU96/ajFY4H9CsXe5JX1Xm1kXLo2nvQ9JuQv0BSgkd
uagscTWSZ9PaWRyZnNNEu0IRuQvGcm2Ig+1BE4KOOoitU0SMWOHrBpaCHUlNFYxj
6fUdbQI+yLBcA9xISrBXEeLzoy4j+lMlAqvxQqdf6KhSTm8VRIT/aX/uvWWKeCHq
kpN3C0L1r45NP1BBM5i38xDBR8BLkfZ3Qk1o8l8q9Z9QR6aBkyptFT9suq0sQV7Q
gjUTeI1bDCT2wNCL4owjs9Jw5mi3Tql1daUxBZzrfL8D/6P4Xo/awWfFLNJfMX8T
4XwAl7VWhfpbZmZ6HNnZFEjjSdxULHxWAr/qY+Ah4uV41M/+YJTKvXPjUptEX0Fj
6QJA0GzGwhMCNmN2AlvosQwq2ZdK9Ekh99t26aU9U3XgO6RdYIQTTrrDiPM4rTZj
clEV5Kx5T5xuBU+Ok3A4+gXCxvVqldu3SWMmiKLAtvsNuUGNHpCFLKZFM8HIgzgr
eSLxtKeIMCAZrXJl4+RSVzHaKN/GQnS+cMSHoSfHpxPtE0hcg1p4rr8uLSERE1TJ
J3ITP32sCPbGgzLw18aRLZ37TQjBXTvq2sHxrMc0l4e3eJ4ahXBxj95LeZT35nel
9bNrxlk++7I6BMP7bBj8pujpW97ZdB1zi6jJjP7CWtQPNJcK9U2h29BkE/qteYK+
3TxrQZV+4L8/HMvTarjo75g4W+jX646Qw/IullJHCbDuFlLMmEalos+Xd/ibemZK
jdPd56f0p4yuQH9+WGvHZ4r3x2I/R3hfhQrjEk3xKf8NskRTjX09/YmdE+ZTtXmK
7TLGgdjgetmfcDNpMKu91VeWt6E5bdd9oUk6mJWQpJi7gLxd93++NSNvLbHa+HkM
1XVP50Lj4bMzRyxARgLq4pdC6+ph7uIPk7LSHxX5I8j9iboPlf3TlDz+4n3fvhxh
Wqm9b9IJhHp5CLdQOBi1wIr15SRHA/YpVwicPyX8y35qeSDwPVCUH5ldNwjyN75E
fWvSO1QyE5tbseFiEM7ZjDKTHxCUmqp92Z85c+Dif28dKPCwm5UmB8UDY1yPWH92
GYL6AGgJ7/634M60ur8863vuHa/wROKXPmaGflJe/j7mZr0wcqSJKZ9SOb/SJVL4
AgbzqRm2aanWwQHBFwRxN3HWoIqTiHUVGMzKHJ2WeazdJxokhWh0qQViFXuHtFXj
y1ewbEpMYAOS/vqHv3PWB2ICXgqLjCd+A9ufBymStF71kTN9zZlpMKAySDmbGfbu
05TF5EUc1+XbI80+mutD9/5EFTimOOVRZu3nKB6+UcQ73hMJIjQaqr2HKS+X0pU1
z5NIFWCtK0YQ/nE0g7gqRxo45/kWcUFCvBVi1L/N4p5b7IkaV1oZpcBcNP/CvmB6
+Wo+nomcHgIOAYdOnXjDZ7ty5eLngE5GZke+9m9or/1ZPnA43zoHptrg8PvMVArg
0dVQWYc6K7fhndpwYPZ/LYrd/IurZGmBqmUmPoLRpixS75euJOd7cgyda2taje9q
ASMt0wTIZEpnJ1nlTDtcTC/pXQVX9prRAV/c5tlAe92WutJsFaDeZ87Ges4SV3Ss
VPFHyNwXIjADJLTuV3uuq0XzstbBZo99q8zZvXdETMlfb2y5Ot+ywHoDUEjtBrP1
cXsastxVv92vO5Y/0N7CmsIVXNBS6bk1p1mh+y3LgYjLu1NqMnOGLL+29rMZR+X5
JGx3hx+U9CGrEPUADhhxBhRai8bqvv6siQtrxftKUfgcpp4zbfnoA1D6aam+aiF9
nhzuFslcQd+Oyt6/7zhvV1/6ZCPeFiwpNTBjYG3ukZ0OKQKGkXw/9tI15TaPlV++
M7CC51H0xjc3EagsL5hHsqi6qY/4iIW1b2GDbKBVylwSvOA11YJZsnF6q6rfsJb0
En+Ir2A4vhGayknjfwjbXYOVeU79dWIer5Fp4tErwufO7u+Rh9efPsAyVeByGkuP
lc8H0wVKx4nUgtvrq+7oL/EOHzqpzC7RRZEdDzbPKUNIa5srxRohRtOZtPT0CcWQ
xHHqPUUUil8qQpUDeowv4VDeK3Km72MZrLki6VQE4JGvYM9Qp/n7HLj4OMzvkZv2
MTS+Lr/KSueqpjKs4qFmRb0RWO6zniC0v0nSw+UoF3BQd+l29dXKAcj0VsmwAXKF
AFyY8lgWXixkXudywAFgTVcrxFfT7hB5Vs4Rz5z28sjbjC/NWI8+avCTPlN84e5W
AindS1nW+6v6QD91crrGxCghvFX4jGIg9vT2+mRXnVSHMLkhBQ+i0en8UShuEny9
3z/DzgDWcix1Nr2ihNJ8ow62JPYh1ORbOsJ+HXWCiv5UuhWR1jZhI9Wqam5aIrdg
wasvImQMWpo2Fp9jyGXVevgcuwl2bXoZx8drNpDVl9Fq7NvA6K4ph4TzUp1YwKJo
HRMVRJf1JppLwtLWdjKO5jDdRKnUNl3vQ7G03VDMQ9odHVN342XA/CvbPTG6iBT1
rOFxGDfd83rJIyTt5grnMf2WNSrY92lkgnGKAkuXwhkndoPtZc7vDoKQckLp3Xch
KcauuiIoxvRupR7LBkAbx0EPFjoUc6EOydJaJHdgTOcsgJPwwHYOb5mLdyRP4wNy
9zY21NgYvBAIf4VN/2XFORIhDjBoswxTufRm95fJqCLPV4lUdnm5O8s1Mn85j2oo
xQDGsBOep+tzD864vIvmeAFXcBJskYva5BH+A8uTk6qO/wE7yIGG3T3J9O+LBYpe
vWB8ym8WWApmMAoDoKcmzIHXu/l6S3KW904Qzdo7F7EARASyMWT+nbsbFyBPhaCT
n2r8+UOrSHvtJ6ha5yFL5W0uzjSMfbTFMHVMhf89yJ1EB3N+/+FWW52c5LXGMBfz
FlQrLXonwnzQXdynxUQRR40Nwfuj2j1UtJBvxeW5Bal2PklQwZzk2FEeh1tYw+tu
MJSwBNaFA3M5TfwqyK5CQDRMahsAr3RVWr3cENdMxiC2P0HDa7+ZkTieQFbBw5/J
RzmpZXxib0df2INrUiiqXH1QYoMNpvDgDUURrWDkq+h0iL2N1ou1wfOF1U5sAzJg
azfHXKWHhnRO3DUGxfjiqW233PIucD3Y46ck110HMhZ21rYM9uI9B2lEDEyZQBGT
YEbicoOqoIxrq15rjuMJKY4EXqWSxTPWnH7PSXASpOc179MYMUyvQCpvWsFplstj
5Cg3T1biHMcZ237H+7h45NvWoEEuNszJ9b4VZRyRAHyfszR8q0u0PkFEwwxn5dE0
3BxPvtl5fv5ZAm7cdMo52Aq/knzr9zqKVrOr9HKYlZYpZB62AYVU2c4uVn+sZyZd
WQRuAmr6TafRMddKwLyvUabC2Iu+f7YunHik5nXtYFWI1A0Cbcsu64F4jxhpyR9U
MWu4JNjFfuOi/wrzQTAGCkVoqC8HqEr2esW7v90WEVDPWrsTl1T2Em8KUWqP/0ms
7k8vRW5Ezc/CfyZ8dmDcOuhf7YQmeqPCH6e6/LVODMS8EOxfc7YXz3ZqkzUfWVB+
QRTX3r6TCVM5Ik0ouizcy/egsgG9rWKI+YODMD4uwIjFMrRsAWmToYSuUYt1HZV2
RLdCPPWEZLVoVWdhdozY1TUb9rc+ObjzhvkmuX1cpY19XHsN9LcyvDdNHBDFeNYc
Qek1VlyUPyfFT6WHWVIKRw4PtMBP3AtGV8qunN9aVMj66I2omLRk0M1kyI8VyMqk
SnUJXDUwy4JhbcUJBSHoypDzj+sPg+wUaX3zS9aH2jPLrJI7u/k+CIgjMyZnLHWh
j8DgFgA6FJzLIpJkbk1kyFtUxXAJG6Zo0ch2r14PzvWfvsdwODqFDWqlKQT0Evd/
aYWtWdpKmM9T1JDMHAqZjPFMy1Anz+s3Rv0FGKhggBfAzg92RQWdM4SjZCOniC+v
mtJHgghx4NY3+mKyp7WnBtKJRNv3NVYeMI2Qbn9e9vfYwuIKzDw6M1WA+H9Z1HtG
3BIwaXdm33s8DvIzZGLCJTLAWNOXSuPb6wEhVmVLg//c0lAR+RwaHiiAgtZpUE2b
CzpiHztv2W2iPG8M8FI/+ObSMCa1PjzQ/dK0t2oCQNeqVEb8Y3HZ0MbHocip0tBJ
f03FaeJOI+g1dwbjiLjo/Bf/AtpEnkZ9GeQC/aR+5hdCMlhaTComsCBk6TDENkoS
eWkaeTcuh0xvzlnAl/D36YfAX5Yj1YfTqEDva3h1s/mCVxZcz8bp+TYZYO58n99+
eP8MmLrFwWczDBzqfvZ16I63XkNFWvuTLQIuA23oPmbPqgF5PA/qj6vrMBjNcwzb
Wh0QsjKXae+oX2AcRMr/n3E+AQkwgWoWt0heJk8A/rcv9KTTXt+4AQBBN4/RE8If
MdKbnZo4kgz16RE69h8SEBEbRe0qSAkCa80Ra1fQhV8FpguWxU1GY48w3ofbhrc5
ICPCcm0vXCvwreSwya7mZz0BIhE2k10xxxQGf3N+ZcknnRa9WCA6lu6C8IOn9CnO
WM4Fkgq6U6OWPEhU0Ad8DvtB6guTtLqzLFhzoEqAjehf/94o6BrtVt9KtpnlL7Xy
yuCIgqZnNjsm35sbkWSXcInH01gF4T9B7CXATpjlK06kVCZDswt4r1uIA6La61cv
VdanuMMVa5D16IHSvnPnrVLMvQmifq7ttVVFihugHwF9wao5Y8CVHSL3qfb0/Ta+
RhO2UBUMzJ77xN1UngtJbY8kZ33NCyDzOZt/stTO54q0hNKFdAjDEZBDmLeoemj2
+ETOnKj583IQJFbFbEhmzghVgG04n3knIv9SW5R7VSc/H6otCIXf2iUOr6Nx1W6v
7DSiDlocltYdTw5vI7oOL1NsskZ+vvSUF2WgOPyRrcDDTCZk8m4XcviqsaF9M+BQ
cPYiO2aNusN+29/R6NeSkto2CiK0KyUKtGoNFsVilR79GRGStKv9eGQEe7tWhqjj
aLOAaZBczRpzhrM3Hr55xvpe9w1KRrDi4MyGV/iexnGKts3seMjKTbDitXz1HQbL
HckGZcrsEnzaYomtk/5HHowHF6SvGujSIH6YOd4ZoXdEhTtVHa0Sx2dyZsu2P5OR
bmg8HilzyQTmyVtL86yqQ3XYPPUHtUwTUFdhzx8VabKZKiWoGTmaDXA0JxGEK7Ch
YSij1dWr2fCHLX5oQjQW7gbDKMUUqPaeGX1cYEdekMR38rJ88lsUQQl2F/5l+Tn7
7hRZ/xdaEMdZs23NhFs/zSNGlM/rCbFNhjF0e7GiWsNfvdUl5hwcpaiftYnkpDzo
XED7lF8ILoeAWIX3xHBvUkGq846w9R7cLEiHtqSUtcbyjHIWoX1vrOun9vqaMuFR
rgeB6gH9LA1sUmLPHGkaGKgfTr/JqGvCwTHhOR+sg9DYdCpx0v5RBD4v1xXG6U83
sJMPT7pjJg7ifWnZRU2OTDlggdMvFOrznMJmqEl4hzrrBMAL1HiJmu6V3r7pSvrh
LQRCNqmFoJkuigxlVU/+0MsOhzJBLXXw1J8OyyMsvDpRSD+MBkZ2kln6aFVu/cnE
dSqDW728qU3+MwMxcOMCuQVh/Vz9qbDqurdc3TKdbnwwIaeTjse7Em9DCiJe2eWu
U/WnQ0tjwr6lymlmw/4uEeBn3G+AkpEDr7BsaT38mlyRY3DgAaYjdmhsKan7SEis
Y1JvlPMZ9UPNTTvA2Qa1Qib3PDcBxhAuva1InBhQFAjtOfBU5UnnsTKe8lSSB31U
5vlIXiTfZPNnLoaieDL4v5dOnP2H0YqjOQd+sdKLi451Soj8slmVEURT5v1QMVnw
UpKNkrYTG85XtZhtGeJpVE1jLz41pblzWGqg6C0f8ijildn0pzxI7XCKNku2K7vs
NRgsReahfjRGwqP4DcBt1hjxc2VGATjzNHEL072f0v116F3UozDm/UVUzoZGag2d
+ApNGEG9i1rZfH4UxvdVNAx3sEHW14RO7KtifsG0/cECjAUMPmKBcB+a6gOuvdWH
WAt7A8dPBqiDNzRFjDVGXjObCyShjIHRqmUBo7OdbJF82Xk9Nt3kMZ2DQtxB8r/v
0XAzrR+jinKuZd8zArY3bZn6ZEPz7RHzphPqhiCWB7xm4rJaYTg+3+/h2I0svVpH
/Mskue3OX+8MoMjoXNLn0vyf4gYH/QghRkq0fPusfDOkKVLixLDEyZ2JPyZk+Fp3
49sU+jL5afbwA9BKCLsK4Yc4oKEiBg03HXuEs24VUcXynNtbwrL+2bYThmkaerA5
ru+xBphndExwAN+gNr0G+z8/licC3Iu4ZWSPW+akrcUAcoJTmuRAPEqPdtgTDkOc
5LaKrVeIwHgf8qW9xEYa81dTE6THyVf5p3HnrvaV7KuhbdOflnApXKJ2KxUIARZ3
5zQrMimxzjTCmipbGyCQxilveh25XCu72ALniQZwJU2kpXvipJafpMurViy7tEPf
pU4+ttDDAc4LziiFNbg4fn1FpHaeqEwRQU++NImtsKGZY19f4sauxFXipHmYNDm+
xQ0Hr8beAoBeKc+nkad+0HGSuEG4zSvUEa/Zw6rRP6AowNcqnf+mmzMSn7sqeeXS
DkFEk/NKdtcDuLyxz5GuiRDlHeEudfr81Utg/OIKLt7+9M6JkeD+AOJMcVcQjEc0
0X7L/OApwit8AeIx/b19tjbtyg5sQxOusDGr2u0AvceKhJkKe6/6M0cWN9MMIJdL
fyHb0s+FLbHc+Fh1cjrm0lQJxGBRunFB/bck7xId9aop3SBGQJmug2kBG2CNsPfB
barsNhroRqEzV+u7jUPaaYef6L0p2GFGxr/xwELT9bHJuqMhepEdtkiwEvOY2d54
1jcAAzfhO9Pu7KU6F+vGVaBL6fKzqFirooo7biVjsStdNAGWRCemoqJNwR6vz8Dk
7vnKwXes5QrrC9DF4VxWs82z9uKuMbq/6/qtKlPv897hO6oZx0JwxDNh+fX5w1ZO
HPUlrj+XnLAB+VZfWW7eRkBdoSmaYt8uUhgFVDtfuor7fVk1H6OwZ/XDekhzAPrW
2Krw0di14TLF6MkoinHz9ZgfeloATwEg/EbRm8exQx8lxBp8ME0RybHxp2K87xaG
euvz987cQ/M+1BqMaeE0Draagdxe9YGXZ8pSkBaE8cBs8LFIxijjslZi0skew6tn
xfAInU5+RLulHqPgnJR5CCi47HviN77/oTUOnTZzXPpSaK9MAvFd1hBb4RWlX1uO
fIk/V592L5PKXzhQsbaVIhOoWF121zgcD/Cfo1WkRVJ5qxkOpp7fOWF4av0pMC6B
c5gQ2oGHvoSMsbp4zmkT6Ja7BkOze/gaBsa1BIYoqNAHCsyy+K8Gp0m1msiSB8U/
Z9L14sykggRx6vxr9VNIsiU9/gYUd8IbB93wy9WWEw2Y63UzAXlxD1xCVDRex5j4
HCaeyHG5bTchhnRgHMUmsv94+/GbU6YY3xde7Uo7BrMLKP0Psb/GXU+lB5aSNhtn
OhsyjiQTb3SAhssKfa+z9IUPbrzQ5KefUhGxwWbOfE3zn8oKsXrNCmyvYovdmjCK
6l9zARxiLUmTWdRcIJjtDtuT3dEtyhR7tjpJR7g0dgrQDThVMV4HMNznV/RfbPSy
1cPwS4SeiBaJ5o+y7OEsLf4gR9CSbL/SV2b3YqNBQV548zYj4ADu4xYGhdSYszAV
n22+tT/sNrPUssNdA+SEPwmYyVixaEXCpOW98ZmmuAznEdksZoFPTXgqHkNgcO2T
Dt8EyIawzYqm8JlWUK0yHXlH4gzdZZZUUrHSx7uJ4P8b/Xmj7vFfs13HqwB3gJGX
WHOAvuud9tMekqZY9VEFfL9Ff4LgkjVJJ/tc1APg+BRwRESqd/QNM/MNoSN5VV97
Pmp6zzYvrXSWjh7bTSf29K7gcaHTEQO9jqWpYxNDQtMR/UNHQAvtb8ek6TOOn67x
5My0sUAZXWur/q++LXBlRiYzIgh5SKwXOc+n3D7UySayBfEPPYnRcW1QzL91MGtF
eXx+HIGuK6WfIHGZUqG4ykA0nieRilY5ZtQMfICYnO25nqSNAHty6TzSqqjGLZKh
YtMzHO7LFproOXmfLbChxtH8+Kqhf+DlstPlXCJ0g+bmIwi92zNlM9iLWbWovXRw
3F4AO6qx0jeFnmeJVFm5gbv0w9Bxhm+DNORHSW/WWys0fa06aRqZAmH3eweOqh98
zjqG99B746lpxidmQz5NZlGaV4gM9bemEDDCOYEpWSCMZSurfrtoE3c6GLoEqkUZ
Nh/whF9T+kLbnYF5KxFbFXpBLaYWMepwf4yfVSLsmejn1IG0tiCBQlWNlFaD1Mek
D3JP0rnds+RnwsAnY/2ivEUyfJGK2f2C2nRxdEoNukNLtHfn0sF69qwISYa493jh
Dan1vTluqJp8p8FJM2TB7Ll//t0f99962JOCFqZsP3oWtF38bYZbumaaxYcgRIOL
3qfG9ceCbZHyn3acXBe053N9Ylz+gRggZmv3CFLAjVvlttuJHC0ivjIClwRPhEfc
8zCiTi9pwcMvUrRiizJdSla+QboQDd/ACp2JNAbsKzsl1L9Hx/v0q4pyA3eXb2C0
azpau9cXu2/TPFEBRnx6p5oMAmoGzCFpOkI6QVtbVtFH0AzORYAKrNIK9VxFpO9P
HxNvm4QSyfLUCcw7l2VNqLHaO6ALAKloaLTPsx+Xx+KGsxWmLfE7g5nXUaEBKnpW
Vh0iDPY7Vpcr2nL6dCWVNx7tOLGVeMCx2GLWXXE/EtVUByjpNQ3s8FRbznUYW6sk
V4wWcfdE6woJXW/Ij/SnowLJf8eW+z3xhZ6Zd8YSVi39Th4n4nH9gEnfkUltHj5B
FMLk9eYOgYCEE2ekN7aSb+5TaxS6kBjtDDDN/v9XGV5uRmDfz6p+hmAxpbEiPixW
A94VNj/uK0DIpYFnybHZnhSQKIfO1+CtnpMmmTBDrUP3BJzB1nFa98EMp0bMkEsf
/sELfpEA6A7pXfZ5hlqLgLRsJU2+bYYg+S9e6RwNObrRy5lVSiXB3kTPRJcjj9oF
hwOxN+KIYnyqko2GfJ+EHWznhx0XVSQLiaE/6/N8jDQd4NAIBYs8z4/DiLGED70w
pPij9Gq0hkiPnRcsOTPR5Ysa3oMrtCgchF2ZOi7R7WFbFdpDkghci0t5rQX/XYtp
BNbbeRRYQlOcb5ZNp5lIzj+EYIdinHqL3y/ICkMMohGtzQGb+KjCfohcJxKOuHZQ
DCwgDfIRYX7f4R75aoDXt56YQBxSyp7gwXqtcYnBmKrcLNErxShCcSdHd5e721GY
jer+prKk/NBmf71kFNg1heaR/xpG98gAvygyOuCP/OuVWP9yFPhAZoJV6Uj0JIQL
GOJLkOOGNqvU+a3aYE1Hwk2teeURVe0mM1/hPtAOuvvXn/G4y9sSpuH50A7B/b+S
Wsf5qoxieZJvEidVipfMWAQcSfLVLZNXn0Mr1tJwPWNvymLWox87iKWOL4NLZo4m
prB6pAnjbHyxB/s96F2uxRUaaoEIlA4xr8lP1dQaCRbXTqUPLL9UzEsyPpC7iYZy
ggXIEVeYUjAV5Ht0LymZMaI7Z5aEEcogTleuY6HdpZ3vDtYS1YPUVhHFH/blIQcO
ZmEvBbc+KwFTPdn8d+KRaLOOx3j/OJe0VPaJIUsgNB3xaBa0hCdISqFf4KWS1mOe
Xb1cdF5NwjOkCf87/OyDnnOXOAFSXSRluwzWAxd8vWGlYfVo2qSpkrRPhc5QeyW8
C9tJmw2687KE5BrZ/HvLgjDg9FSVc2fsG4z/jvNTo9zJT7lrOBBGk4voewfAiy28
b5BtnpRH1a27o43KrVhKywBJMYIdfbjOdsUmud4j4Wf6aE5Ph1FoEAtik/fmodWQ
ixZZVacfTs4qEfI0YGX0Ieh6ssmFNbRJLRzAwyeZTeCE0Csdmrxm7P8k0TSabpgo
Y4GsRzHVaR29nzmO6G7I8vrFXhrI88bx3rBsPby0FDOWz3i8OaWd1RTLpw9P7h0C
/yCyxsypZ8OURlfURRJpPHI8d4ixQALBSEf87uPlGOBq1BNpTftu+JwClF30S/eh
+msQGb43P486MNxaZi58Ro6w202Rp6o7UpYpoy+uGGIx0tTx3qRnwpVfOhijQ785
NZEtj6Z0jDsWPw+MrR67vhBG3NpUwTOyvRyiT1FJk1O9RJaooOmNOuXcjOhGPHY+
O5ALKydhbuQ8Svg/1OBnGZFRscLy/9s0wxUHPJjPTFsl2hnRLwX/I/jNx7HJ32KB
rGu41x95lKxe9QeKBeR7jVkVc74sXalQnX2DdKbDBsEEEvdlyyK2WJkYee/uLJZ/
gkRPW1mjNgxxhqvMQukMB+lanmVUtUhU3E4PxulCwW+xN0mD680LR3V5B+DUEybr
2/WRknVt0bk4sZF4IKASlYTw6v8T8v2zulR59VI2jsYu3VZiGSN4n/gKBUsE20UA
sQL9MVd+hhTBbFq0n3VRnelR5vpS4UQHVuxZQsd4NbTeXK1CfLYKFGxLw/8o23md
VDMVjNPPQH8kJCQLZnHYCCICAd+pfbT9ndPRJPmExlg5YMAG/LbGACs+yNmmeLrz
bpFt9aJk8W91WESqZRH8qSjZBSzYf1PaOImkfhcdsPxMRvYTYY+ZlZUrdR84JFEJ
1enE+0cWX50q1sXe0Wg4a4ClL0mFW6uSM05TmB2tShtaZE2vjJNGqg7w29CyW37u
4TcvcAr+qvkI6bcD5Tl6axj/60LJyLA0N0uVQfOJeV+RUC+psiWpX3hGQg0pfyB3
2egRls4YFpzN1uPfonlXXcVe+wgWfS6J1KxNUMsxg7IoAk9umB5Mjm4JyZ2neBxD
RXlwPVwhcQM8iFNlD3NuKDxfcpsS5+MPu/H5XWF1xM8PS6kw1pF7TJdi9DMcR7eL
fONy78itM4phFiwonnkQ2jCESzzNeK3J2towwEDJA95aEb2y+SXy6CF/R43YL3bO
z/mkxcrkKnESTwJKGx7EMjT1OP/snvmsyXprHAk2bScOKxImyQUOzM3e904Oy1ge
aCyjeT2xNr0JVH9yZEaF0+Ned/1ZkmvjUoqSFffr9NCAiKk5LyFcisTU77J9OVmf
lcU/yeDLaSgF4dfmEeBdHfSaXdVUHmRqMRXXlXZNutjeVq+pylkCCpe/EHRVExQD
O4MTCi2eCxHDPdMDDZtxCTCqiKlRLiKIufa9v5ATem9GXwA3tM+PMoAsuQ7k+ojE
EQATbW7ylNa8y2ZesrqtYLDcyDEedx6XoLGtHgxKvzrZ4Lc7oUUETru7TshNmv1k
/tb3rqmI45UHbSf7/NqR64bNsr7/AetD3gGjFvKSAKZHZ5lHRnM0OIB0OfvRMa/w
NhqgsInUclOa68pXBDkPPCOmOdtedF2FmdHaiOQ9myto90gylAslf/LH1NOq2XeS
RWui9P/rIhlBbQsfQLwY0XnZryV+IFxdnrAtlrlU4thNZaX/iNWLyeU0qtosAS1e
YUKU7dOwgHnj8F6PJJaABIsVXK0KgjotfpdqhPi/iSs9o3qbxuZRFgNecni0Z9mB
aWy4oKJLZxKmJv7KoMHutmZOHYdbIQEvCENnJWjeQ8kd0LW8tsfcI1Vtt1NJOKPx
imYSYaKojINjT7hJvHvnC9ruQSB9NtNUT/AYO9tLJ4TWEWkCS6gavk490sY5w92z
yplio9VvXe1EmS+ZxMpH8m94S+X00VrhlpmYZh7yG0ywOeDVmOuuSbx4j/vp8JuK
YfPKkHcWP7+U3E6WR4Y3s/MAt8XW8/payYHOR+mzVXSgGh8SZ2IgAqxB5nPwGp8L
9xRiLwXd2hguKuXwiMWW4zW2jS+HZnKPkiizTofmJi3ddqH/aSAQeyIZvEr0hdct
E2/LmNTR9ZeDane47qlHxKBgTtN6LXaVQ57MAvHZS7CTpDvcviQxXCR3txa72sVW
Zp/CylnVykQlqE+SmAtX0l0CGeeaIWNb4v3M/3j11R1T+gGuep4C5x7bi1BleUt1
3U5dPQuad5WEeHQottaPCb9MK7JKegEs63x/al/J4FVO4kYkGLadyw1MchlHjpNG
cP/ZjPHlllSidrgBGHJGWBgVz0iNAUaPQIqLD896iY8/c8Aji9oWh4CZMpms3jhR
op+NeTu3juZNIrFtwOPOEbLRG64M438qDe9s2Rn/p28Z+cOaxH3czsLyRmhuAb8u
FcTsGDALyJKuZd3kh6gL3WEuwCz6KAO1qUVbNuQmf6gDLxRfcgQZc1aaD/PIU0/N
KEnYQRkjciZKzIVY342JLn/CU/rJTdcr7CzWUUTn0xupp3WUWiDhE/QBcCtNbjKQ
RPe3uXnH7Tjtx1A0FqIuUFa103/ozoBRMdZ3Ec8lxyaqVo9hs094ozp8QvhtM1MS
i1vulweTSQlrHtow3U3lfH//8FlFyP/mS+pd26+Z0mpqMuNinstl1FUc8kdVgYDF
r5sZrLeTBvM6fo7AJMpnRgSmQfYjGQ6FkIJfS0Jm6P3X9biF71V823JkKfu73btI
IUDW05ZdpPw0Ytg1kUQHFj6NJ/rVFRDO80kndUOtcMyVnGVawKFfSsJNidhd351U
gsokSHsjOZsLaJnuguuWz4kC1Qdb/F969OrcPViDFlX0sxfjA36cmRTJ8/tPQFhP
i9iQS41ZI1WpqYYd28MsKFBJ8Rr6bOlf0nBVysZceABzHRcO6fA0/i/KLg5cXM6d
MC2lJjIQXlKAmIKKYrMZbwWDoeLAhbMxJyepvj190GbcYb9XZtCtZHSBIZ/OAqFL
rFdUqSV5q5j47hhc11qFX1deYU7eoxnn5HS/o3A/Gt/ox7PEJmsMwsCrHD3Mwtcs
KjhtsLgZGBj/2GM5TMo6ErYJaOQunHYbrSVzdZlzcCKIjhbRsqi0cRW8yJF+yGAV
S2s8fGclRb7ZXPIptbrVEw6zE4XCnWepPxFw4bXZVdOTwEcbKYJUywIxJCm/lTNX
MFV25lAL4hikqS6kpBN7o2TZzJFR77iJTpf2vf5GgtC9Y4fvUk3tCN/En46Oh6R3
hcIXibYIMQOd4CBNTgFTVQ8ft2Z0mysf2Adzi8rXyjyrEh25Tdwmk/gUX5ydCPbQ
eCqKz5G6ywPUnWJh4ouB/9oo8x6IAsOvuXjqmZPD6kxV233aeKIagOPZNzDLkz9y
y9VD72pBjWAqjNAVTBJfptuj1nc/SDpQwOSmWeelWvChhpIMSZ/HZnPBGnPNu7v0
S76P1VTLJPdqlwE296QJe8UkMkiF6OXHCoFNk8CDW47IOpNJexGENCjeWrMWvVMo
xs+QAhTgeGDR9eCeBeQG2927PH8BRruHKpkZDkVlfZ0GSyLxexcEQYmMYl3VtVqq
U4X6d6RjR3T1Qk+k34V1hh1XbjLV+H6rjrWQTGrU1eaRZQKvcXPcbZnu+iEKY6El
jh0H4eze6/Ma3DXSzS1+0VKcTRdj8nmRDUBDwpp5yqLf+ujQWYiSf7ErUpNAsy81
Jzppys23ktCnMJdizVOW6boxUxo2N1643WtA/JZdKrysGVj1XEDjx1Zdh3A5v/b+
1LGoc8aQlEp+idPC31dHPqRAjHSXsPw2VLGqAJYaGq5HfDehPIf5b8EKkdrbF5Dm
mzu/ayKgjPGScJnQsiK5LiyZWbeatcCL1Aw1OX/t19SkWxssVVQMBKSbjWVQcPK9
Kmgg7b3RJtYmu9+8UZiZCHvSONvsQ0OvEzq9yyRjHXXSy7XTtr5A0a3GxmE7GA+z
NmK3c0O4vyjW6gE6h7RWV5BtKj3NtLXHwmclRC95tvQ6IPFZmq5jEqpyOMYA5Vn7
RFi5hENV1nWLnqKUQi6VYsnTV29Wvmzo13tE02DU9oKdmZtB6glQeJUMknAB5pOB
I8eetBTVZoVK5r+TAOhZJvqaPQR29c1WTgNDVBsCuPrt3WE7Rwa2JhBYEhVWE2i2
Co3wZyT1rk04W716QOb6xypGtQVu48/4wqtihAYvZKmbb1R3u8OEfhOaRDKcSfbx
0MdhFx3/6kYYDP7PGzIcDYldhOPuGjWmTBCQTpcHWdaRn1+pQ+vW52Z/GF3+HnT2
Gjg7DxU5mQT1wNd981SJE0bpPP7exE+1qjkaAiWZKPiVgiBLzH0VHQW9iaG9RaEr
bL/7Z9vdvV8C0FtepfyB0hJh+VIbG7QUVqP9u09zI6AD9g1tDWNL9ixG+QYPe7oE
RXrottqCNFi0ly1mVGUdu+kxH2KS2esNcN77TOThPqefUfWRRR2q5KM+z4M8rqmS
9Luu86eWPkFaoAWWp4q5b4NQjGHVEnpBEADnco/yP2+9cAr6CWuNKs0XuXoAXojY
0+a4eIwnL8M4ri1yVCMRvWnPnCCcrRhWvjtC7YMC7nXumW7SmORYdzqBjVI3FXcq
Wfi5386WXHqJKiotMP4j0eWokPO9xrwi74ZILMQV59YiDMo16e6dby1iYvtBrlif
XrRHcaAfDPRda9R8c87NLHriimU7dOI2nnBnlL/Yh12+nYCsy6+aw9t51GX07Rhf
zjSZU0zphnhjZ7hGh/RUbGPXqWSu8icWFZkhPJAdrf1PH96ca3xFA3f8YK7KJEIj
iFtSAelHKxzcQO0rcspNVA2tOWzTyMrdbsByFntyqFhdTgLstgzlMoEB+cpwVMYC
cJqDr8g3HIr67y5CsFNSR9bv4xMnjq6dSJYcS0UsPemvJ45Y2YE6qlT+aTShdt4P
SjysHAYa+cNivd9X126FFHUUWIidAhbdpapYN2xB5ySaK+XkrOdpanjqZnFaaZmj
Q/X0b4lmq2+Xtpt36E5ZUwHz8C/wG1Bi7d8K7DoeRFiaP2tBBnKrkQ9WT+DI/oTL
kk4fabRBVvZwB8Aq8JsCIdmWKzdX5n/CRS5EiEFxtCYyKPf6aVEZqPQqlggvHzTA
yZaXH4TJ93OiGUIez1MuGEidI9kPC5XRMa8dfWIlfnLSSWCWOwk4uy2hziLKg6yM
SQ63REBfEY5pPf+pilTT4hg0a5GPfXbmiCHkIK+WfSEn02SPqCkuxOTWSBrwUHzv
DKUteP0t7pPJ+T2SBDcNq/EemufZTyvhM2oSEyZRgsxnSc2kb/BebgUTencfqBow
GBwb54EDfha2+zgPVE2+fEC2zTwsQKbISvHKHX9MADV4TJThNCLv/QRm28HKxsC2
eeboC4D86622FQt7Oiu9VE4p5h341pWPmxZHm/61Dc9JuC0ehFj7k8Ijzc6P1r85
8aThCdB6+aQ9s9fgptRCcGhXAiYDmNu0WvHa6mNZ0LWrupEZ4TmBz1359ADJxcFi
pxaQp3XiUfQIbdXCHgTGxOHS1JmZy5sT2Uyc5+YUKaKfoVV3eZzzmCsog8luzSXr
kU2SeX/4Wr7iM9gwXsUKxX/IFTN0iowPRyXoRKmXksFYLHK/NWnwB5AZzvIlrM5M
7U/JAbz44DIXjT9lOrBHxIGUPL+L84cS+l3HdGKc9AmaeJlvz4Q+/N16MI6doAeJ
Q6T/Xb8b1ko43jHgDqUs4prlpf8BsDFT+QwEYxw2h7ng1xz18/UC5wdvB9vs8R94
qDftmR6BFyt+2hhBsKDkgMtfml7oUE1ggvkZAqH4430LaEKtpTC5GoanxAoNGxkK
qGg1T6VPTzMpCC93b/0n8zsdKORCNUSl12PEexUzqZfKJcg8DWNkIjOXqlhHRtVT
v+fqqIUUwSs+lTHKfhmTT7UtLF7aoOvdQ+9L78yY+mv+EdtLdbCqh5HAMiIMPFBU
ijmq7sdsK6y0rTkIUX+xO4XhfReCw+wypXigZFRmCzy8QtW0TVcrl4xDooId8dBN
5K2zV9Z0ymKpVlAjb5h7a8HlWngt7YSyUxcuzHxbvEGR4P16aC7IebuergItYDUl
Jo7q/zF1iqW21qd788kUath+WaJP2bqLE2PZ/oGekZHTvDtG72LZxh2lY+xgzy2i
zr2FnfQHJHWBwRLlUhOILvCGdamJShhkKoQN9bb6flVd4F8ngWmAkjOOag7MrcDy
a7ILKSqxFBDPWh+zxvdF3J7nSWKIKCn8c0ZiHI7btH0DkzYrA+4qBqk6j3Uvi0v+
RKrmD9DRWiMb7JFuMIovkK8vTv7+RvTlo0KbOJJQOs7SO9nZRbJh3nOrwcu3itZ2
1X943qNAI4CZyxEcAm6ncKnrw5qRUiai5ij9RnxIc7f/Qq93Zxrfd/QTE2rW5FMY
HWtvXc6ULfNcUuPnFXly8X+RY2ule8FsGo80UILNIs1zoxUTtueiaTLWTzRr/OJQ
QSjAZmWkHF7sTFQuk0QIEHeVBWsgUzopJyokQr5X018cSzu+DlYVOFrr4Dob+l3j
LCREeHtRdNQMl9yw0YhkvbgQGsI4FIDCohclLzpvtKARK1d8L8cf4+zcdUpBFH2C
xAXqW6ymltZ5B77uDN9RwpViqMqqNA4Ca9Yjhd2W5joOjsEiQRCu7mE1blnf8FXD
GVaOt4pqo6TukF3iPEOZ7xalC6Wtiz9ShzHM9owzrQu2V7jpTUwMSURplgwKEXI/
cVJykSMfziR0hOJvv/rFpTwVZ854yWMatYRUU1q47hJMy2A6atnyW4WWSeHZ1aS3
KKxTG1gLbeJ3o2PTRdWegmjfwTsZjmPx3uuXQ9Qtru4Dt9tVCYg9aK8EqdD6Y5SC
la+hrkVSaXfp7/ZlNOT5n7W3eY6Zpuvk5V1b1Sre4E/SgGrFWyLHvq44c26r30Ey
5Zqz1UaggSySaSEgaVROCqgpJAslnlr6n6F7rs+OXIVXVssj7WiBlDkO7u6SZjbi
5yM4T1B5UstL5g4bMhAL6c3GYNccdeMPKG5ntiyDh/2vTQpUUZT0Qo59bPmqsA9c
cF1DMdTirows5AOfA411Lj067+fFAzjGlTyXGAcduzf9FJWIASxShe5dHSYC1HUG
4urCL/5J4f14rqwGO0NqHFD5qEKHxVMz1/ho0iIy3N2QfRxRilAUSRa6G+HWo4f+
lU0h7g7VJvtsKIVFfmelH+ECgSoZn0xZDBPNfhcDW9fpqjYHrRO07VNoiV8QEYCB
87zs794vm2u0fjHtzAdyFmZoSf6g3Ahxi76j4E7fQ3FYrDZ7Q9ch9q5Ui54owe5e
NmiTaerDgcxb71sHK18H/9ZyIjpkmCr7DmR//ReVXLUZSbMhUWig9UYvDfSvyikM
dXKcfWQr/4DY0h8tEiDLZeFn8Amcq29GmYLytI7CERgeYUzugTev3nJqsxi6+96d
jzfHseI/Nmv8dQjmkloB7joy+CwM1CqH2o+wInAfoNoUUN6Xlhf0BxNCbcn2GGew
ZxeDmULNKzMH83dO3OCwhiEoHZGW+4jjWKTvlp+7see+0cIDCPlSpwRFRWWYF7yl
lquugpJzKHCDdh47/MLgkAkyGgReXkRbyd/L4IbOxRn45d4sag8mAbO24YRhAhKX
OLbU+b+Ne4yGGpeQvOLyWJpplQTXnp3PwEXm0FH7osjKulAW+kOorP1gDyfZ4BvV
bBDbqSrPIwJveQWjYvFBb0dMawDQYKJpJCGEW6o6SRekkOWF5m2q54JfsvUxXJG9
EgkWO6zihsutWhMbqfxNBlNyOqKHwRIpZXpGagd9g8KRuuWPqfg7CHh/WNDBDY+O
Vea7slLBFJWmF41RDOsprYahV3I9DpGrGY7l5wm/nUBLpo+N/sCXwQJRYqyN+j0V
zyN9wYeddbuObl7ekO5yzMQriyCj+aC6+v02bmxjm379WyqgcvovoDxsJg1ujrWG
JIaZPTG/PvnLh/2capCiR1sdIcWxv5Sl/nB/WK5DbPJAOGLko8AQj/KPn9APdIVX
LgtGSCE7/F6/iIQOzGEdOO9ieZxR8LfMIPFFvisKhwSnvnFff+vGbNO8QSlE5n1x
fEf9b+vKKucSZMZ/qq7e+6TXS656FLwvHQVhJKp16/91YYauGDjQb84zs7YIZ6oH
Xn69IHsd2Rg8Cf18Zgs+dkQJpsEGgmRhPsFJCR4X5hPrLHT/e3GfKdVqw5maMwOS
2rP4qo0pdONGTKty3sIrsQjTBgp8tzdcigoI4dYBw46pnPDqO6MVI65NhOiTfBHW
3K/ECwomsA8+pF8Dllx35UDL7w8lqIAA7j8nQspxPaauKkvIx9GANBz/OqnEFG75
ZJ0dcHq71WUtou3d/8U7Nz1PRl4ce+4IWN8ZASc/WfF0TOxJZDFrp5634mnZ9e2m
ZP56DKDJ9Qb0c7h4Z4ID+fnjHfR+EGqWSJQ/8k6Y46pxVEr7jWz4JkoBEwJH2MzC
x0cOYcOw9FXnuQaVEOtiM3We+u8uCmyKMShOpzxTFT6G8TF0YURr5GPLMj9tbNVl
dQ8bvWvXvwG7zTfzcsKzxwZOQwNoDC2F+flo92KH1nXG8lceJOEM4zMWSNhjjKuH
ZYVTUXVSI5x5IJCWFSy288kQ7pss0GOzCbJz6bftLkSHVJ9qROmr6nn/glCfD3c7
U6CpJ6z6pQVbxQATtLXbL4IdGxhZUEm0Cy2h3ElbkhIkcTXLiCNE6VijRF5G+DO+
oNfSXFYCK6tc1dCuqvhJbklfBEFC0pEyHJSq8E3J6+zheQMyqTVRRVuk07D7d00e
yHz1/nflaJ/3wOb0jLX2kI9QztuHoROgoN4haFUri3zcPznwL4yMIDEM1rQ3VEto
6OwG/OAtX6CQu0eC8pDKRp9YzyMNN6AQJIClZyHEzJ+ePYLc4b/gE0pJqrngr1Bc
xtRBk9jart1uJRbTbxonQafOv8J4fSREXvkFmyblrvl1DV4Qq3khhKZy1ULj++jD
cUGIF+BywN9M48t8WsSGYdvhGQ0MIwSLwRhjne8aberDvkKnkiizsvY0Vn2Xc1l3
uLkLo32sGaHmykTcU7OcuZwXAhbty5L3LL50w4r7i26rQSn+obtv74P2Axl5NoKE
GNJcqF7p4JWTczCReQWVhGuOfPLUaMtXrRKSeFrKu/PBvAtxN0XsLwGCKcqWnNNZ
E35Cv3q9cfrtno1B/aeZfFLv1YwjIIp3YKurRhbfqTKFLPBTPT70uz/PvSqd6pi8
ECpZEFBYvhO1qHcA44puqaSgJn9iCPNSdeXkGpetsXQy4Fyx+65v2VjDFmNNlMtM
ogEbZmUxyuHpBFQfLMYvpep0KrzR39gg8XcZwChzepZgW3UTCiWjGeVAbE2fKzqR
SZIBTPqJ6Z1YrSRE9aEPXk+rtKvMPhkNKay6blviP5y7qouQmZMfXb3PMxt95DS2
mjRIPZxS3NACYjPc8X0rC5wkB3QUrftHLlCj9EnV6wYIIyDw3k8zDqBuKkgqhZGR
lQ3NpeB2R/DrLWCfT609IPq3ZuWIRrpFK4mdzDy28C3j/SskGe7TpizYAMkCOiNQ
CJQ/C1hkv/k23nqg+IBcveeFU8VnnQxkYqSlRHffmXa2Tz2nK9mlO8zxIWJdie3R
qtHiBpiCs61xuWbwwXlGlYQhIaXtHDqC/KcZSdgq1Pb5VmSRRBJOZgLjbcqBb0e+
UfTVLLrAQGibTCcQsgVZBNMLVfn3z7UDDZRR0nZQsoyvG0XPUXzZKajSwm7M+3SR
HBgTr0gTB/mux8fTYa539p7Lyeb+5M2ZsgEi/sri2udkZ2OGeWr7ro1kGnUmpn2i
m891kw5rDDzbKCI/JFQ+0DUP0AKF6dlVbuVqxk8FQtPpRUEoXGLrHgo4X6zHxW9x
arlaYE+0R4UpdFlp6krJemW4jnkB6JT/Qs7oIqEBtQUiKx1gsPrAHxiZJwZQ4kgm
2juJSQ9R6YukkRwvQFGAamow52owmczL/saCsdQi/2PNBI5ssW6Y6YseFNpmgvg0
Q++EC1xCIbL+pNnnae3sdYkv75BNswGblvzltlo77xZzd/IngSCwDch+xC2fx/xA
I8+a3C2qBCo4WmHwi0zmra67VFhNqW9zWYnvld3uJcSsR+Fq0xkUPV4FdgUF4VEI
42B1+P4jPCpG46Q83W1yqxwLvPh3a7MJb8r/54pI6YDuDxdOsX3fhUH712HkedTx
O3Za7j7VklY0cGQl7bl7dSqxEztUetnAiLZcm2D9Qkw5j9FZJhvm2uzwfiCwP7AB
xKajU2gkboIy4ISrBMeAXRMwF+RZlMUy1iB+ztKdvKUSjtIYuej2/JkjhU4M5D+p
b/kP4E8PzRMImbZoK+QWNwk6C1jkHn2wHrF1/kWgM6CnkVqNWFEZlUduEt50Hpeq
bzzZsarqcJaYbaHE5Lrsv5rWc2SBIM46n4UFxoBFo6CcQ+UYO4WWZaIfzd2f4e84
1Tc4kW2ewxmjaYkgF6GEhMaNuqLsf7DjqVubranUXnKUk8S0WhIF13ynCLRw4H97
So5iZ+4bc9H+B9RShUMR6H9e6q9INYU3s3XKNrbxSkuVQXxozmXP+aBFM1oOzGTZ
sxHuWr08+VwjsINGRGbhbjTCS5u9qKDhevkQySxbD8vlsncsbNFqEPKkG9CfVOS+
EcJNIwDyUSBQs207nG1Z4xLgpn6M1xHivWvauTpRRS2a31MTHeRTp3rkVh+ViISP
E2Z1mo62xW9hNhpduRERWwb/giYWhlx+WT2oqoIG1WeY4eoJobZMIryc29/vDr3A
o/5e6JNF3h3tDTZhfO/EVfzK3yp34HfvfCKeElIWVmxCr80WKvA7GFJom5Pu7fD8
gGoJ6NxuGdbXEBLKSGKjTNqSTy9N5DnwcLFAMlTovHbHHJu6/ycwslOZeN++cVQ/
gFhprhKxCGFuTYqLF0enKSnVUtLiL44+YpNYAso9Utc/N5W/+MbfXypphJFzK/BP
Pw8kZ4PkRw+DjtzSq61w+C7lFTLnb+u5lNxkD2S0RshXuOJGFqqmPmM49295jcnK
8oJmIIfwWEBaOjcDXJwDrXInoDazyCiRK6voaV0aJsJ8i1eGiuqpl6T+QT8BaXcj
2TNYuZdmCzX1EFasaxQmSj+CgbPpvb+YtRIQdFB91ATmMAUxk4a2L/NAdIMVK2YG
ZYosGFmCAXgqgmfXiTM+Pg0BXWFb2r/dpb7mURW9snQE3mYHuvxm8kiWRQo11MD6
0iec41Z442uhDkSqYaH0sat2ruFtHUImWVNen+cpuys14t9j8wCC0UQ6pzpJbkPF
vfY5iUOJpZ7SulG/J7mMXoRx/QKAfrbBCjgBcyabUy5Df37Vy114MSWsWF0axZun
ldlrrqm79u7R+32Undgkg3oeyUChAqEI05P0q1gREsj4ZM8OLfgnjUHtX/b/Ybe4
q0P1g2T76PdUIXRmgxbPk1lP61VEUWF+v2tSGJRdzMplx2EOvfNSTm4fuy9qnOvk
7bHduceRwVRAB2dabMme00JgA/Jc9mQ0kYKpCQRZdAB/6mrlkkARIvR/+5aJK3KI
2tI0W3j3596GKJ/UUZXSbDHgggwYq62wFRna8AxFAjLNLaCE/Ty4LJgyoVraCdsS
6wseBioKiGWC9roHhp7+uMFMNS/e6LL2JZ6Upsolr6kbacr2P72gjc1b4IbX/bbl
/Yc/ctPpnUbO+PYjDtq0u/pM+gDlRDdQi8dqE2ljtT3WaRbLqEHntggTG4f5M4DN
RR0WbYFOJYbXOaQxLlfkmfebZAFvXb4qBkMLf9RLSajR3MiNMJyseWXt3y5PZlPN
dYTlBsU+4YMbSfIHnyLbhcFjkcxedRcS/xnKUJWUhThZENbldZw+k1ZViH2tuHtv
VNRqr3pp+63uKkfhwVMqgeDwte1T0uZVgjIwiZo/QyXj72EgyXSF3eKe9pJj9SFh
SoSZh/151eRFFKCmRZMU2+7d9qw4Dqhu8IV4R/wYCXQ4+ecksFPtEbJGOQgU/zZh
7Y5yyg/2uX5UHjzQvraN2GXFEsBzEYi7N2gwRYN2WgLsNCVHJskswczweO2VnTVN
AA0GkG2kMWpeRjytQ/cZYs+8YtkXSVb0eCyhyHhT+8TXVqnIHlBMGSwRbS9N3vOM
rH1oF+SnfbcvtcGag9A28VHUKROVQoqV4rZxDaVp6BKC3EYlSm34mH/IYIzyuoDH
dBVjZcMDRzY8odDu3asCo1DSJh49xeRXP4NzzJ483NwCXfEYwydEbzycd/A1e7RL
71wmQA5cV0DllBTLFEVwXcb0vl/GlKoTllpREG4ncSmrWViGZrH//uS9D7V3JIv1
zwBhaZvmnF0H+rBymnkrs4L8Ae1X2GKJrvbZa3XRWG+dGsssr4zNTlgwuTGAkub5
vDOKqnlr2UyO6B0SEA45Dbq7AIvQ4JhZAXRaJDCyYEKZSoNfvEU7jjStWMOJ89aG
W+YCwnYOLfYVwcgiCMcBp6TnkQn7T+ycGM9IcuZWHB18JGykGY0akGSOOmoO0hxe
qnnaEXH3O/Ectx8F9cWIki14Wi+JxvH+Aj6FkCFs5bKpiuuZuec9F4ZqUgAd/rZm
CyrqKoJHIXSphbYaG1bZElIsnH4wAH9PTplu0yDCX+QsgUR2jKuZ7zZ5zALQ0w4I
5307FD8cLJCMTo9/46ZwIB3pmUK6F3l+uytall/9iyAotTOraUFFnpk328JM/7AL
3IiARJrk5mAv9RO/aTt9GqnGYQl+ISF8gfH6lQnj0Fv3KdwtXvAsMYka9vNb7lqJ
SvYRFIMcHzsSG8hea/wEklRq+KhHbi5U4qJn9Ytyjk+1UFAi6Tt3xFXFLijUoLD7
vk6FYonGPxhv56SLj4x9K8d+qilCaAaRXye1mSNkUkJ7C9cAGPTDQGzOqQlfAxYW
w7O7Qzk3E9JWTwcN62ZqcmMwC2pgex4xxoJ+4p2Bj3qsX2sJQJTpOGbyXJdleeH0
WQH1qlOK8japusphNkJ9BPxUf13vsVqtYR417rPyhW/4J8Wy5qzN8RjqsmwuENyo
2gSBp6pTQrahxK9vOfz6U0DoZhwVU3v+Orj6ZGLWx6MZbOL5hIQqRnq5REEu/QrE
2IyJAbDDmS3HN5QxMDfSLlcwuoWTRp5zLOHCfcr7hZAEc9l3pasYX2R/fg+LuVoS
ZGeVXuu0fMECODF6UWdDLSoCy8YZEUNlSpFYV37AE/hWW645RINIHCYXje3ux4cl
yE9NtoD1I36H+xA9KHLCcDHrVbyYdjQe9zNpRX7e9ajfUADyX+xuydSEdbBywrER
v8q7hjE1N8SYjKGpyJSHk6mWt3SKr858qFozLpo6pkaGNsekpSxQkN8h7sXT8ZmS
w3iQyelpbbrYqaD3sNn/p2HwLO/RJebj+dzLWG0lMCcnnX7MhNnnqmru4ih42rle
uLmJzR2g4LvrfTMtcWyUQTI0PuP8nlPo3CsKm/sReuvaYJznrsyb27c4FoZt9CUP
ItmffNjGX4y/ZyjtLwlucg4lwvT9aJr2P166LE3TIlnffwh2YVFJZpLpc5nCqbDr
jGotJbNhhMyybzRHYKfEWyJ78sif6x7ne/c/y4jRUX/8IbOA1dHiX9b3w4aOXOCk
VjZyY2gtlElOgw0tX/N5k6TsLTmJeNziFXaXHgRfRa2HDas+cG5oX4xLqcK4qy/B
AiT8CJmZx/M9KN3Lx3fOEoMO7SViG7VdAJIfNR8RCZbAgp8dLvG9sTtTIVQqTeor
QP4jQB9gpHm5wNfx+I6/9krqnIEEuT8gp2UWUD4YfaPEE6k1b0HPGuup6y+sVUkJ
4agY4iCwXX/uC8hBLJ2eqv8Sy/Bdmc02XhEt5fJJ8Syxd6LzCEo4wllWQtM8pV7+
AXWmhQSLx607WDtwqJX9lj1qXt4p6FSZopvUZ8uqwSnch2dqd7hv2QyvNYDH1z61
r0WxwvpGNcF+78TPs/0mgj+kH3y0ZObpyspsX1+Qd57Pqlg/WwniS4mTNRaWJbmf
Iwf4lzCqcwqKRW8E5WXHSpQx+Vf9M64MQkBLmYt1ZowkJIbA9llsA/nbYsns+5ui
gBnX1O60C+7RopByh/Q6sRGhv3R9UU63DWpIjnfoyTgsKCRZf9ln283v9kyVAK+S
b2ZyCf09irks/NbszidsNH3MbtWOqLEAKjTMIiKVAa09pvI/nk89vgE2I3oL8c8S
n8SE497PMJZPgAvhdhQRNodS6KxExsUsTQ66Sq0vXxq/4RWDS5uOlF77S8NVqggh
zm5m78UGl231zoQNMWnynqg2cC68wlV5k/f7MM5EWP8VNbE5Yzo7iFWY1aBUyUDj
NvkOnpQmjoDvKfygekyb2amwQ4i1EnH+G0LDxhtx8cFWss1ObXB62WNAu6Xx1DdS
wEeO5edZtSV2S82oyzcQtlxYJYHa11eEKISVNwrt6pfiukFsZEy5huBCHCM4RVqe
mlQCPt9DD/l1kRHBAi/8dAJzT0Pch6DNyORW+LV400G+1Wi5J8JLVotaau+yPFdC
h9voD66/gIj8RnsY1I3KuZGtXNLGM/IE4EjZluLgwkAhLhmZB8gfvsRRngUVz06v
/aWA7MSVZQ1lhgnfTHHf9IoqPeRA6Gya6oMD0poppw48nIiHphRlPGxuLzBfLSoV
0Kv7u5c5kBCmDyK7sL0+K3TRXVQtKCKaLFd31YHi02CyA+X9Sq/6XwADXL7Vp5cJ
IUgAqiEhf+49JvV6PYpxbInmqL2vSE9N4XBBt8/Yz6M3T8MDwmi9MQMgWMDxbg4P
xHIjoFje2q72knBvcWMG5NC5+xUqATA5ZaczW9PFzZ/FvVrSrLSATc/ofB11R2BU
fPsOFhsCOXOt0KnxPSJFEDdpz1J+OY7PA4E28OnMrzO8u8PNR/Eb+vSsXUW3SE0U
sQhugghastBo4WcIyRoa//69OEs6b63hMVcD6Q3N2UAr/6c6vTgafBDfkfQPE9dn
KcT7G9lEc0CSU45poCPldYWuhuQ4hV8IDL3dEgwy+XlXR1O9SE30iJOM+6FLz0Tk
l3K6QGFsXjaqKIQCE5C4L1/4LZZ8DLVbvuyiRD30/QOOh+xjYIxirTX6IV2O9nvZ
7KXS8pb4PJ5f5ahSr3JQZaXjeWEkzlS3rI3XfHn0UV8+W7yo8WvabCqtHFzmpvN8
ZmclGu02gBRx0pFfmSyYDvhNrv7b6+YNUDrCjg8PEfVGij4lFY3EzWGRy23san6k
U8OvnXWuEwmva+7Upq+NaJa1aa181FbILyp9KCAv4xR62CdCvydXaHKNE0OL+jZT
ZnfcQy4PdRCg5eMF/lWwFAQqmdvPItEMkD/N1KsC4XWoJGtgb6nYed5j0YyjXvbn
r2sX/24L5vRR6q5k3+5LeJx+N5yaabDs/4ljwAu/THqO7+sFvGRBObZHC/4H1tkD
Pxn9OeYXqdFSPic0m9a8aZ1znhgsW6zOwKGI04KQkCop/GVtUmQpdq8VMBXFqyAD
4++L/6JedRp4SptDL0YRVPaUcr1EMvyTyEXtYrUJ9R0AwfAT+9netuvQiIQck0ZH
/XFC+KbGBw9C4VAxKrG/Yt07PpcO8DH0L1i6wOZRmQfMleqIK4+gtnCdxaVJXrg4
qUO2EKpjw3Cw+LJRDRZW+tEwOpcbRpKgSvkvovRh/O79DG5tgzDTHpBjBLtHH7xc
cN66dHZgN8xRx4nBn0sj017xgi6fxAQJb1F24Bkt3uOYBlBvPlXMsyB+cFqhNz+H
aD8OU/kY+uOSsr1pVuIGElkRqf60cvyuyajmSoztvy4BWDvbcJiCCfmqJLcjLPty
jTD6iBWytOTwaK8EnZ5tJDQi/1gTERdWb9hgLtQljHdZ7Ym6fgoPDLCg4P7A1KUk
rsIz2dCR6iM7wn7P/9S4FjG1c28EiKsinSzwxPXKxa2XKlVIK5loKbzuQCXUjPEZ
9dY0/7nR1YXUVLajrN581j6MVIvpEu+4MIwVoImn68PS5JptucwJa/WJv4C64OwN
XP+j+UnBZLp65hI9OLvaQKT4XpZHmToD6kti2Hn6o0yBlYjvfIy1I4P/CSl8+ztz
ev2U48KCKCHy2K6sQdEyr7kPbokkQlINqhy6aOI7VBrgul6O7K9XujLO5euZRgMY
rS2rEUJAxuvAcmaAuwUvtLePFZ0+OD131BjJAxRoni4zFFFGmZ6fxlBVXfWZUHHU
fvTZgx3mwOQjN7fJ285XgMoK/kmRDOYw6dwO1//Zb4uDUtGvTbCA41tSysPCT5m7
vC+JRkfBDaqTyHah2c4qCZ1SDqsLL5Ms3yLwa6oEe/Fz+jxmwj2A/6cPo2HBMBzC
VMMjhYhIpnCLSCNjlFfsrpwFI5OMxwuR7ILZUDiw7D0cuxsYUGYFtIXDzDwyoRk5
QewpeEviwx5zesSURr2e5yng+CKORRx04yNDzwheeKpm+RjZ/or6OVXLlG0tF2ap
A8oB9WuoHeF7spgUtXmoiNSoOXH0KqxhJCbSxAgyYtIu+WY7doiUQC1XpD5PEqpb
Wj5p93hzEU3Aeyb7Y+4yk2HMZtjulbYFYFDXrn9N+qol0QN1NtRhf4yr4wJ6o2h4
TY5UaxnvTU/A/8XBc5Gwcmzds7Jo3yM2YbNJbhgeeiNZ73sZOmzvTVlNE1l8GBby
z6b9JBRU7uTBn/aiReCjzAK8iW6xouOxXZ2HXxEQPc8B//kxMaHLGz33ZvcjcxQZ
ZxJ5vQ4MAOQaEdoBVB0tkrn4FeBKKsKF/ChMHUgCRAEH6+OGheyjiy1hB3vvjXxB
cZ5SMyd/KvAFRlHxzZNbyZEsu6gh5Drc7Oyh7rPHCAMWUFZGezgH23gJTuscB1G0
WEkq8gMfI00LR4heS9BpaylsCPepoD4W6dMqRxHUm/OoVuhy7JSwG/cvMnvCuYcW
tyUn1jwkZwxes0/8AzDuW0YUfwmvYyTx26CI7s1Yo/KOKBVcGkqyW7RN7foPdylg
YYDPCapFIiqkBiKiMKFL3fhNV6xGlfZajzqeGQxUum1Rg1vsWGUGYbuxbLSxQLFF
nq8rQZbvX9XBJ49ZpO3YVFtNmRC8hqpkiLGR0RBDjnGrVQtX7ixQ0eeNVxzhIXcu
LXh9XiCCJ2L/FiUNg4DzkGrprCFQZINCSau7UNzaran5dTylGc91Jrh/fzaTuXoA
tS79fTjOjx9H1hW0KzP5AaqKfxjgyI0bTiKYSpJij4a3BfKGnFA1TdQ5F1FCjPld
7/VE0Xb5ANh//CihH6gmQrU7BKSLT30CkJvop3c90l84bvsL/bGbjFLKVBmVtrqW
3zytuKjT7yqWqGHaDYCXK5tz5SvGjKzNBT9fYVkDtwdcouZWfLj+pFejzGRBsuON
XnZcw+IGKZHvUhC9UX41WWwrprLGXnOVT1R0F7iCXeHlifmK6wlaHwL9A4NuIM1R
eRU8IeHDgWRxVM/fP8YVvR643ZzK1l9/tMTbQ1W66uvvdcuOAemUqR8wwz5Wnnc0
C+/5WlNbajvoASQTe1NAffFm44zyRbjxc+ohFWMelELF+cOVAIeEnDzl6GAEj2QB
vunUz0TTPX4f6SLfsjp8zGHxlyYhsnmQzitoNhHMZcSppHwYCPNzVyMRvDf8uA/S
hRbiz6Oc5GCp/6a38Fiq57v5KpuXiBekRMWqNcmFbBxiV1d2hC2Zr7sxtBP0xE11
irWssWzF4DcFH/GQzXwcBbG4yuo9FfEeyLuVYW1xK+PAkq4zlwIgUvncmPPYIoVj
8kNfqm/T7y5cVE8QBt2r1wMPrSL4uxzkjL0+lCMOvvS1cBHgjp9kBngeh8ZjJPn8
uRmNcin7c6WQzhWyvLFOSCZiJ3xZ3ofrP1t4IUShYPXy0S106iDMYQnenHpeKwDK
gqxcHFKME/eC/soOHCUIGzHHcBm+dMdhpKS2GxEYmU5F1LCT7F5yHoYTOV456kg1
Z2e+Ve4UPs28tWcIDpVGuBYS0c+YDsHBqu/kUyQOf49qzPGIa+zV3ffjqbBu/ZUt
S8SuTnrCDykFzey34X/ya+ZwUnFpzvgHesXc5s45B6bcv9eriKEQj6LOvUUQ3vgS
s/0XxfT8HyX49GacanfdAEYub6qIjNldLxjxvaZjqGeN4exfc4BRuzkr2PXbtN7B
fVUdQLKiVjUPb6x7LpoYyFzadTyvJ7EyAtReX8/dFRgwah0ojl/87EXwLFBncHzE
AMU5aBL6J+M5cuKf3+dt3JofASV52EbVRPY+cQuRgPlyeeEzz0s5byU4+KbineAk
LP393QMwifMzHB673h0g63WrYBAtUJpAPFF581Rjqzoa2SLwREBNW1pjeb6Rh3ZQ
Sxnfd55q8Ro44MOUo0NrCEWtR7iksWEnFXGSY3q9pcX/at4iEFjKWya+nJduBgdP
hflbqf7JTsnx9sZ2FKHuquqeXNGfa3b92wX+pMrHO07FPWuy21NwPmf64b4clhtR
vqMnpvQcvJ7tGBSmCZ5rBE+GNj22cRmiowTRTHrX6Pxy8vwj4UuMEAGUaME1w0nr
T3YWdupahYQD6EqahtpzHO95TliAHOFs0CqyUeDhWnZwaGny8l6CBUqAgrk2snh3
320ORYs2xKbK8dsROIf0dwAaNJwgCMWmN50IXBh2iuLZQN7G31qzva6FLYaD8w+P
0ldAjyw2z8nYzila2pgxpLG/cBNuY9spqsbUZCMuDFGQnxYoO+zLnG1Kx7HXSf2K
2UpczAtNdXDjbqbeaI36f3X/rUBCqOVhfulKVIdjrl/uOs+GgCbR2SSjyIB+z3h6
1aFOZ19MUuyT5lT/bU0RTnZZOjQ7o/CMaBKo4YfthKip9UzBDveq6L6cuijJiKpK
qDo+2PKTwCl8FlOaT7csRl9+6Vqv3dmWvS+GNBzjrCkEZVD0ZhLZD3QuTqLwYdyY
77shinVsjVJODpzhcRIhBD9v+pOKbdkR7OhaOebeFLFXmTsjBOGuye2zd7upYOeQ
XGKdp+wiYIXmrgWLJmuyEOvoareYNAdDKY84NRfVthRxlRmF6Wl+q3Pp2I1eio6j
KCNPL2RzPhkXHTnWjTYtgzQ+bVGYzX4nPK1x6qq9az780Lx4sIIBHgkzJUW6ufPR
xqE83nCh63WWnS89/gWnyJUIjRsB6yvp0+OeW3dPyACTAjX6stlch43gO0IawpR/
5vwEaRroJBG4iDe+RH12o9frjXV4A0InaoRMx7s53P2jUGOZXLduNPvPFm1mxUu+
ky2d5IhMuK0civ3aXEhgYcz2oWYz7/tRGARqUt+pdgQhVIJ63sOlsAyYFRQjGcWj
x0ZS/V8YeqdCiClVEQm0NyCKcCZqlF1hXuKuoP5qsHBfYRLx/WDLVyLGvsS0pgc1
H3FqxLACtmMw3nnInFygjE2BPx3kS5jeWrbO3BdvEbptEpxEdRuciCM5boOx0grU
bJljlHcLvLKGhvY2VL0AifyN5ztNDaDrjuOIxI+lFMvCYHCLKk4aUkezbHrORmVb
5Rxe0EX3taZTHPoHRa/jfZy5B+kEcHRrNeoGwyAQsY5L1qk/yylTAlHW6uwQBvk2
LYXrtXK0RKQmB9ovqQqUjxZODgVvR7Qpuf386bf7Wzn8b2dQYySILYu/wkjk9n1E
Zl5dW2wRWUEkI/TieQlnwHp+x5xrShzhWaNJiHC2MOmCoNpAF1aTh2zrg99JWyf2
KbBOV9V++xqWhSpHTltNSUe6nEHGeGEeDPbxKZzO5GsMEOazY+sQctJJWe009CxS
++quCy4WQVcNlOtF899ZKrXD6Ai/waeTPLJCMEIAOEQudyvn8J74FyGhfNZq1T8r
NXrnbI+PzpVszNV46K6mpOQIbdtOk9wruEYozK1JhNjbgFB9FU7spU3Jcpacew/L
CHt0P2mGjNoVCuS2wt/6SvepaAGSvZCypmUeRR6BK6GysQblVf8gIue/KHNH7rTE
k2Kq016C1FivAikn3hpiCZtR9vji8x0D9tB+EKuDgpn5CvM5Oq8MMRtzFM1KXppT
l72xICkMLKOTWe8qk1ber0ZIvwoF3UDf3o+MEHkcGp2Ocazz1GLimoC5RDHnBncA
sayreOBJ6SpW2F5ac9S5QK/w9YQAHRMZv/XLJsTSve14lNzzGkBc8cvlS3oboY4S
p8ACDbIS/IbqitNhH4DIec1qLhzhY3BtyxYVA2YGPiJc7iAUs2iSuQos6JwORfdr
iSmkBeLhAWn2Fj+pEpornI4sNUs6jV9BSr0iQ/D1CxvwBQfMWLtKUt3Uf+sCZAe9
7SpVEliPoSEkxA0Ul9jD6h1at2M0mdyhkX24JBNMZkfyummxetlGStuXtidilQf5
MFUaqtErjsofWHLlbKMEuM+3KqikqZQtmizC1rQef0cQAKX0sG4KzRZ1xxbBoPao
6FH1Zo9tXb++y3bPYD/ma0GRr2rfmiWhlJUDjSYWxhr4YTYAZzN3o0NdXBippT7U
z3tNWF4vnzeKBMLP2rZSEFbG/jW9QwxfAXflX51ozTfzk7VXdZWnVdYqxVTBHE9m
bV30i5VU0Y2tKfFZL4y3cZ6BOjrOyZWlGqr+XWGmf9n4XOUiiGBVa/tEEtc00Qzf
36zc+J+bCKqbMFxmsdhEvGV+PlhtN5CTUcWV6myG0lAaGnd48sABpFY6eE9Mr0C4
HL4+6DRKRbaTTqII7q+0sD5NsV6iYFMSMXCs3H2wimS2eb6vMSxwvhfQlVXiLkIH
VvFQMEI53Hz0WsL38hHtrnwkU9BmYrGO5PSJ0kaNaEg6LdYDpRXv0Ai5sHzdvIgd
9B5+5Cwium5IQZKqmmgks37eDPTVcV2962jczmMIpZaeHCNZjFTsbxaIt/nl6yiz
mF79DHJnaoLcm5GS1Jg29FjDgHIC/QggWTC1tdjliBlsAKW9iZSi5pg77s7eFA8H
Uu9nM8g5DncI+QgZBALJ/3tmLuAfARy0gmmB80oDCYBe1Zten5eoK26utAbY/WXX
r+wJLUn+uKc+IwGypUtpB6tQknwDyFG+D5nuFetEEXRFhVMjuzcHn2ftrywznDX/
4z4lkAzMN2fLo/ZSQzdfnCYEDvk4+x7dIMg2ltjeksK4FPz6/Zl0Fkwjs6d8LZPX
MkRkz6N1eKvSjTFihZpZaDkE45uXQD0zJc0cnWkJTpe3NV5Lr+9H/YDER5pM9VkU
3Yea+j/k1Sd6OUVdxjVU9lL7kMWWjigetxxnuO5y9FkxSx7FrqKZERaahh9FN2aZ
hGsG9L9tBfinA6+4/irHzT5vPlXsI+DlBWlfZBqjU23hmJ2z7DS82h4l+Owa3Ja3
x8MkCb6IYxqfwSz9Ucwl+EVXP84SSEvoD7hIOFVEOcVa1+b8M5ritqKxRc1y/7OX
Bm2FDTeNEsxESZw3cCS2RA4MNfuPw/4gBR8Z4rCg9p4Qvg19pcMWCGrb2XgjRq6+
LIICT5abwE6lryqy/teJYmHEk9mnhfa54DrCJpA8hM3McCAIm+WQIl6tCXoKl1i6
cYk3XBrTD9JoDhgSrVpjTZ8Z48UetvhsYNgskS+OeDtOtpp70AJ7p8WqJyG8Cfv4
OkKpIiRy7fhbjYwlkH4Aqv0aPHYMRTSLW4tgSuGzdGw4awe8U0nZ4woQ97DC+Az0
rh07TiVpNYWUPt3f8kR/Ly+qsvlZdyJQAqcgj0XJRo+IlIitT8Rrd2WIRBoGXuzo
lFzT9sOugSmG5b8XopFIvu4xOHCg8NpJBsMyNsltbFCTtVNsdX9XfGu0JbHHoNBs
TF83hNIZINGtTgPELfkQ2QdqiZVAkZ0E5b3wVGHfpcTu69I1ydDPsPuxcWiW3tZ1
A0h3bJ9n3zFz45Wi8AFR3CC1ZZLmTC0ocZUrcndZiUkQiiCAH70AAlgPpT4L01yo
uoCaaMoNeVAho8A5g5GSfh0VaBMcccLRkOwQGx47sEGMBcTtQArHbudf6JMqUrEz
KmyxAxtfldLsM/VBKYOLCB3UjjUNbDGqcV4ok1tOt89EbcqfYMpkeG/JCbH0+1Ta
mRJRxrlY+N4Jq6PSxbDhpwArSbeXXuzV0+4Im2J65as3/6ajaapTv6Rhpfq1PO2a
W43jagrC3EQgF+C/JpgUAffEYZNCYQ7ZY2mE0nTpGO/uhhxwApesLmq9Y7lrCtim
4a+YfOpyTOi8Rv6L5MQP+HWJDM6qXo9xfyfXS+zxMeicq258gjvWdhB+PGkKWYS4
ImjdgfyYXPn1zejTLl0lww==
`protect END_PROTECTED