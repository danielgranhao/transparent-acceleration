-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
tUcr7prok7c6eH5d0supXNGHLdh8HPnKO3yIBuR8elm0LGc6mGS1Lth9x5aB7O++cMhdLjaDo35p
MijIbRiK9wPv6u4FFxxR4SQ/TxAdkhkLtc3RIARGR5mJkb97obJUeEVTm/BWVbbZddHgo+36BonV
px8spk3RR+esx5Vc7pjxoIrTTvSS5Q5b/Ulu3x4BuZUujsfMSMQoyJlhgxECDioNT3Sitj3bJjDG
jGpx06ipvEHMUdiywpokCjCIeazMk1VgVdG115R1riJh8SqnwJVB7iY/zHpNDk7GcLxiJRKThnj8
eN7BpZG2SQ39vkAy1/rrOSciWEZUFx0vpwSQ1g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5184)
`protect data_block
8l0ZDKErjr0sPw1eAliTHkK6IJd1LdmuiawuV91HYPNaFd2ZZgu0tUTFJAVFzSHlSWHZfL0Dygjl
1/R9XV760ouk9gGKMYpp2TMoKJj37LApgaBmxsZS4N0XI51HVMpO4wY77zlqFL3Kp7diNw+0d+7g
OYG4O+RjFw9AF1WEEZvvpf9Dn/iZiJpZNia44L3RxG67HXFyWlbHL26rNWv53jfGuImCW1N6OiKF
dtT+lrOGuTvwoXbxQNo8egYkGQciNJcgi1LOIIR7jkh3usmVw1lGfQhqPpj3z/0Nw6eEQu02e8Ho
ttyDTzqlz/pQnO2C1nt8Oh1PdeyZ87lFptsa9tPixpl9TC4CAqKqaT7gygQl6iUSETXKQNlH0qBW
IgPbsZ1IUFJfpjoNSos7PYG/lAGcmkzlwJ08S7cR7CR9malKvnZLF4K4YyBdFMPbM4EiFI17xMLE
mXxfBqJb4m1cgHqf1fbtpQuAbDMOu4trIFVjGHiOTgnLujO+RqJ+iINplF+r2lfMO4lo/5WPz48Q
rKrbkF9+0EhYS0xZHhmFQGVPUtB6Ba3OaQb/cCXMc+7oyDS75ap25Ka0a1fXjHY/glF1X/9MYIiw
u2Si+WEjr5oh9EXWkQP1o1WNRG9jutwNsA0HI+1FuDDXYMEPI9V5C9FyAidA7DFxYEG/U3GxC5kD
igaBqFliMFHU8WjIglFMHg0ZUxsXcSV9H0RFKhJop+Sauo340dEZ3H+lv3oU02GRVtFXVUR530tX
zStaaMzTId+ysqWWpKpI1n8OhS2n4dS5REi7OXkOZ7wQw18twA6u9cgpSV5yCuEQYmTdijZ9NKqR
ypIEiZdzinwp8v72rP+jcivu5mUwLEIeQIkl5OGRUF9X+EA1Xlb5DjK52aNUt5oHCQg4XdVzaYMH
WeWPSU7jI7ON61DtIbwdq6PpufSMZ5WPbkNKH8b4eGvm1lQVy8v+9GD7hAHMEh8zRLRlA94dBsvl
2e1jdzDIK69ZZPbDX8xSkv/rNkE2fMphD7TqysHRR3eKM8qNIFdE74WqXpIJXEprveKK6uaTWEzK
kpYsOf1Ii+zr9dHQ6r8t/R/48zT72E8L+7+XFOmHtpGxUZztGgETiAp8PRwZxrRAxXtH1thlSRqS
uU0Cuu5J10KspfQuITn4ZhRMkH/ipSaWP6D6BkZarTMOxv+ou54fW0UYLKQPx/ZVpE/S/HDOQxgC
kYTm3A2J52gHwg3IFaT6jrBzUDQW8eVp6dE9Xr6qzBvndjHlStCGFuzUXrB/rDZp1ddt4nsc8nEQ
JJp5H9I6keE1YtTjnYS3zJgGIJ2CRaTX6bZ3q3NTku3yeb6AnlBSjfAVAAFHp7TNHsBA6eZIWErw
aZd23WTvcvcHJ8j0XD9g/PqJrROGt2Zqr90bhh+RRsq8UYifhYhXis01xW4XFMfmZckzprTWfYgl
GOOu9IWQMCrkED1eZCLAjGi3IL16eM+EP6bw9t5JlFYSoseU4uv4D9Bjcl2NwB/HVfW/FT68PWKI
hbS9zQv937Jx4rpUIKPpBplGbS21OHeER9HTDYsTz8VI1Yjx6LOvYfygdwESotdOiHI9uMQNji04
raixsyJEWUhWFmjfzUeX7WRNLVvPLVxPXzcKz9Nk5aSLqBVdr0FNjt5MPSxQ88JB98Mo1Oswvqnu
IlTra5XHUFLInvtvZgaDCX+RQPjHB7lTI7RFv/2jb4M7nzIV6pZKviyHJFtJehrfomtxTCbc0e+J
JDZhRlzsce9tXiVIs7PUQGGF/Fkrtg9zZX6LQTc/9EknMIFBfFZwR/cq6IgYnY461sQaDGD9NXH7
Lndijhy2/juhW5NX+XE5d8ZvhY1i4rROTVdSCEQZlNSAjif1DAfD8iVbBzcP769uLAN05j1srOUe
2PpEVGCtTGzK97Ptp7BJWyDEB73OO9OrCQC7xH9EREi9u59Xh1qDphxKKAB9NjSsW0dkNh7PEPUz
nd8fkzNijG5jDn13AIa3NRvPEWkdRUUHnBb0Br7wNgT6Em/1X8pYDbxA+pMZdagjy75AjIPOT+0P
XptiUpBuliP4tDEkxGJGSYw71fRCc/85UpubhHq23CnymbQ5y+8HwrIHsFgNjVzzP2C4B2HP+p6c
KJ6yXBO1UttB6qh3UmOjlIW75r19xzuiQPhaod0QTGBeSpEaYgNBIRTzf13XMP7NwWmrJKXkTypu
aRypMPR4MW0ba2LQOfC1RtzmGvKKBQeF3gbQxa2SGCvLCN/Nm+ZHEffGo3ZkyBLXXn6kZVD4StyN
vgBGXje2uoxlwjn17lH40cIeS9JF+tv0qEMlZodm0B7m/gyAJNVzaj4uSQSvpwQ3DTEGhUxQVBb0
jG3OMeICdzWUQCiWAZSD7klaO10ZWiCtyGT+/YoNXSsrdiyVr6NZPbMsJGDPSvPvY0eS0UHSf/6w
r/jekCX6Toqqg11mlY6+mdvxZO9nB5ogWKWKeS72WiePNqCDVnTkjKUE5Vo2LBijM7wvvpidyr8J
CsAT+WCFUQ1bo7cmlE8pO3iu/cana3HzNjUMDpafMN7oiyjpcmTSBHimtsPNQXEbzAt5DBnPHERD
LKEAJAzdEh5o2SAkYS8DOkYtOUFXpECcr3EcBvVC0vAV5ApzL3pxQH0FVQVSLZhxvliSNZYqG31K
r92vNy1O2NmeOg9TANzJSfjgU9o4Kh2AXwOvtipVvHnHps/L1C0PJTEhXPosMBI/FDnFFySpChC9
YV2ZV6k88lzc5yWGt2DqjhGfUzoWb/Xj7rcohwQYJhDylG1jU0bSYzhplWtWa9QwtzQ6sCLl2Cq/
A6Ok59EgGi/5Kn4YIOfTPg47piJ35uXFLoYDq1QM6yHUUEQHO8V9DfrOht/+M8JlcjauBylW/ZVJ
94lXy8PvWCBTAbSFbFtN89LqRJ4QliT2ksQUx5dSuw5B0l/JS53RK1Keebc36Us7F5cKfGg/whxI
s8yrfgQv5A1wHN4w18bHaOu/zq7g2UaLW5mUPtkguChiUkvD2tpE/KCzF0ra/skefbWneh6C8wWi
6AYqrFj6o6EPw9jNhy21YR5dGJ6WQx7n2S0y3PJEtUL/IxpQ/M2uJdB/exMkNitieXaTy9cTF0h0
Vq/hR2YHEq2JXfMoKH665DHlnxMQNBK4VQ0lZpGVB0+7z/HNC5Jjmj9RmJQVdcDBAOxr/xAYvWeu
B09N57b+S56SdHl/PD1b+kod3Au9WYFjMWIe9goJXkXyhDBwc8p8BPksDBWNugGko1/lkRP76Lox
dbISSdHO2H8nLdSZea/VVlp/rw32Ci9K3XQl4qQ/wR1FfCQx7nfzRzDrwDTTZpnIAl1tGT0UPC37
X4cV+iKcfKRVyoNz2V7QE3IRA7/TeK7mBZynm630J7UxtkN6bD0VLyDhkgTcol6lvUzPmEwe8cZ1
V88ImQ6sRSmT3U2WwyZdx9HkE/dc6Y99ZuCgKErydGprrq6TCjYeutgv2W7Ja/I+RFPMmLikOv3J
wZUOZXiFhIFFgrNtHk89mg6S5DGGEs37qopbX1op71e0gPW/V4NJSh0R/z3wYvGgymQ+tvjDfqNe
BeNehF1J+PfZT8GDZALxxoXKnBCGiIcuZs53c8YMDa7LC9T+e+HB77O+kklK2YmyKuqr2r63G2QJ
mxiISpvxICaa2N/AyKTNpBqr2qESQ4405+w+32jMQcOk9JlP8O03Pun0XY6evcIhg4mOuS8jlxE+
1RaMAiLjFgT2Dr3p5pYAR1OL5+CO3pb6MlgLC+ehK8Tfl/v6n9WJDpf26EepAJmdi7ypABMhupB3
KHAklzoqWzWxtTKjwY27NxchjX0lm6kfrPjkt1wf95ghC7rGjtFMrFV8n0x0JCgzLin2B1QCamv8
Dfo2eFDiv3pdnPmtpxPXWXEzsUQ1eR8aq0nwiUKBnVxVYwd9iKyesx/B3tVi6zT4eIdT/0DcaawF
fwvP45P1qN3QJPtDpqVhQ3HKldfMtZUOXdE7VqBW9U4pA29IWwj9Cj5MKdHgmY/6ZmjEugr143Ln
/1ylO0xnTa5dqmPpDE76RY7xB9HEHlJp2Oy99UcA9grar0K5dqbXBDEkuCHx5scN7i6mfnV9kyl3
uxuIjjOq23s1NXwXng+YJWMb+k8t4hXsHp0Z9ZveALH7D5gMM+OHf3FBeQQnFlGYuMTZyh0Vmf4e
9YgxMUWFCzBjmH6weZAQENPNWeIuC936bxncixteWFgfvS+CYwu5s+BXB35DqmVKxl6f/yWSVJQu
rBZApdfvWXWgaZ8N/qlb2S15F8MuAj6gYXjWMJW7ocQMe/wvvJsPIuSzgYL5IDRrTU/x0SAEf1Ks
+z3YeC6yhmB8xsmKFUvT4Df8RBByo0McWxxbcVSm3J2V+byjuco+GChM2Q+M708dz0cho5aKRrbk
e15bP9Qz1T0vUwXZnSQSg1Y8PmTkHjGEl9g0aW6pu9TvSSapjEVnKGjeyCVYU1282H0D9Kf6t8/Z
b1rxRGwT0mVZ6B+j43u2Qni7RiWuvt5S/bvpFiUcSzyeyIdvk8bT5Hh7vfwErblpspY1kPfk12dv
EDKZKzPSFKtRpnFvxApFuiChzBqMWZbZBbplOEo3ybQtpEn54JG2ufb49gIOsbvO8ssGn0itsxBT
vgNkLimB38SFOcPAFi5g+B7b+egXoVLVd6abecFzgoklmDwLGOgeoVIFZohLK9mM9W37BIqg6X9h
0VrEBuU3yshs37fvk2FLkl81V+Tr++dYMvc2KLkMHsWokVQwvTEijFt4kZLRnfPdbrgocPTuKhGQ
feuAkIwgyvy2FO5JL7OXfaJzdsfoIQLjIahaRlISzvZFkR285zDMeoMFdtmuPe4QHF1NirfbaZtQ
6IqIXU+u71tgAn0KLj5DHQAVHDV7J6aSnC3aCxPm/nN2Pw2J9RnJebXO8WoVPzlR/Td7u9ONIK5E
FUE+KJKFtruf0Qh0F1Op8/CAjXwKhQiyKCO8/PGv4GmsTkEEiAU+uE+Z9qd2I52mx57eNUk0oqub
9JdNDetTqlSFyzdZwHV0ow30vUglU/VJT/bkY4OeQ31ajyDwLk1yOqyjzQj5jdREK4xoQncM8cTI
RfkRF/6Bi16IIUiKru/GhYY+AhFmK71iGrMgIg/wkqs/q9+ijxr7i051nhszDFmiAjdfgyYvMEhG
Q3ZKWC8lDDi7yVsKnaF35kywuXUYNOOrGwasYGdeccywdb+5aCY/7RjRYzi7wFLsx/5O7Q/sC3b/
2llPOwGeVZZlMWqt5C6Rd63B2quEStdeqOw+Lzh2mdPQETJxX+712+/+iQH8qn/US3MbEqmywu/4
sCi26G4dWLVhljO8Tu5ZmvAVCX61SrTJvw3IX6tU8UewAcKeDHwh5yLlWDFTuDTwzdu1GAgsJ43/
w5Ib9hVVbURV05TW+tnxM2n8Ish/QYGk5s/MTvNzb+AO719Y5CZkIGv5T5vVoRvc+5lweHP7zDv3
rb48L6gBvCFTD2BlCp6oA7w738bOWBRjIyaCU+2/ObGCyDbAwZyfLg6A4hwUQ+BcKiRd2yaJATiw
/U/SVTB5VYtjMSqkJD4t2O6NMMm2v1rdIHsSH0XP59kwH9ZEe0TbrYkOiwleI//HFOBhU3BZ8Cin
WvwQCk9J/JKUP74EyCm7KNCX9D7j1G2wocSox7dDMZhY2+H2aWTbZlecdX7a9cIDX5jYtsSKA7wQ
RhPelqLyJY1FjJWbcHncRkg8/+WpBqqwsoTXQYVncUttAwVgkXuJNcjA7TFOZ0D8hQ4zI1D/i6Uy
/VOqqm9rK/0NzaMv5haZ73XoBOgbIAfVVt7SxiIn2U9/Zy3C6Z2HlRa1SPsiu2i67EExp9JaMury
EVA1ufFBeK9ZbxXWlIZKx/UKgvlSMIovSbrprIVr6SELKoJRptfN5S4FxoX/LdRlulioone3284X
sYBRt3yZlgMc8k07ap1VZ/i5JHIAEpGxdDlZUD/sODu503ZIE37r40TzbsJqWcz/HpPp/1/QHoIn
KRnlO+If9vpMMD3ZZ+5wlvACldZgZ7JEpIJtQ2JRPEYDoQei3+NXaDXeAuk+bkHTXJgmhFYtoNEe
GQkYl5+gfMF4Wg+iiZZinke6VEVU9n4BbvrvZJmGPMEFl6JZEWgw3PMBAEIbIggnwRtjKZP3Iobb
zMKCAatYk62tfwYqLlwI5uZBLFn/IlIlruDGiq9FXPpu6vWNBFgGh+DFbQHyYfBsJmLf42KBSD5y
RaQmkuDLa2Hm5oa5gRkKhSEjC3scb2XRHGjEaHOrrjjckmxNztLIenxbqXa9oL7yMmXgHdYmzcTE
Dv1pu9Bre8BXkARBFADkTtqH5qrgb1rQwYGcJ2VNtPFwYDl0EuYLms8SRY4YDhbawwCd9X81vOaA
qGGpJXLmO56UFEDV70p0WS9iiPfFaXdONVl87Eiq3Mft5wUJIqp1g3uxTsVIASy44m8isiG8ebay
tooq4yho5aOld9RiEEla5u4IA2066cQflnT/xGiFYAli4k1kEhnrXeg3cTRbl9FQt3r1LzT9qxEz
HUJoL8fUGGWG+VHA5X6+T83pbv1tyOmp0BqHXF52NQ3EM0fgrNOWgiV1eanoh0mbdNQicLKcrY8W
aGJw/diP1VESJd45GZHXCVMO41aW51RaMEWETTqH34upmusMYVS1q8MeN1H4ujbIA2ieLRKk2/JZ
fW3mNtEotiWkAPVJBgQ7ePrRUBs7YOK/EUstdxsbKI8qg2o2vN3Jcwoo7bsIXLWDfDYL3Yf1vGfr
M4b5+uEbZgIMN0E3owWSsS70qEzlgd1bngiJTYYg81mOuSx3uuK5eYtFBj4AOFiJYDcS1Alf+4v7
exNQvzvnCrXiuF0IyQKaVonD+c8q+c4Lu/Dzm6311nMf8PgThWx6d3DS6C3UTrO22Psg8o7o
`protect end_protected
