-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
--pragma protect begin_protected
--pragma protect key_keyowner=Cadence Design Systems.
--pragma protect key_keyname=CDS_KEY
--pragma protect key_method=RC5
--pragma protect key_block
WzunnCKO/gQXnwqJ5xQHsEGsPAkUtdmzDPFqf2wId3q7EMyS1wFDJAYBHjd3B+EH
LZ9pzOp2AfQlZNDwWJtnYlc5d23pKAu7hXlFGmcAUMDcanD1C4nUp1IrhXt94DpQ
P+Frzq6AOgIPGpanRZBiu9YoFGamerdwiJRwj9jzvXbySEAmNadOUA==
--pragma protect end_key_block
--pragma protect digest_block
7DBy4696uBXTzs5HAZ18YK0BiVs=
--pragma protect end_digest_block
--pragma protect data_block
G66EQM0/cKTIMHnN8hCUcwZnAPYeI2JFsOUYk7MRcKyw8OOpgaCpxfDjpkD0P3/q
4pm1MWS7R2dpO61nhKh1khpUZYWxSMynHzURQ2Od0NI/n/UnMnrq5xnG34Hzd5TG
S2qZRQQtEt9UzDaDJXB9X6Nn03W3ONfPZ1lv2LCF0M9O4ULHfL0PHtbsIz5ny5sP
IonfEkQ4PIfOJmEm5jUtgvT/R3DlUjPv/FDqOh2ty84T05fNXrsLI/dBToR1XL/B
B2+L3LjSRIIi2fPk7zyfHDHDookVFNv9KFZQOKoh756LZDrO+owe5y92sVeQ8I7v
6Z2mtkEjyy0FoApM8PI20hpQ6iqYzNoRagp2F3ZeHwMi/k2vDf9ek9ZBUXOabPvk
GvpTqcGxCvL1cdi9xCVNoB8EejBnyPXtps5A1Ws9hFE9nayVbyspZXi+LuZaMJ1Y
ogxzQ6tT32xDVrLVUhfiybMfXyy2f9o9VvV8VKKBcMop/UcQLHewJ36TC3dEcZtS
aFBMtmb1wuQPI1M24nflLXfvPjG3hg+YU/mF7lNTCZ8u+VN2rJscBWWUHSJzSPgu
8hy80z0T7RNs8T6bjgidpRYyKjz0lsAZ6S54KmE0BmQc1mdLAUkh8ujJhoFad+tx
vro8lJQkxnnJdY7AkCDM/ozloJgGEdzsgtDwsiowLy4+l8bl1Ca4DA+QROKWVk3M
LzIZb9F7/aDqvhj7Uci0g+GH3lG4OsXAl8IxhQPEFxglMBM1Y7QSjj0CDBfiwxuv
TEhkxl64p+/sQxwbCdQ2Tb9P1XEz9Q3kqFmOwv+PZ/1VNXpNzOebWcjWjBUSPMMg
84cNekoKEBviYsl2A/ukkn69RYHPZRINyUqHPGjVKZpBsvGuj7S8QuU+7uSF3dae
cLVpKkYEWiUxpum3GmleA9JRfQhNilCNNrVmug593Nfjy2fNs8Nj8U2YIxQSzvSj
8BPECYAOUrh5EA+CSck7/fCkJ3CnRTvMEsfJHvdLS2pAh37RykUeMt3d/p8m7co8
3lfDRCF1IQvJBwErhhgPU+MBlQ6bOpC9SjZgwCTA644ttsx4TjEw2oT0y3/11uBb
DCsmSUejyLNnMZCmNbtP42tAjEgNVP8ZAty+VF/k10VRp/zcv7kr5KiJxnQYAncc
+CK1xXYIWMKJMFyl+GwboqHnI7PPzIT3D4wCFz9VE0M0iLx4QIV/TKrAZL6E4o1K
1h6n9Xmv8/kfl7HKKTBiMR2WF0/S57o0RJe10nhfYeWvNKrebYOHHq4LkTib+a/T
GwH7tBMmdoqcCUM5N68SeZL6Y/MjZ6mADCE3GbNQ1ZjXhhFxVdf1I1FDTtTzczpm
mfLqA8EiTBIWYEV7kaCFJK7cV1j/hlqrNgZAlkeJttcjuHDZ9laMrbbqLQA7XEGe
6rzlfj6Bm9a16nOgWOvpeK0loaM4Ocgs2DlYxq4DQs8Sry6E91DaYm89NTmbn2Sz
DIqL5POIqL8ATFMu7g8EsKdyFxI1j38st9ipAdyS/vzdc10Ne/KV/Btc/K7JpaYX
bTUEORAwmPH4tbxvNvT24mPPqn/9mGVpvtGT4mi23V5FiAX9hVpmoV40+kJJGwiF
bgCqqZ1Xtr375KkASVaGJRFA5xBPqXFrjApYkETePZdj2pgOin+9EJIJ56DyxHKl
Hdh1gL9x18Ne5DcpEhfaL/CNkeZVbKNVfHgt7MegOAqWVNIIuHVVslMYoeGffDUg
pCZ0QoMi/GpSc+ckbyb6eAnuFfGskM4vvpDKnzDTTjZYhTzgKy17O61JSaIe5PrB
OhLjEHxzP0wxeUGn2aN344tzNDVI1/9RHmUdsiIko/Vf7zuMk29v0yfeDkmHoUDr
c8So1z0P1uiK0olCX0VMIj1aY9lksEh2h0+vikNUmzxY9MzzIkabxqXh5nVuavFa
vZmclH7hrp/3QdVsyf7uNW3fYLfXYjZhik95iafypTTiGiaXY72hK4O9UURvbafX
41RvCj2ygynG2CcRzgLoGLMAFkH1wV1bxvjmOih9R4ouFUXpHYOTOZFoQRDKP6IT
aJHZAw6Rw/v//tSq/CYTgwDxIWyA2Spb+d4T5DBwaCUuoh7b3hIFYWWs39RfOzzq
bpKJoJag6P0P5dHwkeExJ500XDgO+t4SDhYA3JVYYoHZ3Mj5vd7T/av7YylWbtd9
vhJcOtXiECviKUM6BJO+uQJNVji/vF4gZBuSic45wzt278qGTBiGXVo3CjscLf1t
2ir+obcm0BLyr15at4YGEgCsN4bZxmxFW2lJjE0KbtEM4GqOVtRUMjb6+C5mesu4
W9hBdtofVtd3CMnM0mlNIty04J//0yLDS1fvTKHcokYQd7CU51knSzCdkdJS29HW
x1ey6xjYMk1d32jrxdYwhTj8ANAPAwA8boIRntIg8OQGJn9UNvYsXlRlveVmJaCJ
97K6bg+D5dDPITH5xUYKG3ftcwa6jeCpahMoQ7H14jk4xeruGl8vgFevj5XLAQNI
P8JYgPJBRPDuQO9Iax9648Mq0cuP0k6KwuZtNJYKOi1mufOACr9ZcUrFf7BG4W7Q
SKnayxkIhRgDX6NJYMglEfaZM76/eS4I8aFoiECYg8Dftv78WEU/G3QnIFSd1MEz
xfhJ+8UKGbQ/n1ayKbwSoEzMHrr3vW37W1Qjdzhll2kvyixQZcivqYsnOhkMlFxj
Ye6+l183mBFjS0y+o0SYRJc5rAhzm7qlH/Z5evfNOdngyZRXqXiffKcqK84xnzV8
m3+8WZ6VZ5TeTvM1zkDcF+KHVPHm4EzwxQZq3VFmrS17m7vtl2B+L4p4lqbP9DD8
aVxW2GJoqOVRofF00afOeTNakCCAXYG2Gg6vYU55P3H4tGFy7bSVEhsdGl6fjPan
Rf8ygD5834It1zVr11WinDakBS5VNSJ7dm7SAxy1ixpdUD89HAtYynCQ8nILCBTY
iX0OgVMK6cvAsVBW06OOVxm2lYkJdqyr7bj2n0rjp9L3eXa1GafChe/hS/l9vwYi
F8YhyrDEGiExhrKnqtsKku7Bdkkqo5r3Xr4Pxk0Iu90/qxQVPMoH7kmWJiVj9FcY
VCqU4088vxbabgf7PwYxXHqiKg/9HJckvSD15hBkXbWroSYwCP0PrI+qeUN1U1Si
zqanLCcdIczk00toMUS+fVTjAwO6+JFYG3bzSEZ6dNW2osDmqOmGUi2lzZ+rqjMZ
4ivaXtt9bIU3n84vYYGVz6xspQ74sDg1Kt77gdYaHA7WuPqAL1HaC6zIepiEU+94
d9OUOo0lwwN5/arBEvsF6UN0FTYtHJrW7/EhdFzsHDm0zcQn+gw05VI8oJQFvNER
RDXWzwo6LMqAeYc7+f2l52oJammeHxAbNplD7vS4cHh6UWAAJpudLREQWNlyO2zC
YPk/SlFXc9FqJLFwhwXsO4438/bvLrvsg1ALjxIEgR0ThbyO8eNtNKqWjNg5cJor
bFKbS/ufhpaqxd/H6+f8SFEfgstkbT29vg8KyqYIQVGkoGt2y4iwAgANxvntf2ph
JuPp4+FOUQH5irXvciTnhbG3UgyYnkDWdYGJQT68CT75cJP8bIhxxRI+5LPCxN1W
qUOt0UiVhhUPU7haJgtObl2U67iMqR2QtaiAe/WjTsn5IIAgHiOqEYTEili0BY0l
c0EFroGxIA0JB+At7ARiNcw4polWOBB0tDesOLLmrLJEe576L2098K5AhTWgDaZA
RlONmAO2XPfMLHqFS8XXA/fABged/3VinlRgkv/e4KDpdd5fQyO9eXOc04ZetXx+
2CXAFE9dG72M7VDro7Y+jYczMDCgDIrZSd/KSn99h/kBCWZYnVwnEfCl/Rt0LhpC
IOzKgwPTKIFlP0bJYqntFDgL3pm+09HdFmo7vVZoomotgKkztsA8fVcO6NhqLUCz
6JuO/PKITM9PtPo5gImw52M/rXKDys/AtdjafAqEIPM8dm/vBj39uaBTj+hseYGV
3CngPNe3m8WZAv62dMANfJ6+QvetXGTDZGhTmYauQpu3aP5aq0wZX+Jye4vujY6c
qmRARIjbBqwOhZah4hMRK78oySgW+twunwdGsyNGtj+CQN+Wwiq7j8zFSsyL0MXo
8km8EiI+SPhqCKyoer3FKiGXJiRx6fJW/GMfmK8yGbYGju95mt4WEw02r3Y+Brsd
5kwR1vFRVIzY+A8lVm/ZhMEEsNZK3CRjlQs5+2BunMKz641yjcAEG+ZcIcNvWq+m
yGsI3oqjCcnU6fBKparmqjnP4I0M8h1/m/P7H+TWuMtgALYVsZMxQ99A0n8polGh
Tr/87MvVQDnpmB2NFt4Pg71Fil/zt7EGBJNjHIx6u12G7+gA76lRRX6NT1+txEfk
IoCquAfoy/NMeYHq2O2CWQtjVrMVwB7479uFzfL+psbAsDqiV3TJmdvgTb7nGoo8
id0betZonlpm0YFGkqpaYhj5K5FRHejdDFcLlmE/Nt/eBFRCn6nSXooXzNxVxkA6
xRZRI9xMObgdACqrHNk3JvjC2O79uihWO6faZ5b5SwhCVPqWNnuk+GRsNpkvvDbz
xHQMRGN3KC2T9nTxbWXivZ2S7dTclZRq3QjMEokMM8UDa8vdVhvlRfBHca2tuOU5
MYWqk3mM9S8JTYZGas+L05MgMYLi9Wy6KA6Q4TnYvELhHbbmE/Y3/MIxVDdv8QGs
9a8SZ2+rqVQuzjJMnHaxowj91HDdwnFIY17i2dANeLic0fNt5o/9hnfSfA/1WoVs
Zq6m23YuSK3+eYWWYaFZdhOUgubRoLqy24cz2HtVsWiIL5OJ5kNZ9iReg+epgeZd
zsl32+FdYHh/pqXkXeyRcnODVZCQIOlJcz+0dirVWyNeeqOAyJrixu4p6XlnUT1l
DRksntk/3YAw0V89ZVEGeZ3B9Szp3xK5hVvsTMjQESFe7dLwgamAqDYIoJkjg2aa
jyAufZiB6fQbBZ8908Y1Qjdpifq2V7lzYrZO3tghDwSiVWxml+5r0k6kRLMOSQ41
pNOMl8B08Yu0qOBUoxwK4CLaI97WhEr5MSYIj78p929aCRqVCY4JGYw8lE1IONJB
NmGW1Td/eIaKxEJSGmOaZM0yznf2TCguD/jN74NXKu+ZQ0F8claoMLguMvnkiJ4A
8j81BSvZL6hEBSLvAqY47zkebj2YIXbhtbIsSaVqbsgDFxGX766jDn0jUISA6koT
kXM1NMLUb+i4+CJHAHCsQqX7tuEeR3R9Vfdspkc8hEW9YVP8I6xOoTEOaowhxx9f
21uL9ioGvBMGMLcmiXjMyKiO/09e3pxyDyTTnQ4MbulCDWzLb5eFzvGBrOIcKY4d
bQnvCpm7xj2lCZNjCgWUXEnepvsA6+kNBT07ETHPYJs8JhDnRhgJjsPT8TqwqoFH
mdmTKuAPpvh5j/66Bp5BToYmC9Qx4u5Hhc+z9PBkVPZhNLTwHasvJa+tv4DT7fIK
B2pUyR7aB/xo2il97gH8d2ba6vAYPtDMbCQNVK8XtWa3/yalBBMPMTN5fhaGjnfX
0qT5yHezHSCxbzETQJcQjN977E3tjN8p8ylvDNDSpoFKgGxZVtzq47Jhr6Zkt9uO
S1fuU1ccL/yn9nYtKP5nlMxYRp+kMCKlXNEP0pWZNCoGtOYrf+yicSnU4coiQaJ0
Dp9s1iz5yHwf/2dFP6An3lgn6eikTHSmD7Unmj0PQdZ9fNaVZLsmO+12OLFgd5CC
JFj+qnmHpB/if64nRCJ5EieAR+W5exGOOXcLONU4E4TcC4rkO65D4lzi3HrJVdKs
E/IUjPmvhdHft+Kq+xT+tTIf1N9UIc1hhnrH7Jy7s4G+vYI8hsuq0Zhy9upskHi4
t91r84YRy+CScdk1B2735taf3qMv3NAjGKcqfx6EebQu8iEjzR8AdTNh/59NoqVw
4wKQ2Os7kSRq6pOJrh4Thh/cH/z6kUrYb6BjglJnLO5+jAYgnxKkJoHLqzb1rj5d
9zKUwU5p1MSmJ6oK1lEWDYKyblzkbtugTm9n3Yto/MdfQ2GbaC/Y82+rV33LUzyj
i24PVxzIa/dsD5aiudQjHWmA46AOk6z+zyHJmfZJpxpw6RebEdO8Vk/uA6jaJl1b
KaGzPAUmL00Fazucdg2T5bNPCgVTaB9Trpjdm6QdwTsdlVj7y9DkT39eAHlZZrfr
hdYhem+TjNsAlLEI+JbQUQAvq0bmnaOka4OcdZGzezw16s/vYrBSBLzQbqz3Qn3l
Z+8qZRLD2/FvCg86LB7LiAcdBUxD2nHIHzb4k6WdA2BzS4gVqB4Tz+ZhhCkJAgGB
95NV4GsMauDMg6vjP0biR1QwPDZptW0MigHhMykPUgA4/XdKUpsbTW636lcAgfF6
fLpmWRV9IYihHUCPtm48gMLUDBAWDyYmivGRSxtB/t4ErUwUxM/gA5dB1DKz0Tq7
ylQvggpVs/CGpOxbwFAXK54b2ZhyZ9g8+pfK2O5ftlrEnCSOJnYeDmq0awXk0LgM
otSXWQpsYRq+hiXpzN0kOzRuoq5jGpb1EiArvKaIlLkybohrImprsnUJwIwRPZKM
qzKEXqbKipRraakmm2hiqJ/rsMlCViuy8+bbU2kKYHKuepsWs9dLukNHhBEEvxsv
67Pi/Uik29vQG7+aQyfPVl337+uH9aTqpMoX065RhaHKXg+lyy4koMU2BaYJ9mmu
mY1EW7fMYmCiOIXE+6LozuwX+AD8V9RqK9112LuVnAg4/70IoVLeFt+BbG9SCEVp
r6oq18QbUJeBLr1ssBddgtkxfPn4tagT5gkC3GKKR70MEzAr7W3n4JyjG1cjR6Xm
iqB+YF6+3iWHEifnlADc79QXCuNVRbEhcygcSSJlUS4MRL4ZXuZa4U3qggn1sUpc
fnBr2OnqSweqhI5cqmVmRgbyGSh06CKEzYqnKN8sZdPARgTqy4Ij63N5DWMQ6Qsh
YB8Bv5ukarlYjy0trgGOpPW+PM5erdOSJS355jKOkrZqFwhvm5nDq5DGWFfYurVr
HlHWywEy+HpxfAJSTcMMk7iMjcjKQBEAal+DQbJ3MfOTlY91Ea2mvHjGUIjD6w/y
x72Y0ej/J4SoDYDhA1IGiSeAkq+omaD6WNcrVkOR/Ip8JnPtJXB99MY3OlIWkWN1
BVEMfmlmyO09fmENRY158EderTakV7EJG1TibzFg/2cdeljvqcY48c4tmM5JmW9s
1yHXFhco2dwaoXSD1pfnillCI4v6ptWNNDCJKMStXVptXlvRo8Ag/sYfqGZwZsU7
Ahw2m9aDRV+iySISha5/TxC3/y+c98s4qFsFX3W5m/izwks9Iwp/2gkVkoPnnUGh
pVsWVkCiqa3EZuPbVuIHrB0VECntdkVtcSr6hAWgt05iOQbZ0owF6+aJmXu3Ruzh
uw/ujGmySI0VmRim1Hzc7QqWfqTyjzxEnWX7OoJBGW5Pez9EXLTyrerKai5j2Ogc
hZuyUotnthr97qs11QoeW9H1gyOyhrPIKkDn7NmcxRpYgga2VMBXWx5mjHPfXP0P
AUAE8LjaCqk1epja7Q4py1cYYQZCeaFjq7pjPctjB3eMAhK4oXYclVPcRewUe1Kx
fHVvZ2DoCtpT1JCf2HNfns2sL6bAgFB+gd6n05NthGTQr7CA3d0Wz45Z7allJ59u
MzntXIjqaKMlyy2mmlmUKZJzyphRuYpsTK29EbaqTxqF5CN92ob0BtJR9ALBwhh6
9OtuYd2KutNbosGvqcjvtxaU2ye/if55DD5U9nHgXZprQ+ioezCb0ROdmMwby3eA
SkINgKfYsaYqQ/Z0Hsxo6vHhmdcxXvaoEY6cM3mkoe0ZZ1bp9zODe7ZilGFti3Q+
sU5OcuSzpfGcow42Y42EWT4R/nt0wWvKj56JCe2ZoyZ8DC51+GW8M9+o3XMb1YC+
2TDttnAHsRH33nNqvGmn5d4yW/mmXBnsGtepQp18tRNiAzXg1ApOG77+rXBl3aIU
ICsdB0a3RtB4I6hbqJxWWZyuxdH7WtIzqIOL3UocY07NuLo5Tz0mrgQwdCXB7zuf
dGVEbO46NV7qvqAG3VMzrFhJV4aqK9xGiyxhi+SHO4FMTAWPGuJTwewsVkBCncnS
3GQTzbrcZ3YJvD+eYf/EjDP27I5tZov5KlogUx6C+OQNVYJirs4hzZE1Lgezw2t5
NPidQKSujmMux/0M48hvEbu4ofvie3d8qJt7+h82/KshAYcikxbRXRvhwbeQcU/d
Fiyz6VqyaSNWRflRKSjKi5ldoPRrUYCHhY3XryKbkQtlyqAlYFDscBe3HB3SKe7E
kUAOHG+cXFql+WKXE2/shPmfw9fVjxVEgyEIBtYqgWgORi21w8GjRtxFiGc1EmSO
Xb7hq6AYnFwQOkE0ziq4dvftO0pBJrl84d4X9sUZkpghOHlvPFEvTlxKVzNzq6oZ
JItRFeczy+C40k1YGoix65yCX+QuK10P0E8+FVf+KRySLsa9rBVj2sCFIIfnKSgi
ImDRwCEF/V6ZOWw0dNxQX7KsIndjeuh3cUQIySP2yxG1GZdM8e+h/7vZQfGpbYE6
uoJs93Ied2HbGF0ZtQ03GAg4Uj8w8aE/krfMa0Jb1BJIGEw8a+z6b74qRyg+nBBh
g2XkX/vsp8aUiJZJZpU1tpCbVMuchUh0x2GJa+NbNVx/eX7r5VNZg0ENawseBnf4
YNPJZdGyb4gY4NEiOUnZGtENG/P1bbAihgYLksNFu6JCuaWwhKJ57I42WU9HMPry
t6jcgOf+fUmn2yzO/fBvNY+ccb+LXGMs3s+H0Kr/3Mhrwm0z/4zdTGw2iPwB9MNY
H0udOSyVfGX6HcAYGjObv+fc7u3459NB2K1Ycm6nxNaMXRULUMTqZpLhAzCy+Qtx
Lru6H+YVCpW/8IY8DZg1+hj/YR25XtHgGtgqKPZtVyH+fP+E3REt+Y/qh4CNeML/
pCxwAgJex3mPRRlkGR9xIfT4ExoFHKXQyGSYBQvZ8vtqzsaZZbhWbaGmDjPbTPSb
KCHai55VPaVccV18rO9w5w/SLKhpqMwDTaiXaY4EMfvOro8uOWiv9Nu147DOKOM6
aV4DZEqBQLwWyWj05KlLqV0nuCKzZ39Oguk911CVGNb9ux9n72BlZ9OijLv9zv9q
P6RQDXmzVW8zatlI2qqCusEPYohOuU1xjUhcnmJbO0TipDdabmyVXj4+FxcexGna
wW1r6oh5MTLtj8Z1h7ONK0nRfkiGkOwx0RXDumVBlgyC8Z2TMFcLA+B0fjGqDydS
g4xkxuolzNg+NI8VfCXJN39lWDV1MQqnmxcngCFYnhdN8YYPJBUc7dv6z0jRCQFQ
GP5OixJUpywPFO0f6CsaTu69Rwez5R3cvFy4w6kYTYO7+irbNBUvkLqqjBON7d5j
ETME3JGq4voeWWdZ1LRaqfGXs7b4QHBpa/p+GjokiHts8jPfjQRSduU/GqZ5r+pC
eXXrzAeGjLx4H7TwvOgUNUEyZ/9bZG5Y0BgPgw+gJkJWNj4WSr3nQk4Vv3pTOpfo
iANbh39MUtFejzrJo8IOEpbkFKTFjHwIEAS3S2NCcrFV/kS9KbWJrq2gFKLWt1l7
FjzD0c5Qgut03IVqFlpSHKcrsTfDFfUFXISt9K0z0CfgvSX6a68Mf+oltP8YWrnl
DqYIbL1pE7hR0mNzyCy1NAAsZz9BBI+r0yho6m2ODQJ2nONUU1eDa92O5l9cVVMT
eMQHpm5dBkJedIc6OxfhuGHsnZPifMA0m1aqQ1bH2UZ6IdfSqOa+gfgy8mZ+pOui
bvCvdjZBwwiXFgQAvXyxfVZsgTEJdZh97sHrKXT7YurpJB5v7V9Q7xmas+v3sA8Z
McNamcPS4pfJ+HQpACifLDyx00ObIJLGbFbdRIW3MIt+hO1IcBVtUtv8gNT01ybb
Yb4Yxwm+QWoz+fEi1xFgg9Qtm7YLH2TEUUUJpzDHGBgEuVdhmgtqDJReoMQNc041
kLWuTpRuY652ez3kj/qhCZHyPpfq9Qaf2q4JdzMcf0s4dgA2fes5SEtmtXNWHyg8
q1RNDeuvhSRYJJXKOWF9HwwLxtqTX6yISOM6x16a2GTvE5I3mZ7lg+Jr40Xddswu
IdTWToCxg4eyxYlLDyVyKjFoMGWvlGL3inHDpxUSeg4r6HSlVJ1/kRHqoMwIQMBt
9J15+RXQ0remBgnw6cGNI+NtbQqiUGgKBCiUQ7pUIZihW60uCk1/9paZPCZvESA5
X27aG+qsTK+pEovthgCLvtRoGeoB58fx6+a75sVxanp3zTE+UfbWkhprdLPjM4Nn
46rX18Ci4UZ4469Q6o8jgWzyiDY6RXYIBJtL8ah9+cj1r/5myhWNSgnul/w5GuiI
TdaqaE4M+x2LR4Gqhs/cd4x9P8MLmqxrHs44EMyF57dRBWG/dJ9Pz48kFXRCDWE+
WLDnRyfheNhfT8siioqg4Yl0CB+H07auT+tgu1lQXu8=
--pragma protect end_data_block
--pragma protect digest_block
B6zNLx+5fqQ4MdlCpvBtHUe5YxE=
--pragma protect end_digest_block
--pragma protect end_protected
