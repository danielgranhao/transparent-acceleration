-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect BEGIN_PROTECTED
`protect version = 1
`protect author = "Altera"
`protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`protect key_keyowner = "Mentor Graphics Corporation" , key_keyname = "MGC-VERIF-SIM-RSA-1" , key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 128)
`protect KEY_BLOCK
nDMyXII1N6CcrHojWTMJd/OxZ2qtnLlEUaww1qOSMhpnrkuLoJoEV4E7KBMZxOp3
rIAB1qjorhng+ITDa6WxfM+GzwEN6I+vFjQOtnmQkcGT7yh05KOkMcGP6+2VGtgh
O9VkAoUzC2hhT+Irm3igclhMatPoRodxxnIg6fBPJ64=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 64, bytes = 7201)

`protect DATA_BLOCK
8Sv9Wxv7OiUGEcDuTSDWaAuNHp1vmBrGNjZFm1vrqkcSDH3mgTAkfYnAxPKjoo7L
paKq9OwcFb3/bXaR0JEUwk0XGFJscVXkE3P5eSYaDls7q5OYcONElc/4nrMYXi2J
ifdyfR+8X0YbqXWKHHa1ZrTximQFBzjSLHJFN6maGHiWVnzZkzVgkS1AbDTjoQNr
K5509eLlggzRxPJ6raiVZRTZpRqQUUl8k34IgdhTWn1zcTQ1ZgDoudBa0jemCKMC
A66rl9Rgh/F8+m3sUVDbHPOsNn1VCF9eo6wmZQKKhJvIdsuEG3idwdYZkkkSRg43
E77oDjNe1SegZtbXOCvDYa2Rukt2shlItLqlJSFwcDIOKQ5tqcNwOJi1d2s6TRud
T1IMUlXvveB343+8whMOWQQRQJwHN5DDS/fM88FaNtGZlIZ8lLtaYP+uLjX64cq/
/pCP4UTbvPOCW9WBFSF/PuhsOtbFB5BA4P6LwdFGtlsT5pLJ7FGCQE+om8lXGTn2
eoj9d7LhWbEjDU9+dWaCOO54TKrAAZW1QYOYKjVO7sTiAnp4oMsIMliTRJE6DNhB
9LXvnZs+vrzWLZ2YEJUw3DS6HCYpj9i2Ll30H+KAdIX6FxNsRrunRQlgMCZln88p
56KGxn4IdM8U8yhfqZYB2PF57Dj5d1tpqXUpryOMKT43VeQDutXFC0N3EaFhBC6k
56/lsQqpoW9XEjfwsokmneqKvZl9+e2oOtznKn7ujTqfGmeMcPimvWseAYkp9If7
gof3/nRfkFBMxHd9vET3tADtXQoZ26Z2PnvNyl1dymfwqdJQwh/qx74MwhXUKXfY
Qf+I5GNFuo9tKkEVPd1Bmdc30P/uuZ9g+pKfSwC5U0s/hhUcGRP/D4WGiRLrRgGi
CVFOe6TytJxx0nM+Aeg1XBH3CVs75bNk8DOgG7v+1qqeEJlOoqsxm7fRagZKe//K
ZoO4eqJyQ2WwVY3xJsCcnqxrOgSX8uLZGmU4FTC8FViEC3CEYdF+l8DyFWbfTnfW
AGBAUS3CXqAN50JygquMSOskx+8WWn42cQ00gtK0aHkJlA9EgCOx/puPcnZlDKAu
s1PMuJ2gtxPPXAwsltIwjENdv3F4IiGF5o5I7qzTHg1au819WsDL+ad95f7j51WB
vtlGXkGYul87sfGpSMXK55rUdAxYajWNwYT3k9FRkkeHc5DH+N9KPpBLgSAYPp4O
izP2xQ5x+0XMAVbjg5HimoV1hKspIN+xFB3Zz/28JobWW1fMJlr1bxLP65tG5eRZ
Ug3iIj3X5RpIfEFH6T6D3b9now7Qz+4SFJg6/bp4lEFXS30wXkd3OsPZ5OoVbQiL
9ACnp3UVhm74dqx9yQCXad5C3SLo5bno+a7hP21Q4UYJ9BWSgcUdjq58kR3xHJHA
sw6omGCaHVvUw3O+aPXcslQqSJHiJV6OplavSs3OD/QneJuJB52A8RWOO5iXFJvQ
6zHv12tXX7osbDk7h/Z3NnB7xaNVEdsqNVmJ5c5ZI1ng+TQm/wz9ct5DxfLT09fH
r2Xnb7cbed4OVMN/p7chEez4uNLFUTlrOISswaGDL3qbQM7M8ZYWiXaT71jB/5SD
x6Jn9n0O7j135ESprvW1iiLbiD4u7tkr04CBat4AKCZJ9vr3N2Fndz474uqi/gob
4cuNqagPhQ8DlDa2RrpQo0UVuOKvtdEP8xuufO2P3D1dDJLloDGIBeKyAfzMVepl
CqLDDEbtUOdPMgc3jIl3LUvahJpf6BQJ66HqwQxR++Y5TL5lXbGHgkor5Kya8mOU
DxjV+cYecwBhwr0yxpxUl426p9X/qLO/ZENpsJNBhIFZTZDaOhwQsi3AE2F0hnr5
X9Dt2ZgxbmfUKOzAxZIZ0DhjvQLWgMHT6nXf9kZaXKgHonIo2PuOoTIR0DGDMMB7
WhhcCuD8RZFb7gofbII6vI/gmKBqtVbgKwNnXgcjR9wPNh8LD5Q2hSZLAPzivwQk
V1QQkQQDNRUZ5ZzGIPxdDEcC9UNfEZpISzcwZf0yhoQbNgzBmMp6M9THDFp2Vtik
0fjlEZ1JBs9PoWnX7KLfsY2sgO08v/6AGyPPsdnORbhumOBBGuEVIYfJJ1pYvVdx
T8/HdB24TZxctUBVOeWRAEWaK3wOzQBsZZvWEwFjnvNLrDFaJU8XqW0BWDEzSgBL
Bb7ld5A/aoaxy0JOGoVUp0kYpk2QFvAAvp6EJs8Tb+76Is0JCPiGwgzeTHJZ89c6
IWoO3OcDAEXl7VOzPdKj1+/xTD0GV4zAQkEAekgM4lKghFOrkcrGS2AbESzh3zmT
kwJEMz/vd0YmoDY+wO/4iUoqboxPAQeWkcl/dnk/+L4eVXGotUAtm+oa8v3or/ZW
GcMuGtNu68frn5mdfd3yZVLF8XYvsFHQjNU3u1kGDK+r07EjfpYdprMavTItN0wq
xDxDM+UWI6wduifCmZhrfTdjh6c76W9YhYKruVz7ux6EisN9S970ZJM9QoLMAsnA
GGfOz2JqtYpu4FHRJoYT6o58TsCGXBbuLaT1+5nTcH/YieBTARIqUXhjwVHbEDM4
YxB2muVRI9+Uo/JqAdiUdnwezosl9CK31+7Ct2gk6zv3/FbTxJ3zarLag1WEHHwF
C+/w+y4x7OJzALt6qB2Q0NDPsSv2Uh0tLlB+/6W/D6OI8DVQLP28mFCA8HZjb0oo
06ogLQNOgN8iRACjB+ZWw7w+ZV6U7o9XoBfErV2aA8O/8GXzfLx1/jf1Cf6HiaQg
AWkMVLSKG3Yqgxc536OI19xXH4CnM6D7loQ/o7AlfygrtS3CTi/mkLnxjDWlO3Q9
m6WucvT8dRI4hSVMtoQ5EZJzi2MSRDpH2KoADcvi5XUKm29/sUoPObzRzgdh0vSL
nER2AMwAm889iEdiLX+hsRfLlQxxWzBV8PrnOydF6aWsDwRMp8E9QGFXNNABhe91
utEhWc6Xk1GJS2nbyYaKH/E5l+BwFsandcTeonyenIJRN9HHcI3a5pZ1e9Y2BPvd
lwrFBixruVk7aLFqE2qL7lZ80nwzW0x+TXlINw95wWYjq0IPPb9blZQ85uAisfQC
nDeXOPyj6xv5pZgPkorsyOdzJdGSYriAVcPEUUslcJvg1sII6MIjSnZTPogyE53B
KA65CjPeUjkkqKetgNXjXSab7M8pSuJyWU89bgmC5RKUxsO7fnIswu1Mh0nnwG1p
BlfUcfbwcZYMXf7YP/6Yx8haMYIQHnzW1X/pQGXQ1ERnWK4UQ4qf9eZoS6lJACWv
i++pti8RhgigXVNVgSN1sh3BT6W3cElq4JSb+tuvF1gyrVbgXQa18J2fQrEC7yS+
G1bJxrd7NeiPOWyr+smDdngOM0pre8EVd5TEjvv1njbA6jfOgfw+vUo2790H3HKL
Xm/2N7WKpeMb5ZWdWEkU1t7vuwXgMhWIk0d1JgWZ71oNSD627b8V/VQ/c8hpnURO
CvC8A6fsu++lRddVS3QCMYfNq3BuQdiu9FQDZRwOtJOT7jwcCvrhndSpLHBvV+Is
EAsktDpiJ+0hpz29WFcdQkfL4GuR+j6O3PxD8nbaZCVfTK8sYUuBZg1gvX651A58
jpR1beKgInKkbzc/3y+1Akl6vtR5ooWJDitz6DIpYXKxBAyO9SaCMJ7xGHokY2Ti
3dkwrEm/PicWR6s8R5tBNpJgIUYYePrAdUTDZNxww5JEoY5YRMV63y7TBPost6Ca
YT5rBMex5ia7r8dmfNz6xPDUGlccp/kmJ2zJEMt+4RLYXc46FqdXbsV6RpCyF2is
C9qeKfx29O8z3IIhP83egYSxvQpX54Y1g7fR0UQeDrTNmw1ohwWmsAdrQztONREW
1QghBuxnNGqeip/D//fp/3y596IkfHwTqtEIfVI1R8kja464ukIieWxo8rzlj7ZI
rk59UaITHkIuZwyAy3mTGZSsrdRV33OiB/RYGYGJMQTWZayFiw+U4Get86hBO1KR
i7w+5HIRltMIag3KnmFs5EBx4NViL710vImTM0xOpTO9mhqv4slp6ZToMrbLpWdk
tbKYWKPjSYaqaLZcWt16gqu8HDbHLDTMaM9cDfidfsLLyajeCuBacsvJFfTV83K/
hkLaR9UpD/KjINUqrKs7ar10Itq+bOPlafJoBtTkyBB277NhlxRbnnDxtLUWRLTu
zHV4fbw7iCr9hwqI5YImRm9NwLh5E9QWNFhTyGgwOmuGK2CZNJhK4QdjELXxIWnH
7Pa7D0NXSWFl33LFDqwkOCaKzShi3oCyGC8QmcAk6cB5z/NWaJReXlDs5ZjEkUzd
zSbx6+e4HPWjeK2WIvQ+zneLrHQYe3OKNX+FygM7eA1/h+LgAL2/SC6d9grOYdMn
Nl0XvoczDjOIlwyT9TV2YQWsNiij7NybI6OHNwwvqRmgrB7WoqXYHDl7sBRHudyE
oqfwxXDDat+02Qjwxscg3dFXv6/Kg+t8ffHEL6lHxP8SHmnmfe9eHJ1200/560hD
kKmMKBvgUAYUL7e6zHwGecWtZBsDYG4VgRtM8Dyc+FU7hSDHetXU1B64fAONll+Z
Tkqrbn99r5nIL9NdRoAf5yo2qysP8MWxNryYNXXIvZsO0clnxOdf7FOpFb5+bDCe
IkyHk0BnwL4DybIWQF4KJHy6q26a2oWt9rF0AWnHR/lJmOATmoBwAuZI3gQ8yn2M
lGP5gGZ9MCqLZXH+6VtwS5M33tGxL72YS76Q6qKGH2FKQt6NAvdgndnyXH+yKu7t
Dzc/WxzmwPGHCQmX2tjnWbomUEKit0tFifZyBUyFDqM06rUxjj6GbLC5er50ZWjB
TdHUBmJZ1Z7ZZhgPZa1UBo/zV+rCzKcY3s8GpRden4oz0HohJIz2ihSuJQqzrRay
6LzsdUuJmRQzER965JtmSfRJxfVjFrr1KC5l1nwjJxUpZnKs/ftaW/afwv/K55RO
V+2BTakFkgzs7WHTvYeCYK0Ukmb8ermbAbesrWSnBsV9OZq44PKeZyAFKP7qVi7e
8GwSwuBW014jCoqaJiJmCuKj77rd4+3U7xWhBxn4lBBcjjovF32AggBzauqh9L2Z
n8MvhyCYEVVlJGQ5viqLZWkcb5vMJucqbVn3cI8xLd3M/2+lUSpuGSOwvDk6wMnd
1MpSaPuht3rxoucuRRrtQqgtOOexvJS4a7SaokhMlYjdLYVCqk9ghmyfKrLFO8wU
YsrebdmVr+0S59Hmi+DMLaLV9mwSXWNS4NPGnQJyHmdQm0RtuDSei2DZRto+dziP
4tjqo3kLeR53AFcOmbxTARlVa3bouHAb+DDZCDnbN4JHgJt15UFHhRMbF7Q8gTNY
bm8bWTQWu7xjCo8nZU4ZW+xOqC2de+8kMgKGGINfVr5m1QzVAOoibr+0McHIFA86
t9UNGN2i34/TvIJl2jfQGh/QTz1Kk8/8Fq92Za/4TQDUAL7ijWo/KiWBUIkY4Yau
5sGa4VcoQFULNkd9t6R6fu5IGeSOx2lXww4/FPz55C7gGzlhwIKcUIDnp8Og0Zqo
KTF+uDa5qXNJFQjDowKB1sp6gwkoEhqn12CUQXYTb+P9oPCbuxeAhUVbaQloUgev
XbvMM5VGoiVh7ch23ijbH4BREx42Ft9+d7MO5jEwmSoR+JJc7SvV+jAd/Go3WVy6
s0gci5Vq7aJGahOuHaYq7cA60Tza7rsTB5hTzeYMKtk+81efHHng/IKOu57lG4oS
ZkTI4hpMf2G4FTqxPQqHcfrWM+yF9xu8OEIAfPI1wvFt2GVxpLHfjkG8EmTwcUgp
uySAcFGpOlsuE3TjnOubZt9EMdijDf3JX5B0jAUm9Bs9mMvWQeVPAp8ZnDfxRcv9
nAOOC4kbBTEQW9chV5Ljx1zaqzNbIKqSd/+f7eSOOdmJTK3LVF+7NmcTmOdvXoPj
6JvoDXhALMx6DwsIpkeYTn9nN+NNmCd+GqHjLLjtu6tldRkOFvWrlIusfv5U6iQH
v65p3iuQRigbrLUVry5Q0y0yeVcEWvulD86PgsepMy+EqxYWIfd+GflvDaDAJWNO
kwalk/yRHVhiREqdH7Evhe9miyPMCARMGQpLHgrktNq6jjwFDkuU6cJ0O3Rodpnt
o7i6JJasICuyHEVvu24sZI2H5mckI/YixF1CdUX8nxC5295CA/xkRZ0C19AACtMv
UeAtZU8HP1sGMRqad0SXY6yAyGnLVRw35IRKYgvxrNGFcIeHyb9A4+uE1to38y1p
nc4w0/WVHDvIGWly6yCwG+Z1SDRzpQLZ8pzGGZe8X73FhCQery+VItW8EeigJiPI
uJBZ991Ehfvj676e83/EurWNoq8jBDfwSTBQKahtbAWjp2z/SHSwrSdZHKoKIi2j
88zaHOy65l2b5nmGLln73Zmvq1lpHmlIiOrGTd7sxRKSKTG95xYwTF2o45MUGMCi
YMt1R96HoMIM1qTqDTiOfW25gwggyEecPljshIyWoCFy5OuXSWp7VW9ojQ1HsZx+
qLArxtn8WZ7vdIWtK5k1lSpfNTLiN6ejiHUgt9mRyrXLqEDVp+SVFMjFVpskTCWy
Bw4ERtW5ejIQiHb1YbR1s1LHil4l2CjpxTeEC0/eyxcrBbI35+iAfpPHneXmG/B2
eDeer1FUKxBSQnkyBdr/OpkbIOzOG7PFZMYdDbJm80WPw6qUg0CLUB5OTNgYhuvY
8gegRsfwSoTrRutd8e2tdryxzoH5xCKxZbD514Ns2EIfzy5JM7U3JXYx0wLS4O5w
LKkBeiXNEIUosYi4orXgq6BRXa2aF16zYBYA5vrOJfVPJJVJ441nTdzNTlHxQTnx
X+mkHY8WUo5DDG2o0qZQEZ0mxrxbKT8ad7w45txoxdHzDcwedeaQ/zO3qEa69KVm
dUnMwPSHfBEvxFyTTUBJadZ4MsTAOC0tFcYUCaKuZt6rhnlMZQdyiUHR9O5OYN5V
xOLvazglYXljW9ILdjAd4mWS+240Na/ov85Iu7r/b6kCZismDByh1p1WctUpeFlJ
5iJ9ryfJBvdci7f0Csco9j+UBOh3nXd0xPEQgKJb24x2a/cODzxwEI28J0Ffh5Qy
+y3053eNOcmLAnLTQVF4WQfP/O9TN61fxbVdjjlwcERlXFm+wDNRDrR0JNncyefs
nruku+DW1I+wfSHAZH1CHfkmzrYvdGcyRFoBhuHNyx8u06oN/pcoxZYgcgm9xTqT
CXBzNM8Wk/FYPhwhGXJHS/15PV3UhO8YZPU3hCK69wNvzKMU9AAL3SRztpExvCJw
eePIdnjVGY22/YQo6a6p75Evi/DHxu5E8Vv+PYrweGDT30qpDZMUw9M7t6ZitYjC
m2DGgBNlyjNrHe6eGca9rMex7ibksNPima29lzk8pl2MckVJhoMuBLgFSJNcX3uc
AWYBPhx4Aci3emSyxcyjveXDXcQKuv1JKgS/bnkuDAE0/YXgZ/e6z6FEjyYdMvyu
OWT71J3luyW/EmYBDmtjssWRtm+0HkcCCqKbIMS7AetHKBNZatyPND5WHBfs4+xo
0YYpepZLlZKDu46qa7g/eXYk7jMiAjcw012xtLyHYwPXbgjzEf1vbgmsdmceYPk1
MpMEZN/xBJFBEeAfGkU+JpviiHw5TJAM7c4o+iONbrsarrCjcbf8GIzIZtpQnWXq
vbGE6iZ7vhngdRXG8cytzi0LbUN8K7Exe1/B3i9gYYbFpH9u1HGWzBiarW8z3/kX
s6CRhv4zWf2f185dz1ng2N8AQU4hP4drKgHtDTt/2qxSumyiLup70xhx4dyTrGyr
WI71iQhifm9wENxYdhcDrhH6Unzm34WXzBGx9O7uh3pKP4Vl1h2NHeeIXIjGPxDW
h7kk+zy/TXc7cNCbjCMB4WmVxG1gvAgXQv3kZCpVcy2Eg9OdtNK3v/KgSQ8C3+Ur
b7azd5uSgtjkiwPTXO9chefeSb4szx6sEdxddPnzVhwnRFszHCKesbl2PlloVcPv
ssyE8gj9VlBoE6ftLYEi52XB2OMlSx4KNAaRIdEfOytc1s8Xc1VYWKdAOah++iDL
bb8vpqSaHGj8zrLx778xDUhaa5rdn4ExRKNsiHF2DADOFMWrBiJoRWPHtgflKmyR
HHtgwbbq/pi2rIoCe/95ZW5C+is3Kjwv2G8GYL9fbbBHEfYixzovEuna4CwajnSx
cyH1ZmQX4dL2RCJTWDeqZcRK5/vV3AbOPXl2iAaME57oEZVqs4AlFz/GhFTbUgq4
tfLYc77/w8c0RO7EYqh0b2EQr7WVY608OpDKTpU2WeG4fOCr73XnzlqWZAl5wDPm
MUKVMchptT/edt5yjYE3u8id4SVYp1NkkFldY1TKS+Z8mLxueOmkB/tIAVobssdK
ECf4uHu+HiBH4/mqU+zyw4OziYI6XNksRh9oWlLc6/92pZ1r3m0e34z5P437lHEN
FgoM7519XnDMeV8XOYaH5ilyv82p1M0FPP9ZL7EpdNXe/CzQrNiS6m8XwNBOFdPF
EDJJIv50vXVi9zT//Gc6D+N4U8cJQV0who2cxsiGx7zj4kjyFeikpFjAVZqcaYwl
JU5CNBipEyAO+zxQ9PJ+0Qv00+N6mxJyujGD2z7IhzzsR3cteu6z0zPD0x38L+qe
mTm7PFpV7Z1oon3RLareXdssWSY9RuMC7+fr5y/lxe1Ugj5EVFi1xKrCiCHqZz86
t8yyVhwNlPIkWDE9K6GSMNrhvdUqsyKbEWWRgjl8K+KheQQkuj93MzZ/ZAtj1b+P
cOZzTWaDJz2iSO86FLjcoPVsSE2ErNK0quWPwRlMdde7Dqx6J8lS+VZiBUDBUbcT
BAEwG8c/dEyJ8MCj6nG/CS1XuxPzUkUVuhPzZRxn2O+0AAUUboiXYAWa2ktV339b
YsFQ91Nud+0U+KVpR9emZxG8L8UmS+KEXYB+QfyeKyGYasOBM2yyra/ZL0Kg8CgX
q1jaTl/ho3+ZX4bX6Nx2DWb5DnucHxvW2G+OqUzDyo/jbbN/Y3uBdjtj7LmpaqyX
cLmAhH0uxWOxWl+QTwoes+UF6v1dpAcW1JghpvH4PDBky2IQ1Nq+5Xg/vMdzdyYe
GbrjQNfg8ygXh+qQrAJRRoaeiM3HFJmLKyPgAKPllYnorvF9ONOfGnNxfcCLUHbN
5Z/6nMhU/kuuqsimiV8xAlnOaE8eKPW3fwCZMx+qdycyeLsarqsb7Ak3IvoHvits
VDT7MNGZRrrqnYikMGL+EXW0xn2FOOv12FKsVU+ABfkdg0vkxIS9WkxOsEkJkjje
MWPeSixYNxuxSK0tUry3BhkdyrGGQmCIwGCOv1M4DlinQctro6lka2pKx2s1mCTZ
wC55hsTh3Hm6KJIvaGhfHGB02EMVFOCA5lIuxcOM4TfxZT7NWCw6gHJpusUw/AHJ
M5y50dWi+Hwe4lLczTTYx/DhMru65d6FRB/YZqBp266isWisGOo+LU42Zx1H3UVc
JDBaJwugpVqI2MmtPkeZZ/x+sJhkoWACfdpOTsw9dwifux5ED9RWOVwSbmAvO18E
LwFSJ5v+QwSIkC4tkxNOJCL8EN7gahitfSYr1MvZ1551rFwudZXCRUtsgzVNR90r
jV1RQ15Qq7HExO9IO1Wmnq2T16PfXZOlli7Wf/QA2bvNMGp0xUAfRCZWxA72NCvr
QOaxKkqTLQeU8F2Tuf+G1/kW/mr179do+eh9YPbQW+U=
`protect END_PROTECTED