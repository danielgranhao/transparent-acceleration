-- (C) 2001-2016 Altera Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Altera and is being provided
-- in accordance with and subject to the protections of the
-- applicable Altera Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Altera
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Altera Program License Subscription
-- Agreement, Altera MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Altera and sold
-- by Altera or its authorized distributors. Please refer to the
-- applicable agreement for further details. Altera products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Altera assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.0
`protect begin_protected
`protect version = 1
`protect encrypt_agent = "VCS"
`protect encrypt_agent_info = "J-2014.12-SP1 -- Feb 26, 2015"
`protect key_keyowner = "Synopsys"
`protect key_keyname = "SNPS-VCS-RSA-1"
`protect key_method = "rsa"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 128)
`protect key_block
l+3tm4o5lp2PzC2i/UtNk3OSNd8vxK0Vu0gEqQWurm3BcrCz5afvR5wdfxZkblEn
1G6iVl9wb5/yiCICOvHj75VuUMfUNt8Y38j8IMwNKHIGIWvAVuxA/UaiYaZmobI0
FWOS/txT2J0Edr2sBsuYu4Aji5EL8HFD5o2cnAmHtaQ=
`protect data_method = "aes128-cbc"
`protect encoding = (enctype = "base64", line_length = 76, bytes = 20608)
`protect data_block
r1DCnL3SsWcKwOBAkteDoN7k+36tl6Zh71T9ZbREM1iIa8Ltdw/ug8PeYooJc9+q
eExSRHlVuE1pFWS+kE7sIfqcC/gNnlwQqRc0W640+UraaQv2LdGbJ2eCvcTvh2f4
eGcgQrNte5bL+RG2amwZ7CvGY6FQ8pGeAcqpi9PWNywzAPh3wjrWj8z4lyVRYMnP
r+Gke6SyruJWOo8WatomakGPbN8h6RNQSaERAcOdMAjRSea2VeKbzzTT5qr6z7Ws
3E404dW3rSPwrAYjoDVHDXpu+MHi1F/Ekuc8DuYKeluLINEhtw+fD/Qapa/N8MJN
P0bMSYSqT+BKp4dDGJce2bR4xjJjnbsJrTJqKfUjzZysnRK/KUWWfp5FTJ4gcKCQ
hFzLzNhwkHzNaiQoM71K9xs9BFoJWi8lAf2R5QKVwHHipqNhhIB9+3UWqx26kdk6
ivKqEDgV+gocQqZ24RT9jNC+JP37L4+7qAkqsVaN2JK/qlIGg7UULO3Pbe6aPlib
K1Gm9OICdXDeRwY/L/qs1a8KYeXK1Hi0iJjDPDQJ0g292cEw+XZPBsMvzTe0Hf+j
bYoG+v+Tst7D5suy4kLbcRFDeUjTQqeq6oCfw5ziikf7s3XlKn/HC7iSYqDDomrd
38Cu9I5uryPpZHRcYohWyyAVqPoyNrKWmhxCWzt4MqKx2yoA0lMWUcGQUzC2zHVc
KA74k/BmP4DthUz1dZHPLAWFe0bDzdYWJkGUSE1l1GFOwawDx0Psdnxwe6ghb9vx
joMK7P1KEPMhqO8yzislnB/T2nBrknxxZDWvc2OW4QjFQDSBaDegu/Eh/gZmAq9f
dGti4Mmvnz1wyKvWPytSSbbHmynysULpLOUUv+m4grh/Lt6OKfg3Aq0i/cDA355B
pYIfh3/LzenmeeKacYwMOJGI8B5gjc5t0kGorPFQaP51XzG/MTIhdDtm/S+AEeDv
txtoeOvcmCiHHKGBHlmiXnyEQW+UifYC9lSODgK9j+whOfN3sqK9YHJ7fUBLWbZi
B2tej3u+aQi++FToDN5szNdERKYLe+Aehq1Ife3tJzjW8bUH/bg0J1gFPSAwJgCg
otXv0L+12iZhwYte67E/laIurYN6RHIp+HBVkaGcYcfgfU0x0e/Gjn0VJx4PZAQw
4iq4GDQ/qgBet0DSpIiU71Fos91sb/GRhI+924EUWxG6fmoBRPFIMwLD35NO7ZNZ
Fi25HiTs0/6uXF/Y3AhbxNmXqeBHX67rKHU1fA4g7nFtujvwKsZZcvT3Fh/oI5Gz
UyM3JI1jFKV4TZfLJEA+kdm+orA7r99empJx96nwzXaf92xqyRuPHpgMa761xgnr
iOGDoC+6YYJtX/sAaTsOxwGuPTnyrTZ+2w2LjmJV1JipzGuAFc2BHUL5kQ4DXqRY
CdC7ApR6IjFpdg0EIcwNTSSdywBnuLtQuPQOrQA0sVeaLEgluVVfBfpDUxoWVILZ
4DH5T0HCNF1WQ2ZJNyJz3ZlLNns8g/Z0ABzRSkoBsTx9OgDqCyBDp86l6oIHuriD
2BPKzMXlOB49tnXJYSIewCRxmb6pgIV9zJqkgDaiDcfJVA98nn2De35esmQrpQjc
O5AqUr/TtaaCCYFDbjS6enjZAmssPI0Sc3bSpcf/sFYLUalqLCwljxAPew4tkZyY
lw+E/KbRFdh7Ul54uTX1+hg2D2usWdk34ARur7ybDmP6KBLa4mOV+hrOdo9w/jC/
wanPsUFFdj1Vero/FFRbRfz15KmGCEEMFEnt9FM2bvyzgXRyyPNo6ahwQXjyqvr2
UALQpu5wHdGup6WjYwQ3NaMcPh42vWjMIQ54yzp8f3TtqBPxnsuRGk/gJ1Qa/4eM
8zhwqtPV30glkffHG5jexmpiUsB9qiQ2P6pwAcA7VFGXTcGsRrx3a7w1odhFPQpl
2i//4aH+mw3nwPoqskgbtCcI7XbNDIbXnBcLzt+0NnArWPiWxUcZ2GlcXgk8UacX
K6qS2X0hugteGd5DjN12/fuZjCrQCGVhahZnrFIEz6We8SFCnihgPCBNSrnKyA5c
7EYcJkCD66CqUheSZ76dfOtD2B9qIJksVYnyiW/+6MgjEk3Zoh1huAjAiAqxPQfh
dHE6nHTisWdhqh2F4V1CQHXI1h14rm53DT9PZ12NQov2Xxn8SaMoyb4PPnNJmQIu
0sxulY2QOmQMh9SEQHU3olOilWywRpxN/yLny5JFlTwNu1t8Jjmfw6uNQooSaLo9
TE+JvVObAd1Ynd6IKNgoLNdRKVPSc6rTDYZG3bDHxZBxnImRebxRrXrH0G1/r4B4
JsqiyZ5OerORb8c0tArGzQ/QoKcJZa83AQ/dUZTK84wnegqqL7XdCxm8WU47Srhl
aYZ8mdtZSTAYuQjjCnsvVO7x0FBAI8GAeBrRuuRvyL1VQ+tC3P3t3gRZxkU2NwFt
qAQXdSGo8MiwC3bpKgi7C3Txeb5LqicNFmyMtDQl0GUomXjQSeFKjwt1DVMKiDOa
Uap32gIdyQ8GUybVzUDBCX+ph1ggJ2MkN0q1L2qd7E/h+1e0uanlojrCeAZetwoj
Kg3OR3SFCVK4cZ0XjVgvJGnI4Dv4GVHkEIJzID+vc31T7oIXjFfc8AzSYbBz0EcY
gbDgYidY+F2llYqxVdNRuXH/0M3/MLBbBFAoXpmVKVHytSWMqz0cVRnrbMRwDfXs
yFgl+yXL6qQpjmtFWWZrBL1k9t49Tg0w2SbUIGhAAzsTjZWmNCbVr/A+JibDJfmY
QumM0nFn8PHUMsh0RAzbTSG5ckir+KldbOVUL7ctY5Bl5iP9zdxqBtbjIh7EfAjv
tjCwdxQ0TDMVv5Mg0NtAI8c+cVQjxbCHbbHaf1L79mg5k02VsJD6EbOyWUGg0CRx
yQ+1EjTm2fFROr767aCgKfGrrs2GKBQVMn5CBdHchK/m6RbIISLTvI6N5wvPwgmX
ywKLogYtqQvsLiwScI3ZSk/GPeO2MYBCOaKNSMx8kjC8MOsOvI0hh8+exaezwIEq
dCxZ71Q0xiQew7emy6CUsDYOSIquAvyH/q0SwILkE4luaxuveEfxopKhvZTSX+ra
4oPfZdGswihCNcG6jgKoT7tE2sM5od7vrV/jOK1bdtwU+Sqj7V3IUle06UlBlGsU
Na1ihdOkwnCTgjTuZ+dvEbXi/LsD3vbEiPb1hwflMqC7OKvWY6SpTToU+XXEIofb
kLbH3ZsABhYX4Kt1CjKhdpeh5SFOoKPxNfPgrgJvgnGa0cJskNAK1+3M3Wyp9Sz7
L2vR6I5oJy1CGZThHxasEbMm78Nxua43hKe+Ud+Ebt71Ld+R973U+hqODClfYikj
X0AR96GpeEXeu1vHaiZwSKfdtu+7c2YM1wJZJpkej+O5sKtnTbnrc8M0Ar2LsCS0
AIAYmMnytsEQPtK5RGcV1BqAN2e7YpOF3ojAnX1u1nSfG3pgUmga4QBRiOUC7N98
5KnvjXvZChSbjONVXFnKQKP90d5ZtKuM3Zj4iDl7w7dm1TU3dpFpOExEmax/kciK
MyzJVRfxN60UEjOOtkYLHha1CRo/cKViJdm6IZDBTjC3gVDjw8QdGnzdBQws419E
SmweEjogfXPWQLenbDqkS0Ijmu57UNsXLAEj7l6ZRHFNnO6o6v+uwO7JodRBiVgQ
TTn1u4/Pzuzl/SEp3Hgegk5M7mMxEbs+XJOGSAM68exzdFX2FCY1H/YApojkE+oL
Vz+k5A6I4ibKZnBlSFOipBMdzlqkZmgen6Gz4LQGXjceIrUHGlRhikLsQ+4/MCtc
eLkgrg5FyMnGGKFNRo4mUE60bpMbIOyPAgLLkkw8tQwMwDmUbVpBRp7i44aVVX5l
SQO1e6KLIJTzECD8Zgc7TIqPyeMTFyWnLe/nV2GTfdfVSRhShEJqpYniMtAq0xRc
CJcoYeCI14SAWGUq0LdtcRPPcaRlCVNsuSIJ1QB5K7pVsWmsWAsIpDQl5AhsrHs2
8iFvmn/xMDgavKpc7J9tVJbltwFiJKO9m21DnLbWWI9mao/fj0wbDa4MBv1c5qLU
Rt6vUCv8YgbnILqX+dNN5cYEKxFZVL61zh6waSJb9sg/WDTusuePKyrbEbza3Ih4
uq42GPI3wI1Lq1q1CfiFXy8MgVmx8y+pUUako4KHZFGH9QrF1i6KJHH6Eo1EG9gM
sTanWHCnYY5ZjrboKQCMIyTCIvDBeazV1MHa5P3HE6B+UrfoDGBiclP4tJ1LEUtU
7jWJ/LSFg+oCdps1m+c0dYjbyLcYvtpaHnPdjupZh4WOhy2nRwyj/NJyufNfoRQq
+JftHxxY/NpQLqM0wOD5scizhMNCLfO30f+X28e3p3TxlRIwyFLeJQuoixL5SCEI
grOC86mwK3TeAYAQzsjOWaUpkf7nmmzRukcj3vT3XIrnkqW6hrNfLWD+cQYNez8B
55ZMNDMrsFK7nPJxt2wXTFoTsyOzWyHCHQgEhJErJ1ypkWfBZ26xkV9JYWlb4fO2
nbpqNDnWdr6FoXe02/rVjC9paHfVIeZ5ezVKUeu0OTqGEnazZPG300lT+XAtXUk3
2wJvWRoVenVeXCDdxhdjepKC+H9tQukKFjjCwWy8uLCXZ3Dex3ypSLITy6hd4HsW
RyHn+pcF9D79R73OW8WcUcMdASEwdgBhzdBxJNElxtm3x1fL980OPPJ/KuLao3A9
PW/GPNZEoCKFVAFvGzKofLkxqygAmwoBK9CrMNqDXWQPQnnXavAfq9I+OB9Kp2cp
IJPvx3n60Vy/PkQcCPPeIm3u3ztP+TQMqo/mgvEoTLN8GrDiT4tLy61/02kwe+Q+
D99kEgjMu8jg8m07KmppNCRJB+p8+NGanOU7DInXUIzTzz8whHKLBrb40OpEupaW
IbUNjPK1Wizwzw5/y/OetCc9tD4OclmuyGpIuFDDNyJyhyAVdxcuJMYVZbipifEu
a+suuUqP8MmmGHkNA1bGvdWeCC6Deauf2P4lFvyZOZgOzJy7rN4NhZK6xj/odeIB
OwPqWInBr6vlAQOrPY1qg9g4Z+nOFEyPHJ2T64kqGbxEnZr8xfF59ipfmeYJjbwo
crz8biSCfDtTfYbW+0y49e35YpsURmCILBn761/vw+4qe7wh436SzlAeM/yj5l2r
B0P4sr+a4Oc0DLOM/yeAjVaszGkMD/0D6soNgdMlXtezEROjSGKScL1ddizFbWKI
VwP8rGKPv9xraZwd3tqcQVfc0mEfcYMQRbsRpJpstE2XV2OZeDKcITFJr19G0VOg
PqXMFEtBiBGGIukQ/j/Mo3kC7RPZSkHn2PtTMckhvhf6Vy4O2SWwTHlKH7Axlbzw
/7v1Vd4DkAIng2WPLdF6/UIRIHzwaRScxMn8t5vDFOqjzlQe49niKSk+Z2mK5vMW
61oP46sPEyVHL0xyZNU6tjRsJLU7/yZMb4eB3dXvFNq4AlQJTkOPGkKzqZZY2d97
cq9Hg0X9vZls2OBFDF28JgCk9e1UxeU/JdNcf/9cmsxNA4vWnNIQ8L/nh+0UW549
zHEBqj2XWmw5tc+AIikfiXbYVNVmIIMpFr9BoTaLA2fkSdsIJ4GVUT/x80LXubD0
aeMxw+stLqxguhh/UD+HtNMfYGzXMwqqobhFOtr3sSEOzbRu9SoXoe66BZKeM2kZ
JTb+5TCLIVADpYrvGB71+ODIB6wQ9B3U6i1uOSNPLhuGkB3XzbH9cKu1f352vtEG
AstDAUVDeyJIdvkzwpOWl4x+2Ci6UkvdO0pHJevKMAmy2pRMjNV8EjrCrUsOrY8G
yawB88QKCX3gM8CjYsiVRbVBECjSxY4LUFliIyiPW7vr8M21TSsgw3yo/nTBRG6q
wpEw8iaJSzYFw/eQ5u2k59cEyip7ecqKeSB01kW+q/4/4AmfJBMBnycMoc0/mzEA
N+utPpwIquS4LDUGKcTAIfMMwL1+EcalUnPjJ+xEPTQYYKlfDf0D8wcSVRB1ebmG
IaBSRUDAKqkQBhoX/Z94Z5HIVIoi9vjlmC9lYIvZzREvfZAkgPGn8dC7e0dC5o7+
6UrOzZoH7RSuj20MBshn7e+p/LT35xiqAn/aVb9roQ7WX2FFxOyAvn7eg6VSCOej
d0kDVIDTb7wvQB36DnGpO1kZxMUi9xMi9rkqc+e1y9z6Ptvc7IawkcXFm2f8XeG7
3eO2FUjGWXBBaBTVlATwPaIilqw1UroKfYcx8jtT72pHd8PbqKuRjSYq+NC1Yzdo
leFJ7z5YjI7oMlQOLsK1gnV8zuzyu1eM9pe8TTOf190MCsTnB5Gn3JHk0eVdtn1m
bSy5b2I/RHOSuOjA6PUFzRSkQOiyjVtd4wZF5uG3N2KOODF3/6aKfPFbOP79ubUu
jhz8KjC57fEukcNVVjrNFuC9pZM8Ej+8+3DJXAE68UauASRu0g8R8NZ2S2scBBr8
mjSx3d/9M2tRervWTQ+gGxqth2LKDsFtQqnHHD/Ir3zU1sU/kmYpd3UYRU/4NnXa
btQTn3odQTDu0TXUE2zqjkvcFV7iRLanPMi/H3D/dnJW0oqAuZL3B9h5MBPMxpPP
FJ90v2lN9h9Tj6JIYLvGWCtQxGK6l7xP5CfKwsZ9QnhbrH/dCu5oqEq5R2VP86lj
GTscTQYmzo8ro2MDIY28nk1XQUmTEAAjvejhF7geIk+/n+z8sc8G4tJC3bXwVWi9
WxQ4R+J63Bo+zJm6d8/7Q4WUPTwcSSPQzVI4g8bpoVFy+nw1/Dnqgg1R80aGlBHn
uGJA8G04DYQ+yDlNNLQokFWCh6VHmFTY/FU0GfeNPMStShQWqbKlbGd6KSB0A9DK
BoygNTgxIdrO0XdzjXtHfZd39jdCpJ+klluTUZCA9bsNpc4S84gzxeQsZSy9wxvx
U7QnCQ29G70taCOE2hQvDECfLg5S4AzhbebhIqo7ogM3jgCbYnte1hL6yikHu73J
Kgg76/QzqIxbHiQ42+/e0rER53rdYkpEgoRO8QnOINhFKrWwhoZca6VWxMiU/C2t
kE2c6Blv8iAP1tnkN871URHpVHtKYdvQtjVv4h6pkNdaE7pYSXRwSpWtLJxiFut3
sHq8FGCQRh3opO4AjZ6fVd/DScJvqfdJr2TLImFoE6cEAoa7Ln4WkuxAWx6D1MJE
Bdyn06JZeRhkOYxN9DBLyaHRCtiDPH89bLiWvvV3ihkAtxPw2a7jU/eZgcikwEeB
WnllzwQUEM8giP+sTWQeeR5V4Z7gffjVb9Mq8LxBEpgcjilkJF8DzBNyMrNYFodp
C9Yce4ApmgjnXny70d8htxMrt7ZMuZQHDOBsasLRUZ1lFSsSCvddo/Q3acwsiIn4
C9fzyE8b5g08HgWJLziidsvgAdfyoxagG6+3JMZWAUG5yaPqOnRuu59Fhc8HiVsE
narVSejImjIMJYtXI4FRflldm0a3r1FI6C4f6xTLhqXx4rQBkSMA/h8cv8ECMYXj
XYcWbBYt9cQCxBp7kreHp2DB4KVOw+w2lKqJqjRL+Sr/MiryXc93mSV8aGx9D4NT
QxWvCHaSrg5z+TkOVKtJxB7OMMSSB1GiJY/tky/8uxVkRwolNr0wH0lEgp9Tl6hC
g42VIgjYXt0JEUKt5U1KupHhCfo+nZLEDFycQ8Nu/uUmf12QiW56/bCDUOSeN859
AAuZWQQSlGAfKy+O3ENNTpglNfkTxWzoLAXjU9xntVtq8YrFVC2mTOGVdZ/JO+6Y
TEpiGGjupdRGivqINFKsEC0iIv0k5Q72YO4GU0cgl07PTHr/jhanbh10WqaHLoxa
A5z8WZ4LtULCxjOFWEaAa9AN2oWvWF6RkNs3vf4Y/U+nIRC+ljvBwgW6HghHhMBM
Vr4wKd0CSc9fP1Smq2ouAC1k27RbFzuq0gfsrkJ5U3P9i/ey+JNDMm7aZ2fY1xfd
zzOX8rXUz71WJeGCXpQUlravxDlzurQEMgiUhIIiSE6k1cUQa69F6PnnK4kbnXdr
PsETpXoBpHTr89pgm8yZjSHPA4g6WC+Tq/d0urP1fjlPr4HihqL3aNBR7X3zTobi
iSewtU2HRHuh0Rgj7FOnzshb2ZtnEWZSEodYZCIWHiEd+5s0/7LKcfLnkG7qsF1C
SzAR4dI5qyksBzMfGtTZOXNbJSIqXEZu37m7BWxpSUQ5OrTrioVvCNzMXJO/Bf+r
PAh7q5rWYaji7MvBjFYeaiHtd9JZse9aW3nL7jnz6zdVzftWe8EuKWrk44WXvTpv
sqk0qIWjLvVAmxZ1jfekGuTiqOs/vpkUPYg7G7Qekr1Q/gr97BCFHwJ3HNnCmKC1
hEG5nBpb4z5u2bAcmoCBC/y1YT2A/kt3oM/USU0DFRbnlae8nLRUXEHs2PZP8mDl
dqW7R4ALpEZOIGewCWIsnOQaldrdPQCLvIks3o0NDJnjC5KF7nu0s5lOWzoXvJrv
rL/sIVDspNhiQcEZBDLA5WSBUV2dcWMn/94lvnjfjeTq8f9E470YtCWn2EHwktk1
PLWOHFrj8CNKMBJXDodrZq+83wFU8Z8mEZ7JV4/xwpDmGzPdoM1QEgsxZbHvax53
rI4yCZuXOk3GXZc66dbdXMtYd51tDx/GDze/lJK1Yhz37zNxPABFGnQ2OcM3/YuT
1ONlwo2UpshmGsTp4wDJxmCtpAI5fClYsasSB/Rmlbu+WsMO9+eqvSnNJTiiGg2a
QDHIPAGjHKmZbtYX20NVNpceylZEHvvW4v/t+vdtN9ipPExuYPQ85V/yxX40qlIz
6vHcRjartx4PHA8utSF6NfySiD2aLaREmC6JE1J7ZZpxDust2Oqxptrh++9Vx4r1
Buq5T4BD0jQLM7NQuQyjY+eUDYSLNiY8vFshkJJgmtZUMatUha+JydM+JBT0Tojb
hWXyIw76MMZPFUda8Rjbdt5ViDgIYNjrBU3g1253LqVlKZShKvIyVH+OrvlZ/UTQ
qmMOtT5Gry0a+VOOd+eIEd+TGEzMmR/tr3IQXlVeGAI6iQWAOxJSTLky3RXIrFdm
wfOBGBng4gFj2piggSV306W0nVuokUC5jpvKsd9WHLOs8/GiWJIt6W8u84ZkGf7i
Em/te6RTv70XVASNsh8r4+WLQOHQEg6oeyw3z8A/dQOCy5Z2kgrwBNRbGQKPQIga
OwG7o/tbk2/V5rV9lIYa/zDsnawhXMvLfPeAZKlbLOjra8s9rD7b3KQm0u/5NOYF
GxbuzkQiDiS05KFguB9LquM3tWcEO4LlJRwfEf7VZvPnQwzW84rLVSyY94wbycFY
/8fpTEapl0QIWcWQkn1ZSRMuJv540mh4H/xrh8ERqHGxkF+qkacllYkwmYG3tQtQ
zZI7Lg7C5es1TI8Vl+bw5Ngn2v/SzWs9KMRdlyj2OX45Fq9aJ8GnYDp4x5rrWRxw
EO/tdIuGIaAxxAT5b557zCDxvtL6JqgqJZ4WsL8qFC0/zWEcZnqNAU2Lo+wXeyAA
smWePSrvk2B2IvStf7ZAAkpZVLPaaO1Vypk8Ks3MF6ki36f3dCl24sYYK8X+K+DT
ohjnsoFbFqkRSbq9U0D/vnnod4pVljpjhazLmI9SHtQuRQy5Z+G2ll/vk+kH7wzM
QKZnef93dMxxnfOTdSEA9bWCnopiKkPZr1wkEV0T/4Y37w/yWwW9ZYBPaazB3Vq0
5/orsSe/VoAPNRZgt1tLFf6YTfLKwnHGEy1KRuzgyk9B1vgkKAg0EoZWzhXlyJvR
ROKJfN0t+U6ReuX3hHzYWIcOVcQYIxUoImEiPhX+LF0sAHXyBa7ZZ2l9qpofKxx+
KFUY+K0vE5ereFMIh8xdU3WIYI6v3xCmEDRDo/1oszRg3hchN7ZdNkE2rfm1DkCo
3n/OjcBT+9Rlb2NNsWCL80pfNHuItxwlMLkpJURTFlCCWXUvo78zuPBQp95SD17f
G7uCgnTcLArPKVyhS0uAEDH/zb5gULbdt1Xnb7MUqFy+8L5hAouRf3SpzAgEnkUb
ips1y8jMeLLmyfCAAHDXvMJR0p2rGNveN0E0BOKQUjqmu+qB+T0aIiLumGbqFykb
JAvJWvPyrQ2P52ejMzormiiNzrk0CXytr2JPkQR+wKJFAaY4qmx5xKYwWqTlQiDJ
ghi30jcwLhwg0aXbLaPmfP88DWBedvY14CucpSmiiZmdRFPa/UrfXAQrXod71pYZ
i9FFGfNno2wsXIsr3aEiVji+MvRaKbKibfIz2y/5vR3QRk446K2O2csNKffCbXOZ
3jjzYU9AgXjHY26q29o4u9nXq/7o1KmE246fLa2LmWUcCFLkxQjduCchtkdReyQN
AmxM0ekorWyQ2bRM09JqBJBocNqP1FgkIzNOVh5oc8UnJcTwJtojqkEVsy1FCPOv
ATRcJLM7AgsUM55ToXp/1n1VU5N7QGPDgaljZkQxVPE52p6WRyKJFpYwXy21b6Ck
PrCeMapL2iFyzuByC69dqBpsGmCTYu3ijfVnFsMw9G59LZaRzeF1J5i5FetDZG2y
pcAusjJOopQesB5EXQg0w+j9xgvBuDlaNpWnSJie6YgADW17eudpNPft5/7YSHdP
mVk6aSqnhK13P1V1R3QLb8Y09SF8U5t1+xPtJZr2SY3fjVrCiEraBcEHkhrvUNUn
tZXMUzfkOMBSAHsveG3qrEeLa4JManSgrBC5D6uJIgo0FYsm17YXAC3X9Ic+zV1A
ezEL+yuiWQBK7S45IIUOdFituk/z+AdxSJtvxZHQnU0rgZGwLjTaD+4mYloXWMWt
IqtZ2RtrcMbsNLHKHWJvwgleH5nBR9o2NjsGux28+6cEgKpo1liLkF6Wbu1vSJwE
s09FPt6zld1hTfe1WmMfQXRKneic0bFho6jUes9u72aT2wzR0B7mnySV7UaqBS4L
oLOVNkW7HrLIzx7zVQtfyKEUQ6AmZVbYqDYUn4suarN40nzygaY67qlPCPhQx5Pz
nBzHqx7oIpAlYr7dQc9N8g81srd1iW5AJGlPa9wCrWpWynOns4bj9Q5D0OZxGjsv
pW9zOXh8FgQbeCQqp8cJ23n5/5nNLWbGYW5eFWeqayDQqWU2GcVydMDWlNZiiPHb
/OjBGtTzlYx4PPbR3V3KRzWR7FVqDKacJS8//OwqkMZ0ObK/eMr/H2TU76QDVYlZ
lGGeb/Q4ncAOsGyLZ44HLMgzDyXgNx1V9MIon9C0/59clLY2wyPm/hJYwnQY9QoH
Ai2hXgSua/3aiV8Cgy+gMDoxjReDQUL/9cJCQjNSP11WM05neCEYtV/i98tQ2HRS
t7V4WxsD+A6Ax0nB7SlLCvHLSZuh9Q2+gwxvv7l5Myr+geax2Zp516tncFwAKZt4
nDxtP1mLpyJ9NWfybwbqM3BSmNwa01yPXTKAfJTdbCQR0JHQkELDMUIvWXPK52wu
5kr6H46tqJGNFNfD0+fd6BENwrRxcs28qmmAD4koQVrEoPRjBY5xitPaBOWkcjdY
ZZgktED595ksAiyaqHFGP3Jw45pnhIWYeBCuPkq+lmM5AhLqfv5VYBPyDoDWB9Bf
yYOtOROHZibAZbaI3fh4TIPQubbReYNd6pTBnB/gejHQzdyHl1kSIYBReXQN2mqs
GZjA5gWxXv+yQALCFJoHsRqfy7ql4+oJUUePOP+PKt85QDQDdK4UmDS49qaDC/u5
5WPBEywTfJgiloaJDJWfBTSzmCRLobNivJde28AaPXVOht8w0gOb/E8bQHyaGhWe
BLTHczfGAIGsv+eOc6i3ZoAm3m01q8lLMqKh1GS5CcgVw+eQeslSYj6Fcy8BoW3H
gL17PV7qhrbguSsfM8y4KqiT5jih9q9Ynhvw8ayr+k9D+YACQ43J43I63ks2KA+q
xUlHMFhROoQ/3QYXbMuFKlzclPCJzUXHaUBj44M+dJhnOoI+LJrYHM28XxwM04jM
s38NXGb7erWTsMZ1WMueZ2zaKIcJar4mmpuQn1MiHL6/74jarX2cozGrgaO5pNUQ
fuYy8upJW3iAq31sa4k+94F45mpmD+8jyZZdWHz3L3iGkNz1lpEddt69PHQ9eyRX
qkijTS4sVAG1+RoObJnNYDUm5i3+oALKW5GctPmdspRDQzJC+JqeKT5lXbRtUDlp
fod0lnTi3bOxBP8Wq81hRrGBwO7PqQ93AgRFaBD8fCaLkf75f9Wbt8aftkkZ8anR
KBBWdVyDAYTQ/1STz5HhncBzdJBdb6bRKQjM4UJOHOzvL5+XgOCv3zbcX7SAxP0W
zrV7jdmGezRCljiCgbyDnF6jj9CHViLmgo5ONi2etI2MCvFk6x7lNyfoQO2dwAMj
Iht0b5t8uH3R2LY788FA7kcwJp+bp77478osXNqPk/UsZPJzcFQIkUhTR0BEowm+
4+/zg1meEX4oQ6cTdDP05TqrNXAUP8Zv7TSK850qV1VAXy2y+MrAa7A7J7jTj/eM
Nf9JxDUEzFNTBABMeEVQNnfaFTzomIc5NbpLZoJL0nlmsaSkkGUkmOLt8zJm4+y9
N4uC8ZmNtapKPea1C1RaEfgfAiiInHgpitamXYlkJDC4xMQv9taIlzcEDvbtNJAo
8AL2sopMCsl93N4a0dMm0qRpv6tlnLwXzQotT6UAqQaff5D4tEyqhCn95wYr+Tnv
wb0RTfzjNrWmXb4tOPUvKZ1PNwunKXcEFNZ0wcwk5z3nn7bM6R0hv9CCjt4HIgOj
aK5D2CtNw80yXDdS6S0auJ0M6QCib5fNLcTzn5c0Emk3XN1JnZfx6qPcQSuXr4sR
365lGn5JOol93v/lT7BjyztP3Szp5ksPeoA3MGhYHmFft6a/sfTPJNzh63DeXak/
yeZ/co2M/Kn2+BSddOlKKYONk0Hy9d+ksG9iLuPBnpnkv/IAj5kMqULap/3yKwB5
ygKoW+d/MJWLIC+gYyJuN1KSHj1tKv2H+2R6v19jOAghT8c+f92cRz6lKmDjHV8H
3Lh0UjKUqxETOCXqGt2tVIW/8mCnJelBXcvvx98+Z1DPMxlj0PCZZQ6r+RalHkvX
1S6USrhl04t1djsNJ09fTeg2qXwL0HsfWcqnLL8eWZ826rJjuSNp+b678cW9P0YL
Vc7CwFUfb7GzQY3N5DSFYD7sJGpnrSU2/qkrBBTXO1X6yjrofT02N8e0GUpFaE8t
XhJTtnAMn/t2+eIwDZVD7ZptwDKn+wDkdKY5mdwO2nWGiLuFbW7qaleOU0IZC2Fw
2gUVai9ZsnMw5H4g02lsYvcYfBGa8OtY1usIjYosAIFy3nD4DbudWGIambaM3rIJ
8rXZeXZWt2JY5vf1UXKu6rk3Y6Xu0Dy+wg45Y2bDhbvuApO40MDog3xTgMeBa1Ev
KdcECkt3aAZpqBV9vhTzYhhEcq2uFZnMnqwsbE1cZm0SKvrOWW32ckA5kbgVo8Om
E/iwMEqahGfTCVbJjKLZfaXNBLKS5Nd9pSdluxS+pskgHC5Rfc3m8Imt2ALLX027
+kqZwXzMuQsiLqceEqHQbQCTT81tf78jBKhYSaT6LkO25MRv7t6LwCDCWUqs/+lk
bPvD4BSVtuA+MByndfoBWDEwFBbwm1p52XJDf9APU5IsDUA61eMyLpVfaDzyIeEZ
spHWOFl2QdLt6XIjDbi5oH62agN5T5qUKTFB2seapjvGueBk73FeWM5ITb5Dl5i1
7dlx7ahiaasTmPNdtKErt/zJMJCTTgvyzDyootvAPCbva9YjtDHlcg+Zz01uK4Hm
KwfGknT8WWs/sroAv2m64EtDQc7l2xcBC9ed/lEQXK7Q+j9fJF2ksHQ19Q0JAj+h
/2kx+puUwcajvWf2hSHeMuCxiMidxSON/lgCYKZyv7RmEnbzPXoH4pewBHa5IieF
b2T4W157MIdNvXg928CMClclNj81F3mBHT+qgjiqe4wZlKOPDmfo/qwBXA1EIfbD
ZkwwHkuXhfdIBXtyT3bzEkUnlY2weMn0UxWkrBoAcYEx/xZUWd1ZoZbKlWbBSD+e
GjOP7xLH1WgdMZhuTJdQdKlVQiB+zFAiygGybgNrQ3Jfl6b7b9vFSGAz1e7JpZa8
75IbKt6jheyedaZxE1S1iPbOu97+t5zOi+Nf4A4lEdp/JFFU6c2kWBWGK4pyxa4c
pCg3WjcJgowBfZYHgaK4OxeuI0mffiBzCcr2D4V7BGJ4jjiByyyrf8Y08ZIzu4/1
rW7t/G2lwMO9H37emfuoHa+ul0RA7edNqAPv+BKfsOU8lc2Z+u29lhXvzk3X8Y8f
alINQFcpvCITCGrepmRS80Q0IvpNgRWo4dFkT1k5NgAj64KGbtLkz0ilr1d02YSr
wBALtvQNYZT8mo3Kh/LqD7ubfHbV0B5XZu8I7nxPlTYUjZSmWkRmbqKdQSNStvHZ
1zAElMFABtJeD9SQb42gPO82GLmnQc9DdlgQkQRNLTpDUCr0kmPNN3JPWyKsh0my
IlgjwKgj1kyxzCoKMDYYpW7lYQpWF3EH3wF7YqMa1pIzMS/+7tvCtyCp9S4tLodz
Zmb8sCTpSwZZji6BBhIqcTRDSnn1XwnP3n4P+aLjzxlq9oJrFje2VmrlWnjsl6rL
HvIKxc9IoIzFJi6LzmYQVie8tQP2HMMFrKIU11Gsivb96eK/SU7en5A7UwduuZjz
Cd9rzMoTDEULTczmMymxBtoxFWQbfnQpsJ4YSO+eV/vY049U4j6Hk4vk+xlAouQU
VMsXnKTid/6jGkkLMub5j8NUq8p/WYNsQz56zFtm62oG9qe7EwXwF6byPfKPzJA5
cQhkOQemJv74Ad09c+7RWbtUn0mn5u/120zyC1JIOONpHLSXTuopeAdHQJI8XyZ4
LZBCxB61onDHs6P/VZEshqqvy2j6bc+v2Bktm1mQenypCYUVwkpl1p7a5hyxxCle
ild3WWuSC1wo/ld3v4HNETiCNnGID7X6RCV+USU4hGAxDvYiuItN8HsLdymFa8/v
SHtjv+VclX5CcmNRUyykkB827MhbqzFalwzYT2LfRmiDq0RlXmvgaH65wYXwhm1F
VHu5lJb6m4wE4nIv/S0eydvxOYgb0FpbEuwHbplPQAoMIJ29SSykidcNjU2f80ma
l6wxaMtbkF2HX9jnZQXY6GbY+wTcKEEdEWiu1t/NaY2GMRcl/MIMfHdBJao8es7K
mgONpjLOE5pU3gqmVs1/s7MBtEHNQL6jDGsbEytCuE0YQZpKzZkg708s92yNqXKk
ZYKUfDWAFo4yhw4OcFBMEb6ICz93LD84dJ8x6rMaiisU9CGX+UiWbl5efcLZlXn9
2MdleZ4Bp+s1qG32SS1tImGQ3V7w3q2z6nR9syWKUQHUzjDGrfaavRFJxWvFLCAs
ShVq3U/dB+tzVpvMpRxe7ULgL6hNO4dEmA+pK3b7JtJj4l9d32rY5b4GiYyx0HiT
qD6eYUMvOEVz3KecgrNpSl5enGz6UPWysUhO2d6gYqVkrCd9ujUIkiY464XasUQx
ars1HCOL/rM/wi7pPyH9xLSD/x/uO7tOzRx8xl5mIPeyr48XPxWv0n8Iosp3EeQJ
Th5PuXoKUt8fRfVyQYBqi/sOcPWMyefWzCXvrYvF6iQrG4y+mFDyMTp6OpqtBqca
uOB8dIimyiltt2PhdyqDNbTb+5YcDeUP3Chd7POK8ck5qROYqYBb98BDyGbv4TcK
OdLKjz7BrpdE0ASCzOmLBg3cTLS+noj7lft5v1FLRPdMpnGG99k/KIm8DSiVUv+3
CH8Xb1vMkMQmAeRYK1vjlfeBZVUq4WyaNZortnb46ij7Em5XXlMkbtSbJDVsbs3k
aD8Z3udihffSNCZOIHmbV1N030MoJ6J1cSwzC+4tPhJ8NqB4G13U7QmI1/rYRYCR
J6WhEu7yX3O4kqaZvlNZGeDlFGkqn5x1ZJvEcDBsQFQ4vpHHtS+TlRrbxQx/lCiU
SKNDXXH/mw+Vj0RDlFMKdLScR9ImIIZ8wSydZIrpc/AfILWtRwvC4hX6JVALLEUf
9RxRvL34QFrsHWN3dNNUbuB60RbXUFI4809j4EJ8DZ6PK9XGaXFPmeDRs5VhNeO8
dy+AoVfVdjXIoK8NdcaiW175/TTglbTkuebeG9GMCfij+nmGeRSs+MoG+vpYDSHd
StLvyQQEr59nwpARPh3OdHy1RQasnwltu5mNGrzPS22JAywESRZQOkIiU0lRU/Ca
W5xokR2VTnDzXHDsCYJQauQltC8Dwma0lbQymgU5bK2wPglt8xc0oQCNKiZyHT/l
dQk5PNkYy43pIqueDv1wgczMvrqD4SvPhGNDMpqQCG4H0emlMLMJ6GUwAhK+/AVX
qLAADA7xGdiTKmmS6DS8q0MOIZY0GgN8msH8h7g1B0SzZ3zXpf1MRpKe9ZancnQb
orpXB9yLLQFEHNN1W4SlhdjkoY0yKStUWhPS5UkZMFah4fBKpTC3A/F5z4mLkKfq
YgLen3cVwxXYvXCMUcA/QDSADwAa5fOdLLRtvu2WTg+roQS6NffbjMNS7hkTAAbU
cB+SUewk31IYhRW/0OutK5VNICiegkwHFymHjk31bakhxyxqqpxalvB+cAffm0UA
kmMwItRK7lIYIlp+2I/LbKfeG+MB40bU9I74LvWm5U6dbl7YNHTdb9YdtGJPaFHG
Izx4EKPGHEcpqS/VRFSISBqeCHIBYM/BMYDUOC+uBWstWayY5/Svl9M73u5iljNx
wpl9SWIM4AetSyzKP9IQitz+for8Vmknt7P48rDhQYIgRn/S2YlWQFqiywSPxZbg
a9tAQnbb7MHejNaCH9BYjb1gmdLTjsF5Bw3xMr4O3Cm9JH4LIS+BgS9ALvDKfViV
asY9yXgT6jCoWJDBACbsCdzNp/xhQ/VzS/EUB2GeHZtkQX081roJorVSLe94ThPZ
/4uwMaBcJsn+nq8BjBGLRGZZR47hU0s6erfuAcFUv0C6jeChvap8B5yO/1nGRVwM
TZziNbEBDNX+4yTwtibW44EBg04v4wbVJ+pktQzgnBrtNhgPyZWHb8w3O5zOkt7G
AZo82GMA9Qu6bvrVSi++oEQzorVN0iP5+Cxt5kmebq5qGwzJdNalbowpwa0o6aB2
besnUXcZ5o8INv/LNZV4FJ2O67ALq8tUJhRAIYVLROc8WY+zrvnbiIkMutWP+noK
xF0eV2rZseMeoD6bHE4d5YQpAPev7zIVBAtrkgkH+cFbFFrhBqbUSUlaewlkDcGt
Y7Jr1PpeNQ6FmoOCl2Xm8o10BUT7GUo7mjpK9sWscMenrOOi2WBr4lHP3OcPwbjC
F4hw3eFhkjSxUYuChehWjnwR5/np0A4uJGCdApLP9k0HoHvF6F9VhWQTBJO8gpdr
6HfdmZOXdYRXdY3McQaxtr6yz7uqB2Nd0lcuswnAT6Sp1lRgYKtI5w0L4gshPlbg
vT1KaDfVU2W0hmZLZ7j4OyPw+nYYEaxzRS/jVkzdcEcn4N2IjJgLb7LPcnNC5v70
qVcu8FwjIhatjK6fmysV1K7ni16af/fjTVev/lYZIzz+OnO+eqdHi15th+08q/Vu
1/rRZL+WoRe5j9impkWNh/kXT5hztAA/3S0fbwYZ3HPb6Drm4Ql2UPmIiQpAl3To
SBMYmJSuqdZWz3iZkaICa6lNlZeKkSjUcgOIm6GMkqD71OnkvQyrBD4auSKRqsey
9hwg6ZLx4iOW4vEg6fZ1HOWGZA1tCxrZbrfaX5UBb5kBxa/G4t/IvheqbpGCPCG1
A7gVk2l8XJZXkCGAndGUYRjcgYyYeiILz618fX+cN92WjnCKSQ2quycdZrhmIl5S
iPRyMrlk0Qe8woQAJb64Ulc9yzWBUHTw6p/Qw5CocWcaD+bZn1LvYRbZGoqB8iMR
Gpit5mymK//kZkk0X/1+RcnD7+fQAHbsM+B6rZmTHwSuSlyuevtTpeSnV6P41yy6
pv+mwxOE5iHcKIA++tFY7SfFILdqvNYjRSNiwPLQ9NUQv0VpwgEmhrNZCrYH3kBT
OF6WrKAMp9Z9wAqLf9fOV1uc37tEQizFDO+MV0czEjzfsN/Z/7qRN2bPeAXLa9Df
T6J8J1GL8UZx6inZ6wkDpFAP3lHCNO3aY0OX02hWgQmKj4ZRRRuF+NBiqvHFwB4l
e28gS2OBPwm1dNjuWrCHSMFe2CBr3cevU3SpYxRsCLpgxAthi+ZrEA8P26SSatFi
DAkt6+t/hMU3pe/jHJfFrcCzbd/JZMNsLBiqjQEoyC0o4wy0U178uCf7cOa6m0eQ
Dr42lNFVBOofvsWvtIgfBPvROYoQx+jXiyN1Lj3wpLe8g8ZG/pII3+ZtbcSpySfo
RLB45yM7iN1xlo98NPho+WjzEw0KMd808sFjShuKL3bFfgQnYXzsMSjnkI7tIsLR
VEGIC8Jb0zKwoGaOCi9LEDdS0gMaSIiJuRlTcG1WBnP58MEbQlTjPflGe9C4dy3z
YCKgoHQ7/KYHDBGEo7v9hFMYi0IsbBfoPMvykWM77ncxl8i/Zp19cFq1B3G7CwcG
lQGMVa8BmsqtLK3mtb7sYHA5h1nHgUv+edsn7e5bTGJ7RQ7bsYAikcueploM9XLU
srN/vDrIt12por6NTShB5Y2u39f9UzCBFOui1rK6/yf0VcFf+BUVRpwDFk3cMihN
ud9t8MlIboz/B9KJA0ArFI5jYa73l56epNEujUs5TBgszS2badsCAUmEjhq59R+y
gSgewVcj7MQqxDx2XxESx0eDA7ix0N9soTRZlGhSdjeFuImLMw8Oxy45Dq6z7xVP
mP+3JwH02J7SI2WscTPbIxF4gJzi8TOkRbUSGeBtoWa9sOiFJlA6+IEcwZO6biFb
P2ufU99kp+lxLFef1i2wsNCh089vNXBihZTP7AGYCOKZHanTPX9mvNHp1ho1mmm4
RHDSMQE2rCO9FaHv4yrmrpoECUZw9SYb7XBEn5BdB95Cq2jkDhXWJRK2BrllpsJ+
L3yIk1sVofWp28nh2PVZ1KujHmI+XcNxdt2FSyXKvsxjDYNRk9YJpswm/MdojWt2
4H6f8LxuUFAIGky/EvUAGGbAhlRI1WIFumuVffL/+9Dqu/xQnjtJRFxnpgwh+tzd
E0jj0ptG4RntG8IDQi973AHlSzAwhauDp9O6SjtrgNW6NQ9H371TuOZhz3MHoHwk
aFuxsylvjN6sSOgYJIKKQcHcopwlyj8EV8nHntaEU1n9YAZSVsWv50OT9KRrPMuC
thf+OWLo3fMcWqK0dPE/OHVzmKweRZyDDLthuuO743dSTdr19y/l3XKLFnrWJd9I
iAjogmb7mKwyyy7WpUbkawOn7dTmjVixctkFPiSDr1QQQOkXL3RYdjRN+1pWt+Ir
+fHesfXdJSJEzljkbaveKLllHeQYXWlcp/4jhhJlHnlNeCVs4x6cvqPMSREDiwqV
337hY3WZkW9jCyadVzSlF/DkgOzb8JyMt+O9y3qAVR3f2izWLO9RRVH/fU0I8ByM
K3YMofapNJB6CCOac4S0C+IKSqIAVj2JRz1zPpdrGXy2b56C5CHGSUkZ8k8pZJ1i
PWwyxlE7crjWQZr1NblYtfvRwPAxfnZNjaKowMLvbBHvku2+k73eRFo4YgAw35nD
RjhI7jsHoIC7xnUm4Ol42nCE+8LMpwTscdnOKEHkEKuCryvqED0we7QeQBq5sqd6
RsmWOH6MiImTHatqTqFCTVpPcbrJpLZkgp8t0TtvYfZcV4sw6mkaIjpfUM7J0ZS8
U0nMnfqecM4ik/xQ/pNJ5T1YF1bAzoyd6S96M0QuKni/N2pISXyRV2indn8szK0I
TkMB61j3ZOJ6cgFQNcQV2nIaHZPJFIGpfS9bKg/WG/IcCCrOBDegkATCb4QiTxvG
wavPI/JKyYrmEPB6MZWalYpTDfwC3hrJLwUACz9eaQX/hhUkJ8t3lMI0dlp+MKLW
x9UV8uVgcAeKBtJID0PNuvurKYTTCxIxP4TuSXvqKwBTA/Xq8USZTlAR0xy0DXUo
8CT2YnoJaRamZK919Yt/MXTjFKG3dpZLusGp3S6qqEgpWjNqgPw4JZfOBYCpsNAt
TCGSWvTzafv5uZu8TyQk5M8UkS+BUMWBrmc8A0FUOKfE2NvKjL5stjsENgWnLZMF
0F2lpqKHFHpmEhWiqBFIl6vp+3iHNoqeuY8zeqPSnNmvC9XtLIm8EFrNHD9fcoyq
NcePyCq2EE+5sWK+2xsTHtU21tJLY1O7vciPldwn6WJ4sxDUbJv19JIGHdqF144n
qh7GaOB/McHN9zEruKucBciFPIoYXFrCd58sqXcqraX5cL9MiclTq1wnOy0XFMu5
qSvDNHSrfJGapUa0iX9a8gSkSHtYAC9BYhplitQ4tBuu+PWf1Ybh5vuOeYLVQalV
8twZcU9WYMCDAPo3lCoWMwQi18gcVJyiRfOa81sZTmwZUBovPgKbHmJt+iNk7t+K
AFOH7MrQ0BGpSCmg9PNHiLM4Cw5XLqJRCzs8EBaE0evzMQOh5cZqeTGIhXgD6Iz4
DAEOLYAMgi6PAa34SDrxGhe1Ct6l2/0L5MFrxBu6s09mb5/5THRtvdyUNWAsVP/K
cUmVgJ7czYTeMCQSUwu37+n8/xdU1wWKlDhVsPt7tCp5Jq/53bZgGRiJjwJFkCtK
hbGjsR+u2gYuljACvHXcfqBKjddpumRrmb75sQt2n99x4lHmC898K4GcgtZ0KkaF
8R5qRjPsta60hw7ccBSM9MNnNpa0Az6qvmX1VgMNstrreH1p5HnsBe1oamewWhFE
v8GYH6BtAvmkbUShkaR4pP1/tsFiVQjSqU+kj3spaOs+cPQHaIbpBMKj/XyuWw7X
4vLtyJtaLCh5oK6sB9VaJNPSRkCQr59ZSI6mupmDZPWoglGd9YJJtf9YBU4p5oBG
H4jUHccVIUOZIoX6AGwgVnqKsXDWTTBJWq+lU+lP8Cak5hCqnaxlTudhs8YXa0Qk
+9QtKLTSUkOW97c5/yoEz0UqyybY10pmCDctr/xQAWy5xlesM2UPmiLsjWM4GynF
RWjKV+/6rWXAHXmOMQ3BjsiZzSgUmcvuJW2NIsNCr7XcI28sMQ7FOkHBkoB8eqDD
BqKE3Kb485i8NVKhuM/MacCyNdLdShqSZsCMTzN7qcpMC4cefRbKtnPrCdhntrqI
GFYkHAmMo1Lfz0AV6UuNKITFWlrywo0L1GykOQxQ9KQrCUxiRefvI2zOBOH+Zxyn
H6MqlhXiahqANYNvbnC9iy4k3KmF8xqg0aHPA6o7Ejpu1v+6WkgvcDN09tPSDVUM
Pybsh/74n1PUUHMYw44BoK86SbHRUxKPCctlQduZASKBlmwL7tE1MBM+eF5qrAhh
H0Mme0HzLNuQX5MjRhroKgC/8DcN+CxLYNE5rlkcjcp2riwOFWvBmI3xWQRBAltO
BjGKVR3aTHHD7RVfCkfqgpYiSSnyHhzoIkkmuqsCu4ch4WcsvGEufomnRBa6QNL4
K6K/hP3S0UPEL0niabJw4Y3osDUBLudq3IKRWZG4jv5Rh/9OM7o8Da5RaKtK0XR5
RwNvwCCki251nHDzJY0Sz182SQFDVJKVz2mcliMviqM4d4emm9y9H3pxb088ng0J
5NoLkIcaT75dnBtCcecpfCoWlw9P59B7yCYRVfDx2CaMk+MLAWlg28PeOHCZM2bn
JM6EACpHqaCQcbG92i7jmJr1IazHZzYfVBKQ2EJsgtWUTyP+z4Wo7OG5r5vTD6jZ
6Q9Mr9vMSYa8kHQDRleXPBxdZykxnEcxbCFuv+utq6YzxYDQRcRlKw2OkCroGM7M
b1kNyALuq7FyEwEqRSSoeW7rBQnH23IoOE+XXliFtjj+YMAnd3IKboFzzW7r84+r
wb0JYUFReP+dMwM07znFTVcvPyxlrqNkA7f0nrdtUMlILIUDEbNedrYIrZM4ubLX
mKRBw97JhJ5aGZyBqJ8oldoJe3b7EXJKCoPuWDrRzXvqkyivaJfKHQjS4eotJqkK
K86zo+wMep0TBfK0Usf7PF/NJ99iRrMYBO7CV7MqkB/NljqniFR3Duq5DxzyThMa
bbVtDSxB16YN8UqfNKd4eMTJTaaNYGanHUZpxfnW5WeqfO96lJ2xPhq+XaH7hI5C
67cogUq/jMg9oR52aqocVxLRWa40FwRrOUf4CLHNJ3HkVqaLs4n7O0yQ0t266uFH
x3j7MYL7pBVrG5pP45MPB+IVP+rCGsnIAFU1CwAZQmX9EdslbmYt5i5shcFU/WuY
dD8hGprFhssoxZawtZUkpDTbfUeb9jGPaUHyK+1SCVhSzpwU4WuyYz1CAMSbeOJ7
+AS8OLdcAarHT8IfCS6M3Ls1ApQMlA9nfTIjToefBUNFKanm0pH3NKlCynFTV5KH
0QgUSiltfGryxXNhx+kNSqP7Wn5Egz21qU1idM68+waYwvI2Y02SAmfJ7QWAf7TJ
YQZgBob3mAiXFFAagNHbOKMc3G/c94vrO/hAqu6szqX9EVmSflGf45D9jT+lMDgs
ggJc+BjZ3be4zNp2fR1KVqs8/jrNIuIMCIAGKz/FPujLJOrTb9bpwpnmZOehjmcp
rm0JZjBuiPloEuA0whAqku/o+gJx0yv/PdzvwHkqOxWdWqMce3b86un7Dw51gk4O
uKL/LBODF842aWPtX+sAlzwBkNmymI6bQI0ltxhUMq0XHE/8qNMShWKg258zJuQa
PG8vY4ttB2tHQ3mbY/Ji1NTDHIJyo6Xad4ECmaysXMlf4ALnmk0YiRed/HnjXEqD
IVz7blHjDiTj6b91WwwQbd0VwjjYts0E6IVLYzGOhyW86nt+E8D3o28dmaaCKBm8
RzX4feBXoATU5VFc8zzjWi2Vrts3pA07oOhkj/RGqFSu8Z2Hg2nlzj/FBiaAEObB
r2Z9qsM6Oezk1irKZbLYbN8k9dfFRjgK86qjMKnUL4AvmAsugF7nIJy1It0nQLCa
xyjVCazeDfITBIPePCyQSmqFfbZQiZA1eBJHFnx2MzFgEGyNKaQEadnOhdY4IKP1
BxGH1HjNiJ9T/HGNtcUSUZV7JpefKoIzCxZRxREMzbo1Lg4jbL3jgTVCBivymMuZ
Qw8c7t9JOCHYSnNy44Mr/4cWApn5460eYVrhfjK8cFMFxW438B2rT5MYPBgdpDCr
sTxdSnCNvuaUs+BZniDuEuUW5g7xh0Ylm4Iar1i6pmddRvxWEuFCxhbVr3nJYxh1
hPsyIxB16F0HvFtDUHpfoNcuIHnfIaTM1j/HQv+HnMuCC3Z8wELBrLQPLBxWBCiP
92ls5L8O/lYKFHznF/AxHScb/CRyg4FLbOjMWCcFigF6OrgZG59CJccf1oALiz4Q
vYxNbMKSZDFmX8XpJykBUR3/P6XSUnh7r9MJb5TXNMqp2csOzC2+rzsoyBrnIg2d
7+zaxYE4fj+88AqKJWmsALvYQQxlHw4ZP+qWx2Kyw8xmk4ogmSuWxXgS+q7+sSAr
TpOXTD0mfpAtL62gES+vjJWJz2qx5Pr6bGkMLdgrt+iDLFHGyBqNzd4D4f7ApTVo
3iIwL5q6K7oGJ6Iv6qLnOMV0Di7d3ynwntuQrDJ/UdYBH8gaHDCWOA3KvtFSAQIE
9ESD5gs1PS7z2+XmI6OvKIfZSp2zf/c7sr77fsUCjuFsip/qsZZstvVHnav1Vi+q
lNS9Cdu/GvBlVdaKipE5gov+uWmExua658gvX6sfrxKqWw5AQxQA0owckGd2CtVR
JMQhG65d/nCTOp2+bPw6wtLewcogFAr6xnSwRMA7W2mTC85r0GgOJ/B+meu38+h0
y5yYCtVTkc1a0B1zSZD/x3Mp8H8LTYx5/18YEDATaxjjB4ZhP1ZEdKR8lDzqIo3g
+cfVTgZPAC1tAKtt17VjQ8CwRB/bGjMlhVFHejHONMawvlwdgIKNpJ6YfHo3lMHT
uK8gQUCmk4DX4oMpgy/zJCJWsEcUY2Xwm512hoSn2XbkvZd+w8wDbNGAxN/ps7tr
syyRT/7mf/cA93JfRbh8GRcV99sBFzrZpczHnxQqPjLUR/D4RBceHwY1LScMX4ub
ZMQZyzxkK0YgAx/x/U8tKZL5vowNk53x5M6+dBB+hj5KlQB1QYGE6E/ew7ql5U2V
BE4aRA2jeO57/3y3/IYGxuudT6e2c2hS+0vcejJA5UTPBRy3dNWi6/KYZhqneU+H
8sqklJQcOudHYO07uunqLCFfl1EvJOcdCDdZATQT8U6+P1qjcHbOUe8/XUI+48Np
7iKhWsaENhMF7feMDLmGHD6v5RCEratbLZKwpvcnrbsUIT0Pbaa4S41uOYoq13DQ
Xnda9rJFN6GER31462QK4LHszCaEIxlSKY9L1zQePxg2BnqFHYVZgXXd1oxtXJmR
aS5DOhthlNi3sgcukWrjpB2tcZ4Z/W0+v84p0qfjnr6Z7IBmoJ9q9n568HgjJ5BI
Qj7S6jDhXz9tPf39ZJ//SQyaAWUZx2Y4+vnlddJqkWP+tprAFQ8ja/vJmv11b4Hj
FztQnjREm/QX1RIbkTSq+w0GmhL54WdhSy1Jmh4Sr0ADTdzCelNe7lEcCtSAX0xe
OQAEyDjDmzTe7UsrtOyuQhOKwr514dg3DgWOUudD7VmFx9F98xj3y94hkx0aizUp
bvQ80r0MWveTv8YR2E6Vq49i9H9V7PcegszJH7sJ711MF50cACqfPlSnnNvRIcA+
IJDgCciozzz1b0vt4gxxUtUrRjz2piZkIuMg5colETBectHnMJze3xtG7uxKLzxn
FwqhWN3W8sygm/ylTYWmTO2hnMtZgtzXCqFB2HhS+IthMazEBmUbbKUBbmkqma4x
7n1xB5UIEEGRY5GVJpcHgfg8XDbg71UPzEk87q11mzq8ZHKo3EBdZKTPavBvAp2I
kKwjvbJ8hGL6lENZzICVH0+TqYZEsmL4hSVsqoAUkeJJbf2G/xFo/rtN+mOhp7/i
EWMRqIPbwFxYXm32OFlcxth4qThviFDmh5gym8+ooIb6GvyXi2JCn8CPIea9oqDr
x19TNGhNGObXsIh4QYjDMbgBEho4LOe5KS+hODSgrMH/eKrfCHvnQ//FGdFfOR3Y
ATmwF5CwfzPmxPfZhvTJNxadW2XUe96ND+6arGMmZHhQDXfaaxZi5CBs5wMlywdS
5Bw/xnqEHn3x//85s40paRvvU/I7ObhPeenyjUqlEL/XKip0VeLyz2KxbI0iK7Ey
kElhL6V1phnLwQaAk8d2dZVbor5Y16jeiygBrwpJzCSnaK1D1cHvkrGyKBjIJrLJ
Z4xcwHfDffcB86rO2hCAdbOnaEPH5QMF4jEFsPElm0+1oUEdfiLqiARSHcVpD4V2
F+SKuDSC2kuxo9EYc6Zv0G9PY+bG6fLKUhTvQpkuIv9YmqAjRwptCRaDPYTlth61
rRbEOgHl9HtVlvZ4b9iUwqltWRvbcxCUB6q/9X+Y+0Qxkuixtq3MVi+ss1y18wT6
2fu4D4KgiWV5Ok7viIv8wYvudkB0Eb8AEUNybeYPr6YPxTLtKLwcuSq2wTfJGT/Y
e6TSSSkf3fXkj1KepJB1LPTcxBthIe/DpqWb85eEPFZss0kT2tI2fxAIeMUBlu0T
YjsjAKw16X804PBI9QXS2FgiDrAHIlnVRwd6mdQ/GW27I9EWoU09fyVNtgvUyycU
7VlHe+oGdq6SWXw0UxMajmR5akHCsgrKeBUDTCmB5GMTvOD1DLEoUoCJn7yN1cD9
n+pN3Y6Cid/JpcsPTcX+6OU2q2BIhVkzDuyiV3m9gtLdP7y1dUNP/IStMFI5wyIi
8/R61dSRTpthPGXjl6WEAL2+SHVovVHafXVFp3d/GxHF73hhW1URaGoJ315diHj6
fJVT25VoqqDdOYSgAiCR/TzaRE9+8eMUOBtNaHYLn93QJSbcgPrMEpogcQAl1e5c
a4n9drvDqv/YJR+PpN8aEKbVQhRdzs70vAIwhjwAsCP2l/GFt+yJCZQFBezot1/u
L8xc2vy4hi2GIUWpmTbrHWEbDJFcg7ahfoxvVQsiXbjyUrk1Q+/UbRficUOYX9V0
9QFDmdUWyNGUgAiVskHB7eaUVhiVv0NzZSBsq0W3eno/Ze9k7niunmz7ngZlgM91
d4JOF1Yy5tchPVOSufHdN/fKjWMI8lFi4m0H0O74Ue/ZCaFBbRAO5KcwZ5Li/8CA
xZj71Mm0E4+V8q8EjJj2/RrtSipk5Xqez4qKRo/K39FTPvs+YYjY74RT9J9A73to
3T3MjlOqydudVIp/FB72xOV1vCVP96F6aODRVjd+tA+8O+KIoBRDD+jUujvx7foY
M+xEIMZrgFH6imLCl5ACv8kd/en94qMVczsVX+k+AUgS22Y8ImPBiZcoBTK0i9mL
y6cgc4DvOo/bq/lkJhntMY3gxuqzuuym3gXXYG4u/H+/vZPH0k0s/K4ijr56oEiP
16j9hGPkUY8CI6qyhS9KQwKa0BGHKynchn69532rNXnBJZbmHBvDkB+a2IBEEl5X
OlPXQHALPC2aRN2HmNdmPWabD+zGrGcqS+6k5k5lZ8t3TUWK53Y+DHD6P5wPqmll
3CnmXRJyD3eukatmD1BCSBoPbJA7Cuijl4kZ+TMl+02zgiS4K+0nG1J/XurX1GCg
OxIKsMbvv46SBNyYIgx+IYiLYqpfF6gaEH57uZpGrRp60Ey05m957MokWN3knyRy
QiTdM0K4EHPi5bR0CImDBy5DFgZ49Emy59aYezTBMIyaPwKl8dCdVSTP8MztuFtD
f3QkiLnlEcFJFmuhRzWDmPb+fnmv53+1K7PFElBLhTBSGjYlaUb59k1gtkzOwKsK
Bn1ZOxgOIoZUywV7h7oLQkOYjJfQL4ltC+/DLN79dQnBiBriQUjqOABbqvkeEO+y
X2n7UTyqeHHD1yrz1fLxlWxy8EqmvLyFE79QlAPFdOx2HvSDSUpN7jnk+IpVnsld
NDYTaGIbhb+kP2d0/FlbhByEt9yN0dawKEZWXxkRozZsd0ArN675knWYainP7oJh
NP0fiEaFLRkKvpKhC3lkP9WTi/22EmLDUAEQJwVCrR2ZcXCeryL0NdOIc91N7q6Y
MEfz3n4D+zQUaKRyqXgI37lP/LU0taznVOhUxStPP8qeyo0bmYfeE3CCBvQUpUQ5
E0z0Om4JRkyNMPRVHu4Uuy14g28/GTYCs6PFkvcJz8upmZ7EXXYbEKZ6oRp2k+iU
6gjck+aPE2/IZ39td9dpYBfWGgzecaFbbWBj7ZbsUD8+/hjduK+Zn/d/Y6/rTql2
I3epiCg7YN1UGVFb/KorIyf5/dRIWCxo+6XS7D2f2TK01S9yS+2QpRqxBHEOmLEY
Mily+9z2M3NlOUqDJ4F6tAsDJW/fuyHd+qYj+fVs9uHsyO4grWBxpVG1uoIXMyY3
52UfENGYVsfEEv4jPRuJeMw0nqxsvlgQSKD33AvdqDmbuMKrIJvz85uSD92J9Hxe
aEaWHbyhzsEYP9qteAipNdapxdAAhgrM8OQLwE2vsIctOSWK8FRJ6xNuAXMx8WzV
N0SraDz5jQ455OWZMj5wMr3KSAggxm1LIrC2XLiKSt3k9XtddhB/52EjNhztiGIT
rb4h3Tde5zA73NLSvj+1xhudqmxtSdCWMPcM12/hH7a0L0Nnkiy9X0ZKxRtp07Uc
EbMA8IfVdNBS7lGylQ0BRA==
`protect end_protected
